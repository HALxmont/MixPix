magic
tech sky130B
magscale 1 2
timestamp 1662760421
<< metal1 >>
rect 157334 700680 157340 700732
rect 157392 700720 157398 700732
rect 202782 700720 202788 700732
rect 157392 700692 202788 700720
rect 157392 700680 157398 700692
rect 202782 700680 202788 700692
rect 202840 700680 202846 700732
rect 89162 700612 89168 700664
rect 89220 700652 89226 700664
rect 160738 700652 160744 700664
rect 89220 700624 160744 700652
rect 89220 700612 89226 700624
rect 160738 700612 160744 700624
rect 160796 700612 160802 700664
rect 72970 700544 72976 700596
rect 73028 700584 73034 700596
rect 160094 700584 160100 700596
rect 73028 700556 160100 700584
rect 73028 700544 73034 700556
rect 160094 700544 160100 700556
rect 160152 700544 160158 700596
rect 157242 700476 157248 700528
rect 157300 700516 157306 700528
rect 283834 700516 283840 700528
rect 157300 700488 283840 700516
rect 157300 700476 157306 700488
rect 283834 700476 283840 700488
rect 283892 700476 283898 700528
rect 8110 700408 8116 700460
rect 8168 700448 8174 700460
rect 162118 700448 162124 700460
rect 8168 700420 162124 700448
rect 8168 700408 8174 700420
rect 162118 700408 162124 700420
rect 162176 700408 162182 700460
rect 153194 700340 153200 700392
rect 153252 700380 153258 700392
rect 332502 700380 332508 700392
rect 153252 700352 332508 700380
rect 153252 700340 153258 700352
rect 332502 700340 332508 700352
rect 332560 700340 332566 700392
rect 525058 700340 525064 700392
rect 525116 700380 525122 700392
rect 559650 700380 559656 700392
rect 525116 700352 559656 700380
rect 525116 700340 525122 700352
rect 559650 700340 559656 700352
rect 559708 700340 559714 700392
rect 149698 700272 149704 700324
rect 149756 700312 149762 700324
rect 543458 700312 543464 700324
rect 149756 700284 543464 700312
rect 149756 700272 149762 700284
rect 543458 700272 543464 700284
rect 543516 700272 543522 700324
rect 24302 699660 24308 699712
rect 24360 699700 24366 699712
rect 25498 699700 25504 699712
rect 24360 699672 25504 699700
rect 24360 699660 24366 699672
rect 25498 699660 25504 699672
rect 25556 699660 25562 699712
rect 105446 699660 105452 699712
rect 105504 699700 105510 699712
rect 106918 699700 106924 699712
rect 105504 699672 106924 699700
rect 105504 699660 105510 699672
rect 106918 699660 106924 699672
rect 106976 699660 106982 699712
rect 137830 699660 137836 699712
rect 137888 699700 137894 699712
rect 140038 699700 140044 699712
rect 137888 699672 140044 699700
rect 137888 699660 137894 699672
rect 140038 699660 140044 699672
rect 140096 699660 140102 699712
rect 265618 699660 265624 699712
rect 265676 699700 265682 699712
rect 267642 699700 267648 699712
rect 265676 699672 267648 699700
rect 265676 699660 265682 699672
rect 267642 699660 267648 699672
rect 267700 699660 267706 699712
rect 396718 699660 396724 699712
rect 396776 699700 396782 699712
rect 397454 699700 397460 699712
rect 396776 699672 397460 699700
rect 396776 699660 396782 699672
rect 397454 699660 397460 699672
rect 397512 699660 397518 699712
rect 428458 699660 428464 699712
rect 428516 699700 428522 699712
rect 429838 699700 429844 699712
rect 428516 699672 429844 699700
rect 428516 699660 428522 699672
rect 429838 699660 429844 699672
rect 429896 699660 429902 699712
rect 146570 696940 146576 696992
rect 146628 696980 146634 696992
rect 580166 696980 580172 696992
rect 146628 696952 580172 696980
rect 146628 696940 146634 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 148318 683136 148324 683188
rect 148376 683176 148382 683188
rect 580166 683176 580172 683188
rect 148376 683148 580172 683176
rect 148376 683136 148382 683148
rect 580166 683136 580172 683148
rect 580224 683136 580230 683188
rect 3326 670760 3332 670812
rect 3384 670800 3390 670812
rect 164878 670800 164884 670812
rect 3384 670772 164884 670800
rect 3384 670760 3390 670772
rect 164878 670760 164884 670772
rect 164936 670760 164942 670812
rect 146938 670692 146944 670744
rect 146996 670732 147002 670744
rect 580166 670732 580172 670744
rect 146996 670704 580172 670732
rect 146996 670692 147002 670704
rect 580166 670692 580172 670704
rect 580224 670692 580230 670744
rect 3510 658112 3516 658164
rect 3568 658152 3574 658164
rect 7558 658152 7564 658164
rect 3568 658124 7564 658152
rect 3568 658112 3574 658124
rect 7558 658112 7564 658124
rect 7616 658112 7622 658164
rect 144914 643084 144920 643136
rect 144972 643124 144978 643136
rect 580166 643124 580172 643136
rect 144972 643096 580172 643124
rect 144972 643084 144978 643096
rect 580166 643084 580172 643096
rect 580224 643084 580230 643136
rect 3510 632068 3516 632120
rect 3568 632108 3574 632120
rect 164234 632108 164240 632120
rect 3568 632080 164240 632108
rect 3568 632068 3574 632080
rect 164234 632068 164240 632080
rect 164292 632068 164298 632120
rect 147030 630640 147036 630692
rect 147088 630680 147094 630692
rect 580166 630680 580172 630692
rect 147088 630652 580172 630680
rect 147088 630640 147094 630652
rect 580166 630640 580172 630652
rect 580224 630640 580230 630692
rect 3510 618264 3516 618316
rect 3568 618304 3574 618316
rect 166258 618304 166264 618316
rect 3568 618276 166264 618304
rect 3568 618264 3574 618276
rect 166258 618264 166264 618276
rect 166316 618264 166322 618316
rect 145558 616836 145564 616888
rect 145616 616876 145622 616888
rect 580166 616876 580172 616888
rect 145616 616848 580172 616876
rect 145616 616836 145622 616848
rect 580166 616836 580172 616848
rect 580224 616836 580230 616888
rect 3510 605820 3516 605872
rect 3568 605860 3574 605872
rect 166350 605860 166356 605872
rect 3568 605832 166356 605860
rect 3568 605820 3574 605832
rect 166350 605820 166356 605832
rect 166408 605820 166414 605872
rect 157610 605072 157616 605124
rect 157668 605112 157674 605124
rect 169754 605112 169760 605124
rect 157668 605084 169760 605112
rect 157668 605072 157674 605084
rect 169754 605072 169760 605084
rect 169812 605072 169818 605124
rect 143718 590656 143724 590708
rect 143776 590696 143782 590708
rect 579798 590696 579804 590708
rect 143776 590668 579804 590696
rect 143776 590656 143782 590668
rect 579798 590656 579804 590668
rect 579856 590656 579862 590708
rect 3326 579640 3332 579692
rect 3384 579680 3390 579692
rect 165614 579680 165620 579692
rect 3384 579652 165620 579680
rect 3384 579640 3390 579652
rect 165614 579640 165620 579652
rect 165672 579640 165678 579692
rect 143810 576852 143816 576904
rect 143868 576892 143874 576904
rect 580166 576892 580172 576904
rect 143868 576864 580172 576892
rect 143868 576852 143874 576864
rect 580166 576852 580172 576864
rect 580224 576852 580230 576904
rect 3234 565836 3240 565888
rect 3292 565876 3298 565888
rect 167638 565876 167644 565888
rect 3292 565848 167644 565876
rect 3292 565836 3298 565848
rect 167638 565836 167644 565848
rect 167696 565836 167702 565888
rect 144178 563048 144184 563100
rect 144236 563088 144242 563100
rect 579798 563088 579804 563100
rect 144236 563060 579804 563088
rect 144236 563048 144242 563060
rect 579798 563048 579804 563060
rect 579856 563048 579862 563100
rect 3326 553392 3332 553444
rect 3384 553432 3390 553444
rect 167730 553432 167736 553444
rect 3384 553404 167736 553432
rect 3384 553392 3390 553404
rect 167730 553392 167736 553404
rect 167788 553392 167794 553444
rect 142154 536800 142160 536852
rect 142212 536840 142218 536852
rect 580166 536840 580172 536852
rect 142212 536812 580172 536840
rect 142212 536800 142218 536812
rect 580166 536800 580172 536812
rect 580224 536800 580230 536852
rect 2774 527144 2780 527196
rect 2832 527184 2838 527196
rect 4798 527184 4804 527196
rect 2832 527156 4804 527184
rect 2832 527144 2838 527156
rect 4798 527144 4804 527156
rect 4856 527144 4862 527196
rect 142246 524424 142252 524476
rect 142304 524464 142310 524476
rect 580166 524464 580172 524476
rect 142304 524436 580172 524464
rect 142304 524424 142310 524436
rect 580166 524424 580172 524436
rect 580224 524424 580230 524476
rect 3510 514768 3516 514820
rect 3568 514808 3574 514820
rect 10318 514808 10324 514820
rect 3568 514780 10324 514808
rect 3568 514768 3574 514780
rect 10318 514768 10324 514780
rect 10376 514768 10382 514820
rect 180058 510620 180064 510672
rect 180116 510660 180122 510672
rect 580166 510660 580172 510672
rect 180116 510632 580172 510660
rect 180116 510620 180122 510632
rect 580166 510620 580172 510632
rect 580224 510620 580230 510672
rect 3050 500964 3056 501016
rect 3108 501004 3114 501016
rect 152458 501004 152464 501016
rect 3108 500976 152464 501004
rect 3108 500964 3114 500976
rect 152458 500964 152464 500976
rect 152516 500964 152522 501016
rect 181438 484372 181444 484424
rect 181496 484412 181502 484424
rect 580166 484412 580172 484424
rect 181496 484384 580172 484412
rect 181496 484372 181502 484384
rect 580166 484372 580172 484384
rect 580224 484372 580230 484424
rect 3050 474716 3056 474768
rect 3108 474756 3114 474768
rect 169754 474756 169760 474768
rect 3108 474728 169760 474756
rect 3108 474716 3114 474728
rect 169754 474716 169760 474728
rect 169812 474716 169818 474768
rect 192478 470568 192484 470620
rect 192536 470608 192542 470620
rect 579982 470608 579988 470620
rect 192536 470580 579988 470608
rect 192536 470568 192542 470580
rect 579982 470568 579988 470580
rect 580040 470568 580046 470620
rect 3510 462340 3516 462392
rect 3568 462380 3574 462392
rect 171778 462380 171784 462392
rect 3568 462352 171784 462380
rect 3568 462340 3574 462352
rect 171778 462340 171784 462352
rect 171836 462340 171842 462392
rect 178678 456764 178684 456816
rect 178736 456804 178742 456816
rect 580166 456804 580172 456816
rect 178736 456776 580172 456804
rect 178736 456764 178742 456776
rect 580166 456764 580172 456776
rect 580224 456764 580230 456816
rect 3142 448536 3148 448588
rect 3200 448576 3206 448588
rect 170398 448576 170404 448588
rect 3200 448548 170404 448576
rect 3200 448536 3206 448548
rect 170398 448536 170404 448548
rect 170456 448536 170462 448588
rect 138014 430584 138020 430636
rect 138072 430624 138078 430636
rect 580166 430624 580172 430636
rect 138072 430596 580172 430624
rect 138072 430584 138078 430596
rect 580166 430584 580172 430596
rect 580224 430584 580230 430636
rect 3510 422288 3516 422340
rect 3568 422328 3574 422340
rect 171134 422328 171140 422340
rect 3568 422300 171140 422328
rect 3568 422288 3574 422300
rect 171134 422288 171140 422300
rect 171192 422288 171198 422340
rect 140130 418140 140136 418192
rect 140188 418180 140194 418192
rect 580166 418180 580172 418192
rect 140188 418152 580172 418180
rect 140188 418140 140194 418152
rect 580166 418140 580172 418152
rect 580224 418140 580230 418192
rect 2866 409844 2872 409896
rect 2924 409884 2930 409896
rect 13078 409884 13084 409896
rect 2924 409856 13084 409884
rect 2924 409844 2930 409856
rect 13078 409844 13084 409856
rect 13136 409844 13142 409896
rect 138658 404336 138664 404388
rect 138716 404376 138722 404388
rect 580166 404376 580172 404388
rect 138716 404348 580172 404376
rect 138716 404336 138722 404348
rect 580166 404336 580172 404348
rect 580224 404336 580230 404388
rect 3510 397468 3516 397520
rect 3568 397508 3574 397520
rect 171870 397508 171876 397520
rect 3568 397480 171876 397508
rect 3568 397468 3574 397480
rect 171870 397468 171876 397480
rect 171928 397468 171934 397520
rect 185578 378156 185584 378208
rect 185636 378196 185642 378208
rect 580166 378196 580172 378208
rect 185636 378168 580172 378196
rect 185636 378156 185642 378168
rect 580166 378156 580172 378168
rect 580224 378156 580230 378208
rect 3510 371288 3516 371340
rect 3568 371328 3574 371340
rect 8938 371328 8944 371340
rect 3568 371300 8944 371328
rect 3568 371288 3574 371300
rect 8938 371288 8944 371300
rect 8996 371288 9002 371340
rect 3142 357416 3148 357468
rect 3200 357456 3206 357468
rect 174538 357456 174544 357468
rect 3200 357428 174544 357456
rect 3200 357416 3206 357428
rect 174538 357416 174544 357428
rect 174596 357416 174602 357468
rect 140222 351908 140228 351960
rect 140280 351948 140286 351960
rect 580166 351948 580172 351960
rect 140280 351920 580172 351948
rect 140280 351908 140286 351920
rect 580166 351908 580172 351920
rect 580224 351908 580230 351960
rect 3326 345040 3332 345092
rect 3384 345080 3390 345092
rect 173894 345080 173900 345092
rect 3384 345052 173900 345080
rect 3384 345040 3390 345052
rect 173894 345040 173900 345052
rect 173952 345040 173958 345092
rect 135530 324300 135536 324352
rect 135588 324340 135594 324352
rect 580166 324340 580172 324352
rect 135588 324312 580172 324340
rect 135588 324300 135594 324312
rect 580166 324300 580172 324312
rect 580224 324300 580230 324352
rect 3326 318792 3332 318844
rect 3384 318832 3390 318844
rect 173986 318832 173992 318844
rect 3384 318804 173992 318832
rect 3384 318792 3390 318804
rect 173986 318792 173992 318804
rect 174044 318792 174050 318844
rect 135898 311856 135904 311908
rect 135956 311896 135962 311908
rect 579982 311896 579988 311908
rect 135956 311868 579988 311896
rect 135956 311856 135962 311868
rect 579982 311856 579988 311868
rect 580040 311856 580046 311908
rect 3510 304988 3516 305040
rect 3568 305028 3574 305040
rect 175918 305028 175924 305040
rect 3568 305000 175924 305028
rect 3568 304988 3574 305000
rect 175918 304988 175924 305000
rect 175976 304988 175982 305040
rect 135990 298120 135996 298172
rect 136048 298160 136054 298172
rect 580166 298160 580172 298172
rect 136048 298132 580172 298160
rect 136048 298120 136054 298132
rect 580166 298120 580172 298132
rect 580224 298120 580230 298172
rect 3510 292544 3516 292596
rect 3568 292584 3574 292596
rect 176010 292584 176016 292596
rect 3568 292556 176016 292584
rect 3568 292544 3574 292556
rect 176010 292544 176016 292556
rect 176068 292544 176074 292596
rect 13078 286288 13084 286340
rect 13136 286328 13142 286340
rect 173158 286328 173164 286340
rect 13136 286300 173164 286328
rect 13136 286288 13142 286300
rect 173158 286288 173164 286300
rect 173216 286288 173222 286340
rect 25498 284928 25504 284980
rect 25556 284968 25562 284980
rect 163498 284968 163504 284980
rect 25556 284940 163504 284968
rect 25556 284928 25562 284940
rect 163498 284928 163504 284940
rect 163556 284928 163562 284980
rect 141418 283568 141424 283620
rect 141476 283608 141482 283620
rect 192478 283608 192484 283620
rect 141476 283580 192484 283608
rect 141476 283568 141482 283580
rect 192478 283568 192484 283580
rect 192536 283568 192542 283620
rect 137278 282140 137284 282192
rect 137336 282180 137342 282192
rect 185578 282180 185584 282192
rect 137336 282152 185584 282180
rect 137336 282140 137342 282152
rect 185578 282140 185584 282152
rect 185636 282140 185642 282192
rect 186406 280780 186412 280832
rect 186464 280820 186470 280832
rect 396718 280820 396724 280832
rect 186464 280792 396724 280820
rect 186464 280780 186470 280792
rect 396718 280780 396724 280792
rect 396776 280780 396782 280832
rect 151814 280168 151820 280220
rect 151872 280208 151878 280220
rect 186406 280208 186412 280220
rect 151872 280180 186412 280208
rect 151872 280168 151878 280180
rect 186406 280168 186412 280180
rect 186464 280168 186470 280220
rect 151078 279420 151084 279472
rect 151136 279460 151142 279472
rect 462314 279460 462320 279472
rect 151136 279432 462320 279460
rect 151136 279420 151142 279432
rect 462314 279420 462320 279432
rect 462372 279420 462378 279472
rect 149238 277992 149244 278044
rect 149296 278032 149302 278044
rect 527174 278032 527180 278044
rect 149296 278004 527180 278032
rect 149296 277992 149302 278004
rect 527174 277992 527180 278004
rect 527232 277992 527238 278044
rect 40034 276632 40040 276684
rect 40092 276672 40098 276684
rect 161474 276672 161480 276684
rect 40092 276644 161480 276672
rect 40092 276632 40098 276644
rect 161474 276632 161480 276644
rect 161532 276632 161538 276684
rect 10318 275272 10324 275324
rect 10376 275312 10382 275324
rect 169110 275312 169116 275324
rect 10376 275284 169116 275312
rect 10376 275272 10382 275284
rect 169110 275272 169116 275284
rect 169168 275272 169174 275324
rect 186682 275272 186688 275324
rect 186740 275312 186746 275324
rect 364334 275312 364340 275324
rect 186740 275284 364340 275312
rect 186740 275272 186746 275284
rect 364334 275272 364340 275284
rect 364392 275272 364398 275324
rect 153378 274660 153384 274712
rect 153436 274700 153442 274712
rect 186498 274700 186504 274712
rect 153436 274672 186504 274700
rect 153436 274660 153442 274672
rect 186498 274660 186504 274672
rect 186556 274700 186562 274712
rect 186682 274700 186688 274712
rect 186556 274672 186688 274700
rect 186556 274660 186562 274672
rect 186682 274660 186688 274672
rect 186740 274660 186746 274712
rect 7558 273912 7564 273964
rect 7616 273952 7622 273964
rect 163590 273952 163596 273964
rect 7616 273924 163596 273952
rect 7616 273912 7622 273924
rect 163590 273912 163596 273924
rect 163648 273912 163654 273964
rect 187694 273912 187700 273964
rect 187752 273952 187758 273964
rect 234614 273952 234620 273964
rect 187752 273924 234620 273952
rect 187752 273912 187758 273924
rect 234614 273912 234620 273924
rect 234672 273912 234678 273964
rect 155954 273232 155960 273284
rect 156012 273272 156018 273284
rect 187694 273272 187700 273284
rect 156012 273244 187700 273272
rect 156012 273232 156018 273244
rect 187694 273232 187700 273244
rect 187752 273232 187758 273284
rect 152458 272484 152464 272536
rect 152516 272524 152522 272536
rect 169018 272524 169024 272536
rect 152516 272496 169024 272524
rect 152516 272484 152522 272496
rect 169018 272484 169024 272496
rect 169076 272484 169082 272536
rect 134518 271872 134524 271924
rect 134576 271912 134582 271924
rect 580166 271912 580172 271924
rect 134576 271884 580172 271912
rect 134576 271872 134582 271884
rect 580166 271872 580172 271884
rect 580224 271872 580230 271924
rect 140038 271124 140044 271176
rect 140096 271164 140102 271176
rect 158714 271164 158720 271176
rect 140096 271136 158720 271164
rect 140096 271124 140102 271136
rect 158714 271124 158720 271136
rect 158772 271124 158778 271176
rect 8938 269832 8944 269884
rect 8996 269872 9002 269884
rect 172514 269872 172520 269884
rect 8996 269844 172520 269872
rect 8996 269832 9002 269844
rect 172514 269832 172520 269844
rect 172572 269832 172578 269884
rect 149146 269764 149152 269816
rect 149204 269804 149210 269816
rect 494054 269804 494060 269816
rect 149204 269776 494060 269804
rect 149204 269764 149210 269776
rect 494054 269764 494060 269776
rect 494112 269764 494118 269816
rect 106918 268404 106924 268456
rect 106976 268444 106982 268456
rect 160186 268444 160192 268456
rect 106976 268416 160192 268444
rect 106976 268404 106982 268416
rect 160186 268404 160192 268416
rect 160244 268404 160250 268456
rect 147674 268336 147680 268388
rect 147732 268376 147738 268388
rect 525058 268376 525064 268388
rect 147732 268348 525064 268376
rect 147732 268336 147738 268348
rect 525058 268336 525064 268348
rect 525116 268336 525122 268388
rect 141050 266976 141056 267028
rect 141108 267016 141114 267028
rect 181438 267016 181444 267028
rect 141108 266988 181444 267016
rect 141108 266976 141114 266988
rect 181438 266976 181444 266988
rect 181496 266976 181502 267028
rect 3050 266364 3056 266416
rect 3108 266404 3114 266416
rect 176654 266404 176660 266416
rect 3108 266376 176660 266404
rect 3108 266364 3114 266376
rect 176654 266364 176660 266376
rect 176712 266364 176718 266416
rect 171686 265752 171692 265804
rect 171744 265792 171750 265804
rect 176102 265792 176108 265804
rect 171744 265764 176108 265792
rect 171744 265752 171750 265764
rect 176102 265752 176108 265764
rect 176160 265752 176166 265804
rect 141602 265684 141608 265736
rect 141660 265724 141666 265736
rect 180058 265724 180064 265736
rect 141660 265696 180064 265724
rect 141660 265684 141666 265696
rect 180058 265684 180064 265696
rect 180116 265684 180122 265736
rect 3418 265616 3424 265668
rect 3476 265656 3482 265668
rect 163498 265656 163504 265668
rect 3476 265628 163504 265656
rect 3476 265616 3482 265628
rect 163498 265616 163504 265628
rect 163556 265616 163562 265668
rect 176010 265616 176016 265668
rect 176068 265656 176074 265668
rect 192294 265656 192300 265668
rect 176068 265628 192300 265656
rect 176068 265616 176074 265628
rect 192294 265616 192300 265628
rect 192352 265616 192358 265668
rect 175918 265548 175924 265600
rect 175976 265588 175982 265600
rect 196434 265588 196440 265600
rect 175976 265560 196440 265588
rect 175976 265548 175982 265560
rect 196434 265548 196440 265560
rect 196492 265548 196498 265600
rect 171962 265480 171968 265532
rect 172020 265520 172026 265532
rect 193858 265520 193864 265532
rect 172020 265492 193864 265520
rect 172020 265480 172026 265492
rect 193858 265480 193864 265492
rect 193916 265480 193922 265532
rect 173158 265412 173164 265464
rect 173216 265452 173222 265464
rect 196250 265452 196256 265464
rect 173216 265424 196256 265452
rect 173216 265412 173222 265424
rect 196250 265412 196256 265424
rect 196308 265412 196314 265464
rect 174538 265344 174544 265396
rect 174596 265384 174602 265396
rect 197722 265384 197728 265396
rect 174596 265356 197728 265384
rect 174596 265344 174602 265356
rect 197722 265344 197728 265356
rect 197780 265344 197786 265396
rect 169110 265276 169116 265328
rect 169168 265316 169174 265328
rect 169570 265316 169576 265328
rect 169168 265288 169576 265316
rect 169168 265276 169174 265288
rect 169570 265276 169576 265288
rect 169628 265316 169634 265328
rect 193582 265316 193588 265328
rect 169628 265288 193588 265316
rect 169628 265276 169634 265288
rect 193582 265276 193588 265288
rect 193640 265276 193646 265328
rect 175826 265208 175832 265260
rect 175884 265248 175890 265260
rect 176010 265248 176016 265260
rect 175884 265220 176016 265248
rect 175884 265208 175890 265220
rect 176010 265208 176016 265220
rect 176068 265208 176074 265260
rect 176102 265208 176108 265260
rect 176160 265248 176166 265260
rect 197630 265248 197636 265260
rect 176160 265220 197636 265248
rect 176160 265208 176166 265220
rect 197630 265208 197636 265220
rect 197688 265208 197694 265260
rect 164878 265140 164884 265192
rect 164936 265180 164942 265192
rect 195146 265180 195152 265192
rect 164936 265152 195152 265180
rect 164936 265140 164942 265152
rect 195146 265140 195152 265152
rect 195204 265140 195210 265192
rect 153286 265072 153292 265124
rect 153344 265112 153350 265124
rect 158806 265112 158812 265124
rect 153344 265084 158812 265112
rect 153344 265072 153350 265084
rect 158806 265072 158812 265084
rect 158864 265072 158870 265124
rect 160738 265072 160744 265124
rect 160796 265112 160802 265124
rect 161290 265112 161296 265124
rect 160796 265084 161296 265112
rect 160796 265072 160802 265084
rect 161290 265072 161296 265084
rect 161348 265112 161354 265124
rect 193214 265112 193220 265124
rect 161348 265084 193220 265112
rect 161348 265072 161354 265084
rect 193214 265072 193220 265084
rect 193272 265072 193278 265124
rect 190454 265044 190460 265056
rect 157260 265016 190460 265044
rect 157260 264988 157288 265016
rect 190454 265004 190460 265016
rect 190512 265004 190518 265056
rect 114278 264936 114284 264988
rect 114336 264976 114342 264988
rect 135898 264976 135904 264988
rect 114336 264948 135904 264976
rect 114336 264936 114342 264948
rect 135898 264936 135904 264948
rect 135956 264936 135962 264988
rect 156322 264936 156328 264988
rect 156380 264976 156386 264988
rect 157242 264976 157248 264988
rect 156380 264948 157248 264976
rect 156380 264936 156386 264948
rect 157242 264936 157248 264948
rect 157300 264936 157306 264988
rect 158806 264936 158812 264988
rect 158864 264976 158870 264988
rect 159634 264976 159640 264988
rect 158864 264948 159640 264976
rect 158864 264936 158870 264948
rect 159634 264936 159640 264948
rect 159692 264976 159698 264988
rect 193766 264976 193772 264988
rect 159692 264948 193772 264976
rect 159692 264936 159698 264948
rect 193766 264936 193772 264948
rect 193824 264936 193830 264988
rect 119154 264392 119160 264444
rect 119212 264432 119218 264444
rect 145558 264432 145564 264444
rect 119212 264404 145564 264432
rect 119212 264392 119218 264404
rect 145558 264392 145564 264404
rect 145616 264392 145622 264444
rect 139762 264324 139768 264376
rect 139820 264364 139826 264376
rect 139820 264336 142154 264364
rect 139820 264324 139826 264336
rect 118142 264256 118148 264308
rect 118200 264296 118206 264308
rect 137186 264296 137192 264308
rect 118200 264268 137192 264296
rect 118200 264256 118206 264268
rect 137186 264256 137192 264268
rect 137244 264256 137250 264308
rect 142126 264296 142154 264336
rect 178678 264296 178684 264308
rect 142126 264268 178684 264296
rect 178678 264256 178684 264268
rect 178736 264256 178742 264308
rect 4798 264188 4804 264240
rect 4856 264228 4862 264240
rect 168374 264228 168380 264240
rect 4856 264200 168380 264228
rect 4856 264188 4862 264200
rect 168374 264188 168380 264200
rect 168432 264188 168438 264240
rect 188246 264188 188252 264240
rect 188304 264228 188310 264240
rect 299474 264228 299480 264240
rect 188304 264200 299480 264228
rect 188304 264188 188310 264200
rect 299474 264188 299480 264200
rect 299532 264188 299538 264240
rect 117130 264120 117136 264172
rect 117188 264160 117194 264172
rect 133966 264160 133972 264172
rect 117188 264132 133972 264160
rect 117188 264120 117194 264132
rect 133966 264120 133972 264132
rect 134024 264160 134030 264172
rect 134518 264160 134524 264172
rect 134024 264132 134524 264160
rect 134024 264120 134030 264132
rect 134518 264120 134524 264132
rect 134576 264120 134582 264172
rect 119798 264052 119804 264104
rect 119856 264092 119862 264104
rect 138658 264092 138664 264104
rect 119856 264064 138664 264092
rect 119856 264052 119862 264064
rect 138658 264052 138664 264064
rect 138716 264052 138722 264104
rect 117038 263984 117044 264036
rect 117096 264024 117102 264036
rect 135346 264024 135352 264036
rect 117096 263996 135352 264024
rect 117096 263984 117102 263996
rect 135346 263984 135352 263996
rect 135404 264024 135410 264036
rect 135990 264024 135996 264036
rect 135404 263996 135996 264024
rect 135404 263984 135410 263996
rect 135990 263984 135996 263996
rect 136048 263984 136054 264036
rect 137094 263984 137100 264036
rect 137152 264024 137158 264036
rect 141050 264024 141056 264036
rect 137152 263996 141056 264024
rect 137152 263984 137158 263996
rect 141050 263984 141056 263996
rect 141108 263984 141114 264036
rect 119614 263916 119620 263968
rect 119672 263956 119678 263968
rect 141602 263956 141608 263968
rect 119672 263928 141608 263956
rect 119672 263916 119678 263928
rect 141602 263916 141608 263928
rect 141660 263916 141666 263968
rect 114186 263848 114192 263900
rect 114244 263888 114250 263900
rect 137278 263888 137284 263900
rect 114244 263860 137284 263888
rect 114244 263848 114250 263860
rect 137278 263848 137284 263860
rect 137336 263848 137342 263900
rect 120994 263780 121000 263832
rect 121052 263820 121058 263832
rect 143626 263820 143632 263832
rect 121052 263792 143632 263820
rect 121052 263780 121058 263792
rect 143626 263780 143632 263792
rect 143684 263820 143690 263832
rect 144178 263820 144184 263832
rect 143684 263792 144184 263820
rect 143684 263780 143690 263792
rect 144178 263780 144184 263792
rect 144236 263780 144242 263832
rect 118326 263712 118332 263764
rect 118384 263752 118390 263764
rect 137094 263752 137100 263764
rect 118384 263724 137100 263752
rect 118384 263712 118390 263724
rect 137094 263712 137100 263724
rect 137152 263712 137158 263764
rect 137186 263712 137192 263764
rect 137244 263752 137250 263764
rect 140222 263752 140228 263764
rect 137244 263724 140228 263752
rect 137244 263712 137250 263724
rect 140222 263712 140228 263724
rect 140280 263712 140286 263764
rect 176654 263712 176660 263764
rect 176712 263752 176718 263764
rect 190914 263752 190920 263764
rect 176712 263724 190920 263752
rect 176712 263712 176718 263724
rect 190914 263712 190920 263724
rect 190972 263712 190978 263764
rect 121086 263644 121092 263696
rect 121144 263684 121150 263696
rect 139762 263684 139768 263696
rect 121144 263656 139768 263684
rect 121144 263644 121150 263656
rect 139762 263644 139768 263656
rect 139820 263684 139826 263696
rect 140314 263684 140320 263696
rect 139820 263656 140320 263684
rect 139820 263644 139826 263656
rect 140314 263644 140320 263656
rect 140372 263644 140378 263696
rect 168374 263644 168380 263696
rect 168432 263684 168438 263696
rect 189258 263684 189264 263696
rect 168432 263656 189264 263684
rect 168432 263644 168438 263656
rect 189258 263644 189264 263656
rect 189316 263644 189322 263696
rect 120902 263576 120908 263628
rect 120960 263616 120966 263628
rect 149146 263616 149152 263628
rect 120960 263588 149152 263616
rect 120960 263576 120966 263588
rect 149146 263576 149152 263588
rect 149204 263616 149210 263628
rect 149974 263616 149980 263628
rect 149204 263588 149980 263616
rect 149204 263576 149210 263588
rect 149974 263576 149980 263588
rect 150032 263576 150038 263628
rect 155218 263576 155224 263628
rect 155276 263616 155282 263628
rect 188246 263616 188252 263628
rect 155276 263588 188252 263616
rect 155276 263576 155282 263588
rect 188246 263576 188252 263588
rect 188304 263576 188310 263628
rect 138290 263508 138296 263560
rect 138348 263548 138354 263560
rect 580258 263548 580264 263560
rect 138348 263520 580264 263548
rect 138348 263508 138354 263520
rect 580258 263508 580264 263520
rect 580316 263508 580322 263560
rect 151814 263440 151820 263492
rect 151872 263480 151878 263492
rect 152182 263480 152188 263492
rect 151872 263452 152188 263480
rect 151872 263440 151878 263452
rect 152182 263440 152188 263452
rect 152240 263440 152246 263492
rect 187970 263440 187976 263492
rect 188028 263480 188034 263492
rect 347774 263480 347780 263492
rect 188028 263452 347780 263480
rect 188028 263440 188034 263452
rect 347774 263440 347780 263452
rect 347832 263440 347838 263492
rect 146386 263168 146392 263220
rect 146444 263208 146450 263220
rect 147030 263208 147036 263220
rect 146444 263180 147036 263208
rect 146444 263168 146450 263180
rect 147030 263168 147036 263180
rect 147088 263168 147094 263220
rect 112438 263032 112444 263084
rect 112496 263072 112502 263084
rect 131206 263072 131212 263084
rect 112496 263044 131212 263072
rect 112496 263032 112502 263044
rect 131206 263032 131212 263044
rect 131264 263032 131270 263084
rect 133690 263032 133696 263084
rect 133748 263072 133754 263084
rect 580350 263072 580356 263084
rect 133748 263044 580356 263072
rect 133748 263032 133754 263044
rect 580350 263032 580356 263044
rect 580408 263032 580414 263084
rect 115198 262964 115204 263016
rect 115256 263004 115262 263016
rect 132586 263004 132592 263016
rect 115256 262976 132592 263004
rect 115256 262964 115262 262976
rect 132586 262964 132592 262976
rect 132644 263004 132650 263016
rect 133782 263004 133788 263016
rect 132644 262976 133788 263004
rect 132644 262964 132650 262976
rect 133782 262964 133788 262976
rect 133840 262964 133846 263016
rect 3418 262896 3424 262948
rect 3476 262936 3482 262948
rect 178770 262936 178776 262948
rect 3476 262908 178776 262936
rect 3476 262896 3482 262908
rect 178770 262896 178776 262908
rect 178828 262896 178834 262948
rect 180426 262896 180432 262948
rect 180484 262936 180490 262948
rect 187142 262936 187148 262948
rect 180484 262908 187148 262936
rect 180484 262896 180490 262908
rect 187142 262896 187148 262908
rect 187200 262896 187206 262948
rect 118050 262828 118056 262880
rect 118108 262868 118114 262880
rect 133138 262868 133144 262880
rect 118108 262840 133144 262868
rect 118108 262828 118114 262840
rect 133138 262828 133144 262840
rect 133196 262828 133202 262880
rect 178126 262828 178132 262880
rect 178184 262868 178190 262880
rect 189626 262868 189632 262880
rect 178184 262840 189632 262868
rect 178184 262828 178190 262840
rect 189626 262828 189632 262840
rect 189684 262828 189690 262880
rect 191742 262828 191748 262880
rect 191800 262868 191806 262880
rect 218054 262868 218060 262880
rect 191800 262840 218060 262868
rect 191800 262828 191806 262840
rect 218054 262828 218060 262840
rect 218112 262828 218118 262880
rect 111058 262760 111064 262812
rect 111116 262800 111122 262812
rect 129734 262800 129740 262812
rect 111116 262772 129740 262800
rect 111116 262760 111122 262772
rect 129734 262760 129740 262772
rect 129792 262760 129798 262812
rect 133782 262760 133788 262812
rect 133840 262800 133846 262812
rect 580442 262800 580448 262812
rect 133840 262772 580448 262800
rect 133840 262760 133846 262772
rect 580442 262760 580448 262772
rect 580500 262760 580506 262812
rect 116946 262692 116952 262744
rect 117004 262732 117010 262744
rect 128446 262732 128452 262744
rect 117004 262704 128452 262732
rect 117004 262692 117010 262704
rect 128446 262692 128452 262704
rect 128504 262692 128510 262744
rect 170398 262692 170404 262744
rect 170456 262732 170462 262744
rect 192478 262732 192484 262744
rect 170456 262704 192484 262732
rect 170456 262692 170462 262704
rect 192478 262692 192484 262704
rect 192536 262692 192542 262744
rect 117958 262624 117964 262676
rect 118016 262664 118022 262676
rect 146386 262664 146392 262676
rect 118016 262636 146392 262664
rect 118016 262624 118022 262636
rect 146386 262624 146392 262636
rect 146444 262624 146450 262676
rect 169018 262624 169024 262676
rect 169076 262664 169082 262676
rect 193674 262664 193680 262676
rect 169076 262636 193680 262664
rect 169076 262624 169082 262636
rect 193674 262624 193680 262636
rect 193732 262624 193738 262676
rect 120626 262556 120632 262608
rect 120684 262596 120690 262608
rect 150434 262596 150440 262608
rect 120684 262568 150440 262596
rect 120684 262556 120690 262568
rect 150434 262556 150440 262568
rect 150492 262556 150498 262608
rect 158346 262556 158352 262608
rect 158404 262596 158410 262608
rect 190822 262596 190828 262608
rect 158404 262568 190828 262596
rect 158404 262556 158410 262568
rect 190822 262556 190828 262568
rect 190880 262596 190886 262608
rect 191742 262596 191748 262608
rect 190880 262568 191748 262596
rect 190880 262556 190886 262568
rect 191742 262556 191748 262568
rect 191800 262556 191806 262608
rect 119430 262488 119436 262540
rect 119488 262528 119494 262540
rect 149698 262528 149704 262540
rect 119488 262500 149704 262528
rect 119488 262488 119494 262500
rect 149698 262488 149704 262500
rect 149756 262488 149762 262540
rect 155034 262488 155040 262540
rect 155092 262528 155098 262540
rect 187970 262528 187976 262540
rect 155092 262500 187976 262528
rect 155092 262488 155098 262500
rect 187970 262488 187976 262500
rect 188028 262488 188034 262540
rect 3510 262420 3516 262472
rect 3568 262460 3574 262472
rect 177758 262460 177764 262472
rect 3568 262432 177764 262460
rect 3568 262420 3574 262432
rect 177758 262420 177764 262432
rect 177816 262420 177822 262472
rect 180610 262420 180616 262472
rect 180668 262460 180674 262472
rect 192202 262460 192208 262472
rect 180668 262432 192208 262460
rect 180668 262420 180674 262432
rect 192202 262420 192208 262432
rect 192260 262420 192266 262472
rect 117866 262352 117872 262404
rect 117924 262392 117930 262404
rect 130102 262392 130108 262404
rect 117924 262364 130108 262392
rect 117924 262352 117930 262364
rect 130102 262352 130108 262364
rect 130160 262352 130166 262404
rect 183186 262352 183192 262404
rect 183244 262392 183250 262404
rect 196526 262392 196532 262404
rect 183244 262364 196532 262392
rect 183244 262352 183250 262364
rect 196526 262352 196532 262364
rect 196584 262352 196590 262404
rect 119522 262284 119528 262336
rect 119580 262324 119586 262336
rect 125134 262324 125140 262336
rect 119580 262296 125140 262324
rect 119580 262284 119586 262296
rect 125134 262284 125140 262296
rect 125192 262284 125198 262336
rect 121178 262216 121184 262268
rect 121236 262256 121242 262268
rect 126974 262256 126980 262268
rect 121236 262228 126980 262256
rect 121236 262216 121242 262228
rect 126974 262216 126980 262228
rect 127032 262216 127038 262268
rect 182082 262216 182088 262268
rect 182140 262256 182146 262268
rect 187050 262256 187056 262268
rect 182140 262228 187056 262256
rect 182140 262216 182146 262228
rect 187050 262216 187056 262228
rect 187108 262216 187114 262268
rect 181530 261332 181536 261384
rect 181588 261372 181594 261384
rect 192662 261372 192668 261384
rect 181588 261344 192668 261372
rect 181588 261332 181594 261344
rect 192662 261332 192668 261344
rect 192720 261332 192726 261384
rect 133138 261264 133144 261316
rect 133196 261304 133202 261316
rect 133690 261304 133696 261316
rect 133196 261276 133696 261304
rect 133196 261264 133202 261276
rect 133690 261264 133696 261276
rect 133748 261304 133754 261316
rect 472618 261304 472624 261316
rect 133748 261276 472624 261304
rect 133748 261264 133754 261276
rect 472618 261264 472624 261276
rect 472676 261264 472682 261316
rect 4798 261196 4804 261248
rect 4856 261236 4862 261248
rect 178126 261236 178132 261248
rect 4856 261208 178132 261236
rect 4856 261196 4862 261208
rect 178126 261196 178132 261208
rect 178184 261196 178190 261248
rect 192570 261236 192576 261248
rect 180766 261208 192576 261236
rect 116762 261128 116768 261180
rect 116820 261168 116826 261180
rect 131114 261168 131120 261180
rect 116820 261140 131120 261168
rect 116820 261128 116826 261140
rect 131114 261128 131120 261140
rect 131172 261128 131178 261180
rect 178678 261128 178684 261180
rect 178736 261168 178742 261180
rect 180766 261168 180794 261208
rect 192570 261196 192576 261208
rect 192628 261196 192634 261248
rect 178736 261140 180794 261168
rect 178736 261128 178742 261140
rect 112346 261060 112352 261112
rect 112404 261100 112410 261112
rect 135162 261100 135168 261112
rect 112404 261072 135168 261100
rect 112404 261060 112410 261072
rect 135162 261060 135168 261072
rect 135220 261100 135226 261112
rect 187786 261100 187792 261112
rect 135220 261072 187792 261100
rect 135220 261060 135226 261072
rect 187786 261060 187792 261072
rect 187844 261060 187850 261112
rect 120534 260992 120540 261044
rect 120592 261032 120598 261044
rect 178678 261032 178684 261044
rect 120592 261004 178684 261032
rect 120592 260992 120598 261004
rect 178678 260992 178684 261004
rect 178736 260992 178742 261044
rect 178770 260992 178776 261044
rect 178828 261032 178834 261044
rect 179506 261032 179512 261044
rect 178828 261004 179512 261032
rect 178828 260992 178834 261004
rect 179506 260992 179512 261004
rect 179564 261032 179570 261044
rect 196618 261032 196624 261044
rect 179564 261004 196624 261032
rect 179564 260992 179570 261004
rect 196618 260992 196624 261004
rect 196676 260992 196682 261044
rect 177758 260924 177764 260976
rect 177816 260964 177822 260976
rect 196710 260964 196716 260976
rect 177816 260936 196716 260964
rect 177816 260924 177822 260936
rect 196710 260924 196716 260936
rect 196768 260924 196774 260976
rect 113818 260856 113824 260908
rect 113876 260896 113882 260908
rect 130654 260896 130660 260908
rect 113876 260868 130660 260896
rect 113876 260856 113882 260868
rect 130654 260856 130660 260868
rect 130712 260856 130718 260908
rect 184842 260856 184848 260908
rect 184900 260896 184906 260908
rect 196342 260896 196348 260908
rect 184900 260868 196348 260896
rect 184900 260856 184906 260868
rect 196342 260856 196348 260868
rect 196400 260856 196406 260908
rect 175182 260448 175188 260500
rect 175240 260488 175246 260500
rect 189534 260488 189540 260500
rect 175240 260460 189540 260488
rect 175240 260448 175246 260460
rect 189534 260448 189540 260460
rect 189592 260448 189598 260500
rect 157334 260380 157340 260432
rect 157392 260420 157398 260432
rect 191098 260420 191104 260432
rect 157392 260392 191104 260420
rect 157392 260380 157398 260392
rect 191098 260380 191104 260392
rect 191156 260380 191162 260432
rect 7558 260312 7564 260364
rect 7616 260352 7622 260364
rect 177022 260352 177028 260364
rect 7616 260324 177028 260352
rect 7616 260312 7622 260324
rect 177022 260312 177028 260324
rect 177080 260312 177086 260364
rect 182634 260312 182640 260364
rect 182692 260352 182698 260364
rect 192386 260352 192392 260364
rect 182692 260324 192392 260352
rect 182692 260312 182698 260324
rect 192386 260312 192392 260324
rect 192444 260312 192450 260364
rect 131114 260244 131120 260296
rect 131172 260284 131178 260296
rect 132034 260284 132040 260296
rect 131172 260256 132040 260284
rect 131172 260244 131178 260256
rect 132034 260244 132040 260256
rect 132092 260284 132098 260296
rect 471238 260284 471244 260296
rect 132092 260256 471244 260284
rect 132092 260244 132098 260256
rect 471238 260244 471244 260256
rect 471296 260244 471302 260296
rect 146570 260176 146576 260228
rect 146628 260216 146634 260228
rect 147536 260216 147542 260228
rect 146628 260188 147542 260216
rect 146628 260176 146634 260188
rect 147536 260176 147542 260188
rect 147594 260176 147600 260228
rect 147674 260176 147680 260228
rect 147732 260216 147738 260228
rect 148640 260216 148646 260228
rect 147732 260188 148646 260216
rect 147732 260176 147738 260188
rect 148640 260176 148646 260188
rect 148698 260176 148704 260228
rect 153194 260176 153200 260228
rect 153252 260216 153258 260228
rect 154160 260216 154166 260228
rect 153252 260188 154166 260216
rect 153252 260176 153258 260188
rect 154160 260176 154166 260188
rect 154218 260176 154224 260228
rect 157610 260176 157616 260228
rect 157668 260216 157674 260228
rect 158576 260216 158582 260228
rect 157668 260188 158582 260216
rect 157668 260176 157674 260188
rect 158576 260176 158582 260188
rect 158634 260176 158640 260228
rect 165614 260176 165620 260228
rect 165672 260216 165678 260228
rect 166856 260216 166862 260228
rect 165672 260188 166862 260216
rect 165672 260176 165678 260188
rect 166856 260176 166862 260188
rect 166914 260176 166920 260228
rect 170168 260176 170174 260228
rect 170226 260216 170232 260228
rect 189442 260216 189448 260228
rect 170226 260188 189448 260216
rect 170226 260176 170232 260188
rect 189442 260176 189448 260188
rect 189500 260176 189506 260228
rect 171134 260108 171140 260160
rect 171192 260148 171198 260160
rect 171824 260148 171830 260160
rect 171192 260120 171830 260148
rect 171192 260108 171198 260120
rect 171824 260108 171830 260120
rect 171882 260108 171888 260160
rect 172514 260108 172520 260160
rect 172572 260148 172578 260160
rect 173480 260148 173486 260160
rect 172572 260120 173486 260148
rect 172572 260108 172578 260120
rect 173480 260108 173486 260120
rect 173538 260108 173544 260160
rect 173986 260108 173992 260160
rect 174044 260148 174050 260160
rect 175136 260148 175142 260160
rect 174044 260120 175142 260148
rect 174044 260108 174050 260120
rect 175136 260108 175142 260120
rect 175194 260108 175200 260160
rect 186958 260148 186964 260160
rect 175568 260120 186964 260148
rect 123478 260040 123484 260092
rect 123536 260080 123542 260092
rect 123536 260052 128354 260080
rect 123536 260040 123542 260052
rect 116578 259972 116584 260024
rect 116636 260012 116642 260024
rect 116636 259984 127572 260012
rect 116636 259972 116642 259984
rect 113910 259904 113916 259956
rect 113968 259944 113974 259956
rect 127342 259944 127348 259956
rect 113968 259916 127348 259944
rect 113968 259904 113974 259916
rect 127342 259904 127348 259916
rect 127400 259904 127406 259956
rect 115382 259836 115388 259888
rect 115440 259876 115446 259888
rect 123478 259876 123484 259888
rect 115440 259848 123484 259876
rect 115440 259836 115446 259848
rect 123478 259836 123484 259848
rect 123536 259836 123542 259888
rect 116670 259768 116676 259820
rect 116728 259808 116734 259820
rect 124214 259808 124220 259820
rect 116728 259780 124220 259808
rect 116728 259768 116734 259780
rect 124214 259768 124220 259780
rect 124272 259768 124278 259820
rect 127544 259808 127572 259984
rect 128326 259944 128354 260052
rect 171842 259944 171870 260108
rect 173498 260080 173526 260108
rect 175568 260080 175596 260120
rect 186958 260108 186964 260120
rect 187016 260108 187022 260160
rect 173498 260052 175596 260080
rect 184934 259972 184940 260024
rect 184992 260012 184998 260024
rect 189810 260012 189816 260024
rect 184992 259984 189816 260012
rect 184992 259972 184998 259984
rect 189810 259972 189816 259984
rect 189868 259972 189874 260024
rect 187878 259944 187884 259956
rect 128326 259916 132494 259944
rect 171842 259916 187884 259944
rect 132466 259876 132494 259916
rect 187878 259904 187884 259916
rect 187936 259904 187942 259956
rect 135530 259876 135536 259888
rect 132466 259848 135536 259876
rect 135530 259836 135536 259848
rect 135588 259836 135594 259888
rect 166994 259836 167000 259888
rect 167052 259876 167058 259888
rect 186682 259876 186688 259888
rect 167052 259848 186688 259876
rect 167052 259836 167058 259848
rect 186682 259836 186688 259848
rect 186740 259836 186746 259888
rect 142154 259808 142160 259820
rect 127544 259780 142160 259808
rect 142154 259768 142160 259780
rect 142212 259768 142218 259820
rect 160554 259768 160560 259820
rect 160612 259808 160618 259820
rect 186774 259808 186780 259820
rect 160612 259780 186780 259808
rect 160612 259768 160618 259780
rect 186774 259768 186780 259780
rect 186832 259768 186838 259820
rect 118234 259700 118240 259752
rect 118292 259740 118298 259752
rect 146570 259740 146576 259752
rect 118292 259712 146576 259740
rect 118292 259700 118298 259712
rect 146570 259700 146576 259712
rect 146628 259700 146634 259752
rect 158714 259700 158720 259752
rect 158772 259740 158778 259752
rect 188062 259740 188068 259752
rect 158772 259712 188068 259740
rect 158772 259700 158778 259712
rect 188062 259700 188068 259712
rect 188120 259700 188126 259752
rect 119338 259632 119344 259684
rect 119396 259672 119402 259684
rect 147674 259672 147680 259684
rect 119396 259644 147680 259672
rect 119396 259632 119402 259644
rect 147674 259632 147680 259644
rect 147732 259632 147738 259684
rect 159450 259632 159456 259684
rect 159508 259672 159514 259684
rect 191006 259672 191012 259684
rect 159508 259644 191012 259672
rect 159508 259632 159514 259644
rect 191006 259632 191012 259644
rect 191064 259632 191070 259684
rect 119246 259564 119252 259616
rect 119304 259604 119310 259616
rect 153194 259604 153200 259616
rect 119304 259576 153200 259604
rect 119304 259564 119310 259576
rect 153194 259564 153200 259576
rect 153252 259564 153258 259616
rect 174354 259564 174360 259616
rect 174412 259604 174418 259616
rect 184934 259604 184940 259616
rect 174412 259576 184940 259604
rect 174412 259564 174418 259576
rect 184934 259564 184940 259576
rect 184992 259564 184998 259616
rect 189902 259604 189908 259616
rect 185228 259576 189908 259604
rect 115290 259496 115296 259548
rect 115348 259536 115354 259548
rect 124582 259536 124588 259548
rect 115348 259508 124588 259536
rect 115348 259496 115354 259508
rect 124582 259496 124588 259508
rect 124640 259496 124646 259548
rect 177666 259496 177672 259548
rect 177724 259536 177730 259548
rect 185228 259536 185256 259576
rect 189902 259564 189908 259576
rect 189960 259564 189966 259616
rect 177724 259508 185256 259536
rect 177724 259496 177730 259508
rect 185302 259496 185308 259548
rect 185360 259536 185366 259548
rect 187234 259536 187240 259548
rect 185360 259508 187240 259536
rect 185360 259496 185366 259508
rect 187234 259496 187240 259508
rect 187292 259496 187298 259548
rect 115106 259428 115112 259480
rect 115164 259468 115170 259480
rect 128998 259468 129004 259480
rect 115164 259440 129004 259468
rect 115164 259428 115170 259440
rect 128998 259428 129004 259440
rect 129056 259428 129062 259480
rect 184290 259428 184296 259480
rect 184348 259468 184354 259480
rect 195054 259468 195060 259480
rect 184348 259440 195060 259468
rect 184348 259428 184354 259440
rect 195054 259428 195060 259440
rect 195112 259428 195118 259480
rect 120810 259360 120816 259412
rect 120868 259400 120874 259412
rect 123478 259400 123484 259412
rect 120868 259372 123484 259400
rect 120868 259360 120874 259372
rect 123478 259360 123484 259372
rect 123536 259360 123542 259412
rect 187786 259360 187792 259412
rect 187844 259400 187850 259412
rect 580166 259400 580172 259412
rect 187844 259372 580172 259400
rect 187844 259360 187850 259372
rect 580166 259360 580172 259372
rect 580224 259360 580230 259412
rect 183646 259292 183652 259344
rect 183704 259332 183710 259344
rect 188246 259332 188252 259344
rect 183704 259304 188252 259332
rect 183704 259292 183710 259304
rect 188246 259292 188252 259304
rect 188304 259292 188310 259344
rect 187786 259224 187792 259276
rect 187844 259264 187850 259276
rect 188338 259264 188344 259276
rect 187844 259236 188344 259264
rect 187844 259224 187850 259236
rect 188338 259224 188344 259236
rect 188396 259224 188402 259276
rect 472618 245556 472624 245608
rect 472676 245596 472682 245608
rect 580166 245596 580172 245608
rect 472676 245568 580172 245596
rect 472676 245556 472682 245568
rect 580166 245556 580172 245568
rect 580224 245556 580230 245608
rect 3510 241068 3516 241120
rect 3568 241108 3574 241120
rect 7558 241108 7564 241120
rect 3568 241080 7564 241108
rect 3568 241068 3574 241080
rect 7558 241068 7564 241080
rect 7616 241068 7622 241120
rect 2774 215228 2780 215280
rect 2832 215268 2838 215280
rect 4798 215268 4804 215280
rect 2832 215240 4804 215268
rect 2832 215228 2838 215240
rect 4798 215228 4804 215240
rect 4856 215228 4862 215280
rect 471238 206932 471244 206984
rect 471296 206972 471302 206984
rect 579798 206972 579804 206984
rect 471296 206944 579804 206972
rect 471296 206932 471302 206944
rect 579798 206932 579804 206944
rect 579856 206932 579862 206984
rect 106918 199860 106924 199912
rect 106976 199900 106982 199912
rect 131298 199900 131304 199912
rect 106976 199872 131304 199900
rect 106976 199860 106982 199872
rect 131298 199860 131304 199872
rect 131356 199860 131362 199912
rect 132034 199860 132040 199912
rect 132092 199900 132098 199912
rect 132540 199900 132546 199912
rect 132092 199872 132546 199900
rect 132092 199860 132098 199872
rect 132540 199860 132546 199872
rect 132598 199860 132604 199912
rect 134104 199860 134110 199912
rect 134162 199900 134168 199912
rect 134162 199860 134196 199900
rect 134288 199860 134294 199912
rect 134346 199860 134352 199912
rect 135024 199860 135030 199912
rect 135082 199900 135088 199912
rect 135082 199872 135162 199900
rect 135082 199860 135088 199872
rect 131942 199792 131948 199844
rect 132000 199832 132006 199844
rect 132816 199832 132822 199844
rect 132000 199804 132822 199832
rect 132000 199792 132006 199804
rect 132816 199792 132822 199804
rect 132874 199792 132880 199844
rect 133828 199792 133834 199844
rect 133886 199832 133892 199844
rect 133886 199804 133966 199832
rect 133886 199792 133892 199804
rect 133644 199724 133650 199776
rect 133702 199724 133708 199776
rect 133736 199724 133742 199776
rect 133794 199764 133800 199776
rect 133794 199736 133874 199764
rect 133794 199724 133800 199736
rect 131666 199656 131672 199708
rect 131724 199696 131730 199708
rect 133662 199696 133690 199724
rect 131724 199668 133690 199696
rect 131724 199656 131730 199668
rect 133846 199640 133874 199736
rect 133414 199628 133420 199640
rect 129706 199600 133420 199628
rect 104434 199452 104440 199504
rect 104492 199492 104498 199504
rect 129706 199492 129734 199600
rect 133414 199588 133420 199600
rect 133472 199588 133478 199640
rect 133782 199588 133788 199640
rect 133840 199600 133874 199640
rect 133840 199588 133846 199600
rect 133938 199572 133966 199804
rect 134012 199792 134018 199844
rect 134070 199832 134076 199844
rect 134070 199792 134104 199832
rect 134076 199708 134104 199792
rect 134058 199656 134064 199708
rect 134116 199656 134122 199708
rect 133874 199520 133880 199572
rect 133932 199532 133966 199572
rect 133932 199520 133938 199532
rect 104492 199464 129734 199492
rect 104492 199452 104498 199464
rect 133598 199452 133604 199504
rect 133656 199492 133662 199504
rect 134168 199492 134196 199860
rect 133656 199464 134196 199492
rect 134306 199504 134334 199860
rect 134840 199724 134846 199776
rect 134898 199764 134904 199776
rect 134898 199736 135070 199764
rect 134898 199724 134904 199736
rect 135042 199640 135070 199736
rect 135134 199696 135162 199872
rect 135208 199860 135214 199912
rect 135266 199900 135272 199912
rect 135266 199860 135300 199900
rect 135484 199860 135490 199912
rect 135542 199860 135548 199912
rect 135576 199860 135582 199912
rect 135634 199860 135640 199912
rect 135668 199860 135674 199912
rect 135726 199860 135732 199912
rect 135944 199860 135950 199912
rect 136002 199860 136008 199912
rect 136404 199860 136410 199912
rect 136462 199860 136468 199912
rect 136496 199860 136502 199912
rect 136554 199860 136560 199912
rect 136864 199860 136870 199912
rect 136922 199860 136928 199912
rect 136956 199860 136962 199912
rect 137014 199860 137020 199912
rect 137048 199860 137054 199912
rect 137106 199900 137112 199912
rect 137106 199860 137140 199900
rect 137232 199860 137238 199912
rect 137290 199860 137296 199912
rect 137600 199900 137606 199912
rect 137342 199872 137606 199900
rect 135272 199776 135300 199860
rect 135392 199832 135398 199844
rect 135364 199792 135398 199832
rect 135450 199792 135456 199844
rect 135254 199724 135260 199776
rect 135312 199724 135318 199776
rect 135134 199668 135300 199696
rect 135272 199640 135300 199668
rect 135042 199600 135076 199640
rect 135070 199588 135076 199600
rect 135128 199588 135134 199640
rect 135254 199588 135260 199640
rect 135312 199588 135318 199640
rect 135364 199560 135392 199792
rect 135502 199764 135530 199860
rect 135456 199736 135530 199764
rect 135456 199708 135484 199736
rect 135594 199708 135622 199860
rect 135438 199656 135444 199708
rect 135496 199656 135502 199708
rect 135530 199656 135536 199708
rect 135588 199668 135622 199708
rect 135588 199656 135594 199668
rect 135686 199640 135714 199860
rect 135760 199792 135766 199844
rect 135818 199832 135824 199844
rect 135818 199792 135852 199832
rect 135824 199708 135852 199792
rect 135806 199656 135812 199708
rect 135864 199656 135870 199708
rect 135962 199640 135990 199860
rect 136128 199792 136134 199844
rect 136186 199792 136192 199844
rect 136220 199792 136226 199844
rect 136278 199792 136284 199844
rect 136312 199792 136318 199844
rect 136370 199792 136376 199844
rect 136146 199640 136174 199792
rect 135686 199600 135720 199640
rect 135714 199588 135720 199600
rect 135772 199588 135778 199640
rect 135962 199600 135996 199640
rect 135990 199588 135996 199600
rect 136048 199588 136054 199640
rect 136082 199588 136088 199640
rect 136140 199600 136174 199640
rect 136140 199588 136146 199600
rect 136238 199572 136266 199792
rect 135898 199560 135904 199572
rect 135364 199532 135904 199560
rect 135898 199520 135904 199532
rect 135956 199520 135962 199572
rect 136174 199520 136180 199572
rect 136232 199532 136266 199572
rect 136232 199520 136238 199532
rect 134306 199464 134340 199504
rect 133656 199452 133662 199464
rect 134334 199452 134340 199464
rect 134392 199452 134398 199504
rect 136330 199492 136358 199792
rect 136422 199708 136450 199860
rect 136514 199776 136542 199860
rect 136772 199792 136778 199844
rect 136830 199792 136836 199844
rect 136514 199736 136548 199776
rect 136542 199724 136548 199736
rect 136600 199724 136606 199776
rect 136422 199668 136456 199708
rect 136450 199656 136456 199668
rect 136508 199656 136514 199708
rect 136790 199640 136818 199792
rect 136882 199776 136910 199860
rect 136974 199832 137002 199860
rect 136974 199804 137048 199832
rect 136882 199736 136916 199776
rect 136910 199724 136916 199736
rect 136968 199724 136974 199776
rect 137020 199640 137048 199804
rect 137112 199708 137140 199860
rect 137094 199656 137100 199708
rect 137152 199656 137158 199708
rect 137250 199696 137278 199860
rect 137342 199776 137370 199872
rect 137600 199860 137606 199872
rect 137658 199860 137664 199912
rect 137784 199860 137790 199912
rect 137842 199860 137848 199912
rect 137968 199860 137974 199912
rect 138026 199860 138032 199912
rect 138244 199860 138250 199912
rect 138302 199860 138308 199912
rect 138336 199860 138342 199912
rect 138394 199860 138400 199912
rect 138704 199860 138710 199912
rect 138762 199860 138768 199912
rect 139256 199860 139262 199912
rect 139314 199860 139320 199912
rect 139624 199900 139630 199912
rect 139412 199872 139630 199900
rect 137324 199724 137330 199776
rect 137382 199724 137388 199776
rect 137204 199668 137278 199696
rect 136726 199588 136732 199640
rect 136784 199600 136818 199640
rect 136784 199588 136790 199600
rect 137002 199588 137008 199640
rect 137060 199588 137066 199640
rect 137204 199560 137232 199668
rect 137278 199588 137284 199640
rect 137336 199628 137342 199640
rect 137802 199628 137830 199860
rect 137986 199764 138014 199860
rect 137940 199736 138014 199764
rect 137940 199708 137968 199736
rect 137922 199656 137928 199708
rect 137980 199656 137986 199708
rect 138014 199656 138020 199708
rect 138072 199696 138078 199708
rect 138262 199696 138290 199860
rect 138072 199668 138290 199696
rect 138072 199656 138078 199668
rect 138354 199640 138382 199860
rect 137336 199600 137830 199628
rect 137336 199588 137342 199600
rect 138290 199588 138296 199640
rect 138348 199600 138382 199640
rect 138348 199588 138354 199600
rect 137204 199532 138060 199560
rect 138032 199504 138060 199532
rect 138382 199520 138388 199572
rect 138440 199560 138446 199572
rect 138722 199560 138750 199860
rect 139274 199640 139302 199860
rect 139412 199764 139440 199872
rect 139624 199860 139630 199872
rect 139682 199860 139688 199912
rect 139900 199860 139906 199912
rect 139958 199860 139964 199912
rect 140820 199860 140826 199912
rect 140878 199860 140884 199912
rect 141096 199860 141102 199912
rect 141154 199860 141160 199912
rect 141556 199860 141562 199912
rect 141614 199860 141620 199912
rect 141648 199860 141654 199912
rect 141706 199860 141712 199912
rect 141832 199860 141838 199912
rect 141890 199860 141896 199912
rect 142200 199900 142206 199912
rect 141942 199872 142206 199900
rect 139578 199764 139584 199776
rect 139412 199736 139584 199764
rect 139578 199724 139584 199736
rect 139636 199724 139642 199776
rect 139918 199640 139946 199860
rect 140838 199776 140866 199860
rect 140774 199724 140780 199776
rect 140832 199736 140866 199776
rect 140832 199724 140838 199736
rect 141114 199696 141142 199860
rect 139210 199588 139216 199640
rect 139268 199600 139302 199640
rect 139268 199588 139274 199600
rect 139854 199588 139860 199640
rect 139912 199600 139946 199640
rect 140608 199668 141142 199696
rect 141574 199708 141602 199860
rect 141666 199764 141694 199860
rect 141666 199736 141740 199764
rect 141574 199668 141608 199708
rect 139912 199588 139918 199600
rect 138440 199532 138750 199560
rect 138440 199520 138446 199532
rect 136450 199492 136456 199504
rect 136330 199464 136456 199492
rect 136450 199452 136456 199464
rect 136508 199452 136514 199504
rect 136634 199452 136640 199504
rect 136692 199492 136698 199504
rect 137462 199492 137468 199504
rect 136692 199464 137468 199492
rect 136692 199452 136698 199464
rect 137462 199452 137468 199464
rect 137520 199452 137526 199504
rect 138014 199452 138020 199504
rect 138072 199452 138078 199504
rect 140038 199452 140044 199504
rect 140096 199492 140102 199504
rect 140608 199492 140636 199668
rect 141602 199656 141608 199668
rect 141660 199656 141666 199708
rect 141712 199640 141740 199736
rect 141694 199588 141700 199640
rect 141752 199588 141758 199640
rect 140682 199520 140688 199572
rect 140740 199560 140746 199572
rect 141850 199560 141878 199860
rect 140740 199532 141878 199560
rect 140740 199520 140746 199532
rect 140866 199492 140872 199504
rect 140096 199464 140544 199492
rect 140608 199464 140872 199492
rect 140096 199452 140102 199464
rect 136358 199384 136364 199436
rect 136416 199424 136422 199436
rect 140406 199424 140412 199436
rect 136416 199396 140412 199424
rect 136416 199384 136422 199396
rect 140406 199384 140412 199396
rect 140464 199384 140470 199436
rect 140516 199424 140544 199464
rect 140866 199452 140872 199464
rect 140924 199452 140930 199504
rect 141786 199452 141792 199504
rect 141844 199492 141850 199504
rect 141942 199492 141970 199872
rect 142200 199860 142206 199872
rect 142258 199860 142264 199912
rect 142384 199860 142390 199912
rect 142442 199900 142448 199912
rect 142442 199860 142476 199900
rect 142752 199860 142758 199912
rect 142810 199860 142816 199912
rect 143120 199900 143126 199912
rect 142862 199872 143126 199900
rect 142448 199708 142476 199860
rect 142770 199776 142798 199860
rect 142706 199724 142712 199776
rect 142764 199736 142798 199776
rect 142764 199724 142770 199736
rect 142430 199656 142436 199708
rect 142488 199656 142494 199708
rect 142246 199588 142252 199640
rect 142304 199628 142310 199640
rect 142862 199628 142890 199872
rect 143120 199860 143126 199872
rect 143178 199860 143184 199912
rect 143212 199860 143218 199912
rect 143270 199860 143276 199912
rect 143396 199860 143402 199912
rect 143454 199860 143460 199912
rect 143488 199860 143494 199912
rect 143546 199860 143552 199912
rect 143672 199860 143678 199912
rect 143730 199860 143736 199912
rect 144040 199860 144046 199912
rect 144098 199860 144104 199912
rect 144224 199860 144230 199912
rect 144282 199860 144288 199912
rect 144316 199860 144322 199912
rect 144374 199860 144380 199912
rect 144868 199860 144874 199912
rect 144926 199860 144932 199912
rect 145420 199900 145426 199912
rect 144978 199872 145426 199900
rect 143230 199776 143258 199860
rect 143166 199724 143172 199776
rect 143224 199736 143258 199776
rect 143224 199724 143230 199736
rect 143414 199640 143442 199860
rect 142304 199600 142890 199628
rect 142304 199588 142310 199600
rect 143350 199588 143356 199640
rect 143408 199600 143442 199640
rect 143408 199588 143414 199600
rect 143506 199572 143534 199860
rect 143690 199640 143718 199860
rect 143626 199588 143632 199640
rect 143684 199600 143718 199640
rect 143684 199588 143690 199600
rect 143442 199520 143448 199572
rect 143500 199532 143534 199572
rect 143500 199520 143506 199532
rect 144058 199504 144086 199860
rect 144242 199764 144270 199860
rect 144196 199736 144270 199764
rect 144196 199640 144224 199736
rect 144334 199708 144362 199860
rect 144886 199764 144914 199860
rect 144270 199656 144276 199708
rect 144328 199668 144362 199708
rect 144472 199736 144914 199764
rect 144328 199656 144334 199668
rect 144178 199588 144184 199640
rect 144236 199588 144242 199640
rect 144472 199628 144500 199736
rect 144472 199600 144592 199628
rect 144564 199572 144592 199600
rect 144822 199588 144828 199640
rect 144880 199628 144886 199640
rect 144978 199628 145006 199872
rect 145420 199860 145426 199872
rect 145478 199860 145484 199912
rect 145512 199860 145518 199912
rect 145570 199860 145576 199912
rect 145788 199860 145794 199912
rect 145846 199860 145852 199912
rect 145972 199860 145978 199912
rect 146030 199860 146036 199912
rect 147352 199900 147358 199912
rect 146266 199872 147358 199900
rect 145236 199792 145242 199844
rect 145294 199792 145300 199844
rect 145328 199792 145334 199844
rect 145386 199832 145392 199844
rect 145386 199792 145420 199832
rect 145254 199708 145282 199792
rect 145392 199708 145420 199792
rect 145254 199668 145288 199708
rect 145282 199656 145288 199668
rect 145340 199656 145346 199708
rect 145374 199656 145380 199708
rect 145432 199656 145438 199708
rect 145530 199696 145558 199860
rect 145806 199776 145834 199860
rect 145742 199724 145748 199776
rect 145800 199736 145834 199776
rect 145800 199724 145806 199736
rect 145530 199668 145604 199696
rect 145576 199640 145604 199668
rect 144880 199600 145006 199628
rect 144880 199588 144886 199600
rect 145558 199588 145564 199640
rect 145616 199588 145622 199640
rect 144546 199520 144552 199572
rect 144604 199520 144610 199572
rect 141844 199464 141970 199492
rect 141844 199452 141850 199464
rect 143994 199452 144000 199504
rect 144052 199464 144086 199504
rect 144052 199452 144058 199464
rect 145990 199424 146018 199860
rect 140516 199396 146018 199424
rect 112990 199316 112996 199368
rect 113048 199356 113054 199368
rect 113048 199328 141648 199356
rect 113048 199316 113054 199328
rect 115750 199248 115756 199300
rect 115808 199288 115814 199300
rect 140038 199288 140044 199300
rect 115808 199260 140044 199288
rect 115808 199248 115814 199260
rect 140038 199248 140044 199260
rect 140096 199248 140102 199300
rect 141620 199288 141648 199328
rect 146266 199288 146294 199872
rect 147352 199860 147358 199872
rect 147410 199860 147416 199912
rect 147536 199860 147542 199912
rect 147594 199860 147600 199912
rect 148088 199860 148094 199912
rect 148146 199860 148152 199912
rect 148272 199860 148278 199912
rect 148330 199860 148336 199912
rect 148640 199900 148646 199912
rect 148382 199872 148646 199900
rect 147554 199832 147582 199860
rect 147232 199804 147582 199832
rect 147232 199492 147260 199804
rect 148106 199776 148134 199860
rect 148106 199736 148140 199776
rect 148134 199724 148140 199736
rect 148192 199724 148198 199776
rect 147674 199588 147680 199640
rect 147732 199628 147738 199640
rect 148290 199628 148318 199860
rect 147732 199600 148318 199628
rect 147732 199588 147738 199600
rect 148226 199520 148232 199572
rect 148284 199560 148290 199572
rect 148382 199560 148410 199872
rect 148640 199860 148646 199872
rect 148698 199860 148704 199912
rect 148732 199860 148738 199912
rect 148790 199860 148796 199912
rect 148824 199860 148830 199912
rect 148882 199860 148888 199912
rect 148916 199860 148922 199912
rect 148974 199860 148980 199912
rect 149100 199900 149106 199912
rect 149072 199860 149106 199900
rect 149158 199860 149164 199912
rect 149192 199860 149198 199912
rect 149250 199860 149256 199912
rect 149376 199860 149382 199912
rect 149434 199860 149440 199912
rect 149652 199860 149658 199912
rect 149710 199860 149716 199912
rect 150020 199900 150026 199912
rect 149946 199872 150026 199900
rect 148750 199832 148778 199860
rect 148704 199804 148778 199832
rect 148704 199776 148732 199804
rect 148842 199776 148870 199860
rect 148686 199724 148692 199776
rect 148744 199724 148750 199776
rect 148778 199724 148784 199776
rect 148836 199736 148870 199776
rect 148836 199724 148842 199736
rect 148934 199708 148962 199860
rect 149072 199776 149100 199860
rect 149210 199832 149238 199860
rect 149164 199804 149238 199832
rect 149164 199776 149192 199804
rect 149054 199724 149060 199776
rect 149112 199724 149118 199776
rect 149146 199724 149152 199776
rect 149204 199724 149210 199776
rect 149238 199724 149244 199776
rect 149296 199764 149302 199776
rect 149394 199764 149422 199860
rect 149296 199736 149422 199764
rect 149296 199724 149302 199736
rect 148870 199656 148876 199708
rect 148928 199668 148962 199708
rect 148928 199656 148934 199668
rect 149330 199656 149336 199708
rect 149388 199696 149394 199708
rect 149670 199696 149698 199860
rect 149388 199668 149698 199696
rect 149388 199656 149394 199668
rect 149836 199656 149842 199708
rect 149894 199656 149900 199708
rect 149514 199588 149520 199640
rect 149572 199628 149578 199640
rect 149854 199628 149882 199656
rect 149572 199600 149882 199628
rect 149572 199588 149578 199600
rect 148284 199532 148410 199560
rect 148284 199520 148290 199532
rect 149946 199504 149974 199872
rect 150020 199860 150026 199872
rect 150078 199860 150084 199912
rect 150112 199860 150118 199912
rect 150170 199860 150176 199912
rect 150756 199860 150762 199912
rect 150814 199860 150820 199912
rect 151216 199860 151222 199912
rect 151274 199860 151280 199912
rect 151400 199860 151406 199912
rect 151458 199860 151464 199912
rect 151584 199860 151590 199912
rect 151642 199860 151648 199912
rect 151676 199860 151682 199912
rect 151734 199860 151740 199912
rect 151952 199860 151958 199912
rect 152010 199860 152016 199912
rect 152044 199860 152050 199912
rect 152102 199860 152108 199912
rect 152412 199860 152418 199912
rect 152470 199860 152476 199912
rect 152596 199860 152602 199912
rect 152654 199860 152660 199912
rect 152964 199860 152970 199912
rect 153022 199860 153028 199912
rect 153240 199860 153246 199912
rect 153298 199900 153304 199912
rect 153298 199872 153470 199900
rect 153298 199860 153304 199872
rect 150130 199708 150158 199860
rect 150388 199724 150394 199776
rect 150446 199724 150452 199776
rect 150066 199656 150072 199708
rect 150124 199668 150158 199708
rect 150406 199696 150434 199724
rect 150360 199668 150434 199696
rect 150774 199696 150802 199860
rect 151234 199776 151262 199860
rect 151170 199724 151176 199776
rect 151228 199736 151262 199776
rect 151228 199724 151234 199736
rect 151418 199696 151446 199860
rect 150774 199668 150848 199696
rect 150124 199656 150130 199668
rect 150360 199640 150388 199668
rect 150820 199640 150848 199668
rect 151004 199668 151446 199696
rect 151602 199708 151630 199860
rect 151694 199764 151722 199860
rect 151694 199736 151768 199764
rect 151602 199668 151636 199708
rect 150342 199588 150348 199640
rect 150400 199588 150406 199640
rect 150802 199588 150808 199640
rect 150860 199588 150866 199640
rect 151004 199560 151032 199668
rect 151630 199656 151636 199668
rect 151688 199656 151694 199708
rect 151078 199588 151084 199640
rect 151136 199628 151142 199640
rect 151740 199628 151768 199736
rect 151136 199600 151768 199628
rect 151136 199588 151142 199600
rect 151446 199560 151452 199572
rect 151004 199532 151452 199560
rect 151446 199520 151452 199532
rect 151504 199520 151510 199572
rect 151538 199520 151544 199572
rect 151596 199560 151602 199572
rect 151970 199560 151998 199860
rect 151596 199532 151998 199560
rect 151596 199520 151602 199532
rect 147490 199492 147496 199504
rect 147232 199464 147496 199492
rect 147490 199452 147496 199464
rect 147548 199452 147554 199504
rect 149882 199452 149888 199504
rect 149940 199464 149974 199504
rect 152062 199492 152090 199860
rect 152430 199640 152458 199860
rect 152430 199600 152464 199640
rect 152458 199588 152464 199600
rect 152516 199588 152522 199640
rect 152182 199492 152188 199504
rect 152062 199464 152188 199492
rect 149940 199452 149946 199464
rect 152182 199452 152188 199464
rect 152240 199452 152246 199504
rect 152614 199492 152642 199860
rect 152826 199520 152832 199572
rect 152884 199560 152890 199572
rect 152982 199560 153010 199860
rect 153332 199792 153338 199844
rect 153390 199792 153396 199844
rect 152884 199532 153010 199560
rect 152884 199520 152890 199532
rect 153350 199504 153378 199792
rect 153194 199492 153200 199504
rect 152614 199464 153200 199492
rect 153194 199452 153200 199464
rect 153252 199452 153258 199504
rect 153286 199452 153292 199504
rect 153344 199464 153378 199504
rect 153344 199452 153350 199464
rect 153442 199436 153470 199872
rect 153516 199860 153522 199912
rect 153574 199860 153580 199912
rect 153608 199860 153614 199912
rect 153666 199860 153672 199912
rect 153976 199860 153982 199912
rect 154034 199860 154040 199912
rect 154068 199860 154074 199912
rect 154126 199860 154132 199912
rect 154160 199860 154166 199912
rect 154218 199860 154224 199912
rect 154252 199860 154258 199912
rect 154310 199900 154316 199912
rect 154310 199860 154344 199900
rect 154528 199860 154534 199912
rect 154586 199860 154592 199912
rect 154620 199860 154626 199912
rect 154678 199860 154684 199912
rect 154896 199860 154902 199912
rect 154954 199860 154960 199912
rect 155080 199860 155086 199912
rect 155138 199860 155144 199912
rect 155172 199860 155178 199912
rect 155230 199860 155236 199912
rect 155264 199860 155270 199912
rect 155322 199900 155328 199912
rect 155322 199872 155448 199900
rect 155322 199860 155328 199872
rect 153534 199776 153562 199860
rect 153626 199832 153654 199860
rect 153626 199804 153700 199832
rect 153534 199736 153568 199776
rect 153562 199724 153568 199736
rect 153620 199724 153626 199776
rect 153672 199640 153700 199804
rect 153994 199708 154022 199860
rect 154086 199776 154114 199860
rect 154178 199832 154206 199860
rect 154178 199804 154252 199832
rect 154224 199776 154252 199804
rect 154086 199736 154120 199776
rect 154114 199724 154120 199736
rect 154172 199724 154178 199776
rect 154206 199724 154212 199776
rect 154264 199724 154270 199776
rect 153994 199668 154028 199708
rect 154022 199656 154028 199668
rect 154080 199656 154086 199708
rect 154316 199640 154344 199860
rect 154546 199832 154574 199860
rect 154500 199804 154574 199832
rect 154500 199776 154528 199804
rect 154638 199776 154666 199860
rect 154482 199724 154488 199776
rect 154540 199724 154546 199776
rect 154574 199724 154580 199776
rect 154632 199736 154666 199776
rect 154632 199724 154638 199736
rect 153654 199588 153660 199640
rect 153712 199588 153718 199640
rect 154298 199588 154304 199640
rect 154356 199588 154362 199640
rect 154914 199628 154942 199860
rect 155098 199776 155126 199860
rect 155190 199832 155218 199860
rect 155190 199804 155264 199832
rect 155236 199776 155264 199804
rect 155098 199736 155132 199776
rect 155126 199724 155132 199736
rect 155184 199724 155190 199776
rect 155218 199724 155224 199776
rect 155276 199724 155282 199776
rect 155034 199628 155040 199640
rect 154914 199600 155040 199628
rect 155034 199588 155040 199600
rect 155092 199588 155098 199640
rect 155420 199572 155448 199872
rect 155540 199860 155546 199912
rect 155598 199860 155604 199912
rect 156184 199860 156190 199912
rect 156242 199860 156248 199912
rect 156276 199860 156282 199912
rect 156334 199860 156340 199912
rect 156368 199860 156374 199912
rect 156426 199900 156432 199912
rect 156426 199860 156460 199900
rect 156736 199860 156742 199912
rect 156794 199860 156800 199912
rect 157012 199900 157018 199912
rect 156984 199860 157018 199900
rect 157070 199860 157076 199912
rect 157104 199860 157110 199912
rect 157162 199860 157168 199912
rect 157380 199860 157386 199912
rect 157438 199860 157444 199912
rect 157564 199860 157570 199912
rect 157622 199860 157628 199912
rect 157656 199860 157662 199912
rect 157714 199860 157720 199912
rect 157748 199860 157754 199912
rect 157806 199860 157812 199912
rect 157932 199860 157938 199912
rect 157990 199860 157996 199912
rect 158392 199860 158398 199912
rect 158450 199860 158456 199912
rect 158760 199860 158766 199912
rect 158818 199860 158824 199912
rect 158944 199860 158950 199912
rect 159002 199860 159008 199912
rect 159404 199900 159410 199912
rect 159376 199860 159410 199900
rect 159462 199860 159468 199912
rect 159496 199860 159502 199912
rect 159554 199860 159560 199912
rect 160324 199860 160330 199912
rect 160382 199860 160388 199912
rect 160416 199860 160422 199912
rect 160474 199860 160480 199912
rect 160600 199860 160606 199912
rect 160658 199860 160664 199912
rect 161888 199900 161894 199912
rect 160848 199872 161894 199900
rect 155558 199572 155586 199860
rect 156202 199776 156230 199860
rect 156294 199832 156322 199860
rect 156294 199804 156368 199832
rect 156340 199776 156368 199804
rect 156202 199736 156236 199776
rect 156230 199724 156236 199736
rect 156288 199724 156294 199776
rect 156322 199724 156328 199776
rect 156380 199724 156386 199776
rect 156432 199708 156460 199860
rect 156414 199656 156420 199708
rect 156472 199656 156478 199708
rect 156754 199640 156782 199860
rect 156984 199696 157012 199860
rect 157122 199776 157150 199860
rect 157058 199724 157064 199776
rect 157116 199736 157150 199776
rect 157116 199724 157122 199736
rect 157150 199696 157156 199708
rect 156984 199668 157156 199696
rect 157150 199656 157156 199668
rect 157208 199656 157214 199708
rect 156690 199588 156696 199640
rect 156748 199600 156782 199640
rect 156748 199588 156754 199600
rect 155402 199520 155408 199572
rect 155460 199520 155466 199572
rect 155558 199532 155592 199572
rect 155586 199520 155592 199532
rect 155644 199520 155650 199572
rect 153378 199384 153384 199436
rect 153436 199396 153470 199436
rect 153436 199384 153442 199396
rect 157398 199356 157426 199860
rect 157582 199492 157610 199860
rect 157674 199708 157702 199860
rect 157766 199764 157794 199860
rect 157766 199736 157840 199764
rect 157674 199668 157708 199708
rect 157702 199656 157708 199668
rect 157760 199656 157766 199708
rect 157812 199560 157840 199736
rect 157950 199640 157978 199860
rect 158410 199776 158438 199860
rect 158346 199724 158352 199776
rect 158404 199736 158438 199776
rect 158404 199724 158410 199736
rect 157886 199588 157892 199640
rect 157944 199600 157978 199640
rect 157944 199588 157950 199600
rect 158778 199572 158806 199860
rect 158962 199696 158990 199860
rect 158916 199668 158990 199696
rect 158916 199640 158944 199668
rect 158898 199588 158904 199640
rect 158956 199588 158962 199640
rect 158254 199560 158260 199572
rect 157812 199532 158260 199560
rect 158254 199520 158260 199532
rect 158312 199520 158318 199572
rect 158778 199532 158812 199572
rect 158806 199520 158812 199532
rect 158864 199520 158870 199572
rect 159174 199520 159180 199572
rect 159232 199560 159238 199572
rect 159376 199560 159404 199860
rect 159514 199832 159542 199860
rect 159468 199804 159542 199832
rect 159468 199776 159496 199804
rect 160232 199792 160238 199844
rect 160290 199792 160296 199844
rect 159450 199724 159456 199776
rect 159508 199724 159514 199776
rect 160250 199708 160278 199792
rect 160186 199656 160192 199708
rect 160244 199668 160278 199708
rect 160244 199656 160250 199668
rect 160342 199640 160370 199860
rect 160278 199588 160284 199640
rect 160336 199600 160370 199640
rect 160434 199640 160462 199860
rect 160434 199600 160468 199640
rect 160336 199588 160342 199600
rect 160462 199588 160468 199600
rect 160520 199588 160526 199640
rect 159232 199532 159404 199560
rect 159232 199520 159238 199532
rect 157702 199492 157708 199504
rect 157582 199464 157708 199492
rect 157702 199452 157708 199464
rect 157760 199452 157766 199504
rect 158530 199356 158536 199368
rect 157398 199328 158536 199356
rect 158530 199316 158536 199328
rect 158588 199316 158594 199368
rect 160618 199356 160646 199860
rect 160848 199572 160876 199872
rect 161888 199860 161894 199872
rect 161946 199860 161952 199912
rect 161980 199860 161986 199912
rect 162038 199860 162044 199912
rect 162164 199900 162170 199912
rect 162136 199860 162170 199900
rect 162222 199860 162228 199912
rect 162256 199860 162262 199912
rect 162314 199860 162320 199912
rect 162348 199860 162354 199912
rect 162406 199860 162412 199912
rect 162440 199860 162446 199912
rect 162498 199860 162504 199912
rect 162532 199860 162538 199912
rect 162590 199860 162596 199912
rect 162808 199860 162814 199912
rect 162866 199900 162872 199912
rect 162866 199872 163314 199900
rect 162866 199860 162872 199872
rect 160968 199832 160974 199844
rect 160940 199792 160974 199832
rect 161026 199792 161032 199844
rect 161520 199792 161526 199844
rect 161578 199792 161584 199844
rect 161998 199832 162026 199860
rect 161952 199804 162026 199832
rect 160940 199708 160968 199792
rect 161152 199724 161158 199776
rect 161210 199724 161216 199776
rect 161244 199724 161250 199776
rect 161302 199724 161308 199776
rect 160922 199656 160928 199708
rect 160980 199656 160986 199708
rect 160830 199520 160836 199572
rect 160888 199520 160894 199572
rect 161170 199424 161198 199724
rect 161262 199572 161290 199724
rect 161538 199572 161566 199792
rect 161952 199776 161980 199804
rect 161934 199724 161940 199776
rect 161992 199724 161998 199776
rect 162136 199640 162164 199860
rect 162274 199832 162302 199860
rect 162228 199804 162302 199832
rect 162228 199708 162256 199804
rect 162366 199708 162394 199860
rect 162210 199656 162216 199708
rect 162268 199656 162274 199708
rect 162302 199656 162308 199708
rect 162360 199668 162394 199708
rect 162458 199708 162486 199860
rect 162550 199776 162578 199860
rect 163084 199832 163090 199844
rect 163056 199792 163090 199832
rect 163142 199792 163148 199844
rect 163176 199792 163182 199844
rect 163234 199792 163240 199844
rect 162550 199736 162584 199776
rect 162578 199724 162584 199736
rect 162636 199724 162642 199776
rect 162900 199724 162906 199776
rect 162958 199764 162964 199776
rect 162958 199724 162992 199764
rect 162458 199668 162492 199708
rect 162360 199656 162366 199668
rect 162486 199656 162492 199668
rect 162544 199656 162550 199708
rect 162118 199588 162124 199640
rect 162176 199588 162182 199640
rect 162964 199572 162992 199724
rect 163056 199640 163084 199792
rect 163194 199708 163222 199792
rect 163130 199656 163136 199708
rect 163188 199668 163222 199708
rect 163188 199656 163194 199668
rect 163038 199588 163044 199640
rect 163096 199588 163102 199640
rect 163286 199572 163314 199872
rect 163360 199860 163366 199912
rect 163418 199860 163424 199912
rect 163544 199860 163550 199912
rect 163602 199860 163608 199912
rect 163636 199860 163642 199912
rect 163694 199860 163700 199912
rect 164004 199900 164010 199912
rect 163930 199872 164010 199900
rect 163378 199708 163406 199860
rect 163378 199668 163412 199708
rect 163406 199656 163412 199668
rect 163464 199656 163470 199708
rect 163562 199640 163590 199860
rect 163654 199776 163682 199860
rect 163820 199792 163826 199844
rect 163878 199792 163884 199844
rect 163654 199736 163688 199776
rect 163682 199724 163688 199736
rect 163740 199724 163746 199776
rect 163498 199588 163504 199640
rect 163556 199600 163590 199640
rect 163556 199588 163562 199600
rect 161262 199532 161296 199572
rect 161290 199520 161296 199532
rect 161348 199520 161354 199572
rect 161474 199520 161480 199572
rect 161532 199532 161566 199572
rect 161532 199520 161538 199532
rect 162946 199520 162952 199572
rect 163004 199520 163010 199572
rect 163286 199532 163320 199572
rect 163314 199520 163320 199532
rect 163372 199520 163378 199572
rect 163590 199520 163596 199572
rect 163648 199560 163654 199572
rect 163838 199560 163866 199792
rect 163648 199532 163866 199560
rect 163648 199520 163654 199532
rect 163930 199504 163958 199872
rect 164004 199860 164010 199872
rect 164062 199860 164068 199912
rect 164096 199860 164102 199912
rect 164154 199860 164160 199912
rect 164188 199860 164194 199912
rect 164246 199860 164252 199912
rect 164280 199860 164286 199912
rect 164338 199860 164344 199912
rect 164372 199860 164378 199912
rect 164430 199860 164436 199912
rect 164464 199860 164470 199912
rect 164522 199900 164528 199912
rect 164832 199900 164838 199912
rect 164522 199872 164694 199900
rect 164522 199860 164528 199872
rect 164114 199832 164142 199860
rect 164068 199804 164142 199832
rect 164068 199708 164096 199804
rect 164206 199708 164234 199860
rect 164050 199656 164056 199708
rect 164108 199656 164114 199708
rect 164142 199656 164148 199708
rect 164200 199668 164234 199708
rect 164200 199656 164206 199668
rect 164298 199640 164326 199860
rect 164390 199708 164418 199860
rect 164556 199832 164562 199844
rect 164528 199792 164562 199832
rect 164614 199792 164620 199844
rect 164528 199708 164556 199792
rect 164390 199668 164424 199708
rect 164418 199656 164424 199668
rect 164476 199656 164482 199708
rect 164510 199656 164516 199708
rect 164568 199656 164574 199708
rect 164234 199588 164240 199640
rect 164292 199600 164326 199640
rect 164292 199588 164298 199600
rect 164666 199572 164694 199872
rect 164804 199860 164838 199900
rect 164890 199860 164896 199912
rect 164924 199860 164930 199912
rect 164982 199860 164988 199912
rect 165016 199860 165022 199912
rect 165074 199860 165080 199912
rect 165108 199860 165114 199912
rect 165166 199860 165172 199912
rect 165476 199860 165482 199912
rect 165534 199860 165540 199912
rect 165844 199860 165850 199912
rect 165902 199860 165908 199912
rect 166028 199900 166034 199912
rect 166000 199860 166034 199900
rect 166086 199860 166092 199912
rect 166120 199860 166126 199912
rect 166178 199860 166184 199912
rect 166212 199860 166218 199912
rect 166270 199860 166276 199912
rect 166304 199860 166310 199912
rect 166362 199860 166368 199912
rect 166488 199860 166494 199912
rect 166546 199860 166552 199912
rect 166856 199860 166862 199912
rect 166914 199860 166920 199912
rect 167224 199860 167230 199912
rect 167282 199860 167288 199912
rect 167408 199860 167414 199912
rect 167466 199860 167472 199912
rect 167500 199860 167506 199912
rect 167558 199860 167564 199912
rect 167592 199860 167598 199912
rect 167650 199900 167656 199912
rect 167960 199900 167966 199912
rect 167650 199872 167868 199900
rect 167650 199860 167656 199872
rect 164804 199776 164832 199860
rect 164942 199832 164970 199860
rect 164896 199804 164970 199832
rect 164786 199724 164792 199776
rect 164844 199724 164850 199776
rect 164896 199708 164924 199804
rect 165034 199764 165062 199860
rect 164988 199736 165062 199764
rect 164988 199708 165016 199736
rect 165126 199708 165154 199860
rect 164878 199656 164884 199708
rect 164936 199656 164942 199708
rect 164970 199656 164976 199708
rect 165028 199656 165034 199708
rect 165062 199656 165068 199708
rect 165120 199668 165154 199708
rect 165120 199656 165126 199668
rect 165494 199640 165522 199860
rect 165660 199792 165666 199844
rect 165718 199792 165724 199844
rect 165678 199640 165706 199792
rect 165476 199588 165482 199640
rect 165534 199588 165540 199640
rect 165678 199600 165712 199640
rect 165706 199588 165712 199600
rect 165764 199588 165770 199640
rect 164666 199532 164700 199572
rect 164694 199520 164700 199532
rect 164752 199520 164758 199572
rect 165862 199560 165890 199860
rect 166000 199640 166028 199860
rect 166138 199764 166166 199860
rect 166092 199736 166166 199764
rect 166092 199708 166120 199736
rect 166230 199708 166258 199860
rect 166074 199656 166080 199708
rect 166132 199656 166138 199708
rect 166166 199656 166172 199708
rect 166224 199668 166258 199708
rect 166224 199656 166230 199668
rect 166322 199640 166350 199860
rect 165982 199588 165988 199640
rect 166040 199588 166046 199640
rect 166322 199600 166356 199640
rect 166350 199588 166356 199600
rect 166408 199588 166414 199640
rect 166506 199572 166534 199860
rect 166672 199792 166678 199844
rect 166730 199792 166736 199844
rect 166764 199792 166770 199844
rect 166822 199792 166828 199844
rect 166690 199640 166718 199792
rect 166782 199708 166810 199792
rect 166874 199776 166902 199860
rect 167132 199792 167138 199844
rect 167190 199792 167196 199844
rect 166874 199736 166908 199776
rect 166902 199724 166908 199736
rect 166960 199724 166966 199776
rect 166782 199668 166816 199708
rect 166810 199656 166816 199668
rect 166868 199656 166874 199708
rect 166690 199600 166724 199640
rect 166718 199588 166724 199600
rect 166776 199588 166782 199640
rect 167150 199572 167178 199792
rect 167242 199640 167270 199860
rect 167242 199600 167276 199640
rect 167270 199588 167276 199600
rect 167328 199588 167334 199640
rect 167426 199628 167454 199860
rect 167518 199832 167546 199860
rect 167518 199804 167592 199832
rect 167564 199696 167592 199804
rect 167564 199668 167638 199696
rect 167380 199600 167454 199628
rect 166258 199560 166264 199572
rect 165862 199532 166264 199560
rect 166258 199520 166264 199532
rect 166316 199520 166322 199572
rect 166506 199532 166540 199572
rect 166534 199520 166540 199532
rect 166592 199520 166598 199572
rect 167150 199532 167184 199572
rect 167178 199520 167184 199532
rect 167236 199520 167242 199572
rect 163866 199452 163872 199504
rect 163924 199464 163958 199504
rect 163924 199452 163930 199464
rect 165430 199424 165436 199436
rect 161170 199396 165436 199424
rect 165430 199384 165436 199396
rect 165488 199384 165494 199436
rect 166258 199356 166264 199368
rect 160618 199328 166264 199356
rect 166258 199316 166264 199328
rect 166316 199316 166322 199368
rect 167380 199356 167408 199600
rect 167454 199520 167460 199572
rect 167512 199560 167518 199572
rect 167610 199560 167638 199668
rect 167512 199532 167638 199560
rect 167512 199520 167518 199532
rect 167840 199424 167868 199872
rect 167932 199860 167966 199900
rect 168018 199860 168024 199912
rect 168328 199860 168334 199912
rect 168386 199860 168392 199912
rect 168512 199860 168518 199912
rect 168570 199860 168576 199912
rect 168696 199860 168702 199912
rect 168754 199860 168760 199912
rect 168972 199860 168978 199912
rect 169030 199860 169036 199912
rect 169064 199860 169070 199912
rect 169122 199860 169128 199912
rect 169156 199860 169162 199912
rect 169214 199860 169220 199912
rect 169340 199860 169346 199912
rect 169398 199860 169404 199912
rect 169432 199860 169438 199912
rect 169490 199860 169496 199912
rect 169984 199900 169990 199912
rect 169680 199872 169990 199900
rect 167932 199492 167960 199860
rect 168144 199832 168150 199844
rect 168024 199804 168150 199832
rect 168024 199628 168052 199804
rect 168144 199792 168150 199804
rect 168202 199792 168208 199844
rect 168346 199708 168374 199860
rect 168282 199656 168288 199708
rect 168340 199668 168374 199708
rect 168340 199656 168346 199668
rect 168190 199628 168196 199640
rect 168024 199600 168196 199628
rect 168190 199588 168196 199600
rect 168248 199588 168254 199640
rect 168530 199628 168558 199860
rect 168714 199696 168742 199860
rect 168990 199708 169018 199860
rect 168714 199668 168880 199696
rect 168742 199628 168748 199640
rect 168530 199600 168748 199628
rect 168742 199588 168748 199600
rect 168800 199588 168806 199640
rect 168466 199520 168472 199572
rect 168524 199560 168530 199572
rect 168852 199560 168880 199668
rect 168926 199656 168932 199708
rect 168984 199668 169018 199708
rect 168984 199656 168990 199668
rect 168524 199532 168880 199560
rect 169082 199572 169110 199860
rect 169174 199764 169202 199860
rect 169174 199736 169248 199764
rect 169220 199640 169248 199736
rect 169358 199696 169386 199860
rect 169312 199668 169386 199696
rect 169312 199640 169340 199668
rect 169202 199588 169208 199640
rect 169260 199588 169266 199640
rect 169294 199588 169300 199640
rect 169352 199588 169358 199640
rect 169450 199572 169478 199860
rect 169680 199640 169708 199872
rect 169984 199860 169990 199872
rect 170042 199860 170048 199912
rect 170076 199860 170082 199912
rect 170134 199860 170140 199912
rect 170168 199860 170174 199912
rect 170226 199860 170232 199912
rect 170260 199860 170266 199912
rect 170318 199860 170324 199912
rect 170444 199860 170450 199912
rect 170502 199860 170508 199912
rect 170720 199900 170726 199912
rect 170600 199872 170726 199900
rect 169800 199792 169806 199844
rect 169858 199792 169864 199844
rect 170094 199832 170122 199860
rect 169956 199804 170122 199832
rect 169662 199588 169668 199640
rect 169720 199588 169726 199640
rect 169082 199532 169116 199572
rect 168524 199520 168530 199532
rect 169110 199520 169116 199532
rect 169168 199520 169174 199572
rect 169386 199520 169392 199572
rect 169444 199532 169478 199572
rect 169818 199560 169846 199792
rect 169956 199628 169984 199804
rect 170030 199656 170036 199708
rect 170088 199696 170094 199708
rect 170186 199696 170214 199860
rect 170088 199668 170214 199696
rect 170088 199656 170094 199668
rect 170278 199640 170306 199860
rect 170122 199628 170128 199640
rect 169956 199600 170128 199628
rect 170122 199588 170128 199600
rect 170180 199588 170186 199640
rect 170214 199588 170220 199640
rect 170272 199600 170306 199640
rect 170272 199588 170278 199600
rect 169938 199560 169944 199572
rect 169818 199532 169944 199560
rect 169444 199520 169450 199532
rect 169938 199520 169944 199532
rect 169996 199520 170002 199572
rect 170462 199560 170490 199860
rect 170600 199640 170628 199872
rect 170720 199860 170726 199872
rect 170778 199860 170784 199912
rect 170812 199860 170818 199912
rect 170870 199860 170876 199912
rect 170904 199860 170910 199912
rect 170962 199860 170968 199912
rect 171088 199900 171094 199912
rect 171060 199860 171094 199900
rect 171146 199900 171152 199912
rect 171146 199872 171193 199900
rect 171146 199860 171152 199872
rect 171272 199860 171278 199912
rect 171330 199860 171336 199912
rect 171364 199860 171370 199912
rect 171422 199860 171428 199912
rect 171456 199860 171462 199912
rect 171514 199860 171520 199912
rect 171640 199860 171646 199912
rect 171698 199860 171704 199912
rect 171732 199860 171738 199912
rect 171790 199860 171796 199912
rect 171824 199860 171830 199912
rect 171882 199860 171888 199912
rect 171916 199860 171922 199912
rect 171974 199860 171980 199912
rect 172008 199860 172014 199912
rect 172066 199860 172072 199912
rect 172192 199900 172198 199912
rect 172164 199860 172198 199900
rect 172250 199860 172256 199912
rect 172376 199860 172382 199912
rect 172434 199860 172440 199912
rect 172560 199860 172566 199912
rect 172618 199860 172624 199912
rect 172652 199860 172658 199912
rect 172710 199860 172716 199912
rect 172744 199860 172750 199912
rect 172802 199860 172808 199912
rect 172928 199860 172934 199912
rect 172986 199860 172992 199912
rect 173020 199860 173026 199912
rect 173078 199860 173084 199912
rect 173112 199860 173118 199912
rect 173170 199900 173176 199912
rect 173296 199900 173302 199912
rect 173170 199860 173204 199900
rect 170830 199776 170858 199860
rect 170766 199724 170772 199776
rect 170824 199736 170858 199776
rect 170824 199724 170830 199736
rect 170582 199588 170588 199640
rect 170640 199588 170646 199640
rect 170674 199560 170680 199572
rect 170462 199532 170680 199560
rect 170674 199520 170680 199532
rect 170732 199520 170738 199572
rect 167932 199464 168052 199492
rect 167914 199424 167920 199436
rect 167840 199396 167920 199424
rect 167914 199384 167920 199396
rect 167972 199384 167978 199436
rect 167638 199356 167644 199368
rect 167380 199328 167644 199356
rect 167638 199316 167644 199328
rect 167696 199316 167702 199368
rect 141620 199260 146294 199288
rect 151354 199248 151360 199300
rect 151412 199288 151418 199300
rect 162394 199288 162400 199300
rect 151412 199260 162400 199288
rect 151412 199248 151418 199260
rect 162394 199248 162400 199260
rect 162452 199248 162458 199300
rect 167546 199248 167552 199300
rect 167604 199288 167610 199300
rect 168024 199288 168052 199464
rect 170030 199452 170036 199504
rect 170088 199492 170094 199504
rect 170922 199492 170950 199860
rect 171060 199776 171088 199860
rect 171290 199832 171318 199860
rect 171244 199804 171318 199832
rect 171042 199724 171048 199776
rect 171100 199724 171106 199776
rect 171244 199640 171272 199804
rect 171382 199764 171410 199860
rect 171336 199736 171410 199764
rect 171336 199708 171364 199736
rect 171474 199708 171502 199860
rect 171658 199776 171686 199860
rect 171594 199724 171600 199776
rect 171652 199736 171686 199776
rect 171652 199724 171658 199736
rect 171318 199656 171324 199708
rect 171376 199656 171382 199708
rect 171410 199656 171416 199708
rect 171468 199668 171502 199708
rect 171468 199656 171474 199668
rect 171750 199640 171778 199860
rect 171842 199708 171870 199860
rect 171934 199764 171962 199860
rect 172026 199832 172054 199860
rect 172026 199804 172100 199832
rect 171934 199736 172008 199764
rect 171980 199708 172008 199736
rect 171842 199668 171876 199708
rect 171870 199656 171876 199668
rect 171928 199656 171934 199708
rect 171962 199656 171968 199708
rect 172020 199656 172026 199708
rect 171226 199588 171232 199640
rect 171284 199588 171290 199640
rect 171686 199588 171692 199640
rect 171744 199600 171778 199640
rect 171744 199588 171750 199600
rect 171778 199520 171784 199572
rect 171836 199560 171842 199572
rect 172072 199560 172100 199804
rect 172164 199640 172192 199860
rect 172394 199832 172422 199860
rect 172256 199804 172422 199832
rect 172256 199640 172284 199804
rect 172578 199708 172606 199860
rect 172670 199764 172698 199860
rect 172762 199832 172790 199860
rect 172762 199804 172836 199832
rect 172670 199736 172744 199764
rect 172716 199708 172744 199736
rect 172578 199668 172612 199708
rect 172606 199656 172612 199668
rect 172664 199656 172670 199708
rect 172698 199656 172704 199708
rect 172756 199656 172762 199708
rect 172146 199588 172152 199640
rect 172204 199588 172210 199640
rect 172238 199588 172244 199640
rect 172296 199588 172302 199640
rect 171836 199532 172100 199560
rect 171836 199520 171842 199532
rect 170088 199464 170950 199492
rect 172808 199492 172836 199804
rect 172946 199696 172974 199860
rect 173038 199776 173066 199860
rect 173176 199776 173204 199860
rect 173268 199860 173302 199900
rect 173354 199860 173360 199912
rect 173572 199900 173578 199912
rect 173544 199860 173578 199900
rect 173630 199860 173636 199912
rect 173664 199860 173670 199912
rect 173722 199860 173728 199912
rect 173848 199860 173854 199912
rect 173906 199860 173912 199912
rect 173940 199860 173946 199912
rect 173998 199860 174004 199912
rect 174400 199860 174406 199912
rect 174458 199860 174464 199912
rect 174584 199860 174590 199912
rect 174642 199860 174648 199912
rect 174768 199860 174774 199912
rect 174826 199860 174832 199912
rect 175136 199860 175142 199912
rect 175194 199860 175200 199912
rect 175228 199860 175234 199912
rect 175286 199900 175292 199912
rect 175286 199872 175412 199900
rect 175286 199860 175292 199872
rect 173038 199736 173072 199776
rect 173066 199724 173072 199736
rect 173124 199724 173130 199776
rect 173158 199724 173164 199776
rect 173216 199724 173222 199776
rect 172946 199668 173158 199696
rect 172882 199588 172888 199640
rect 172940 199628 172946 199640
rect 172940 199600 173020 199628
rect 172940 199588 172946 199600
rect 172992 199572 173020 199600
rect 172974 199520 172980 199572
rect 173032 199520 173038 199572
rect 172882 199492 172888 199504
rect 172808 199464 172888 199492
rect 170088 199452 170094 199464
rect 172882 199452 172888 199464
rect 172940 199452 172946 199504
rect 173130 199436 173158 199668
rect 173268 199628 173296 199860
rect 173342 199628 173348 199640
rect 173268 199600 173348 199628
rect 173342 199588 173348 199600
rect 173400 199588 173406 199640
rect 169754 199384 169760 199436
rect 169812 199424 169818 199436
rect 171502 199424 171508 199436
rect 169812 199396 171508 199424
rect 169812 199384 169818 199396
rect 171502 199384 171508 199396
rect 171560 199384 171566 199436
rect 173130 199396 173164 199436
rect 173158 199384 173164 199396
rect 173216 199384 173222 199436
rect 167604 199260 168052 199288
rect 173544 199288 173572 199860
rect 173682 199776 173710 199860
rect 173618 199724 173624 199776
rect 173676 199736 173710 199776
rect 173866 199764 173894 199860
rect 173820 199736 173894 199764
rect 173676 199724 173682 199736
rect 173820 199628 173848 199736
rect 173958 199708 173986 199860
rect 173894 199656 173900 199708
rect 173952 199668 173986 199708
rect 173952 199656 173958 199668
rect 174262 199628 174268 199640
rect 173820 199600 174268 199628
rect 174262 199588 174268 199600
rect 174320 199588 174326 199640
rect 174418 199492 174446 199860
rect 174602 199560 174630 199860
rect 174786 199628 174814 199860
rect 175154 199776 175182 199860
rect 175154 199736 175188 199776
rect 175182 199724 175188 199736
rect 175240 199724 175246 199776
rect 174906 199628 174912 199640
rect 174786 199600 174912 199628
rect 174906 199588 174912 199600
rect 174964 199588 174970 199640
rect 175274 199588 175280 199640
rect 175332 199588 175338 199640
rect 174602 199532 175228 199560
rect 174630 199492 174636 199504
rect 174418 199464 174636 199492
rect 174630 199452 174636 199464
rect 174688 199452 174694 199504
rect 174538 199384 174544 199436
rect 174596 199424 174602 199436
rect 175200 199424 175228 199532
rect 174596 199396 175228 199424
rect 175292 199424 175320 199588
rect 175384 199492 175412 199872
rect 175780 199860 175786 199912
rect 175838 199860 175844 199912
rect 176056 199860 176062 199912
rect 176114 199860 176120 199912
rect 176148 199860 176154 199912
rect 176206 199860 176212 199912
rect 176240 199860 176246 199912
rect 176298 199860 176304 199912
rect 176424 199860 176430 199912
rect 176482 199860 176488 199912
rect 176700 199860 176706 199912
rect 176758 199860 176764 199912
rect 176792 199860 176798 199912
rect 176850 199860 176856 199912
rect 176976 199860 176982 199912
rect 177034 199860 177040 199912
rect 177160 199860 177166 199912
rect 177218 199860 177224 199912
rect 177344 199860 177350 199912
rect 177402 199860 177408 199912
rect 177620 199860 177626 199912
rect 177678 199900 177684 199912
rect 177758 199900 177764 199912
rect 177678 199872 177764 199900
rect 177678 199860 177684 199872
rect 177758 199860 177764 199872
rect 177816 199860 177822 199912
rect 175688 199832 175694 199844
rect 175660 199792 175694 199832
rect 175746 199792 175752 199844
rect 175660 199572 175688 199792
rect 175798 199708 175826 199860
rect 176074 199708 176102 199860
rect 175734 199656 175740 199708
rect 175792 199668 175826 199708
rect 175792 199656 175798 199668
rect 176010 199656 176016 199708
rect 176068 199668 176102 199708
rect 176166 199708 176194 199860
rect 176258 199776 176286 199860
rect 176258 199736 176292 199776
rect 176286 199724 176292 199736
rect 176344 199724 176350 199776
rect 176442 199708 176470 199860
rect 176166 199668 176200 199708
rect 176068 199656 176074 199668
rect 176194 199656 176200 199668
rect 176252 199656 176258 199708
rect 176378 199656 176384 199708
rect 176436 199668 176470 199708
rect 176436 199656 176442 199668
rect 176718 199628 176746 199860
rect 176810 199776 176838 199860
rect 176810 199736 176844 199776
rect 176838 199724 176844 199736
rect 176896 199724 176902 199776
rect 176994 199708 177022 199860
rect 177178 199764 177206 199860
rect 177362 199832 177390 199860
rect 177850 199832 177856 199844
rect 177362 199804 177856 199832
rect 177850 199792 177856 199804
rect 177908 199792 177914 199844
rect 187234 199764 187240 199776
rect 177178 199736 187240 199764
rect 187234 199724 187240 199736
rect 187292 199724 187298 199776
rect 176930 199656 176936 199708
rect 176988 199668 177022 199708
rect 176988 199656 176994 199668
rect 179046 199628 179052 199640
rect 176718 199600 179052 199628
rect 179046 199588 179052 199600
rect 179104 199588 179110 199640
rect 175642 199520 175648 199572
rect 175700 199520 175706 199572
rect 201494 199492 201500 199504
rect 175384 199464 201500 199492
rect 201494 199452 201500 199464
rect 201552 199452 201558 199504
rect 175550 199424 175556 199436
rect 175292 199396 175556 199424
rect 174596 199384 174602 199396
rect 175550 199384 175556 199396
rect 175608 199384 175614 199436
rect 178954 199384 178960 199436
rect 179012 199424 179018 199436
rect 187142 199424 187148 199436
rect 179012 199396 187148 199424
rect 179012 199384 179018 199396
rect 187142 199384 187148 199396
rect 187200 199384 187206 199436
rect 174078 199316 174084 199368
rect 174136 199356 174142 199368
rect 183186 199356 183192 199368
rect 174136 199328 183192 199356
rect 174136 199316 174142 199328
rect 183186 199316 183192 199328
rect 183244 199316 183250 199368
rect 195606 199288 195612 199300
rect 173544 199260 195612 199288
rect 167604 199248 167610 199260
rect 195606 199248 195612 199260
rect 195664 199248 195670 199300
rect 118418 199180 118424 199232
rect 118476 199220 118482 199232
rect 148686 199220 148692 199232
rect 118476 199192 148692 199220
rect 118476 199180 118482 199192
rect 148686 199180 148692 199192
rect 148744 199180 148750 199232
rect 173802 199180 173808 199232
rect 173860 199220 173866 199232
rect 208578 199220 208584 199232
rect 173860 199192 208584 199220
rect 173860 199180 173866 199192
rect 208578 199180 208584 199192
rect 208636 199180 208642 199232
rect 117222 199112 117228 199164
rect 117280 199152 117286 199164
rect 117280 199124 141280 199152
rect 117280 199112 117286 199124
rect 114462 199044 114468 199096
rect 114520 199084 114526 199096
rect 141252 199084 141280 199124
rect 141326 199112 141332 199164
rect 141384 199152 141390 199164
rect 143902 199152 143908 199164
rect 141384 199124 143908 199152
rect 141384 199112 141390 199124
rect 143902 199112 143908 199124
rect 143960 199112 143966 199164
rect 158622 199112 158628 199164
rect 158680 199152 158686 199164
rect 180242 199152 180248 199164
rect 158680 199124 180248 199152
rect 158680 199112 158686 199124
rect 180242 199112 180248 199124
rect 180300 199112 180306 199164
rect 180794 199112 180800 199164
rect 180852 199152 180858 199164
rect 187050 199152 187056 199164
rect 180852 199124 187056 199152
rect 180852 199112 180858 199124
rect 187050 199112 187056 199124
rect 187108 199112 187114 199164
rect 148410 199084 148416 199096
rect 114520 199056 140912 199084
rect 141252 199056 148416 199084
rect 114520 199044 114526 199056
rect 111610 198976 111616 199028
rect 111668 199016 111674 199028
rect 140884 199016 140912 199056
rect 148410 199044 148416 199056
rect 148468 199044 148474 199096
rect 144822 199016 144828 199028
rect 111668 198988 140222 199016
rect 140884 198988 144828 199016
rect 111668 198976 111674 198988
rect 113082 198908 113088 198960
rect 113140 198948 113146 198960
rect 140194 198948 140222 198988
rect 144822 198976 144828 198988
rect 144880 198976 144886 199028
rect 169938 198976 169944 199028
rect 169996 199016 170002 199028
rect 174078 199016 174084 199028
rect 169996 198988 174084 199016
rect 169996 198976 170002 198988
rect 174078 198976 174084 198988
rect 174136 198976 174142 199028
rect 174722 198976 174728 199028
rect 174780 199016 174786 199028
rect 202414 199016 202420 199028
rect 174780 198988 202420 199016
rect 174780 198976 174786 198988
rect 202414 198976 202420 198988
rect 202472 198976 202478 199028
rect 142430 198948 142436 198960
rect 113140 198920 140130 198948
rect 140194 198920 142436 198948
rect 113140 198908 113146 198920
rect 136358 198840 136364 198892
rect 136416 198880 136422 198892
rect 136634 198880 136640 198892
rect 136416 198852 136640 198880
rect 136416 198840 136422 198852
rect 136634 198840 136640 198852
rect 136692 198840 136698 198892
rect 137830 198840 137836 198892
rect 137888 198880 137894 198892
rect 138934 198880 138940 198892
rect 137888 198852 138940 198880
rect 137888 198840 137894 198852
rect 138934 198840 138940 198852
rect 138992 198840 138998 198892
rect 140102 198880 140130 198920
rect 142430 198908 142436 198920
rect 142488 198908 142494 198960
rect 150710 198908 150716 198960
rect 150768 198948 150774 198960
rect 173802 198948 173808 198960
rect 150768 198920 173808 198948
rect 150768 198908 150774 198920
rect 173802 198908 173808 198920
rect 173860 198908 173866 198960
rect 142614 198880 142620 198892
rect 140102 198852 142620 198880
rect 142614 198840 142620 198852
rect 142672 198840 142678 198892
rect 167178 198840 167184 198892
rect 167236 198880 167242 198892
rect 208486 198880 208492 198892
rect 167236 198852 208492 198880
rect 167236 198840 167242 198852
rect 208486 198840 208492 198852
rect 208544 198840 208550 198892
rect 126238 198772 126244 198824
rect 126296 198812 126302 198824
rect 145558 198812 145564 198824
rect 126296 198784 145564 198812
rect 126296 198772 126302 198784
rect 145558 198772 145564 198784
rect 145616 198772 145622 198824
rect 153194 198772 153200 198824
rect 153252 198812 153258 198824
rect 208394 198812 208400 198824
rect 153252 198784 208400 198812
rect 153252 198772 153258 198784
rect 208394 198772 208400 198784
rect 208452 198772 208458 198824
rect 182818 198704 182824 198756
rect 182876 198744 182882 198756
rect 188246 198744 188252 198756
rect 182876 198716 188252 198744
rect 182876 198704 182882 198716
rect 188246 198704 188252 198716
rect 188304 198704 188310 198756
rect 155126 198568 155132 198620
rect 155184 198608 155190 198620
rect 174814 198608 174820 198620
rect 155184 198580 174820 198608
rect 155184 198568 155190 198580
rect 174814 198568 174820 198580
rect 174872 198568 174878 198620
rect 132310 198500 132316 198552
rect 132368 198540 132374 198552
rect 150802 198540 150808 198552
rect 132368 198512 150808 198540
rect 132368 198500 132374 198512
rect 150802 198500 150808 198512
rect 150860 198500 150866 198552
rect 122742 198228 122748 198280
rect 122800 198268 122806 198280
rect 149146 198268 149152 198280
rect 122800 198240 149152 198268
rect 122800 198228 122806 198240
rect 149146 198228 149152 198240
rect 149204 198228 149210 198280
rect 162854 198160 162860 198212
rect 162912 198200 162918 198212
rect 163314 198200 163320 198212
rect 162912 198172 163320 198200
rect 162912 198160 162918 198172
rect 163314 198160 163320 198172
rect 163372 198160 163378 198212
rect 167914 198200 167920 198212
rect 167656 198172 167920 198200
rect 167656 198144 167684 198172
rect 167914 198160 167920 198172
rect 167972 198160 167978 198212
rect 169662 198160 169668 198212
rect 169720 198200 169726 198212
rect 197998 198200 198004 198212
rect 169720 198172 198004 198200
rect 169720 198160 169726 198172
rect 197998 198160 198004 198172
rect 198056 198160 198062 198212
rect 167638 198092 167644 198144
rect 167696 198092 167702 198144
rect 171042 198092 171048 198144
rect 171100 198132 171106 198144
rect 199654 198132 199660 198144
rect 171100 198104 199660 198132
rect 171100 198092 171106 198104
rect 199654 198092 199660 198104
rect 199712 198092 199718 198144
rect 132034 198024 132040 198076
rect 132092 198064 132098 198076
rect 132494 198064 132500 198076
rect 132092 198036 132500 198064
rect 132092 198024 132098 198036
rect 132494 198024 132500 198036
rect 132552 198024 132558 198076
rect 136082 198024 136088 198076
rect 136140 198064 136146 198076
rect 136266 198064 136272 198076
rect 136140 198036 136272 198064
rect 136140 198024 136146 198036
rect 136266 198024 136272 198036
rect 136324 198024 136330 198076
rect 173434 198024 173440 198076
rect 173492 198064 173498 198076
rect 198826 198064 198832 198076
rect 173492 198036 198832 198064
rect 173492 198024 173498 198036
rect 198826 198024 198832 198036
rect 198884 198024 198890 198076
rect 131942 197956 131948 198008
rect 132000 197996 132006 198008
rect 132862 197996 132868 198008
rect 132000 197968 132868 197996
rect 132000 197956 132006 197968
rect 132862 197956 132868 197968
rect 132920 197956 132926 198008
rect 183186 197956 183192 198008
rect 183244 197996 183250 198008
rect 203150 197996 203156 198008
rect 183244 197968 203156 197996
rect 183244 197956 183250 197968
rect 203150 197956 203156 197968
rect 203208 197956 203214 198008
rect 129642 197888 129648 197940
rect 129700 197928 129706 197940
rect 150066 197928 150072 197940
rect 129700 197900 150072 197928
rect 129700 197888 129706 197900
rect 150066 197888 150072 197900
rect 150124 197888 150130 197940
rect 133966 197752 133972 197804
rect 134024 197792 134030 197804
rect 134426 197792 134432 197804
rect 134024 197764 134432 197792
rect 134024 197752 134030 197764
rect 134426 197752 134432 197764
rect 134484 197752 134490 197804
rect 163222 197752 163228 197804
rect 163280 197792 163286 197804
rect 163590 197792 163596 197804
rect 163280 197764 163596 197792
rect 163280 197752 163286 197764
rect 163590 197752 163596 197764
rect 163648 197752 163654 197804
rect 115658 197616 115664 197668
rect 115716 197656 115722 197668
rect 142338 197656 142344 197668
rect 115716 197628 142344 197656
rect 115716 197616 115722 197628
rect 142338 197616 142344 197628
rect 142396 197616 142402 197668
rect 155310 197548 155316 197600
rect 155368 197588 155374 197600
rect 173434 197588 173440 197600
rect 155368 197560 173440 197588
rect 155368 197548 155374 197560
rect 173434 197548 173440 197560
rect 173492 197548 173498 197600
rect 134518 197480 134524 197532
rect 134576 197520 134582 197532
rect 134886 197520 134892 197532
rect 134576 197492 134892 197520
rect 134576 197480 134582 197492
rect 134886 197480 134892 197492
rect 134944 197480 134950 197532
rect 163038 197276 163044 197328
rect 163096 197316 163102 197328
rect 197538 197316 197544 197328
rect 163096 197288 197544 197316
rect 163096 197276 163102 197288
rect 197538 197276 197544 197288
rect 197596 197276 197602 197328
rect 154482 197208 154488 197260
rect 154540 197248 154546 197260
rect 187050 197248 187056 197260
rect 154540 197220 187056 197248
rect 154540 197208 154546 197220
rect 187050 197208 187056 197220
rect 187108 197208 187114 197260
rect 156690 197140 156696 197192
rect 156748 197180 156754 197192
rect 190546 197180 190552 197192
rect 156748 197152 190552 197180
rect 156748 197140 156754 197152
rect 190546 197140 190552 197152
rect 190604 197140 190610 197192
rect 162210 197072 162216 197124
rect 162268 197112 162274 197124
rect 196066 197112 196072 197124
rect 162268 197084 196072 197112
rect 162268 197072 162274 197084
rect 196066 197072 196072 197084
rect 196124 197072 196130 197124
rect 118234 197004 118240 197056
rect 118292 197044 118298 197056
rect 145190 197044 145196 197056
rect 118292 197016 145196 197044
rect 118292 197004 118298 197016
rect 145190 197004 145196 197016
rect 145248 197004 145254 197056
rect 166258 197004 166264 197056
rect 166316 197044 166322 197056
rect 194686 197044 194692 197056
rect 166316 197016 194692 197044
rect 166316 197004 166322 197016
rect 194686 197004 194692 197016
rect 194744 197004 194750 197056
rect 157978 196936 157984 196988
rect 158036 196976 158042 196988
rect 191926 196976 191932 196988
rect 158036 196948 191932 196976
rect 158036 196936 158042 196948
rect 191926 196936 191932 196948
rect 191984 196936 191990 196988
rect 111426 196868 111432 196920
rect 111484 196908 111490 196920
rect 142890 196908 142896 196920
rect 111484 196880 142896 196908
rect 111484 196868 111490 196880
rect 142890 196868 142896 196880
rect 142948 196868 142954 196920
rect 163682 196868 163688 196920
rect 163740 196908 163746 196920
rect 197446 196908 197452 196920
rect 163740 196880 197452 196908
rect 163740 196868 163746 196880
rect 197446 196868 197452 196880
rect 197504 196868 197510 196920
rect 110138 196800 110144 196852
rect 110196 196840 110202 196852
rect 144638 196840 144644 196852
rect 110196 196812 144644 196840
rect 110196 196800 110202 196812
rect 144638 196800 144644 196812
rect 144696 196800 144702 196852
rect 160278 196800 160284 196852
rect 160336 196840 160342 196852
rect 194870 196840 194876 196852
rect 160336 196812 194876 196840
rect 160336 196800 160342 196812
rect 194870 196800 194876 196812
rect 194928 196800 194934 196852
rect 105906 196732 105912 196784
rect 105964 196772 105970 196784
rect 131022 196772 131028 196784
rect 105964 196744 131028 196772
rect 105964 196732 105970 196744
rect 131022 196732 131028 196744
rect 131080 196732 131086 196784
rect 159450 196732 159456 196784
rect 159508 196772 159514 196784
rect 193398 196772 193404 196784
rect 159508 196744 193404 196772
rect 159508 196732 159514 196744
rect 193398 196732 193404 196744
rect 193456 196732 193462 196784
rect 115474 196664 115480 196716
rect 115532 196704 115538 196716
rect 149514 196704 149520 196716
rect 115532 196676 149520 196704
rect 115532 196664 115538 196676
rect 149514 196664 149520 196676
rect 149572 196664 149578 196716
rect 161934 196664 161940 196716
rect 161992 196704 161998 196716
rect 196158 196704 196164 196716
rect 161992 196676 196164 196704
rect 161992 196664 161998 196676
rect 196158 196664 196164 196676
rect 196216 196664 196222 196716
rect 112622 196596 112628 196648
rect 112680 196636 112686 196648
rect 147582 196636 147588 196648
rect 112680 196608 147588 196636
rect 112680 196596 112686 196608
rect 147582 196596 147588 196608
rect 147640 196596 147646 196648
rect 157702 196596 157708 196648
rect 157760 196636 157766 196648
rect 192110 196636 192116 196648
rect 157760 196608 192116 196636
rect 157760 196596 157766 196608
rect 192110 196596 192116 196608
rect 192168 196596 192174 196648
rect 158898 196528 158904 196580
rect 158956 196568 158962 196580
rect 193490 196568 193496 196580
rect 158956 196540 193496 196568
rect 158956 196528 158962 196540
rect 193490 196528 193496 196540
rect 193548 196528 193554 196580
rect 154758 196460 154764 196512
rect 154816 196500 154822 196512
rect 189718 196500 189724 196512
rect 154816 196472 189724 196500
rect 154816 196460 154822 196472
rect 189718 196460 189724 196472
rect 189776 196460 189782 196512
rect 169938 196052 169944 196104
rect 169996 196092 170002 196104
rect 183094 196092 183100 196104
rect 169996 196064 183100 196092
rect 169996 196052 170002 196064
rect 183094 196052 183100 196064
rect 183152 196052 183158 196104
rect 166994 195916 167000 195968
rect 167052 195956 167058 195968
rect 182910 195956 182916 195968
rect 167052 195928 182916 195956
rect 167052 195916 167058 195928
rect 182910 195916 182916 195928
rect 182968 195916 182974 195968
rect 119890 195848 119896 195900
rect 119948 195888 119954 195900
rect 150342 195888 150348 195900
rect 119948 195860 150348 195888
rect 119948 195848 119954 195860
rect 150342 195848 150348 195860
rect 150400 195848 150406 195900
rect 156230 195848 156236 195900
rect 156288 195888 156294 195900
rect 190730 195888 190736 195900
rect 156288 195860 190736 195888
rect 156288 195848 156294 195860
rect 190730 195848 190736 195860
rect 190788 195848 190794 195900
rect 159634 195780 159640 195832
rect 159692 195820 159698 195832
rect 180150 195820 180156 195832
rect 159692 195792 180156 195820
rect 159692 195780 159698 195792
rect 180150 195780 180156 195792
rect 180208 195780 180214 195832
rect 111242 195712 111248 195764
rect 111300 195752 111306 195764
rect 120350 195752 120356 195764
rect 111300 195724 120356 195752
rect 111300 195712 111306 195724
rect 120350 195712 120356 195724
rect 120408 195712 120414 195764
rect 159266 195712 159272 195764
rect 159324 195752 159330 195764
rect 194134 195752 194140 195764
rect 159324 195724 194140 195752
rect 159324 195712 159330 195724
rect 194134 195712 194140 195724
rect 194192 195712 194198 195764
rect 111150 195644 111156 195696
rect 111208 195684 111214 195696
rect 143166 195684 143172 195696
rect 111208 195656 143172 195684
rect 111208 195644 111214 195656
rect 143166 195644 143172 195656
rect 143224 195644 143230 195696
rect 180058 195684 180064 195696
rect 178328 195656 180064 195684
rect 110230 195576 110236 195628
rect 110288 195616 110294 195628
rect 142246 195616 142252 195628
rect 110288 195588 142252 195616
rect 110288 195576 110294 195588
rect 142246 195576 142252 195588
rect 142304 195576 142310 195628
rect 157334 195576 157340 195628
rect 157392 195616 157398 195628
rect 178328 195616 178356 195656
rect 180058 195644 180064 195656
rect 180116 195644 180122 195696
rect 157392 195588 178356 195616
rect 157392 195576 157398 195588
rect 105998 195508 106004 195560
rect 106056 195548 106062 195560
rect 138658 195548 138664 195560
rect 106056 195520 138664 195548
rect 106056 195508 106062 195520
rect 138658 195508 138664 195520
rect 138716 195508 138722 195560
rect 161566 195508 161572 195560
rect 161624 195548 161630 195560
rect 194594 195548 194600 195560
rect 161624 195520 194600 195548
rect 161624 195508 161630 195520
rect 194594 195508 194600 195520
rect 194652 195508 194658 195560
rect 105722 195440 105728 195492
rect 105780 195480 105786 195492
rect 139118 195480 139124 195492
rect 105780 195452 139124 195480
rect 105780 195440 105786 195452
rect 139118 195440 139124 195452
rect 139176 195440 139182 195492
rect 160094 195440 160100 195492
rect 160152 195480 160158 195492
rect 193306 195480 193312 195492
rect 160152 195452 193312 195480
rect 160152 195440 160158 195452
rect 193306 195440 193312 195452
rect 193364 195440 193370 195492
rect 109770 195372 109776 195424
rect 109828 195412 109834 195424
rect 142522 195412 142528 195424
rect 109828 195384 142528 195412
rect 109828 195372 109834 195384
rect 142522 195372 142528 195384
rect 142580 195372 142586 195424
rect 160370 195372 160376 195424
rect 160428 195412 160434 195424
rect 190638 195412 190644 195424
rect 160428 195384 190644 195412
rect 160428 195372 160434 195384
rect 190638 195372 190644 195384
rect 190696 195372 190702 195424
rect 106826 195304 106832 195356
rect 106884 195344 106890 195356
rect 137830 195344 137836 195356
rect 106884 195316 137836 195344
rect 106884 195304 106890 195316
rect 137830 195304 137836 195316
rect 137888 195304 137894 195356
rect 158346 195304 158352 195356
rect 158404 195344 158410 195356
rect 191834 195344 191840 195356
rect 158404 195316 191840 195344
rect 158404 195304 158410 195316
rect 191834 195304 191840 195316
rect 191892 195304 191898 195356
rect 105538 195236 105544 195288
rect 105596 195276 105602 195288
rect 139578 195276 139584 195288
rect 105596 195248 139584 195276
rect 105596 195236 105602 195248
rect 139578 195236 139584 195248
rect 139636 195236 139642 195288
rect 158070 195236 158076 195288
rect 158128 195276 158134 195288
rect 192018 195276 192024 195288
rect 158128 195248 192024 195276
rect 158128 195236 158134 195248
rect 192018 195236 192024 195248
rect 192076 195236 192082 195288
rect 176626 195044 182174 195072
rect 173434 194964 173440 195016
rect 173492 195004 173498 195016
rect 176626 195004 176654 195044
rect 173492 194976 176654 195004
rect 182146 195004 182174 195044
rect 189166 195004 189172 195016
rect 182146 194976 189172 195004
rect 173492 194964 173498 194976
rect 189166 194964 189172 194976
rect 189224 194964 189230 195016
rect 153470 194896 153476 194948
rect 153528 194936 153534 194948
rect 188246 194936 188252 194948
rect 153528 194908 188252 194936
rect 153528 194896 153534 194908
rect 188246 194896 188252 194908
rect 188304 194896 188310 194948
rect 174814 194828 174820 194880
rect 174872 194868 174878 194880
rect 189074 194868 189080 194880
rect 174872 194840 189080 194868
rect 174872 194828 174878 194840
rect 189074 194828 189080 194840
rect 189132 194828 189138 194880
rect 128262 194692 128268 194744
rect 128320 194732 128326 194744
rect 138750 194732 138756 194744
rect 128320 194704 138756 194732
rect 128320 194692 128326 194704
rect 138750 194692 138756 194704
rect 138808 194692 138814 194744
rect 127894 194488 127900 194540
rect 127952 194528 127958 194540
rect 153286 194528 153292 194540
rect 127952 194500 153292 194528
rect 127952 194488 127958 194500
rect 153286 194488 153292 194500
rect 153344 194488 153350 194540
rect 100662 194352 100668 194404
rect 100720 194392 100726 194404
rect 104434 194392 104440 194404
rect 100720 194364 104440 194392
rect 100720 194352 100726 194364
rect 104434 194352 104440 194364
rect 104492 194352 104498 194404
rect 115842 194284 115848 194336
rect 115900 194324 115906 194336
rect 148226 194324 148232 194336
rect 115900 194296 148232 194324
rect 115900 194284 115906 194296
rect 148226 194284 148232 194296
rect 148284 194284 148290 194336
rect 112806 194216 112812 194268
rect 112864 194256 112870 194268
rect 145834 194256 145840 194268
rect 112864 194228 145840 194256
rect 112864 194216 112870 194228
rect 145834 194216 145840 194228
rect 145892 194216 145898 194268
rect 114094 194148 114100 194200
rect 114152 194188 114158 194200
rect 146938 194188 146944 194200
rect 114152 194160 146944 194188
rect 114152 194148 114158 194160
rect 146938 194148 146944 194160
rect 146996 194148 147002 194200
rect 174170 194148 174176 194200
rect 174228 194188 174234 194200
rect 200758 194188 200764 194200
rect 174228 194160 200764 194188
rect 174228 194148 174234 194160
rect 200758 194148 200764 194160
rect 200816 194148 200822 194200
rect 112714 194080 112720 194132
rect 112772 194120 112778 194132
rect 145006 194120 145012 194132
rect 112772 194092 145012 194120
rect 112772 194080 112778 194092
rect 145006 194080 145012 194092
rect 145064 194080 145070 194132
rect 114002 194012 114008 194064
rect 114060 194052 114066 194064
rect 146386 194052 146392 194064
rect 114060 194024 146392 194052
rect 114060 194012 114066 194024
rect 146386 194012 146392 194024
rect 146444 194012 146450 194064
rect 174354 194012 174360 194064
rect 174412 194052 174418 194064
rect 174722 194052 174728 194064
rect 174412 194024 174728 194052
rect 174412 194012 174418 194024
rect 174722 194012 174728 194024
rect 174780 194012 174786 194064
rect 177114 194012 177120 194064
rect 177172 194052 177178 194064
rect 207014 194052 207020 194064
rect 177172 194024 207020 194052
rect 177172 194012 177178 194024
rect 207014 194012 207020 194024
rect 207072 194012 207078 194064
rect 102042 193944 102048 193996
rect 102100 193984 102106 193996
rect 135254 193984 135260 193996
rect 102100 193956 135260 193984
rect 102100 193944 102106 193956
rect 135254 193944 135260 193956
rect 135312 193944 135318 193996
rect 169938 193944 169944 193996
rect 169996 193984 170002 193996
rect 202874 193984 202880 193996
rect 169996 193956 202880 193984
rect 169996 193944 170002 193956
rect 202874 193944 202880 193956
rect 202932 193944 202938 193996
rect 118510 193876 118516 193928
rect 118568 193916 118574 193928
rect 151538 193916 151544 193928
rect 118568 193888 151544 193916
rect 118568 193876 118574 193888
rect 151538 193876 151544 193888
rect 151596 193876 151602 193928
rect 167822 193876 167828 193928
rect 167880 193916 167886 193928
rect 202506 193916 202512 193928
rect 167880 193888 202512 193916
rect 167880 193876 167886 193888
rect 202506 193876 202512 193888
rect 202564 193876 202570 193928
rect 106090 193808 106096 193860
rect 106148 193848 106154 193860
rect 140222 193848 140228 193860
rect 106148 193820 140228 193848
rect 106148 193808 106154 193820
rect 140222 193808 140228 193820
rect 140280 193808 140286 193860
rect 166718 193808 166724 193860
rect 166776 193848 166782 193860
rect 200114 193848 200120 193860
rect 166776 193820 200120 193848
rect 166776 193808 166782 193820
rect 200114 193808 200120 193820
rect 200172 193808 200178 193860
rect 108942 193672 108948 193724
rect 109000 193712 109006 193724
rect 128262 193712 128268 193724
rect 109000 193684 128268 193712
rect 109000 193672 109006 193684
rect 128262 193672 128268 193684
rect 128320 193672 128326 193724
rect 131942 193672 131948 193724
rect 132000 193712 132006 193724
rect 154666 193712 154672 193724
rect 132000 193684 154672 193712
rect 132000 193672 132006 193684
rect 154666 193672 154672 193684
rect 154724 193672 154730 193724
rect 130470 193604 130476 193656
rect 130528 193644 130534 193656
rect 150618 193644 150624 193656
rect 130528 193616 150624 193644
rect 130528 193604 130534 193616
rect 150618 193604 150624 193616
rect 150676 193604 150682 193656
rect 162578 193264 162584 193316
rect 162636 193304 162642 193316
rect 183462 193304 183468 193316
rect 162636 193276 183468 193304
rect 162636 193264 162642 193276
rect 183462 193264 183468 193276
rect 183520 193264 183526 193316
rect 164694 193196 164700 193248
rect 164752 193236 164758 193248
rect 184106 193236 184112 193248
rect 164752 193208 184112 193236
rect 164752 193196 164758 193208
rect 184106 193196 184112 193208
rect 184164 193196 184170 193248
rect 156138 193128 156144 193180
rect 156196 193168 156202 193180
rect 181530 193168 181536 193180
rect 156196 193140 181536 193168
rect 156196 193128 156202 193140
rect 181530 193128 181536 193140
rect 181588 193128 181594 193180
rect 188430 193128 188436 193180
rect 188488 193168 188494 193180
rect 580166 193168 580172 193180
rect 188488 193140 580172 193168
rect 188488 193128 188494 193140
rect 580166 193128 580172 193140
rect 580224 193128 580230 193180
rect 171962 193060 171968 193112
rect 172020 193100 172026 193112
rect 205634 193100 205640 193112
rect 172020 193072 205640 193100
rect 172020 193060 172026 193072
rect 205634 193060 205640 193072
rect 205692 193060 205698 193112
rect 164970 192992 164976 193044
rect 165028 193032 165034 193044
rect 194778 193032 194784 193044
rect 165028 193004 194784 193032
rect 165028 192992 165034 193004
rect 194778 192992 194784 193004
rect 194836 192992 194842 193044
rect 110966 192924 110972 192976
rect 111024 192964 111030 192976
rect 140682 192964 140688 192976
rect 111024 192936 140688 192964
rect 111024 192924 111030 192936
rect 140682 192924 140688 192936
rect 140740 192924 140746 192976
rect 173986 192924 173992 192976
rect 174044 192964 174050 192976
rect 204346 192964 204352 192976
rect 174044 192936 204352 192964
rect 174044 192924 174050 192936
rect 204346 192924 204352 192936
rect 204404 192924 204410 192976
rect 108666 192856 108672 192908
rect 108724 192896 108730 192908
rect 138658 192896 138664 192908
rect 108724 192868 138664 192896
rect 108724 192856 108730 192868
rect 138658 192856 138664 192868
rect 138716 192856 138722 192908
rect 176838 192856 176844 192908
rect 176896 192896 176902 192908
rect 207106 192896 207112 192908
rect 176896 192868 207112 192896
rect 176896 192856 176902 192868
rect 207106 192856 207112 192868
rect 207164 192856 207170 192908
rect 168742 192788 168748 192840
rect 168800 192828 168806 192840
rect 180334 192828 180340 192840
rect 168800 192800 180340 192828
rect 168800 192788 168806 192800
rect 180334 192788 180340 192800
rect 180392 192788 180398 192840
rect 183094 192788 183100 192840
rect 183152 192828 183158 192840
rect 203058 192828 203064 192840
rect 183152 192800 203064 192828
rect 183152 192788 183158 192800
rect 203058 192788 203064 192800
rect 203116 192788 203122 192840
rect 167454 192720 167460 192772
rect 167512 192760 167518 192772
rect 201770 192760 201776 192772
rect 167512 192732 201776 192760
rect 167512 192720 167518 192732
rect 201770 192720 201776 192732
rect 201828 192720 201834 192772
rect 103330 192652 103336 192704
rect 103388 192692 103394 192704
rect 135806 192692 135812 192704
rect 103388 192664 135812 192692
rect 103388 192652 103394 192664
rect 135806 192652 135812 192664
rect 135864 192652 135870 192704
rect 169202 192652 169208 192704
rect 169260 192692 169266 192704
rect 202966 192692 202972 192704
rect 169260 192664 202972 192692
rect 169260 192652 169266 192664
rect 202966 192652 202972 192664
rect 203024 192652 203030 192704
rect 104066 192584 104072 192636
rect 104124 192624 104130 192636
rect 137646 192624 137652 192636
rect 104124 192596 137652 192624
rect 104124 192584 104130 192596
rect 137646 192584 137652 192596
rect 137704 192584 137710 192636
rect 103054 192516 103060 192568
rect 103112 192556 103118 192568
rect 138014 192556 138020 192568
rect 103112 192528 138020 192556
rect 103112 192516 103118 192528
rect 138014 192516 138020 192528
rect 138072 192516 138078 192568
rect 164142 192516 164148 192568
rect 164200 192556 164206 192568
rect 197354 192556 197360 192568
rect 164200 192528 197360 192556
rect 164200 192516 164206 192528
rect 197354 192516 197360 192528
rect 197412 192516 197418 192568
rect 103146 192448 103152 192500
rect 103204 192488 103210 192500
rect 137462 192488 137468 192500
rect 103204 192460 137468 192488
rect 103204 192448 103210 192460
rect 137462 192448 137468 192460
rect 137520 192448 137526 192500
rect 153378 192448 153384 192500
rect 153436 192488 153442 192500
rect 162210 192488 162216 192500
rect 153436 192460 162216 192488
rect 153436 192448 153442 192460
rect 162210 192448 162216 192460
rect 162268 192448 162274 192500
rect 174078 192448 174084 192500
rect 174136 192488 174142 192500
rect 174906 192488 174912 192500
rect 174136 192460 174912 192488
rect 174136 192448 174142 192460
rect 174906 192448 174912 192460
rect 174964 192448 174970 192500
rect 183462 192448 183468 192500
rect 183520 192488 183526 192500
rect 195974 192488 195980 192500
rect 183520 192460 195980 192488
rect 183520 192448 183526 192460
rect 195974 192448 195980 192460
rect 196032 192448 196038 192500
rect 116854 192380 116860 192432
rect 116912 192420 116918 192432
rect 144546 192420 144552 192432
rect 116912 192392 144552 192420
rect 116912 192380 116918 192392
rect 144546 192380 144552 192392
rect 144604 192380 144610 192432
rect 173986 192380 173992 192432
rect 174044 192420 174050 192432
rect 174998 192420 175004 192432
rect 174044 192392 175004 192420
rect 174044 192380 174050 192392
rect 174998 192380 175004 192392
rect 175056 192380 175062 192432
rect 184106 192380 184112 192432
rect 184164 192420 184170 192432
rect 199102 192420 199108 192432
rect 184164 192392 199108 192420
rect 184164 192380 184170 192392
rect 199102 192380 199108 192392
rect 199160 192380 199166 192432
rect 110322 192312 110328 192364
rect 110380 192352 110386 192364
rect 138014 192352 138020 192364
rect 110380 192324 138020 192352
rect 110380 192312 110386 192324
rect 138014 192312 138020 192324
rect 138072 192312 138078 192364
rect 200206 192352 200212 192364
rect 175522 192324 200212 192352
rect 125042 192244 125048 192296
rect 125100 192284 125106 192296
rect 141694 192284 141700 192296
rect 125100 192256 141700 192284
rect 125100 192244 125106 192256
rect 141694 192244 141700 192256
rect 141752 192244 141758 192296
rect 166074 192244 166080 192296
rect 166132 192284 166138 192296
rect 175522 192284 175550 192324
rect 200206 192312 200212 192324
rect 200264 192312 200270 192364
rect 185578 192284 185584 192296
rect 166132 192256 175550 192284
rect 184906 192256 185584 192284
rect 166132 192244 166138 192256
rect 168282 192176 168288 192228
rect 168340 192216 168346 192228
rect 184906 192216 184934 192256
rect 185578 192244 185584 192256
rect 185636 192244 185642 192296
rect 168340 192188 184934 192216
rect 168340 192176 168346 192188
rect 166442 192040 166448 192092
rect 166500 192080 166506 192092
rect 183002 192080 183008 192092
rect 166500 192052 183008 192080
rect 166500 192040 166506 192052
rect 183002 192040 183008 192052
rect 183060 192040 183066 192092
rect 161382 191632 161388 191684
rect 161440 191672 161446 191684
rect 183094 191672 183100 191684
rect 161440 191644 183100 191672
rect 161440 191632 161446 191644
rect 183094 191632 183100 191644
rect 183152 191632 183158 191684
rect 122098 191360 122104 191412
rect 122156 191400 122162 191412
rect 139854 191400 139860 191412
rect 122156 191372 139860 191400
rect 122156 191360 122162 191372
rect 139854 191360 139860 191372
rect 139912 191360 139918 191412
rect 111334 191292 111340 191344
rect 111392 191332 111398 191344
rect 143074 191332 143080 191344
rect 111392 191304 143080 191332
rect 111392 191292 111398 191304
rect 143074 191292 143080 191304
rect 143132 191292 143138 191344
rect 101950 191224 101956 191276
rect 102008 191264 102014 191276
rect 134334 191264 134340 191276
rect 102008 191236 134340 191264
rect 102008 191224 102014 191236
rect 134334 191224 134340 191236
rect 134392 191224 134398 191276
rect 141326 191264 141332 191276
rect 135916 191236 141332 191264
rect 109862 191156 109868 191208
rect 109920 191196 109926 191208
rect 135916 191196 135944 191236
rect 141326 191224 141332 191236
rect 141384 191224 141390 191276
rect 109920 191168 135944 191196
rect 109920 191156 109926 191168
rect 109678 191088 109684 191140
rect 109736 191128 109742 191140
rect 144178 191128 144184 191140
rect 109736 191100 144184 191128
rect 109736 191088 109742 191100
rect 144178 191088 144184 191100
rect 144236 191088 144242 191140
rect 131758 190952 131764 191004
rect 131816 190992 131822 191004
rect 138934 190992 138940 191004
rect 131816 190964 138940 190992
rect 131816 190952 131822 190964
rect 138934 190952 138940 190964
rect 138992 190952 138998 191004
rect 123570 190884 123576 190936
rect 123628 190924 123634 190936
rect 145282 190924 145288 190936
rect 123628 190896 145288 190924
rect 123628 190884 123634 190896
rect 145282 190884 145288 190896
rect 145340 190884 145346 190936
rect 127710 190680 127716 190732
rect 127768 190720 127774 190732
rect 143994 190720 144000 190732
rect 127768 190692 144000 190720
rect 127768 190680 127774 190692
rect 143994 190680 144000 190692
rect 144052 190680 144058 190732
rect 168098 190680 168104 190732
rect 168156 190720 168162 190732
rect 178862 190720 178868 190732
rect 168156 190692 178868 190720
rect 168156 190680 168162 190692
rect 178862 190680 178868 190692
rect 178920 190680 178926 190732
rect 110046 190408 110052 190460
rect 110104 190448 110110 190460
rect 141418 190448 141424 190460
rect 110104 190420 141424 190448
rect 110104 190408 110110 190420
rect 141418 190408 141424 190420
rect 141476 190408 141482 190460
rect 110874 190340 110880 190392
rect 110932 190380 110938 190392
rect 141878 190380 141884 190392
rect 110932 190352 141884 190380
rect 110932 190340 110938 190352
rect 141878 190340 141884 190352
rect 141936 190340 141942 190392
rect 107562 190272 107568 190324
rect 107620 190312 107626 190324
rect 139946 190312 139952 190324
rect 107620 190284 139952 190312
rect 107620 190272 107626 190284
rect 139946 190272 139952 190284
rect 140004 190272 140010 190324
rect 106182 190204 106188 190256
rect 106240 190244 106246 190256
rect 138290 190244 138296 190256
rect 106240 190216 138296 190244
rect 106240 190204 106246 190216
rect 138290 190204 138296 190216
rect 138348 190204 138354 190256
rect 100570 190136 100576 190188
rect 100628 190176 100634 190188
rect 133782 190176 133788 190188
rect 100628 190148 133788 190176
rect 100628 190136 100634 190148
rect 133782 190136 133788 190148
rect 133840 190136 133846 190188
rect 101858 190068 101864 190120
rect 101916 190108 101922 190120
rect 134794 190108 134800 190120
rect 101916 190080 134800 190108
rect 101916 190068 101922 190080
rect 134794 190068 134800 190080
rect 134852 190068 134858 190120
rect 111518 190000 111524 190052
rect 111576 190040 111582 190052
rect 139394 190040 139400 190052
rect 111576 190012 139400 190040
rect 111576 190000 111582 190012
rect 139394 190000 139400 190012
rect 139452 190000 139458 190052
rect 101582 189932 101588 189984
rect 101640 189972 101646 189984
rect 104802 189972 104808 189984
rect 101640 189944 104808 189972
rect 101640 189932 101646 189944
rect 104802 189932 104808 189944
rect 104860 189932 104866 189984
rect 101766 189864 101772 189916
rect 101824 189904 101830 189916
rect 133966 189904 133972 189916
rect 101824 189876 133972 189904
rect 101824 189864 101830 189876
rect 133966 189864 133972 189876
rect 134024 189864 134030 189916
rect 101674 189796 101680 189848
rect 101732 189836 101738 189848
rect 133598 189836 133604 189848
rect 101732 189808 133604 189836
rect 101732 189796 101738 189808
rect 133598 189796 133604 189808
rect 133656 189796 133662 189848
rect 104802 189728 104808 189780
rect 104860 189768 104866 189780
rect 138842 189768 138848 189780
rect 104860 189740 138848 189768
rect 104860 189728 104866 189740
rect 138842 189728 138848 189740
rect 138900 189728 138906 189780
rect 107378 189660 107384 189712
rect 107436 189700 107442 189712
rect 138566 189700 138572 189712
rect 107436 189672 138572 189700
rect 107436 189660 107442 189672
rect 138566 189660 138572 189672
rect 138624 189660 138630 189712
rect 108850 189592 108856 189644
rect 108908 189632 108914 189644
rect 138934 189632 138940 189644
rect 108908 189604 138940 189632
rect 108908 189592 108914 189604
rect 138934 189592 138940 189604
rect 138992 189592 138998 189644
rect 112530 189524 112536 189576
rect 112588 189564 112594 189576
rect 120166 189564 120172 189576
rect 112588 189536 120172 189564
rect 112588 189524 112594 189536
rect 120166 189524 120172 189536
rect 120224 189524 120230 189576
rect 165614 189048 165620 189100
rect 165672 189088 165678 189100
rect 178770 189088 178776 189100
rect 165672 189060 178776 189088
rect 165672 189048 165678 189060
rect 178770 189048 178776 189060
rect 178828 189048 178834 189100
rect 3418 188980 3424 189032
rect 3476 189020 3482 189032
rect 120534 189020 120540 189032
rect 3476 188992 120540 189020
rect 3476 188980 3482 188992
rect 120534 188980 120540 188992
rect 120592 188980 120598 189032
rect 131850 188912 131856 188964
rect 131908 188952 131914 188964
rect 140774 188952 140780 188964
rect 131908 188924 140780 188952
rect 131908 188912 131914 188924
rect 140774 188912 140780 188924
rect 140832 188912 140838 188964
rect 126330 188844 126336 188896
rect 126388 188884 126394 188896
rect 146018 188884 146024 188896
rect 126388 188856 146024 188884
rect 126388 188844 126394 188856
rect 146018 188844 146024 188856
rect 146076 188844 146082 188896
rect 127618 187960 127624 188012
rect 127676 188000 127682 188012
rect 143718 188000 143724 188012
rect 127676 187972 143724 188000
rect 127676 187960 127682 187972
rect 143718 187960 143724 187972
rect 143776 187960 143782 188012
rect 130378 187416 130384 187468
rect 130436 187456 130442 187468
rect 142798 187456 142804 187468
rect 130436 187428 142804 187456
rect 130436 187416 130442 187428
rect 142798 187416 142804 187428
rect 142856 187416 142862 187468
rect 163958 187280 163964 187332
rect 164016 187320 164022 187332
rect 181438 187320 181444 187332
rect 164016 187292 181444 187320
rect 164016 187280 164022 187292
rect 181438 187280 181444 187292
rect 181496 187280 181502 187332
rect 102778 186940 102784 186992
rect 102836 186980 102842 186992
rect 135530 186980 135536 186992
rect 102836 186952 135536 186980
rect 102836 186940 102842 186952
rect 135530 186940 135536 186952
rect 135588 186940 135594 186992
rect 163406 186940 163412 186992
rect 163464 186980 163470 186992
rect 178678 186980 178684 186992
rect 163464 186952 178684 186980
rect 163464 186940 163470 186952
rect 178678 186940 178684 186952
rect 178736 186940 178742 186992
rect 124122 186872 124128 186924
rect 124180 186912 124186 186924
rect 148318 186912 148324 186924
rect 124180 186884 148324 186912
rect 124180 186872 124186 186884
rect 148318 186872 148324 186884
rect 148376 186872 148382 186924
rect 171318 186668 171324 186720
rect 171376 186708 171382 186720
rect 195238 186708 195244 186720
rect 171376 186680 195244 186708
rect 171376 186668 171382 186680
rect 195238 186668 195244 186680
rect 195296 186668 195302 186720
rect 160002 186600 160008 186652
rect 160060 186640 160066 186652
rect 171226 186640 171232 186652
rect 160060 186612 171232 186640
rect 160060 186600 160066 186612
rect 171226 186600 171232 186612
rect 171284 186600 171290 186652
rect 171594 186600 171600 186652
rect 171652 186640 171658 186652
rect 199010 186640 199016 186652
rect 171652 186612 199016 186640
rect 171652 186600 171658 186612
rect 199010 186600 199016 186612
rect 199068 186600 199074 186652
rect 172882 186464 172888 186516
rect 172940 186504 172946 186516
rect 199194 186504 199200 186516
rect 172940 186476 199200 186504
rect 172940 186464 172946 186476
rect 199194 186464 199200 186476
rect 199252 186464 199258 186516
rect 154850 186396 154856 186448
rect 154908 186436 154914 186448
rect 155494 186436 155500 186448
rect 154908 186408 155500 186436
rect 154908 186396 154914 186408
rect 155494 186396 155500 186408
rect 155552 186396 155558 186448
rect 174262 186396 174268 186448
rect 174320 186436 174326 186448
rect 198734 186436 198740 186448
rect 174320 186408 198740 186436
rect 174320 186396 174326 186408
rect 198734 186396 198740 186408
rect 198792 186396 198798 186448
rect 172790 186328 172796 186380
rect 172848 186368 172854 186380
rect 205726 186368 205732 186380
rect 172848 186340 205732 186368
rect 172848 186328 172854 186340
rect 205726 186328 205732 186340
rect 205784 186328 205790 186380
rect 136542 186260 136548 186312
rect 136600 186300 136606 186312
rect 137186 186300 137192 186312
rect 136600 186272 137192 186300
rect 136600 186260 136606 186272
rect 137186 186260 137192 186272
rect 137244 186260 137250 186312
rect 158898 186260 158904 186312
rect 158956 186300 158962 186312
rect 159542 186300 159548 186312
rect 158956 186272 159548 186300
rect 158956 186260 158962 186272
rect 159542 186260 159548 186272
rect 159600 186260 159606 186312
rect 161566 186260 161572 186312
rect 161624 186300 161630 186312
rect 162026 186300 162032 186312
rect 161624 186272 162032 186300
rect 161624 186260 161630 186272
rect 162026 186260 162032 186272
rect 162084 186260 162090 186312
rect 169846 186260 169852 186312
rect 169904 186300 169910 186312
rect 170858 186300 170864 186312
rect 169904 186272 170864 186300
rect 169904 186260 169910 186272
rect 170858 186260 170864 186272
rect 170916 186260 170922 186312
rect 171042 186260 171048 186312
rect 171100 186300 171106 186312
rect 171502 186300 171508 186312
rect 171100 186272 171508 186300
rect 171100 186260 171106 186272
rect 171502 186260 171508 186272
rect 171560 186260 171566 186312
rect 176838 186260 176844 186312
rect 176896 186300 176902 186312
rect 177206 186300 177212 186312
rect 176896 186272 177212 186300
rect 176896 186260 176902 186272
rect 177206 186260 177212 186272
rect 177264 186260 177270 186312
rect 107286 186192 107292 186244
rect 107344 186232 107350 186244
rect 136450 186232 136456 186244
rect 107344 186204 136456 186232
rect 107344 186192 107350 186204
rect 136450 186192 136456 186204
rect 136508 186192 136514 186244
rect 148962 186192 148968 186244
rect 149020 186232 149026 186244
rect 157794 186232 157800 186244
rect 149020 186204 157800 186232
rect 149020 186192 149026 186204
rect 157794 186192 157800 186204
rect 157852 186192 157858 186244
rect 176746 186192 176752 186244
rect 176804 186232 176810 186244
rect 177482 186232 177488 186244
rect 176804 186204 177488 186232
rect 176804 186192 176810 186204
rect 177482 186192 177488 186204
rect 177540 186192 177546 186244
rect 148318 186124 148324 186176
rect 148376 186164 148382 186176
rect 148778 186164 148784 186176
rect 148376 186136 148784 186164
rect 148376 186124 148382 186136
rect 148778 186124 148784 186136
rect 148836 186124 148842 186176
rect 176654 186124 176660 186176
rect 176712 186164 176718 186176
rect 177758 186164 177764 186176
rect 176712 186136 177764 186164
rect 176712 186124 176718 186136
rect 177758 186124 177764 186136
rect 177816 186124 177822 186176
rect 154482 185784 154488 185836
rect 154540 185824 154546 185836
rect 158806 185824 158812 185836
rect 154540 185796 158812 185824
rect 154540 185784 154546 185796
rect 158806 185784 158812 185796
rect 158864 185784 158870 185836
rect 103422 185716 103428 185768
rect 103480 185756 103486 185768
rect 134242 185756 134248 185768
rect 103480 185728 134248 185756
rect 103480 185716 103486 185728
rect 134242 185716 134248 185728
rect 134300 185716 134306 185768
rect 105814 185648 105820 185700
rect 105872 185688 105878 185700
rect 137278 185688 137284 185700
rect 105872 185660 137284 185688
rect 105872 185648 105878 185660
rect 137278 185648 137284 185660
rect 137336 185648 137342 185700
rect 153930 185648 153936 185700
rect 153988 185688 153994 185700
rect 154390 185688 154396 185700
rect 153988 185660 154396 185688
rect 153988 185648 153994 185660
rect 154390 185648 154396 185660
rect 154448 185648 154454 185700
rect 155494 185648 155500 185700
rect 155552 185688 155558 185700
rect 155770 185688 155776 185700
rect 155552 185660 155776 185688
rect 155552 185648 155558 185660
rect 155770 185648 155776 185660
rect 155828 185648 155834 185700
rect 158806 185648 158812 185700
rect 158864 185688 158870 185700
rect 159818 185688 159824 185700
rect 158864 185660 159824 185688
rect 158864 185648 158870 185660
rect 159818 185648 159824 185660
rect 159876 185648 159882 185700
rect 164142 185648 164148 185700
rect 164200 185688 164206 185700
rect 167270 185688 167276 185700
rect 164200 185660 167276 185688
rect 164200 185648 164206 185660
rect 167270 185648 167276 185660
rect 167328 185648 167334 185700
rect 174630 185648 174636 185700
rect 174688 185688 174694 185700
rect 201678 185688 201684 185700
rect 174688 185660 201684 185688
rect 174688 185648 174694 185660
rect 201678 185648 201684 185660
rect 201736 185648 201742 185700
rect 104618 185580 104624 185632
rect 104676 185620 104682 185632
rect 134518 185620 134524 185632
rect 104676 185592 134524 185620
rect 104676 185580 104682 185592
rect 134518 185580 134524 185592
rect 134576 185580 134582 185632
rect 141142 185580 141148 185632
rect 141200 185620 141206 185632
rect 141510 185620 141516 185632
rect 141200 185592 141516 185620
rect 141200 185580 141206 185592
rect 141510 185580 141516 185592
rect 141568 185580 141574 185632
rect 149606 185580 149612 185632
rect 149664 185620 149670 185632
rect 150158 185620 150164 185632
rect 149664 185592 150164 185620
rect 149664 185580 149670 185592
rect 150158 185580 150164 185592
rect 150216 185580 150222 185632
rect 151906 185580 151912 185632
rect 151964 185620 151970 185632
rect 152458 185620 152464 185632
rect 151964 185592 152464 185620
rect 151964 185580 151970 185592
rect 152458 185580 152464 185592
rect 152516 185580 152522 185632
rect 153378 185580 153384 185632
rect 153436 185620 153442 185632
rect 154114 185620 154120 185632
rect 153436 185592 154120 185620
rect 153436 185580 153442 185592
rect 154114 185580 154120 185592
rect 154172 185580 154178 185632
rect 154758 185580 154764 185632
rect 154816 185620 154822 185632
rect 155678 185620 155684 185632
rect 154816 185592 155684 185620
rect 154816 185580 154822 185592
rect 155678 185580 155684 185592
rect 155736 185580 155742 185632
rect 156138 185580 156144 185632
rect 156196 185620 156202 185632
rect 157058 185620 157064 185632
rect 156196 185592 157064 185620
rect 156196 185580 156202 185592
rect 157058 185580 157064 185592
rect 157116 185580 157122 185632
rect 157518 185580 157524 185632
rect 157576 185620 157582 185632
rect 158438 185620 158444 185632
rect 157576 185592 158444 185620
rect 157576 185580 157582 185592
rect 158438 185580 158444 185592
rect 158496 185580 158502 185632
rect 160094 185580 160100 185632
rect 160152 185620 160158 185632
rect 160922 185620 160928 185632
rect 160152 185592 160928 185620
rect 160152 185580 160158 185592
rect 160922 185580 160928 185592
rect 160980 185580 160986 185632
rect 161382 185580 161388 185632
rect 161440 185620 161446 185632
rect 168374 185620 168380 185632
rect 161440 185592 168380 185620
rect 161440 185580 161446 185592
rect 168374 185580 168380 185592
rect 168432 185580 168438 185632
rect 169754 185580 169760 185632
rect 169812 185620 169818 185632
rect 170306 185620 170312 185632
rect 169812 185592 170312 185620
rect 169812 185580 169818 185592
rect 170306 185580 170312 185592
rect 170364 185580 170370 185632
rect 172606 185580 172612 185632
rect 172664 185620 172670 185632
rect 173250 185620 173256 185632
rect 172664 185592 173256 185620
rect 172664 185580 172670 185592
rect 173250 185580 173256 185592
rect 173308 185580 173314 185632
rect 175274 185580 175280 185632
rect 175332 185620 175338 185632
rect 175826 185620 175832 185632
rect 175332 185592 175832 185620
rect 175332 185580 175338 185592
rect 175826 185580 175832 185592
rect 175884 185580 175890 185632
rect 104342 185512 104348 185564
rect 104400 185552 104406 185564
rect 135162 185552 135168 185564
rect 104400 185524 135168 185552
rect 104400 185512 104406 185524
rect 135162 185512 135168 185524
rect 135220 185512 135226 185564
rect 142430 185512 142436 185564
rect 142488 185552 142494 185564
rect 142706 185552 142712 185564
rect 142488 185524 142712 185552
rect 142488 185512 142494 185524
rect 142706 185512 142712 185524
rect 142764 185512 142770 185564
rect 156782 185512 156788 185564
rect 156840 185552 156846 185564
rect 157242 185552 157248 185564
rect 156840 185524 157248 185552
rect 156840 185512 156846 185524
rect 157242 185512 157248 185524
rect 157300 185512 157306 185564
rect 167270 185512 167276 185564
rect 167328 185552 167334 185564
rect 167638 185552 167644 185564
rect 167328 185524 167644 185552
rect 167328 185512 167334 185524
rect 167638 185512 167644 185524
rect 167696 185512 167702 185564
rect 121362 185308 121368 185360
rect 121420 185348 121426 185360
rect 142154 185348 142160 185360
rect 121420 185320 142160 185348
rect 121420 185308 121426 185320
rect 142154 185308 142160 185320
rect 142212 185308 142218 185360
rect 108574 185172 108580 185224
rect 108632 185212 108638 185224
rect 132494 185212 132500 185224
rect 108632 185184 132500 185212
rect 108632 185172 108638 185184
rect 132494 185172 132500 185184
rect 132552 185172 132558 185224
rect 127802 185104 127808 185156
rect 127860 185144 127866 185156
rect 144270 185144 144276 185156
rect 127860 185116 144276 185144
rect 127860 185104 127866 185116
rect 144270 185104 144276 185116
rect 144328 185104 144334 185156
rect 108390 184968 108396 185020
rect 108448 185008 108454 185020
rect 137738 185008 137744 185020
rect 108448 184980 137744 185008
rect 108448 184968 108454 184980
rect 137738 184968 137744 184980
rect 137796 184968 137802 185020
rect 160278 184968 160284 185020
rect 160336 185008 160342 185020
rect 160646 185008 160652 185020
rect 160336 184980 160652 185008
rect 160336 184968 160342 184980
rect 160646 184968 160652 184980
rect 160704 184968 160710 185020
rect 150618 184560 150624 184612
rect 150676 184600 150682 184612
rect 150986 184600 150992 184612
rect 150676 184572 150992 184600
rect 150676 184560 150682 184572
rect 150986 184560 150992 184572
rect 151044 184560 151050 184612
rect 107010 184356 107016 184408
rect 107068 184396 107074 184408
rect 136082 184396 136088 184408
rect 107068 184368 136088 184396
rect 107068 184356 107074 184368
rect 136082 184356 136088 184368
rect 136140 184356 136146 184408
rect 126882 184288 126888 184340
rect 126940 184328 126946 184340
rect 144914 184328 144920 184340
rect 126940 184300 144920 184328
rect 126940 184288 126946 184300
rect 144914 184288 144920 184300
rect 144972 184288 144978 184340
rect 150802 184288 150808 184340
rect 150860 184328 150866 184340
rect 151262 184328 151268 184340
rect 150860 184300 151268 184328
rect 150860 184288 150866 184300
rect 151262 184288 151268 184300
rect 151320 184288 151326 184340
rect 102870 184152 102876 184204
rect 102928 184192 102934 184204
rect 134058 184192 134064 184204
rect 102928 184164 134064 184192
rect 102928 184152 102934 184164
rect 134058 184152 134064 184164
rect 134116 184152 134122 184204
rect 146754 184152 146760 184204
rect 146812 184192 146818 184204
rect 148042 184192 148048 184204
rect 146812 184164 148048 184192
rect 146812 184152 146818 184164
rect 148042 184152 148048 184164
rect 148100 184152 148106 184204
rect 172422 184016 172428 184068
rect 172480 184056 172486 184068
rect 196802 184056 196808 184068
rect 172480 184028 196808 184056
rect 172480 184016 172486 184028
rect 196802 184016 196808 184028
rect 196860 184016 196866 184068
rect 121270 183744 121276 183796
rect 121328 183784 121334 183796
rect 139118 183784 139124 183796
rect 121328 183756 139124 183784
rect 121328 183744 121334 183756
rect 139118 183744 139124 183756
rect 139176 183744 139182 183796
rect 164418 183268 164424 183320
rect 164476 183308 164482 183320
rect 165338 183308 165344 183320
rect 164476 183280 165344 183308
rect 164476 183268 164482 183280
rect 165338 183268 165344 183280
rect 165396 183268 165402 183320
rect 175458 183064 175464 183116
rect 175516 183104 175522 183116
rect 176194 183104 176200 183116
rect 175516 183076 176200 183104
rect 175516 183064 175522 183076
rect 176194 183064 176200 183076
rect 176252 183064 176258 183116
rect 150342 182996 150348 183048
rect 150400 183036 150406 183048
rect 156322 183036 156328 183048
rect 150400 183008 156328 183036
rect 150400 182996 150406 183008
rect 156322 182996 156328 183008
rect 156380 182996 156386 183048
rect 164234 182860 164240 182912
rect 164292 182900 164298 182912
rect 164602 182900 164608 182912
rect 164292 182872 164608 182900
rect 164292 182860 164298 182872
rect 164602 182860 164608 182872
rect 164660 182860 164666 182912
rect 164234 182724 164240 182776
rect 164292 182764 164298 182776
rect 165062 182764 165068 182776
rect 164292 182736 165068 182764
rect 164292 182724 164298 182736
rect 165062 182724 165068 182736
rect 165120 182724 165126 182776
rect 147582 182656 147588 182708
rect 147640 182696 147646 182708
rect 155218 182696 155224 182708
rect 147640 182668 155224 182696
rect 147640 182656 147646 182668
rect 155218 182656 155224 182668
rect 155276 182656 155282 182708
rect 104526 182520 104532 182572
rect 104584 182560 104590 182572
rect 133322 182560 133328 182572
rect 104584 182532 133328 182560
rect 104584 182520 104590 182532
rect 133322 182520 133328 182532
rect 133380 182520 133386 182572
rect 108482 182112 108488 182164
rect 108540 182152 108546 182164
rect 136818 182152 136824 182164
rect 108540 182124 136824 182152
rect 108540 182112 108546 182124
rect 136818 182112 136824 182124
rect 136876 182112 136882 182164
rect 149514 181976 149520 182028
rect 149572 182016 149578 182028
rect 149974 182016 149980 182028
rect 149572 181988 149980 182016
rect 149572 181976 149578 181988
rect 149974 181976 149980 181988
rect 150032 181976 150038 182028
rect 172514 181976 172520 182028
rect 172572 182016 172578 182028
rect 173618 182016 173624 182028
rect 172572 181988 173624 182016
rect 172572 181976 172578 181988
rect 173618 181976 173624 181988
rect 173676 181976 173682 182028
rect 104158 181568 104164 181620
rect 104216 181608 104222 181620
rect 132586 181608 132592 181620
rect 104216 181580 132592 181608
rect 104216 181568 104222 181580
rect 132586 181568 132592 181580
rect 132644 181568 132650 181620
rect 132586 181432 132592 181484
rect 132644 181472 132650 181484
rect 133046 181472 133052 181484
rect 132644 181444 133052 181472
rect 132644 181432 132650 181444
rect 133046 181432 133052 181444
rect 133104 181432 133110 181484
rect 160186 181432 160192 181484
rect 160244 181472 160250 181484
rect 161290 181472 161296 181484
rect 160244 181444 161296 181472
rect 160244 181432 160250 181444
rect 161290 181432 161296 181444
rect 161348 181432 161354 181484
rect 150526 181160 150532 181212
rect 150584 181200 150590 181212
rect 151630 181200 151636 181212
rect 150584 181172 151636 181200
rect 150584 181160 150590 181172
rect 151630 181160 151636 181172
rect 151688 181160 151694 181212
rect 146846 180480 146852 180532
rect 146904 180520 146910 180532
rect 147398 180520 147404 180532
rect 146904 180492 147404 180520
rect 146904 180480 146910 180492
rect 147398 180480 147404 180492
rect 147456 180480 147462 180532
rect 128998 180344 129004 180396
rect 129056 180384 129062 180396
rect 140866 180384 140872 180396
rect 129056 180356 140872 180384
rect 129056 180344 129062 180356
rect 140866 180344 140872 180356
rect 140924 180344 140930 180396
rect 151998 179936 152004 179988
rect 152056 179976 152062 179988
rect 152642 179976 152648 179988
rect 152056 179948 152648 179976
rect 152056 179936 152062 179948
rect 152642 179936 152648 179948
rect 152700 179936 152706 179988
rect 161658 179936 161664 179988
rect 161716 179976 161722 179988
rect 162302 179976 162308 179988
rect 161716 179948 162308 179976
rect 161716 179936 161722 179948
rect 162302 179936 162308 179948
rect 162360 179936 162366 179988
rect 157426 179800 157432 179852
rect 157484 179840 157490 179852
rect 157886 179840 157892 179852
rect 157484 179812 157892 179840
rect 157484 179800 157490 179812
rect 157886 179800 157892 179812
rect 157944 179800 157950 179852
rect 161290 179120 161296 179172
rect 161348 179160 161354 179172
rect 162118 179160 162124 179172
rect 161348 179132 162124 179160
rect 161348 179120 161354 179132
rect 162118 179120 162124 179132
rect 162176 179120 162182 179172
rect 163130 179120 163136 179172
rect 163188 179160 163194 179172
rect 163774 179160 163780 179172
rect 163188 179132 163780 179160
rect 163188 179120 163194 179132
rect 163774 179120 163780 179132
rect 163832 179120 163838 179172
rect 135622 178984 135628 179036
rect 135680 179024 135686 179036
rect 136174 179024 136180 179036
rect 135680 178996 136180 179024
rect 135680 178984 135686 178996
rect 136174 178984 136180 178996
rect 136232 178984 136238 179036
rect 145558 178984 145564 179036
rect 145616 179024 145622 179036
rect 149054 179024 149060 179036
rect 145616 178996 149060 179024
rect 145616 178984 145622 178996
rect 149054 178984 149060 178996
rect 149112 178984 149118 179036
rect 149698 178712 149704 178764
rect 149756 178752 149762 178764
rect 153562 178752 153568 178764
rect 149756 178724 153568 178752
rect 149756 178712 149762 178724
rect 153562 178712 153568 178724
rect 153620 178712 153626 178764
rect 108206 178440 108212 178492
rect 108264 178480 108270 178492
rect 137922 178480 137928 178492
rect 108264 178452 137928 178480
rect 108264 178440 108270 178452
rect 137922 178440 137928 178452
rect 137980 178440 137986 178492
rect 142430 178440 142436 178492
rect 142488 178480 142494 178492
rect 143258 178480 143264 178492
rect 142488 178452 143264 178480
rect 142488 178440 142494 178452
rect 143258 178440 143264 178452
rect 143316 178440 143322 178492
rect 171226 178236 171232 178288
rect 171284 178276 171290 178288
rect 172330 178276 172336 178288
rect 171284 178248 172336 178276
rect 171284 178236 171290 178248
rect 172330 178236 172336 178248
rect 172388 178236 172394 178288
rect 175642 178032 175648 178084
rect 175700 178072 175706 178084
rect 176378 178072 176384 178084
rect 175700 178044 176384 178072
rect 175700 178032 175706 178044
rect 176378 178032 176384 178044
rect 176436 178032 176442 178084
rect 188430 178032 188436 178084
rect 188488 178072 188494 178084
rect 580166 178072 580172 178084
rect 188488 178044 580172 178072
rect 188488 178032 188494 178044
rect 580166 178032 580172 178044
rect 580224 178032 580230 178084
rect 146938 177148 146944 177200
rect 146996 177188 147002 177200
rect 147766 177188 147772 177200
rect 146996 177160 147772 177188
rect 146996 177148 147002 177160
rect 147766 177148 147772 177160
rect 147824 177148 147830 177200
rect 102962 176944 102968 176996
rect 103020 176984 103026 176996
rect 134610 176984 134616 176996
rect 103020 176956 134616 176984
rect 103020 176944 103026 176956
rect 134610 176944 134616 176956
rect 134668 176944 134674 176996
rect 167086 176944 167092 176996
rect 167144 176984 167150 176996
rect 168190 176984 168196 176996
rect 167144 176956 168196 176984
rect 167144 176944 167150 176956
rect 168190 176944 168196 176956
rect 168248 176944 168254 176996
rect 104710 176400 104716 176452
rect 104768 176440 104774 176452
rect 132954 176440 132960 176452
rect 104768 176412 132960 176440
rect 104768 176400 104774 176412
rect 132954 176400 132960 176412
rect 133012 176400 133018 176452
rect 145190 175856 145196 175908
rect 145248 175896 145254 175908
rect 146294 175896 146300 175908
rect 145248 175868 146300 175896
rect 145248 175856 145254 175868
rect 146294 175856 146300 175868
rect 146352 175856 146358 175908
rect 164326 175720 164332 175772
rect 164384 175760 164390 175772
rect 164786 175760 164792 175772
rect 164384 175732 164792 175760
rect 164384 175720 164390 175732
rect 164786 175720 164792 175732
rect 164844 175720 164850 175772
rect 158990 175176 158996 175228
rect 159048 175216 159054 175228
rect 159358 175216 159364 175228
rect 159048 175188 159364 175216
rect 159048 175176 159054 175188
rect 159358 175176 159364 175188
rect 159416 175176 159422 175228
rect 171318 175176 171324 175228
rect 171376 175216 171382 175228
rect 171778 175216 171784 175228
rect 171376 175188 171784 175216
rect 171376 175176 171382 175188
rect 171778 175176 171784 175188
rect 171836 175176 171842 175228
rect 107102 174224 107108 174276
rect 107160 174264 107166 174276
rect 136266 174264 136272 174276
rect 107160 174236 136272 174264
rect 107160 174224 107166 174236
rect 136266 174224 136272 174236
rect 136324 174224 136330 174276
rect 132678 174088 132684 174140
rect 132736 174128 132742 174140
rect 133506 174128 133512 174140
rect 132736 174100 133512 174128
rect 132736 174088 132742 174100
rect 133506 174088 133512 174100
rect 133564 174088 133570 174140
rect 137002 173544 137008 173596
rect 137060 173584 137066 173596
rect 137370 173584 137376 173596
rect 137060 173556 137376 173584
rect 137060 173544 137066 173556
rect 137370 173544 137376 173556
rect 137428 173544 137434 173596
rect 117866 166268 117872 166320
rect 117924 166308 117930 166320
rect 580166 166308 580172 166320
rect 117924 166280 580172 166308
rect 117924 166268 117930 166280
rect 580166 166268 580172 166280
rect 580224 166268 580230 166320
rect 165798 155660 165804 155712
rect 165856 155700 165862 155712
rect 200390 155700 200396 155712
rect 165856 155672 200396 155700
rect 165856 155660 165862 155672
rect 200390 155660 200396 155672
rect 200448 155660 200454 155712
rect 167270 155592 167276 155644
rect 167328 155632 167334 155644
rect 201862 155632 201868 155644
rect 167328 155604 201868 155632
rect 167328 155592 167334 155604
rect 201862 155592 201868 155604
rect 201920 155592 201926 155644
rect 167362 155524 167368 155576
rect 167420 155564 167426 155576
rect 201954 155564 201960 155576
rect 167420 155536 201960 155564
rect 167420 155524 167426 155536
rect 201954 155524 201960 155536
rect 202012 155524 202018 155576
rect 165890 155456 165896 155508
rect 165948 155496 165954 155508
rect 200574 155496 200580 155508
rect 165948 155468 200580 155496
rect 165948 155456 165954 155468
rect 200574 155456 200580 155468
rect 200632 155456 200638 155508
rect 168650 155388 168656 155440
rect 168708 155428 168714 155440
rect 203334 155428 203340 155440
rect 168708 155400 203340 155428
rect 168708 155388 168714 155400
rect 203334 155388 203340 155400
rect 203392 155388 203398 155440
rect 168558 155320 168564 155372
rect 168616 155360 168622 155372
rect 203518 155360 203524 155372
rect 168616 155332 203524 155360
rect 168616 155320 168622 155332
rect 203518 155320 203524 155332
rect 203576 155320 203582 155372
rect 168466 155252 168472 155304
rect 168524 155292 168530 155304
rect 203426 155292 203432 155304
rect 168524 155264 203432 155292
rect 168524 155252 168530 155264
rect 203426 155252 203432 155264
rect 203484 155252 203490 155304
rect 167178 155184 167184 155236
rect 167236 155224 167242 155236
rect 202138 155224 202144 155236
rect 167236 155196 202144 155224
rect 167236 155184 167242 155196
rect 202138 155184 202144 155196
rect 202196 155184 202202 155236
rect 160370 153144 160376 153196
rect 160428 153184 160434 153196
rect 185670 153184 185676 153196
rect 160428 153156 185676 153184
rect 160428 153144 160434 153156
rect 185670 153144 185676 153156
rect 185728 153144 185734 153196
rect 159082 153076 159088 153128
rect 159140 153116 159146 153128
rect 184382 153116 184388 153128
rect 159140 153088 184388 153116
rect 159140 153076 159146 153088
rect 184382 153076 184388 153088
rect 184440 153076 184446 153128
rect 160278 153008 160284 153060
rect 160336 153048 160342 153060
rect 185762 153048 185768 153060
rect 160336 153020 185768 153048
rect 160336 153008 160342 153020
rect 185762 153008 185768 153020
rect 185820 153008 185826 153060
rect 158990 152940 158996 152992
rect 159048 152980 159054 152992
rect 184474 152980 184480 152992
rect 159048 152952 184480 152980
rect 159048 152940 159054 152952
rect 184474 152940 184480 152952
rect 184532 152940 184538 152992
rect 158898 152872 158904 152924
rect 158956 152912 158962 152924
rect 185854 152912 185860 152924
rect 158956 152884 185860 152912
rect 158956 152872 158962 152884
rect 185854 152872 185860 152884
rect 185912 152872 185918 152924
rect 163222 152804 163228 152856
rect 163280 152844 163286 152856
rect 198182 152844 198188 152856
rect 163280 152816 198188 152844
rect 163280 152804 163286 152816
rect 198182 152804 198188 152816
rect 198240 152804 198246 152856
rect 164510 152736 164516 152788
rect 164568 152776 164574 152788
rect 199746 152776 199752 152788
rect 164568 152748 199752 152776
rect 164568 152736 164574 152748
rect 199746 152736 199752 152748
rect 199804 152736 199810 152788
rect 164602 152668 164608 152720
rect 164660 152708 164666 152720
rect 199378 152708 199384 152720
rect 164660 152680 199384 152708
rect 164660 152668 164666 152680
rect 199378 152668 199384 152680
rect 199436 152668 199442 152720
rect 149330 152600 149336 152652
rect 149388 152640 149394 152652
rect 204714 152640 204720 152652
rect 149388 152612 204720 152640
rect 149388 152600 149394 152612
rect 204714 152600 204720 152612
rect 204772 152600 204778 152652
rect 146478 152532 146484 152584
rect 146536 152572 146542 152584
rect 204806 152572 204812 152584
rect 146536 152544 204812 152572
rect 146536 152532 146542 152544
rect 204806 152532 204812 152544
rect 204864 152532 204870 152584
rect 147858 152464 147864 152516
rect 147916 152504 147922 152516
rect 206186 152504 206192 152516
rect 147916 152476 206192 152504
rect 147916 152464 147922 152476
rect 206186 152464 206192 152476
rect 206244 152464 206250 152516
rect 160462 152396 160468 152448
rect 160520 152436 160526 152448
rect 184566 152436 184572 152448
rect 160520 152408 184572 152436
rect 160520 152396 160526 152408
rect 184566 152396 184572 152408
rect 184624 152396 184630 152448
rect 161750 152328 161756 152380
rect 161808 152368 161814 152380
rect 184658 152368 184664 152380
rect 161808 152340 184664 152368
rect 161808 152328 161814 152340
rect 184658 152328 184664 152340
rect 184716 152328 184722 152380
rect 161658 152260 161664 152312
rect 161716 152300 161722 152312
rect 184198 152300 184204 152312
rect 161716 152272 184204 152300
rect 161716 152260 161722 152272
rect 184198 152260 184204 152272
rect 184256 152260 184262 152312
rect 161382 151036 161388 151088
rect 161440 151076 161446 151088
rect 203242 151076 203248 151088
rect 161440 151048 203248 151076
rect 161440 151036 161446 151048
rect 203242 151036 203248 151048
rect 203300 151036 203306 151088
rect 179046 150356 179052 150408
rect 179104 150396 179110 150408
rect 205818 150396 205824 150408
rect 179104 150368 205824 150396
rect 179104 150356 179110 150368
rect 205818 150356 205824 150368
rect 205876 150356 205882 150408
rect 176838 150288 176844 150340
rect 176896 150328 176902 150340
rect 204898 150328 204904 150340
rect 176896 150300 204904 150328
rect 176896 150288 176902 150300
rect 204898 150288 204904 150300
rect 204956 150288 204962 150340
rect 174078 150220 174084 150272
rect 174136 150260 174142 150272
rect 202322 150260 202328 150272
rect 174136 150232 202328 150260
rect 174136 150220 174142 150232
rect 202322 150220 202328 150232
rect 202380 150220 202386 150272
rect 175642 150152 175648 150204
rect 175700 150192 175706 150204
rect 204438 150192 204444 150204
rect 175700 150164 204444 150192
rect 175700 150152 175706 150164
rect 204438 150152 204444 150164
rect 204496 150152 204502 150204
rect 176930 150084 176936 150136
rect 176988 150124 176994 150136
rect 206278 150124 206284 150136
rect 176988 150096 206284 150124
rect 176988 150084 176994 150096
rect 206278 150084 206284 150096
rect 206336 150084 206342 150136
rect 175550 150016 175556 150068
rect 175608 150056 175614 150068
rect 205910 150056 205916 150068
rect 175608 150028 205916 150056
rect 175608 150016 175614 150028
rect 205910 150016 205916 150028
rect 205968 150016 205974 150068
rect 175458 149948 175464 150000
rect 175516 149988 175522 150000
rect 206094 149988 206100 150000
rect 175516 149960 206100 149988
rect 175516 149948 175522 149960
rect 206094 149948 206100 149960
rect 206152 149948 206158 150000
rect 175366 149880 175372 149932
rect 175424 149920 175430 149932
rect 206002 149920 206008 149932
rect 175424 149892 206008 149920
rect 175424 149880 175430 149892
rect 206002 149880 206008 149892
rect 206060 149880 206066 149932
rect 172882 149812 172888 149864
rect 172940 149852 172946 149864
rect 203702 149852 203708 149864
rect 172940 149824 203708 149852
rect 172940 149812 172946 149824
rect 203702 149812 203708 149824
rect 203760 149812 203766 149864
rect 175274 149744 175280 149796
rect 175332 149784 175338 149796
rect 206370 149784 206376 149796
rect 175332 149756 206376 149784
rect 175332 149744 175338 149756
rect 206370 149744 206376 149756
rect 206428 149744 206434 149796
rect 148962 149676 148968 149728
rect 149020 149716 149026 149728
rect 184750 149716 184756 149728
rect 149020 149688 184756 149716
rect 149020 149676 149026 149688
rect 184750 149676 184756 149688
rect 184808 149676 184814 149728
rect 173066 149608 173072 149660
rect 173124 149648 173130 149660
rect 186958 149648 186964 149660
rect 173124 149620 186964 149648
rect 173124 149608 173130 149620
rect 186958 149608 186964 149620
rect 187016 149608 187022 149660
rect 182082 149540 182088 149592
rect 182140 149580 182146 149592
rect 192662 149580 192668 149592
rect 182140 149552 192668 149580
rect 182140 149540 182146 149552
rect 192662 149540 192668 149552
rect 192720 149540 192726 149592
rect 3418 149064 3424 149116
rect 3476 149104 3482 149116
rect 180886 149104 180892 149116
rect 3476 149076 180892 149104
rect 3476 149064 3482 149076
rect 180886 149064 180892 149076
rect 180944 149104 180950 149116
rect 182082 149104 182088 149116
rect 180944 149076 182088 149104
rect 180944 149064 180950 149076
rect 182082 149064 182088 149076
rect 182140 149064 182146 149116
rect 122374 148996 122380 149048
rect 122432 149036 122438 149048
rect 152182 149036 152188 149048
rect 122432 149008 152188 149036
rect 122432 148996 122438 149008
rect 152182 148996 152188 149008
rect 152240 148996 152246 149048
rect 162946 148996 162952 149048
rect 163004 149036 163010 149048
rect 185302 149036 185308 149048
rect 163004 149008 185308 149036
rect 163004 148996 163010 149008
rect 185302 148996 185308 149008
rect 185360 148996 185366 149048
rect 112162 148928 112168 148980
rect 112220 148968 112226 148980
rect 142982 148968 142988 148980
rect 112220 148940 142988 148968
rect 112220 148928 112226 148940
rect 142982 148928 142988 148940
rect 143040 148928 143046 148980
rect 161566 148928 161572 148980
rect 161624 148968 161630 148980
rect 186314 148968 186320 148980
rect 161624 148940 186320 148968
rect 161624 148928 161630 148940
rect 186314 148928 186320 148940
rect 186372 148928 186378 148980
rect 108114 148860 108120 148912
rect 108172 148900 108178 148912
rect 139854 148900 139860 148912
rect 108172 148872 139860 148900
rect 108172 148860 108178 148872
rect 139854 148860 139860 148872
rect 139912 148860 139918 148912
rect 164418 148860 164424 148912
rect 164476 148900 164482 148912
rect 197906 148900 197912 148912
rect 164476 148872 197912 148900
rect 164476 148860 164482 148872
rect 197906 148860 197912 148872
rect 197964 148860 197970 148912
rect 100202 148792 100208 148844
rect 100260 148832 100266 148844
rect 132862 148832 132868 148844
rect 100260 148804 132868 148832
rect 100260 148792 100266 148804
rect 132862 148792 132868 148804
rect 132920 148792 132926 148844
rect 163038 148792 163044 148844
rect 163096 148832 163102 148844
rect 197814 148832 197820 148844
rect 163096 148804 197820 148832
rect 163096 148792 163102 148804
rect 197814 148792 197820 148804
rect 197872 148792 197878 148844
rect 100386 148724 100392 148776
rect 100444 148764 100450 148776
rect 132678 148764 132684 148776
rect 100444 148736 132684 148764
rect 100444 148724 100450 148736
rect 132678 148724 132684 148736
rect 132736 148724 132742 148776
rect 161474 148724 161480 148776
rect 161532 148764 161538 148776
rect 196894 148764 196900 148776
rect 161532 148736 196900 148764
rect 161532 148724 161538 148736
rect 196894 148724 196900 148736
rect 196952 148724 196958 148776
rect 117682 148656 117688 148708
rect 117740 148696 117746 148708
rect 150710 148696 150716 148708
rect 117740 148668 150716 148696
rect 117740 148656 117746 148668
rect 150710 148656 150716 148668
rect 150768 148656 150774 148708
rect 167086 148656 167092 148708
rect 167144 148696 167150 148708
rect 202046 148696 202052 148708
rect 167144 148668 202052 148696
rect 167144 148656 167150 148668
rect 202046 148656 202052 148668
rect 202104 148656 202110 148708
rect 102686 148588 102692 148640
rect 102744 148628 102750 148640
rect 135622 148628 135628 148640
rect 102744 148600 135628 148628
rect 102744 148588 102750 148600
rect 135622 148588 135628 148600
rect 135680 148588 135686 148640
rect 166810 148588 166816 148640
rect 166868 148628 166874 148640
rect 200666 148628 200672 148640
rect 166868 148600 200672 148628
rect 166868 148588 166874 148600
rect 200666 148588 200672 148600
rect 200724 148588 200730 148640
rect 103974 148520 103980 148572
rect 104032 148560 104038 148572
rect 137186 148560 137192 148572
rect 104032 148532 137192 148560
rect 104032 148520 104038 148532
rect 137186 148520 137192 148532
rect 137244 148520 137250 148572
rect 164326 148520 164332 148572
rect 164384 148560 164390 148572
rect 199470 148560 199476 148572
rect 164384 148532 199476 148560
rect 164384 148520 164390 148532
rect 199470 148520 199476 148532
rect 199528 148520 199534 148572
rect 100294 148452 100300 148504
rect 100352 148492 100358 148504
rect 134242 148492 134248 148504
rect 100352 148464 134248 148492
rect 100352 148452 100358 148464
rect 134242 148452 134248 148464
rect 134300 148452 134306 148504
rect 167914 148452 167920 148504
rect 167972 148492 167978 148504
rect 202230 148492 202236 148504
rect 167972 148464 202236 148492
rect 167972 148452 167978 148464
rect 202230 148452 202236 148464
rect 202288 148452 202294 148504
rect 116302 148384 116308 148436
rect 116360 148424 116366 148436
rect 150802 148424 150808 148436
rect 116360 148396 150808 148424
rect 116360 148384 116366 148396
rect 150802 148384 150808 148396
rect 150860 148384 150866 148436
rect 169202 148384 169208 148436
rect 169260 148424 169266 148436
rect 203610 148424 203616 148436
rect 169260 148396 203616 148424
rect 169260 148384 169266 148396
rect 203610 148384 203616 148396
rect 203668 148384 203674 148436
rect 100110 148316 100116 148368
rect 100168 148356 100174 148368
rect 134334 148356 134340 148368
rect 100168 148328 134340 148356
rect 100168 148316 100174 148328
rect 134334 148316 134340 148328
rect 134392 148316 134398 148368
rect 164234 148316 164240 148368
rect 164292 148356 164298 148368
rect 199562 148356 199568 148368
rect 164292 148328 199568 148356
rect 164292 148316 164298 148328
rect 199562 148316 199568 148328
rect 199620 148316 199626 148368
rect 123938 148248 123944 148300
rect 123996 148288 124002 148300
rect 152090 148288 152096 148300
rect 123996 148260 152096 148288
rect 123996 148248 124002 148260
rect 152090 148248 152096 148260
rect 152148 148248 152154 148300
rect 185026 148248 185032 148300
rect 185084 148288 185090 148300
rect 199286 148288 199292 148300
rect 185084 148260 199292 148288
rect 185084 148248 185090 148260
rect 199286 148248 199292 148260
rect 199344 148248 199350 148300
rect 113542 148180 113548 148232
rect 113600 148220 113606 148232
rect 142430 148220 142436 148232
rect 113600 148192 142436 148220
rect 113600 148180 113606 148192
rect 142430 148180 142436 148192
rect 142488 148180 142494 148232
rect 180150 148180 180156 148232
rect 180208 148220 180214 148232
rect 192846 148220 192852 148232
rect 180208 148192 192852 148220
rect 180208 148180 180214 148192
rect 192846 148180 192852 148192
rect 192904 148180 192910 148232
rect 122190 148112 122196 148164
rect 122248 148152 122254 148164
rect 149698 148152 149704 148164
rect 122248 148124 149704 148152
rect 122248 148112 122254 148124
rect 149698 148112 149704 148124
rect 149756 148112 149762 148164
rect 179322 147568 179328 147620
rect 179380 147608 179386 147620
rect 196710 147608 196716 147620
rect 179380 147580 196716 147608
rect 179380 147568 179386 147580
rect 196710 147568 196716 147580
rect 196768 147568 196774 147620
rect 171502 147500 171508 147552
rect 171560 147540 171566 147552
rect 194962 147540 194968 147552
rect 171560 147512 194968 147540
rect 171560 147500 171566 147512
rect 194962 147500 194968 147512
rect 195020 147500 195026 147552
rect 171226 147432 171232 147484
rect 171284 147472 171290 147484
rect 195330 147472 195336 147484
rect 171284 147444 195336 147472
rect 171284 147432 171290 147444
rect 195330 147432 195336 147444
rect 195388 147432 195394 147484
rect 171318 147364 171324 147416
rect 171376 147404 171382 147416
rect 196986 147404 196992 147416
rect 171376 147376 196992 147404
rect 171376 147364 171382 147376
rect 196986 147364 196992 147376
rect 197044 147364 197050 147416
rect 169938 147296 169944 147348
rect 169996 147336 170002 147348
rect 197078 147336 197084 147348
rect 169996 147308 197084 147336
rect 169996 147296 170002 147308
rect 197078 147296 197084 147308
rect 197136 147296 197142 147348
rect 171410 147228 171416 147280
rect 171468 147268 171474 147280
rect 198090 147268 198096 147280
rect 171468 147240 198096 147268
rect 171468 147228 171474 147240
rect 198090 147228 198096 147240
rect 198148 147228 198154 147280
rect 172790 147160 172796 147212
rect 172848 147200 172854 147212
rect 200942 147200 200948 147212
rect 172848 147172 200948 147200
rect 172848 147160 172854 147172
rect 200942 147160 200948 147172
rect 201000 147160 201006 147212
rect 172698 147092 172704 147144
rect 172756 147132 172762 147144
rect 200850 147132 200856 147144
rect 172756 147104 200856 147132
rect 172756 147092 172762 147104
rect 200850 147092 200856 147104
rect 200908 147092 200914 147144
rect 164142 147024 164148 147076
rect 164200 147064 164206 147076
rect 193950 147064 193956 147076
rect 164200 147036 193956 147064
rect 164200 147024 164206 147036
rect 193950 147024 193956 147036
rect 194008 147024 194014 147076
rect 111058 146956 111064 147008
rect 111116 146996 111122 147008
rect 130194 146996 130200 147008
rect 111116 146968 130200 146996
rect 111116 146956 111122 146968
rect 130194 146956 130200 146968
rect 130252 146956 130258 147008
rect 172606 146956 172612 147008
rect 172664 146996 172670 147008
rect 204530 146996 204536 147008
rect 172664 146968 204536 146996
rect 172664 146956 172670 146968
rect 204530 146956 204536 146968
rect 204588 146956 204594 147008
rect 113450 146888 113456 146940
rect 113508 146928 113514 146940
rect 142706 146928 142712 146940
rect 113508 146900 142712 146928
rect 113508 146888 113514 146900
rect 142706 146888 142712 146900
rect 142764 146888 142770 146940
rect 170030 146888 170036 146940
rect 170088 146928 170094 146940
rect 204622 146928 204628 146940
rect 170088 146900 204628 146928
rect 170088 146888 170094 146900
rect 204622 146888 204628 146900
rect 204680 146888 204686 146940
rect 178586 146820 178592 146872
rect 178644 146860 178650 146872
rect 196434 146860 196440 146872
rect 178644 146832 196440 146860
rect 178644 146820 178650 146832
rect 196434 146820 196440 146832
rect 196492 146820 196498 146872
rect 130194 146276 130200 146328
rect 130252 146316 130258 146328
rect 580350 146316 580356 146328
rect 130252 146288 580356 146316
rect 130252 146276 130258 146288
rect 580350 146276 580356 146288
rect 580408 146276 580414 146328
rect 3510 146208 3516 146260
rect 3568 146248 3574 146260
rect 179046 146248 179052 146260
rect 3568 146220 179052 146248
rect 3568 146208 3574 146220
rect 179046 146208 179052 146220
rect 179104 146208 179110 146260
rect 179782 146208 179788 146260
rect 179840 146248 179846 146260
rect 192294 146248 192300 146260
rect 179840 146220 192300 146248
rect 179840 146208 179846 146220
rect 192294 146208 192300 146220
rect 192352 146208 192358 146260
rect 113818 146140 113824 146192
rect 113876 146180 113882 146192
rect 130746 146180 130752 146192
rect 113876 146152 130752 146180
rect 113876 146140 113882 146152
rect 130746 146140 130752 146152
rect 130804 146140 130810 146192
rect 183462 146140 183468 146192
rect 183520 146180 183526 146192
rect 196526 146180 196532 146192
rect 183520 146152 196532 146180
rect 183520 146140 183526 146152
rect 196526 146140 196532 146152
rect 196584 146140 196590 146192
rect 114278 146072 114284 146124
rect 114336 146112 114342 146124
rect 132402 146112 132408 146124
rect 114336 146084 132408 146112
rect 114336 146072 114342 146084
rect 132402 146072 132408 146084
rect 132460 146072 132466 146124
rect 178034 146072 178040 146124
rect 178092 146112 178098 146124
rect 192570 146112 192576 146124
rect 178092 146084 192576 146112
rect 178092 146072 178098 146084
rect 192570 146072 192576 146084
rect 192628 146072 192634 146124
rect 112346 146004 112352 146056
rect 112404 146044 112410 146056
rect 131022 146044 131028 146056
rect 112404 146016 131028 146044
rect 112404 146004 112410 146016
rect 131022 146004 131028 146016
rect 131080 146004 131086 146056
rect 131758 146004 131764 146056
rect 131816 146044 131822 146056
rect 132218 146044 132224 146056
rect 131816 146016 132224 146044
rect 131816 146004 131822 146016
rect 132218 146004 132224 146016
rect 132276 146004 132282 146056
rect 179598 146004 179604 146056
rect 179656 146044 179662 146056
rect 196618 146044 196624 146056
rect 179656 146016 196624 146044
rect 179656 146004 179662 146016
rect 196618 146004 196624 146016
rect 196676 146004 196682 146056
rect 117958 145936 117964 145988
rect 118016 145976 118022 145988
rect 146294 145976 146300 145988
rect 118016 145948 146300 145976
rect 118016 145936 118022 145948
rect 146294 145936 146300 145948
rect 146352 145936 146358 145988
rect 162210 145936 162216 145988
rect 162268 145976 162274 145988
rect 188522 145976 188528 145988
rect 162268 145948 188528 145976
rect 162268 145936 162274 145948
rect 188522 145936 188528 145948
rect 188580 145936 188586 145988
rect 119062 145868 119068 145920
rect 119120 145908 119126 145920
rect 150618 145908 150624 145920
rect 119120 145880 150624 145908
rect 119120 145868 119126 145880
rect 150618 145868 150624 145880
rect 150676 145868 150682 145920
rect 160186 145868 160192 145920
rect 160244 145908 160250 145920
rect 195514 145908 195520 145920
rect 160244 145880 195520 145908
rect 160244 145868 160250 145880
rect 195514 145868 195520 145880
rect 195572 145868 195578 145920
rect 117958 145800 117964 145852
rect 118016 145840 118022 145852
rect 149238 145840 149244 145852
rect 118016 145812 149244 145840
rect 118016 145800 118022 145812
rect 149238 145800 149244 145812
rect 149296 145800 149302 145852
rect 158530 145800 158536 145852
rect 158588 145840 158594 145852
rect 192754 145840 192760 145852
rect 158588 145812 192760 145840
rect 158588 145800 158594 145812
rect 192754 145800 192760 145812
rect 192812 145800 192818 145852
rect 114830 145732 114836 145784
rect 114888 145772 114894 145784
rect 149514 145772 149520 145784
rect 114888 145744 149520 145772
rect 114888 145732 114894 145744
rect 149514 145732 149520 145744
rect 149572 145732 149578 145784
rect 157426 145732 157432 145784
rect 157484 145772 157490 145784
rect 192294 145772 192300 145784
rect 157484 145744 192300 145772
rect 157484 145732 157490 145744
rect 192294 145732 192300 145744
rect 192352 145732 192358 145784
rect 114922 145664 114928 145716
rect 114980 145704 114986 145716
rect 149606 145704 149612 145716
rect 114980 145676 149612 145704
rect 114980 145664 114986 145676
rect 149606 145664 149612 145676
rect 149664 145664 149670 145716
rect 154482 145664 154488 145716
rect 154540 145704 154546 145716
rect 194318 145704 194324 145716
rect 154540 145676 194324 145704
rect 154540 145664 154546 145676
rect 194318 145664 194324 145676
rect 194376 145664 194382 145716
rect 114738 145596 114744 145648
rect 114796 145636 114802 145648
rect 145558 145636 145564 145648
rect 114796 145608 145564 145636
rect 114796 145596 114802 145608
rect 145558 145596 145564 145608
rect 145616 145596 145622 145648
rect 147582 145596 147588 145648
rect 147640 145636 147646 145648
rect 189994 145636 190000 145648
rect 147640 145608 190000 145636
rect 147640 145596 147646 145608
rect 189994 145596 190000 145608
rect 190052 145596 190058 145648
rect 112346 145528 112352 145580
rect 112404 145568 112410 145580
rect 142522 145568 142528 145580
rect 112404 145540 142528 145568
rect 112404 145528 112410 145540
rect 142522 145528 142528 145540
rect 142580 145528 142586 145580
rect 145190 145528 145196 145580
rect 145248 145568 145254 145580
rect 206462 145568 206468 145580
rect 145248 145540 206468 145568
rect 145248 145528 145254 145540
rect 206462 145528 206468 145540
rect 206520 145528 206526 145580
rect 115198 145460 115204 145512
rect 115256 145500 115262 145512
rect 130562 145500 130568 145512
rect 115256 145472 130568 145500
rect 115256 145460 115262 145472
rect 130562 145460 130568 145472
rect 130620 145460 130626 145512
rect 178126 145460 178132 145512
rect 178184 145500 178190 145512
rect 189626 145500 189632 145512
rect 178184 145472 189632 145500
rect 178184 145460 178190 145472
rect 189626 145460 189632 145472
rect 189684 145460 189690 145512
rect 115106 145392 115112 145444
rect 115164 145432 115170 145444
rect 129550 145432 129556 145444
rect 115164 145404 129556 145432
rect 115164 145392 115170 145404
rect 129550 145392 129556 145404
rect 129608 145392 129614 145444
rect 179506 145392 179512 145444
rect 179564 145432 179570 145444
rect 190914 145432 190920 145444
rect 179564 145404 190920 145432
rect 179564 145392 179570 145404
rect 190914 145392 190920 145404
rect 190972 145392 190978 145444
rect 179414 145324 179420 145376
rect 179472 145364 179478 145376
rect 189902 145364 189908 145376
rect 179472 145336 189908 145364
rect 179472 145324 179478 145336
rect 189902 145324 189908 145336
rect 189960 145324 189966 145376
rect 116118 144848 116124 144900
rect 116176 144888 116182 144900
rect 130470 144888 130476 144900
rect 116176 144860 130476 144888
rect 116176 144848 116182 144860
rect 130470 144848 130476 144860
rect 130528 144848 130534 144900
rect 180058 144848 180064 144900
rect 180116 144888 180122 144900
rect 191374 144888 191380 144900
rect 180116 144860 191380 144888
rect 180116 144848 180122 144860
rect 191374 144848 191380 144860
rect 191432 144848 191438 144900
rect 114278 144780 114284 144832
rect 114336 144820 114342 144832
rect 130378 144820 130384 144832
rect 114336 144792 130384 144820
rect 114336 144780 114342 144792
rect 130378 144780 130384 144792
rect 130436 144780 130442 144832
rect 174354 144780 174360 144832
rect 174412 144820 174418 144832
rect 189810 144820 189816 144832
rect 174412 144792 189816 144820
rect 174412 144780 174418 144792
rect 189810 144780 189816 144792
rect 189868 144780 189874 144832
rect 113634 144712 113640 144764
rect 113692 144752 113698 144764
rect 128998 144752 129004 144764
rect 113692 144724 129004 144752
rect 113692 144712 113698 144724
rect 128998 144712 129004 144724
rect 129056 144712 129062 144764
rect 171042 144712 171048 144764
rect 171100 144752 171106 144764
rect 192478 144752 192484 144764
rect 171100 144724 192484 144752
rect 171100 144712 171106 144724
rect 192478 144712 192484 144724
rect 192536 144712 192542 144764
rect 114186 144644 114192 144696
rect 114244 144684 114250 144696
rect 137278 144684 137284 144696
rect 114244 144656 137284 144684
rect 114244 144644 114250 144656
rect 137278 144644 137284 144656
rect 137336 144644 137342 144696
rect 172422 144644 172428 144696
rect 172480 144684 172486 144696
rect 193858 144684 193864 144696
rect 172480 144656 193864 144684
rect 172480 144644 172486 144656
rect 193858 144644 193864 144656
rect 193916 144644 193922 144696
rect 116578 144576 116584 144628
rect 116636 144616 116642 144628
rect 142246 144616 142252 144628
rect 116636 144588 142252 144616
rect 116636 144576 116642 144588
rect 142246 144576 142252 144588
rect 142304 144576 142310 144628
rect 162486 144576 162492 144628
rect 162544 144616 162550 144628
rect 191006 144616 191012 144628
rect 162544 144588 191012 144616
rect 162544 144576 162550 144588
rect 191006 144576 191012 144588
rect 191064 144576 191070 144628
rect 120534 144508 120540 144560
rect 120592 144548 120598 144560
rect 150526 144548 150532 144560
rect 120592 144520 150532 144548
rect 120592 144508 120598 144520
rect 150526 144508 150532 144520
rect 150584 144508 150590 144560
rect 158346 144508 158352 144560
rect 158404 144548 158410 144560
rect 190822 144548 190828 144560
rect 158404 144520 190828 144548
rect 158404 144508 158410 144520
rect 190822 144508 190828 144520
rect 190880 144508 190886 144560
rect 119430 144440 119436 144492
rect 119488 144480 119494 144492
rect 149422 144480 149428 144492
rect 119488 144452 149428 144480
rect 119488 144440 119494 144452
rect 149422 144440 149428 144452
rect 149480 144440 149486 144492
rect 157794 144440 157800 144492
rect 157852 144480 157858 144492
rect 191098 144480 191104 144492
rect 157852 144452 191104 144480
rect 157852 144440 157858 144452
rect 191098 144440 191104 144452
rect 191156 144440 191162 144492
rect 119246 144372 119252 144424
rect 119304 144412 119310 144424
rect 154022 144412 154028 144424
rect 119304 144384 154028 144412
rect 119304 144372 119310 144384
rect 154022 144372 154028 144384
rect 154080 144372 154086 144424
rect 156690 144372 156696 144424
rect 156748 144412 156754 144424
rect 190454 144412 190460 144424
rect 156748 144384 190460 144412
rect 156748 144372 156754 144384
rect 190454 144372 190460 144384
rect 190512 144372 190518 144424
rect 120626 144304 120632 144356
rect 120684 144344 120690 144356
rect 151262 144344 151268 144356
rect 120684 144316 151268 144344
rect 120684 144304 120690 144316
rect 151262 144304 151268 144316
rect 151320 144304 151326 144356
rect 153102 144304 153108 144356
rect 153160 144344 153166 144356
rect 186590 144344 186596 144356
rect 153160 144316 186596 144344
rect 153160 144304 153166 144316
rect 186590 144304 186596 144316
rect 186648 144304 186654 144356
rect 113726 144236 113732 144288
rect 113784 144276 113790 144288
rect 148042 144276 148048 144288
rect 113784 144248 148048 144276
rect 113784 144236 113790 144248
rect 148042 144236 148048 144248
rect 148100 144236 148106 144288
rect 159910 144236 159916 144288
rect 159968 144276 159974 144288
rect 193766 144276 193772 144288
rect 159968 144248 193772 144276
rect 159968 144236 159974 144248
rect 193766 144236 193772 144248
rect 193824 144236 193830 144288
rect 112438 144168 112444 144220
rect 112496 144208 112502 144220
rect 131482 144208 131488 144220
rect 112496 144180 131488 144208
rect 112496 144168 112502 144180
rect 131482 144168 131488 144180
rect 131540 144208 131546 144220
rect 188430 144208 188436 144220
rect 131540 144180 188436 144208
rect 131540 144168 131546 144180
rect 188430 144168 188436 144180
rect 188488 144168 188494 144220
rect 129550 143488 129556 143540
rect 129608 143528 129614 143540
rect 580258 143528 580264 143540
rect 129608 143500 580264 143528
rect 129608 143488 129614 143500
rect 580258 143488 580264 143500
rect 580316 143488 580322 143540
rect 177666 143420 177672 143472
rect 177724 143460 177730 143472
rect 179414 143460 179420 143472
rect 177724 143432 179420 143460
rect 177724 143420 177730 143432
rect 179414 143420 179420 143432
rect 179472 143420 179478 143472
rect 181530 143420 181536 143472
rect 181588 143460 181594 143472
rect 189626 143460 189632 143472
rect 181588 143432 189632 143460
rect 181588 143420 181594 143432
rect 189626 143420 189632 143432
rect 189684 143420 189690 143472
rect 117866 143352 117872 143404
rect 117924 143392 117930 143404
rect 130102 143392 130108 143404
rect 117924 143364 130108 143392
rect 117924 143352 117930 143364
rect 130102 143352 130108 143364
rect 130160 143352 130166 143404
rect 132034 143392 132040 143404
rect 131776 143364 132040 143392
rect 116762 143284 116768 143336
rect 116820 143324 116826 143336
rect 131776 143324 131804 143364
rect 132034 143352 132040 143364
rect 132092 143352 132098 143404
rect 176562 143352 176568 143404
rect 176620 143392 176626 143404
rect 178586 143392 178592 143404
rect 176620 143364 178592 143392
rect 176620 143352 176626 143364
rect 178586 143352 178592 143364
rect 178644 143352 178650 143404
rect 185578 143352 185584 143404
rect 185636 143392 185642 143404
rect 188338 143392 188344 143404
rect 185636 143364 188344 143392
rect 185636 143352 185642 143364
rect 188338 143352 188344 143364
rect 188396 143352 188402 143404
rect 116820 143296 131804 143324
rect 116820 143284 116826 143296
rect 131850 143284 131856 143336
rect 131908 143324 131914 143336
rect 138014 143324 138020 143336
rect 131908 143296 138020 143324
rect 131908 143284 131914 143296
rect 138014 143284 138020 143296
rect 138072 143284 138078 143336
rect 176010 143284 176016 143336
rect 176068 143324 176074 143336
rect 179782 143324 179788 143336
rect 176068 143296 179788 143324
rect 176068 143284 176074 143296
rect 179782 143284 179788 143296
rect 179840 143284 179846 143336
rect 184290 143284 184296 143336
rect 184348 143324 184354 143336
rect 195054 143324 195060 143336
rect 184348 143296 195060 143324
rect 184348 143284 184354 143296
rect 195054 143284 195060 143296
rect 195112 143284 195118 143336
rect 118050 143216 118056 143268
rect 118108 143256 118114 143268
rect 133414 143256 133420 143268
rect 118108 143228 133420 143256
rect 118108 143216 118114 143228
rect 133414 143216 133420 143228
rect 133472 143216 133478 143268
rect 184658 143216 184664 143268
rect 184716 143256 184722 143268
rect 196802 143256 196808 143268
rect 184716 143228 196808 143256
rect 184716 143216 184722 143228
rect 196802 143216 196808 143228
rect 196860 143216 196866 143268
rect 119798 143148 119804 143200
rect 119856 143188 119862 143200
rect 138382 143188 138388 143200
rect 119856 143160 138388 143188
rect 119856 143148 119862 143160
rect 138382 143148 138388 143160
rect 138440 143148 138446 143200
rect 175182 143148 175188 143200
rect 175240 143188 175246 143200
rect 189534 143188 189540 143200
rect 175240 143160 189540 143188
rect 175240 143148 175246 143160
rect 189534 143148 189540 143160
rect 189592 143148 189598 143200
rect 117038 143080 117044 143132
rect 117096 143120 117102 143132
rect 135254 143120 135260 143132
rect 117096 143092 135260 143120
rect 117096 143080 117102 143092
rect 135254 143080 135260 143092
rect 135312 143080 135318 143132
rect 168834 143080 168840 143132
rect 168892 143120 168898 143132
rect 189258 143120 189264 143132
rect 168892 143092 189264 143120
rect 168892 143080 168898 143092
rect 189258 143080 189264 143092
rect 189316 143080 189322 143132
rect 121086 143012 121092 143064
rect 121144 143052 121150 143064
rect 140038 143052 140044 143064
rect 121144 143024 140044 143052
rect 121144 143012 121150 143024
rect 140038 143012 140044 143024
rect 140096 143012 140102 143064
rect 166902 143012 166908 143064
rect 166960 143052 166966 143064
rect 186682 143052 186688 143064
rect 166960 143024 186688 143052
rect 166960 143012 166966 143024
rect 186682 143012 186688 143024
rect 186740 143012 186746 143064
rect 118142 142944 118148 142996
rect 118200 142984 118206 142996
rect 136726 142984 136732 142996
rect 118200 142956 136732 142984
rect 118200 142944 118206 142956
rect 136726 142944 136732 142956
rect 136784 142944 136790 142996
rect 165522 142944 165528 142996
rect 165580 142984 165586 142996
rect 187970 142984 187976 142996
rect 165580 142956 187976 142984
rect 165580 142944 165586 142956
rect 187970 142944 187976 142956
rect 188028 142944 188034 142996
rect 119614 142876 119620 142928
rect 119672 142916 119678 142928
rect 141694 142916 141700 142928
rect 119672 142888 141700 142916
rect 119672 142876 119678 142888
rect 141694 142876 141700 142888
rect 141752 142876 141758 142928
rect 160554 142876 160560 142928
rect 160612 142916 160618 142928
rect 186774 142916 186780 142928
rect 160612 142888 186780 142916
rect 160612 142876 160618 142888
rect 186774 142876 186780 142888
rect 186832 142876 186838 142928
rect 120994 142808 121000 142860
rect 121052 142848 121058 142860
rect 143534 142848 143540 142860
rect 121052 142820 143540 142848
rect 121052 142808 121058 142820
rect 143534 142808 143540 142820
rect 143592 142808 143598 142860
rect 155034 142808 155040 142860
rect 155092 142848 155098 142860
rect 157702 142848 157708 142860
rect 155092 142820 157708 142848
rect 155092 142808 155098 142820
rect 157702 142808 157708 142820
rect 157760 142808 157766 142860
rect 158622 142808 158628 142860
rect 158680 142848 158686 142860
rect 188062 142848 188068 142860
rect 158680 142820 188068 142848
rect 158680 142808 158686 142820
rect 188062 142808 188068 142820
rect 188120 142808 188126 142860
rect 132402 142740 132408 142792
rect 132460 142780 132466 142792
rect 136174 142780 136180 142792
rect 132460 142752 136180 142780
rect 132460 142740 132466 142752
rect 136174 142740 136180 142752
rect 136232 142740 136238 142792
rect 177114 142740 177120 142792
rect 177172 142780 177178 142792
rect 179506 142780 179512 142792
rect 177172 142752 179512 142780
rect 177172 142740 177178 142752
rect 179506 142740 179512 142752
rect 179564 142740 179570 142792
rect 119706 142672 119712 142724
rect 119764 142712 119770 142724
rect 127894 142712 127900 142724
rect 119764 142684 127900 142712
rect 119764 142672 119770 142684
rect 127894 142672 127900 142684
rect 127952 142672 127958 142724
rect 131022 142672 131028 142724
rect 131080 142712 131086 142724
rect 134518 142712 134524 142724
rect 131080 142684 134524 142712
rect 131080 142672 131086 142684
rect 134518 142672 134524 142684
rect 134576 142672 134582 142724
rect 179046 142672 179052 142724
rect 179104 142712 179110 142724
rect 179782 142712 179788 142724
rect 179104 142684 179788 142712
rect 179104 142672 179110 142684
rect 179782 142672 179788 142684
rect 179840 142672 179846 142724
rect 177942 142604 177948 142656
rect 178000 142644 178006 142656
rect 179322 142644 179328 142656
rect 178000 142616 179328 142644
rect 178000 142604 178006 142616
rect 179322 142604 179328 142616
rect 179380 142604 179386 142656
rect 130562 142468 130568 142520
rect 130620 142508 130626 142520
rect 132494 142508 132500 142520
rect 130620 142480 132500 142508
rect 130620 142468 130626 142480
rect 132494 142468 132500 142480
rect 132552 142468 132558 142520
rect 137986 142344 142154 142372
rect 3418 142264 3424 142316
rect 3476 142304 3482 142316
rect 137986 142304 138014 142344
rect 3476 142276 138014 142304
rect 142126 142304 142154 142344
rect 185578 142304 185584 142316
rect 142126 142276 185584 142304
rect 3476 142264 3482 142276
rect 185578 142264 185584 142276
rect 185636 142264 185642 142316
rect 125594 142196 125600 142248
rect 125652 142236 125658 142248
rect 126514 142236 126520 142248
rect 125652 142208 126520 142236
rect 125652 142196 125658 142208
rect 126514 142196 126520 142208
rect 126572 142236 126578 142248
rect 188154 142236 188160 142248
rect 126572 142208 188160 142236
rect 126572 142196 126578 142208
rect 188154 142196 188160 142208
rect 188212 142196 188218 142248
rect 116670 142128 116676 142180
rect 116728 142168 116734 142180
rect 124214 142168 124220 142180
rect 116728 142140 124220 142168
rect 116728 142128 116734 142140
rect 124214 142128 124220 142140
rect 124272 142128 124278 142180
rect 140774 142168 140780 142180
rect 139320 142140 140780 142168
rect 118326 142060 118332 142112
rect 118384 142100 118390 142112
rect 139320 142100 139348 142140
rect 140774 142128 140780 142140
rect 140832 142128 140838 142180
rect 155862 142128 155868 142180
rect 155920 142168 155926 142180
rect 157334 142168 157340 142180
rect 155920 142140 157340 142168
rect 155920 142128 155926 142140
rect 157334 142128 157340 142140
rect 157392 142128 157398 142180
rect 159450 142128 159456 142180
rect 159508 142168 159514 142180
rect 162486 142168 162492 142180
rect 159508 142140 162492 142168
rect 159508 142128 159514 142140
rect 162486 142128 162492 142140
rect 162544 142128 162550 142180
rect 118384 142072 139348 142100
rect 118384 142060 118390 142072
rect 184382 142060 184388 142112
rect 184440 142100 184446 142112
rect 193858 142100 193864 142112
rect 184440 142072 193864 142100
rect 184440 142060 184446 142072
rect 193858 142060 193864 142072
rect 193916 142060 193922 142112
rect 121178 141992 121184 142044
rect 121236 142032 121242 142044
rect 127066 142032 127072 142044
rect 121236 142004 127072 142032
rect 121236 141992 121242 142004
rect 127066 141992 127072 142004
rect 127124 141992 127130 142044
rect 182266 141992 182272 142044
rect 182324 142032 182330 142044
rect 192386 142032 192392 142044
rect 182324 142004 192392 142032
rect 182324 141992 182330 142004
rect 192386 141992 192392 142004
rect 192444 141992 192450 142044
rect 120810 141924 120816 141976
rect 120868 141964 120874 141976
rect 123754 141964 123760 141976
rect 120868 141936 123760 141964
rect 120868 141924 120874 141936
rect 123754 141924 123760 141936
rect 123812 141924 123818 141976
rect 183094 141924 183100 141976
rect 183152 141964 183158 141976
rect 194226 141964 194232 141976
rect 183152 141936 194232 141964
rect 183152 141924 183158 141936
rect 194226 141924 194232 141936
rect 194284 141924 194290 141976
rect 119522 141856 119528 141908
rect 119580 141896 119586 141908
rect 125134 141896 125140 141908
rect 119580 141868 125140 141896
rect 119580 141856 119586 141868
rect 125134 141856 125140 141868
rect 125192 141856 125198 141908
rect 184566 141856 184572 141908
rect 184624 141896 184630 141908
rect 195146 141896 195152 141908
rect 184624 141868 195152 141896
rect 184624 141856 184630 141868
rect 195146 141856 195152 141868
rect 195204 141856 195210 141908
rect 115290 141788 115296 141840
rect 115348 141828 115354 141840
rect 124582 141828 124588 141840
rect 115348 141800 124588 141828
rect 115348 141788 115354 141800
rect 124582 141788 124588 141800
rect 124640 141788 124646 141840
rect 180150 141788 180156 141840
rect 180208 141828 180214 141840
rect 192202 141828 192208 141840
rect 180208 141800 192208 141828
rect 180208 141788 180214 141800
rect 192202 141788 192208 141800
rect 192260 141788 192266 141840
rect 116946 141720 116952 141772
rect 117004 141760 117010 141772
rect 128998 141760 129004 141772
rect 117004 141732 129004 141760
rect 117004 141720 117010 141732
rect 128998 141720 129004 141732
rect 129056 141720 129062 141772
rect 184842 141720 184848 141772
rect 184900 141760 184906 141772
rect 196342 141760 196348 141772
rect 184900 141732 196348 141760
rect 184900 141720 184906 141732
rect 196342 141720 196348 141732
rect 196400 141720 196406 141772
rect 113910 141652 113916 141704
rect 113968 141692 113974 141704
rect 126974 141692 126980 141704
rect 113968 141664 126980 141692
rect 113968 141652 113974 141664
rect 126974 141652 126980 141664
rect 127032 141652 127038 141704
rect 172146 141652 172152 141704
rect 172204 141692 172210 141704
rect 187878 141692 187884 141704
rect 172204 141664 187884 141692
rect 172204 141652 172210 141664
rect 187878 141652 187884 141664
rect 187936 141652 187942 141704
rect 117130 141584 117136 141636
rect 117188 141624 117194 141636
rect 133966 141624 133972 141636
rect 117188 141596 133972 141624
rect 117188 141584 117194 141596
rect 133966 141584 133972 141596
rect 134024 141584 134030 141636
rect 170490 141584 170496 141636
rect 170548 141624 170554 141636
rect 189442 141624 189448 141636
rect 170548 141596 189448 141624
rect 170548 141584 170554 141596
rect 189442 141584 189448 141596
rect 189500 141584 189506 141636
rect 112254 141516 112260 141568
rect 112312 141556 112318 141568
rect 131666 141556 131672 141568
rect 112312 141528 131672 141556
rect 112312 141516 112318 141528
rect 131666 141516 131672 141528
rect 131724 141516 131730 141568
rect 174722 141516 174728 141568
rect 174780 141556 174786 141568
rect 197722 141556 197728 141568
rect 174780 141528 197728 141556
rect 174780 141516 174786 141528
rect 197722 141516 197728 141528
rect 197780 141516 197786 141568
rect 115382 141448 115388 141500
rect 115440 141488 115446 141500
rect 135622 141488 135628 141500
rect 115440 141460 135628 141488
rect 115440 141448 115446 141460
rect 135622 141448 135628 141460
rect 135680 141448 135686 141500
rect 169386 141448 169392 141500
rect 169444 141488 169450 141500
rect 193674 141488 193680 141500
rect 169444 141460 193680 141488
rect 169444 141448 169450 141460
rect 193674 141448 193680 141460
rect 193732 141448 193738 141500
rect 121178 141380 121184 141432
rect 121236 141420 121242 141432
rect 151906 141420 151912 141432
rect 121236 141392 151912 141420
rect 121236 141380 121242 141392
rect 151906 141380 151912 141392
rect 151964 141380 151970 141432
rect 160738 141380 160744 141432
rect 160796 141420 160802 141432
rect 189350 141420 189356 141432
rect 160796 141392 189356 141420
rect 160796 141380 160802 141392
rect 189350 141380 189356 141392
rect 189408 141380 189414 141432
rect 118694 141108 118700 141160
rect 118752 141148 118758 141160
rect 180150 141148 180156 141160
rect 118752 141120 180156 141148
rect 118752 141108 118758 141120
rect 180150 141108 180156 141120
rect 180208 141148 180214 141160
rect 180610 141148 180616 141160
rect 180208 141120 180616 141148
rect 180208 141108 180214 141120
rect 180610 141108 180616 141120
rect 180668 141108 180674 141160
rect 111058 141040 111064 141092
rect 111116 141080 111122 141092
rect 184842 141080 184848 141092
rect 111116 141052 184848 141080
rect 111116 141040 111122 141052
rect 184842 141040 184848 141052
rect 184900 141040 184906 141092
rect 8938 140972 8944 141024
rect 8996 141012 9002 141024
rect 182818 141012 182824 141024
rect 8996 140984 182824 141012
rect 8996 140972 9002 140984
rect 182818 140972 182824 140984
rect 182876 140972 182882 141024
rect 127066 140904 127072 140956
rect 127124 140944 127130 140956
rect 549898 140944 549904 140956
rect 127124 140916 549904 140944
rect 127124 140904 127130 140916
rect 549898 140904 549904 140916
rect 549956 140904 549962 140956
rect 128998 140836 129004 140888
rect 129056 140876 129062 140888
rect 580534 140876 580540 140888
rect 129056 140848 580540 140876
rect 129056 140836 129062 140848
rect 580534 140836 580540 140848
rect 580592 140836 580598 140888
rect 126974 140768 126980 140820
rect 127032 140808 127038 140820
rect 127618 140808 127624 140820
rect 127032 140780 127624 140808
rect 127032 140768 127038 140780
rect 127618 140768 127624 140780
rect 127676 140808 127682 140820
rect 580442 140808 580448 140820
rect 127676 140780 580448 140808
rect 127676 140768 127682 140780
rect 580442 140768 580448 140780
rect 580500 140768 580506 140820
rect 119798 140700 119804 140752
rect 119856 140740 119862 140752
rect 127802 140740 127808 140752
rect 119856 140712 127808 140740
rect 119856 140700 119862 140712
rect 127802 140700 127808 140712
rect 127860 140700 127866 140752
rect 169754 140700 169760 140752
rect 169812 140740 169818 140752
rect 193674 140740 193680 140752
rect 169812 140712 193680 140740
rect 169812 140700 169818 140712
rect 193674 140700 193680 140712
rect 193732 140700 193738 140752
rect 119522 140632 119528 140684
rect 119580 140672 119586 140684
rect 127526 140672 127532 140684
rect 119580 140644 127532 140672
rect 119580 140632 119586 140644
rect 127526 140632 127532 140644
rect 127584 140632 127590 140684
rect 178034 140632 178040 140684
rect 178092 140672 178098 140684
rect 178678 140672 178684 140684
rect 178092 140644 178684 140672
rect 178092 140632 178098 140644
rect 178678 140632 178684 140644
rect 178736 140632 178742 140684
rect 193214 140672 193220 140684
rect 180766 140644 193220 140672
rect 120810 140564 120816 140616
rect 120868 140604 120874 140616
rect 127710 140604 127716 140616
rect 120868 140576 127716 140604
rect 120868 140564 120874 140576
rect 127710 140564 127716 140576
rect 127768 140564 127774 140616
rect 172514 140564 172520 140616
rect 172572 140604 172578 140616
rect 180766 140604 180794 140644
rect 193214 140632 193220 140644
rect 193272 140632 193278 140684
rect 172572 140576 180794 140604
rect 172572 140564 172578 140576
rect 185670 140564 185676 140616
rect 185728 140604 185734 140616
rect 185728 140576 190454 140604
rect 185728 140564 185734 140576
rect 126238 140536 126244 140548
rect 125566 140508 126244 140536
rect 116670 140428 116676 140480
rect 116728 140468 116734 140480
rect 125566 140468 125594 140508
rect 126238 140496 126244 140508
rect 126296 140496 126302 140548
rect 181438 140496 181444 140548
rect 181496 140536 181502 140548
rect 181496 140508 189580 140536
rect 181496 140496 181502 140508
rect 116728 140440 125594 140468
rect 116728 140428 116734 140440
rect 116578 140360 116584 140412
rect 116636 140400 116642 140412
rect 126330 140400 126336 140412
rect 116636 140372 126336 140400
rect 116636 140360 116642 140372
rect 126330 140360 126336 140372
rect 126388 140360 126394 140412
rect 178770 140360 178776 140412
rect 178828 140400 178834 140412
rect 189350 140400 189356 140412
rect 178828 140372 189356 140400
rect 178828 140360 178834 140372
rect 189350 140360 189356 140372
rect 189408 140360 189414 140412
rect 189552 140400 189580 140508
rect 190426 140468 190454 140576
rect 195422 140468 195428 140480
rect 190426 140440 195428 140468
rect 195422 140428 195428 140440
rect 195480 140428 195486 140480
rect 189552 140372 190454 140400
rect 120902 140292 120908 140344
rect 120960 140332 120966 140344
rect 148134 140332 148140 140344
rect 120960 140304 148140 140332
rect 120960 140292 120966 140304
rect 148134 140292 148140 140304
rect 148192 140292 148198 140344
rect 185854 140292 185860 140344
rect 185912 140332 185918 140344
rect 189810 140332 189816 140344
rect 185912 140304 189816 140332
rect 185912 140292 185918 140304
rect 189810 140292 189816 140304
rect 189868 140292 189874 140344
rect 190426 140332 190454 140372
rect 192202 140332 192208 140344
rect 190426 140304 192208 140332
rect 192202 140292 192208 140304
rect 192260 140292 192266 140344
rect 119338 140224 119344 140276
rect 119396 140264 119402 140276
rect 146938 140264 146944 140276
rect 119396 140236 146944 140264
rect 119396 140224 119402 140236
rect 146938 140224 146944 140236
rect 146996 140224 147002 140276
rect 178862 140224 178868 140276
rect 178920 140264 178926 140276
rect 191282 140264 191288 140276
rect 178920 140236 191288 140264
rect 178920 140224 178926 140236
rect 191282 140224 191288 140236
rect 191340 140224 191346 140276
rect 117774 140156 117780 140208
rect 117832 140196 117838 140208
rect 146846 140196 146852 140208
rect 117832 140168 146852 140196
rect 117832 140156 117838 140168
rect 146846 140156 146852 140168
rect 146904 140156 146910 140208
rect 183094 140156 183100 140208
rect 183152 140196 183158 140208
rect 189902 140196 189908 140208
rect 183152 140168 189908 140196
rect 183152 140156 183158 140168
rect 189902 140156 189908 140168
rect 189960 140156 189966 140208
rect 116394 140088 116400 140140
rect 116452 140128 116458 140140
rect 146754 140128 146760 140140
rect 116452 140100 146760 140128
rect 116452 140088 116458 140100
rect 146754 140088 146760 140100
rect 146812 140088 146818 140140
rect 179230 140088 179236 140140
rect 179288 140128 179294 140140
rect 192662 140128 192668 140140
rect 179288 140100 192668 140128
rect 179288 140088 179294 140100
rect 192662 140088 192668 140100
rect 192720 140088 192726 140140
rect 116486 140020 116492 140072
rect 116544 140060 116550 140072
rect 148226 140060 148232 140072
rect 116544 140032 148232 140060
rect 116544 140020 116550 140032
rect 148226 140020 148232 140032
rect 148284 140020 148290 140072
rect 160094 140020 160100 140072
rect 160152 140060 160158 140072
rect 192570 140060 192576 140072
rect 160152 140032 192576 140060
rect 160152 140020 160158 140032
rect 192570 140020 192576 140032
rect 192628 140020 192634 140072
rect 119614 139952 119620 140004
rect 119672 139992 119678 140004
rect 123570 139992 123576 140004
rect 119672 139964 123576 139992
rect 119672 139952 119678 139964
rect 123570 139952 123576 139964
rect 123628 139952 123634 140004
rect 184198 139952 184204 140004
rect 184256 139992 184262 140004
rect 196710 139992 196716 140004
rect 184256 139964 196716 139992
rect 184256 139952 184262 139964
rect 196710 139952 196716 139964
rect 196768 139952 196774 140004
rect 168282 139816 168288 139868
rect 168340 139856 168346 139868
rect 178586 139856 178592 139868
rect 168340 139828 178592 139856
rect 168340 139816 168346 139828
rect 178586 139816 178592 139828
rect 178644 139816 178650 139868
rect 173250 139748 173256 139800
rect 173308 139788 173314 139800
rect 196250 139788 196256 139800
rect 173308 139760 196256 139788
rect 173308 139748 173314 139760
rect 196250 139748 196256 139760
rect 196308 139748 196314 139800
rect 120994 139680 121000 139732
rect 121052 139720 121058 139732
rect 125042 139720 125048 139732
rect 121052 139692 125048 139720
rect 121052 139680 121058 139692
rect 125042 139680 125048 139692
rect 125100 139680 125106 139732
rect 169754 139680 169760 139732
rect 169812 139720 169818 139732
rect 193582 139720 193588 139732
rect 169812 139692 193588 139720
rect 169812 139680 169818 139692
rect 193582 139680 193588 139692
rect 193640 139680 193646 139732
rect 118326 139612 118332 139664
rect 118384 139652 118390 139664
rect 123938 139652 123944 139664
rect 118384 139624 123944 139652
rect 118384 139612 118390 139624
rect 123938 139612 123944 139624
rect 123996 139612 124002 139664
rect 171594 139612 171600 139664
rect 171652 139652 171658 139664
rect 197630 139652 197636 139664
rect 171652 139624 197636 139652
rect 171652 139612 171658 139624
rect 197630 139612 197636 139624
rect 197688 139612 197694 139664
rect 126146 139544 126152 139596
rect 126204 139584 126210 139596
rect 179874 139584 179880 139596
rect 126204 139556 179880 139584
rect 126204 139544 126210 139556
rect 179874 139544 179880 139556
rect 179932 139544 179938 139596
rect 125042 139476 125048 139528
rect 125100 139516 125106 139528
rect 180426 139516 180432 139528
rect 125100 139488 180432 139516
rect 125100 139476 125106 139488
rect 180426 139476 180432 139488
rect 180484 139476 180490 139528
rect 113910 139408 113916 139460
rect 113968 139448 113974 139460
rect 122098 139448 122104 139460
rect 113968 139420 122104 139448
rect 113968 139408 113974 139420
rect 122098 139408 122104 139420
rect 122156 139408 122162 139460
rect 124030 139408 124036 139460
rect 124088 139448 124094 139460
rect 182082 139448 182088 139460
rect 124088 139420 182088 139448
rect 124088 139408 124094 139420
rect 182082 139408 182088 139420
rect 182140 139408 182146 139460
rect 121914 139340 121920 139392
rect 121972 139380 121978 139392
rect 123662 139380 123668 139392
rect 121972 139352 123668 139380
rect 121972 139340 121978 139352
rect 123662 139340 123668 139352
rect 123720 139340 123726 139392
rect 155126 139340 155132 139392
rect 155184 139380 155190 139392
rect 155494 139380 155500 139392
rect 155184 139352 155500 139380
rect 155184 139340 155190 139352
rect 155494 139340 155500 139352
rect 155552 139340 155558 139392
rect 185762 139340 185768 139392
rect 185820 139380 185826 139392
rect 186406 139380 186412 139392
rect 185820 139352 186412 139380
rect 185820 139340 185826 139352
rect 186406 139340 186412 139352
rect 186464 139340 186470 139392
rect 188154 138660 188160 138712
rect 188212 138700 188218 138712
rect 580258 138700 580264 138712
rect 188212 138672 580264 138700
rect 188212 138660 188218 138672
rect 580258 138660 580264 138672
rect 580316 138660 580322 138712
rect 3510 137912 3516 137964
rect 3568 137952 3574 137964
rect 118694 137952 118700 137964
rect 3568 137924 118700 137952
rect 3568 137912 3574 137924
rect 118694 137912 118700 137924
rect 118752 137912 118758 137964
rect 118050 136280 118056 136332
rect 118108 136320 118114 136332
rect 120810 136320 120816 136332
rect 118108 136292 120816 136320
rect 118108 136280 118114 136292
rect 120810 136280 120816 136292
rect 120868 136280 120874 136332
rect 3142 111732 3148 111784
rect 3200 111772 3206 111784
rect 31018 111772 31024 111784
rect 3200 111744 31024 111772
rect 3200 111732 3206 111744
rect 31018 111732 31024 111744
rect 31076 111732 31082 111784
rect 549898 86912 549904 86964
rect 549956 86952 549962 86964
rect 580166 86952 580172 86964
rect 549956 86924 580172 86952
rect 549956 86912 549962 86924
rect 580166 86912 580172 86924
rect 580224 86912 580230 86964
rect 188154 81240 188160 81252
rect 153166 81212 172514 81240
rect 108390 80928 108396 80980
rect 108448 80968 108454 80980
rect 123478 80968 123484 80980
rect 108448 80940 123484 80968
rect 108448 80928 108454 80940
rect 123478 80928 123484 80940
rect 123536 80928 123542 80980
rect 137986 80940 148594 80968
rect 120902 80860 120908 80912
rect 120960 80900 120966 80912
rect 137986 80900 138014 80940
rect 120960 80872 138014 80900
rect 120960 80860 120966 80872
rect 108206 80792 108212 80844
rect 108264 80832 108270 80844
rect 124030 80832 124036 80844
rect 108264 80804 124036 80832
rect 108264 80792 108270 80804
rect 124030 80792 124036 80804
rect 124088 80792 124094 80844
rect 116394 80724 116400 80776
rect 116452 80764 116458 80776
rect 116452 80736 133092 80764
rect 116452 80724 116458 80736
rect 71774 80656 71780 80708
rect 71832 80696 71838 80708
rect 108206 80696 108212 80708
rect 71832 80668 108212 80696
rect 71832 80656 71838 80668
rect 108206 80656 108212 80668
rect 108264 80656 108270 80708
rect 117682 80656 117688 80708
rect 117740 80696 117746 80708
rect 117740 80668 118694 80696
rect 117740 80656 117746 80668
rect 118666 80560 118694 80668
rect 123478 80656 123484 80708
rect 123536 80696 123542 80708
rect 129826 80696 129832 80708
rect 123536 80668 129832 80696
rect 123536 80656 123542 80668
rect 129826 80656 129832 80668
rect 129884 80656 129890 80708
rect 133064 80628 133092 80736
rect 133248 80736 136588 80764
rect 133248 80628 133276 80736
rect 133064 80600 133276 80628
rect 118666 80532 135254 80560
rect 135226 80424 135254 80532
rect 136560 80492 136588 80736
rect 142126 80668 145466 80696
rect 142126 80492 142154 80668
rect 136560 80464 142154 80492
rect 135226 80396 142154 80424
rect 118666 80328 140958 80356
rect 115014 80180 115020 80232
rect 115072 80220 115078 80232
rect 118666 80220 118694 80328
rect 115072 80192 118694 80220
rect 125566 80192 140222 80220
rect 115072 80180 115078 80192
rect 125566 80016 125594 80192
rect 132034 80112 132040 80164
rect 132092 80152 132098 80164
rect 132092 80124 132862 80152
rect 132092 80112 132098 80124
rect 129826 80044 129832 80096
rect 129884 80084 129890 80096
rect 130838 80084 130844 80096
rect 129884 80056 130844 80084
rect 129884 80044 129890 80056
rect 130838 80044 130844 80056
rect 130896 80044 130902 80096
rect 118666 79988 125594 80016
rect 106826 79840 106832 79892
rect 106884 79880 106890 79892
rect 118666 79880 118694 79988
rect 132834 79960 132862 80124
rect 133110 80056 138014 80084
rect 131942 79908 131948 79960
rect 132000 79948 132006 79960
rect 132724 79948 132730 79960
rect 132000 79920 132730 79948
rect 132000 79908 132006 79920
rect 132724 79908 132730 79920
rect 132782 79908 132788 79960
rect 132816 79908 132822 79960
rect 132874 79908 132880 79960
rect 133000 79908 133006 79960
rect 133058 79908 133064 79960
rect 106884 79852 118694 79880
rect 106884 79840 106890 79852
rect 124030 79840 124036 79892
rect 124088 79880 124094 79892
rect 124088 79852 129872 79880
rect 124088 79840 124094 79852
rect 114830 79772 114836 79824
rect 114888 79812 114894 79824
rect 129844 79812 129872 79852
rect 129918 79840 129924 79892
rect 129976 79880 129982 79892
rect 132908 79880 132914 79892
rect 129976 79852 132914 79880
rect 129976 79840 129982 79852
rect 132908 79840 132914 79852
rect 132966 79840 132972 79892
rect 114888 79784 125594 79812
rect 129844 79784 132724 79812
rect 114888 79772 114894 79784
rect 109678 79704 109684 79756
rect 109736 79744 109742 79756
rect 123478 79744 123484 79756
rect 109736 79716 123484 79744
rect 109736 79704 109742 79716
rect 123478 79704 123484 79716
rect 123536 79704 123542 79756
rect 125566 79744 125594 79784
rect 132310 79744 132316 79756
rect 125566 79716 132316 79744
rect 132310 79704 132316 79716
rect 132368 79704 132374 79756
rect 117866 79636 117872 79688
rect 117924 79676 117930 79688
rect 130746 79676 130752 79688
rect 117924 79648 130752 79676
rect 117924 79636 117930 79648
rect 130746 79636 130752 79648
rect 130804 79676 130810 79688
rect 132218 79676 132224 79688
rect 130804 79648 132224 79676
rect 130804 79636 130810 79648
rect 132218 79636 132224 79648
rect 132276 79636 132282 79688
rect 132696 79676 132724 79784
rect 132770 79704 132776 79756
rect 132828 79744 132834 79756
rect 133018 79744 133046 79908
rect 132828 79716 133046 79744
rect 132828 79704 132834 79716
rect 133110 79676 133138 80056
rect 133294 79988 133966 80016
rect 133294 79960 133322 79988
rect 133184 79908 133190 79960
rect 133242 79908 133248 79960
rect 133276 79908 133282 79960
rect 133334 79908 133340 79960
rect 133368 79908 133374 79960
rect 133426 79908 133432 79960
rect 133460 79908 133466 79960
rect 133518 79948 133524 79960
rect 133644 79948 133650 79960
rect 133518 79908 133552 79948
rect 133202 79880 133230 79908
rect 133202 79852 133276 79880
rect 133248 79688 133276 79852
rect 133386 79756 133414 79908
rect 133322 79704 133328 79756
rect 133380 79716 133414 79756
rect 133380 79704 133386 79716
rect 133524 79688 133552 79908
rect 133616 79908 133650 79948
rect 133702 79908 133708 79960
rect 133736 79908 133742 79960
rect 133794 79908 133800 79960
rect 133616 79688 133644 79908
rect 133754 79880 133782 79908
rect 133708 79852 133782 79880
rect 133708 79824 133736 79852
rect 133828 79840 133834 79892
rect 133886 79840 133892 79892
rect 133690 79772 133696 79824
rect 133748 79772 133754 79824
rect 133846 79812 133874 79840
rect 133800 79784 133874 79812
rect 133800 79756 133828 79784
rect 133782 79704 133788 79756
rect 133840 79704 133846 79756
rect 132696 79648 133138 79676
rect 133230 79636 133236 79688
rect 133288 79636 133294 79688
rect 133506 79636 133512 79688
rect 133564 79636 133570 79688
rect 133598 79636 133604 79688
rect 133656 79636 133662 79688
rect 110874 79568 110880 79620
rect 110932 79608 110938 79620
rect 121086 79608 121092 79620
rect 110932 79580 121092 79608
rect 110932 79568 110938 79580
rect 121086 79568 121092 79580
rect 121144 79568 121150 79620
rect 123018 79608 123024 79620
rect 121472 79580 123024 79608
rect 106734 79500 106740 79552
rect 106792 79540 106798 79552
rect 121472 79540 121500 79580
rect 123018 79568 123024 79580
rect 123076 79568 123082 79620
rect 129090 79568 129096 79620
rect 129148 79608 129154 79620
rect 133938 79608 133966 79988
rect 136054 79988 136910 80016
rect 134380 79908 134386 79960
rect 134438 79948 134444 79960
rect 134438 79908 134472 79948
rect 135392 79908 135398 79960
rect 135450 79908 135456 79960
rect 135852 79948 135858 79960
rect 135824 79908 135858 79948
rect 135910 79908 135916 79960
rect 134288 79840 134294 79892
rect 134346 79880 134352 79892
rect 134346 79840 134380 79880
rect 134104 79772 134110 79824
rect 134162 79772 134168 79824
rect 134122 79620 134150 79772
rect 134352 79756 134380 79840
rect 134444 79824 134472 79908
rect 134564 79840 134570 79892
rect 134622 79840 134628 79892
rect 135116 79880 135122 79892
rect 134812 79852 135122 79880
rect 134426 79772 134432 79824
rect 134484 79772 134490 79824
rect 134334 79704 134340 79756
rect 134392 79704 134398 79756
rect 129148 79580 133966 79608
rect 129148 79568 129154 79580
rect 134058 79568 134064 79620
rect 134116 79580 134150 79620
rect 134116 79568 134122 79580
rect 126974 79540 126980 79552
rect 106792 79512 121500 79540
rect 121564 79512 126980 79540
rect 106792 79500 106798 79512
rect 110966 79432 110972 79484
rect 111024 79472 111030 79484
rect 121564 79472 121592 79512
rect 126974 79500 126980 79512
rect 127032 79500 127038 79552
rect 131666 79540 131672 79552
rect 128326 79512 131672 79540
rect 128326 79472 128354 79512
rect 131666 79500 131672 79512
rect 131724 79500 131730 79552
rect 132402 79500 132408 79552
rect 132460 79540 132466 79552
rect 134582 79540 134610 79840
rect 134812 79552 134840 79852
rect 135116 79840 135122 79852
rect 135174 79840 135180 79892
rect 135208 79840 135214 79892
rect 135266 79840 135272 79892
rect 135300 79840 135306 79892
rect 135358 79840 135364 79892
rect 135024 79812 135030 79824
rect 134996 79772 135030 79812
rect 135082 79772 135088 79824
rect 134996 79552 135024 79772
rect 135226 79756 135254 79840
rect 135162 79704 135168 79756
rect 135220 79716 135254 79756
rect 135220 79704 135226 79716
rect 135070 79568 135076 79620
rect 135128 79608 135134 79620
rect 135318 79608 135346 79840
rect 135128 79580 135346 79608
rect 135128 79568 135134 79580
rect 132460 79512 134610 79540
rect 132460 79500 132466 79512
rect 134794 79500 134800 79552
rect 134852 79500 134858 79552
rect 134978 79500 134984 79552
rect 135036 79500 135042 79552
rect 135410 79540 135438 79908
rect 135668 79840 135674 79892
rect 135726 79840 135732 79892
rect 135686 79676 135714 79840
rect 135824 79824 135852 79908
rect 135944 79880 135950 79892
rect 135916 79840 135950 79880
rect 136002 79840 136008 79892
rect 135806 79772 135812 79824
rect 135864 79772 135870 79824
rect 135916 79756 135944 79840
rect 135898 79704 135904 79756
rect 135956 79704 135962 79756
rect 135640 79648 135714 79676
rect 135640 79620 135668 79648
rect 135622 79568 135628 79620
rect 135680 79568 135686 79620
rect 135714 79568 135720 79620
rect 135772 79608 135778 79620
rect 136054 79608 136082 79988
rect 136882 79960 136910 79988
rect 137434 79988 137876 80016
rect 137434 79960 137462 79988
rect 136772 79908 136778 79960
rect 136830 79908 136836 79960
rect 136864 79908 136870 79960
rect 136922 79908 136928 79960
rect 137232 79948 137238 79960
rect 136974 79920 137238 79948
rect 136312 79840 136318 79892
rect 136370 79840 136376 79892
rect 136790 79880 136818 79908
rect 136790 79852 136910 79880
rect 136330 79620 136358 79840
rect 136882 79688 136910 79852
rect 136974 79756 137002 79920
rect 137232 79908 137238 79920
rect 137290 79908 137296 79960
rect 137416 79908 137422 79960
rect 137474 79908 137480 79960
rect 137600 79908 137606 79960
rect 137658 79908 137664 79960
rect 137048 79840 137054 79892
rect 137106 79880 137112 79892
rect 137106 79852 137324 79880
rect 137106 79840 137112 79852
rect 137140 79772 137146 79824
rect 137198 79772 137204 79824
rect 136974 79716 137008 79756
rect 137002 79704 137008 79716
rect 137060 79704 137066 79756
rect 136882 79648 136916 79688
rect 136910 79636 136916 79648
rect 136968 79636 136974 79688
rect 135772 79580 136082 79608
rect 135772 79568 135778 79580
rect 136266 79568 136272 79620
rect 136324 79580 136358 79620
rect 136324 79568 136330 79580
rect 136174 79540 136180 79552
rect 135410 79512 136180 79540
rect 136174 79500 136180 79512
rect 136232 79500 136238 79552
rect 137158 79540 137186 79772
rect 137296 79620 137324 79852
rect 137618 79812 137646 79908
rect 137388 79784 137646 79812
rect 137388 79688 137416 79784
rect 137370 79636 137376 79688
rect 137428 79636 137434 79688
rect 137848 79620 137876 79988
rect 137986 79960 138014 80056
rect 140194 79960 140222 80192
rect 140930 79960 140958 80328
rect 142126 80288 142154 80396
rect 142126 80260 145052 80288
rect 137968 79908 137974 79960
rect 138026 79908 138032 79960
rect 138336 79908 138342 79960
rect 138394 79908 138400 79960
rect 138796 79908 138802 79960
rect 138854 79908 138860 79960
rect 138888 79908 138894 79960
rect 138946 79908 138952 79960
rect 139256 79908 139262 79960
rect 139314 79948 139320 79960
rect 139314 79920 139486 79948
rect 139314 79908 139320 79920
rect 138354 79880 138382 79908
rect 138032 79852 138382 79880
rect 138032 79688 138060 79852
rect 138428 79840 138434 79892
rect 138486 79840 138492 79892
rect 138152 79772 138158 79824
rect 138210 79772 138216 79824
rect 138014 79636 138020 79688
rect 138072 79636 138078 79688
rect 137278 79568 137284 79620
rect 137336 79568 137342 79620
rect 137830 79568 137836 79620
rect 137888 79568 137894 79620
rect 138170 79552 138198 79772
rect 138446 79688 138474 79840
rect 138382 79636 138388 79688
rect 138440 79648 138474 79688
rect 138440 79636 138446 79648
rect 138474 79568 138480 79620
rect 138532 79608 138538 79620
rect 138814 79608 138842 79908
rect 138906 79824 138934 79908
rect 139164 79840 139170 79892
rect 139222 79840 139228 79892
rect 139348 79840 139354 79892
rect 139406 79840 139412 79892
rect 138906 79784 138940 79824
rect 138934 79772 138940 79784
rect 138992 79772 138998 79824
rect 139182 79744 139210 79840
rect 138532 79580 138842 79608
rect 138952 79716 139210 79744
rect 138952 79608 138980 79716
rect 139026 79636 139032 79688
rect 139084 79676 139090 79688
rect 139366 79676 139394 79840
rect 139084 79648 139394 79676
rect 139084 79636 139090 79648
rect 139118 79608 139124 79620
rect 138952 79580 139124 79608
rect 138532 79568 138538 79580
rect 139118 79568 139124 79580
rect 139176 79568 139182 79620
rect 137554 79540 137560 79552
rect 137158 79512 137560 79540
rect 137554 79500 137560 79512
rect 137612 79500 137618 79552
rect 138170 79512 138204 79552
rect 138198 79500 138204 79512
rect 138256 79500 138262 79552
rect 139210 79500 139216 79552
rect 139268 79540 139274 79552
rect 139458 79540 139486 79920
rect 140176 79908 140182 79960
rect 140234 79908 140240 79960
rect 140728 79908 140734 79960
rect 140786 79908 140792 79960
rect 140820 79908 140826 79960
rect 140878 79908 140884 79960
rect 140912 79908 140918 79960
rect 140970 79908 140976 79960
rect 141832 79908 141838 79960
rect 141890 79908 141896 79960
rect 141924 79908 141930 79960
rect 141982 79908 141988 79960
rect 142108 79908 142114 79960
rect 142166 79908 142172 79960
rect 142292 79908 142298 79960
rect 142350 79908 142356 79960
rect 142384 79908 142390 79960
rect 142442 79908 142448 79960
rect 142752 79908 142758 79960
rect 142810 79908 142816 79960
rect 143488 79948 143494 79960
rect 143368 79920 143494 79948
rect 140452 79840 140458 79892
rect 140510 79840 140516 79892
rect 139808 79772 139814 79824
rect 139866 79772 139872 79824
rect 139826 79744 139854 79772
rect 139780 79716 139854 79744
rect 139780 79688 139808 79716
rect 139762 79636 139768 79688
rect 139820 79636 139826 79688
rect 139670 79568 139676 79620
rect 139728 79608 139734 79620
rect 140470 79608 140498 79840
rect 139728 79580 140498 79608
rect 139728 79568 139734 79580
rect 140590 79568 140596 79620
rect 140648 79608 140654 79620
rect 140746 79608 140774 79908
rect 140838 79688 140866 79908
rect 141188 79880 141194 79892
rect 140976 79852 141194 79880
rect 140976 79688 141004 79852
rect 141188 79840 141194 79852
rect 141246 79840 141252 79892
rect 141850 79824 141878 79908
rect 141942 79824 141970 79908
rect 142016 79840 142022 79892
rect 142074 79840 142080 79892
rect 141464 79812 141470 79824
rect 141160 79784 141470 79812
rect 140838 79648 140872 79688
rect 140866 79636 140872 79648
rect 140924 79636 140930 79688
rect 140958 79636 140964 79688
rect 141016 79636 141022 79688
rect 141160 79620 141188 79784
rect 141464 79772 141470 79784
rect 141522 79772 141528 79824
rect 141832 79772 141838 79824
rect 141890 79772 141896 79824
rect 141924 79772 141930 79824
rect 141982 79772 141988 79824
rect 142034 79744 142062 79840
rect 142126 79824 142154 79908
rect 142200 79840 142206 79892
rect 142258 79840 142264 79892
rect 142108 79772 142114 79824
rect 142166 79772 142172 79824
rect 141528 79716 142062 79744
rect 141528 79620 141556 79716
rect 142218 79688 142246 79840
rect 142310 79824 142338 79908
rect 142292 79772 142298 79824
rect 142350 79772 142356 79824
rect 142402 79688 142430 79908
rect 142660 79880 142666 79892
rect 142154 79636 142160 79688
rect 142212 79648 142246 79688
rect 142212 79636 142218 79648
rect 142338 79636 142344 79688
rect 142396 79648 142430 79688
rect 142540 79852 142666 79880
rect 142396 79636 142402 79648
rect 140648 79580 140774 79608
rect 140648 79568 140654 79580
rect 141142 79568 141148 79620
rect 141200 79568 141206 79620
rect 141510 79568 141516 79620
rect 141568 79568 141574 79620
rect 142540 79608 142568 79852
rect 142660 79840 142666 79852
rect 142718 79840 142724 79892
rect 142770 79812 142798 79908
rect 142936 79840 142942 79892
rect 142994 79840 143000 79892
rect 143120 79840 143126 79892
rect 143178 79880 143184 79892
rect 143178 79852 143304 79880
rect 143178 79840 143184 79852
rect 142632 79784 142798 79812
rect 142632 79688 142660 79784
rect 142954 79688 142982 79840
rect 142614 79636 142620 79688
rect 142672 79636 142678 79688
rect 142954 79648 142988 79688
rect 142982 79636 142988 79648
rect 143040 79636 143046 79688
rect 143276 79620 143304 79852
rect 142798 79608 142804 79620
rect 142540 79580 142804 79608
rect 142798 79568 142804 79580
rect 142856 79568 142862 79620
rect 143258 79568 143264 79620
rect 143316 79568 143322 79620
rect 139268 79512 139486 79540
rect 139268 79500 139274 79512
rect 139578 79500 139584 79552
rect 139636 79540 139642 79552
rect 143368 79540 143396 79920
rect 143488 79908 143494 79920
rect 143546 79908 143552 79960
rect 143580 79908 143586 79960
rect 143638 79908 143644 79960
rect 143764 79908 143770 79960
rect 143822 79908 143828 79960
rect 144316 79908 144322 79960
rect 144374 79908 144380 79960
rect 144592 79908 144598 79960
rect 144650 79908 144656 79960
rect 144684 79908 144690 79960
rect 144742 79908 144748 79960
rect 144776 79908 144782 79960
rect 144834 79908 144840 79960
rect 139636 79512 143396 79540
rect 143598 79552 143626 79908
rect 143782 79608 143810 79908
rect 144132 79880 144138 79892
rect 144104 79840 144138 79880
rect 144190 79840 144196 79892
rect 144104 79620 144132 79840
rect 144334 79620 144362 79908
rect 144610 79880 144638 79908
rect 143736 79580 143810 79608
rect 143736 79552 143764 79580
rect 144086 79568 144092 79620
rect 144144 79568 144150 79620
rect 144270 79568 144276 79620
rect 144328 79580 144362 79620
rect 144564 79852 144638 79880
rect 144564 79608 144592 79852
rect 144702 79812 144730 79908
rect 144656 79784 144730 79812
rect 144656 79676 144684 79784
rect 144794 79756 144822 79908
rect 144730 79704 144736 79756
rect 144788 79716 144822 79756
rect 144788 79704 144794 79716
rect 144822 79676 144828 79688
rect 144656 79648 144828 79676
rect 144822 79636 144828 79648
rect 144880 79636 144886 79688
rect 144638 79608 144644 79620
rect 144564 79580 144644 79608
rect 144328 79568 144334 79580
rect 144638 79568 144644 79580
rect 144696 79568 144702 79620
rect 143598 79512 143632 79552
rect 139636 79500 139642 79512
rect 143626 79500 143632 79512
rect 143684 79500 143690 79552
rect 143718 79500 143724 79552
rect 143776 79500 143782 79552
rect 143534 79472 143540 79484
rect 111024 79444 121592 79472
rect 121656 79444 128354 79472
rect 130396 79444 143540 79472
rect 111024 79432 111030 79444
rect 109954 79364 109960 79416
rect 110012 79404 110018 79416
rect 121656 79404 121684 79444
rect 110012 79376 121684 79404
rect 110012 79364 110018 79376
rect 123478 79364 123484 79416
rect 123536 79404 123542 79416
rect 130396 79404 130424 79444
rect 143534 79432 143540 79444
rect 143592 79432 143598 79484
rect 123536 79376 130424 79404
rect 123536 79364 123542 79376
rect 132310 79364 132316 79416
rect 132368 79404 132374 79416
rect 143902 79404 143908 79416
rect 132368 79376 143908 79404
rect 132368 79364 132374 79376
rect 143902 79364 143908 79376
rect 143960 79364 143966 79416
rect 145024 79404 145052 80260
rect 145438 80220 145466 80668
rect 145438 80192 146386 80220
rect 146358 79960 146386 80192
rect 146726 79988 147720 80016
rect 146726 79960 146754 79988
rect 145696 79908 145702 79960
rect 145754 79908 145760 79960
rect 146340 79908 146346 79960
rect 146398 79908 146404 79960
rect 146432 79908 146438 79960
rect 146490 79948 146496 79960
rect 146490 79908 146524 79948
rect 146708 79908 146714 79960
rect 146766 79908 146772 79960
rect 146800 79908 146806 79960
rect 146858 79948 146864 79960
rect 147168 79948 147174 79960
rect 146858 79908 146892 79948
rect 145144 79880 145150 79892
rect 145116 79840 145150 79880
rect 145202 79840 145208 79892
rect 145420 79840 145426 79892
rect 145478 79840 145484 79892
rect 145604 79880 145610 79892
rect 145576 79840 145610 79880
rect 145662 79840 145668 79892
rect 145116 79552 145144 79840
rect 145438 79676 145466 79840
rect 145300 79648 145466 79676
rect 145098 79500 145104 79552
rect 145156 79500 145162 79552
rect 145300 79472 145328 79648
rect 145576 79608 145604 79840
rect 145714 79812 145742 79908
rect 145788 79840 145794 79892
rect 145846 79840 145852 79892
rect 146156 79840 146162 79892
rect 146214 79840 146220 79892
rect 146248 79840 146254 79892
rect 146306 79840 146312 79892
rect 145668 79784 145742 79812
rect 145668 79688 145696 79784
rect 145806 79688 145834 79840
rect 145972 79772 145978 79824
rect 146030 79772 146036 79824
rect 145650 79636 145656 79688
rect 145708 79636 145714 79688
rect 145742 79636 145748 79688
rect 145800 79648 145834 79688
rect 145990 79688 146018 79772
rect 146174 79688 146202 79840
rect 145990 79648 146024 79688
rect 145800 79636 145806 79648
rect 146018 79636 146024 79648
rect 146076 79636 146082 79688
rect 146110 79636 146116 79688
rect 146168 79648 146202 79688
rect 146168 79636 146174 79648
rect 146266 79620 146294 79840
rect 146496 79620 146524 79908
rect 145392 79580 145604 79608
rect 145392 79552 145420 79580
rect 146202 79568 146208 79620
rect 146260 79580 146294 79620
rect 146260 79568 146266 79580
rect 146478 79568 146484 79620
rect 146536 79568 146542 79620
rect 145374 79500 145380 79552
rect 145432 79500 145438 79552
rect 146662 79500 146668 79552
rect 146720 79540 146726 79552
rect 146864 79540 146892 79908
rect 146956 79920 147174 79948
rect 146956 79552 146984 79920
rect 147168 79908 147174 79920
rect 147226 79908 147232 79960
rect 147260 79840 147266 79892
rect 147318 79840 147324 79892
rect 147536 79840 147542 79892
rect 147594 79880 147600 79892
rect 147594 79840 147628 79880
rect 147122 79568 147128 79620
rect 147180 79608 147186 79620
rect 147278 79608 147306 79840
rect 147490 79608 147496 79620
rect 147180 79580 147496 79608
rect 147180 79568 147186 79580
rect 147490 79568 147496 79580
rect 147548 79568 147554 79620
rect 146720 79512 146892 79540
rect 146720 79500 146726 79512
rect 146938 79500 146944 79552
rect 146996 79500 147002 79552
rect 147398 79500 147404 79552
rect 147456 79540 147462 79552
rect 147600 79540 147628 79840
rect 147456 79512 147628 79540
rect 147692 79540 147720 79988
rect 148566 79960 148594 80940
rect 153166 80084 153194 81212
rect 172486 81172 172514 81212
rect 179524 81212 188160 81240
rect 179524 81172 179552 81212
rect 188154 81200 188160 81212
rect 188212 81200 188218 81252
rect 172486 81144 179552 81172
rect 167840 80940 179276 80968
rect 167840 80492 167868 80940
rect 179248 80764 179276 80940
rect 186406 80860 186412 80912
rect 186464 80900 186470 80912
rect 199562 80900 199568 80912
rect 186464 80872 199568 80900
rect 186464 80860 186470 80872
rect 199562 80860 199568 80872
rect 199620 80860 199626 80912
rect 188154 80792 188160 80844
rect 188212 80832 188218 80844
rect 208578 80832 208584 80844
rect 188212 80804 208584 80832
rect 188212 80792 188218 80804
rect 208578 80792 208584 80804
rect 208636 80832 208642 80844
rect 234614 80832 234620 80844
rect 208636 80804 234620 80832
rect 208636 80792 208642 80804
rect 234614 80792 234620 80804
rect 234672 80792 234678 80844
rect 188246 80764 188252 80776
rect 179248 80736 188252 80764
rect 188246 80724 188252 80736
rect 188304 80764 188310 80776
rect 270494 80764 270500 80776
rect 188304 80736 270500 80764
rect 188304 80724 188310 80736
rect 270494 80724 270500 80736
rect 270552 80724 270558 80776
rect 177850 80656 177856 80708
rect 177908 80696 177914 80708
rect 183646 80696 183652 80708
rect 177908 80668 183652 80696
rect 177908 80656 177914 80668
rect 183646 80656 183652 80668
rect 183704 80656 183710 80708
rect 183830 80656 183836 80708
rect 183888 80696 183894 80708
rect 189718 80696 189724 80708
rect 183888 80668 189724 80696
rect 183888 80656 183894 80668
rect 189718 80656 189724 80668
rect 189776 80696 189782 80708
rect 288434 80696 288440 80708
rect 189776 80668 288440 80696
rect 189776 80656 189782 80668
rect 288434 80656 288440 80668
rect 288492 80656 288498 80708
rect 177758 80588 177764 80640
rect 177816 80628 177822 80640
rect 177816 80600 179414 80628
rect 177816 80588 177822 80600
rect 161492 80464 167868 80492
rect 179386 80492 179414 80600
rect 186406 80492 186412 80504
rect 179386 80464 186412 80492
rect 161492 80424 161520 80464
rect 186406 80452 186412 80464
rect 186464 80452 186470 80504
rect 194042 80424 194048 80436
rect 161216 80396 161520 80424
rect 161584 80396 194048 80424
rect 161216 80288 161244 80396
rect 161584 80288 161612 80396
rect 194042 80384 194048 80396
rect 194100 80384 194106 80436
rect 187142 80356 187148 80368
rect 160664 80260 161244 80288
rect 161308 80260 161612 80288
rect 164252 80328 187148 80356
rect 160664 80152 160692 80260
rect 150682 80056 153194 80084
rect 153442 80124 160692 80152
rect 150682 79960 150710 80056
rect 152338 79988 152918 80016
rect 148364 79908 148370 79960
rect 148422 79908 148428 79960
rect 148456 79908 148462 79960
rect 148514 79908 148520 79960
rect 148548 79908 148554 79960
rect 148606 79908 148612 79960
rect 150664 79908 150670 79960
rect 150722 79908 150728 79960
rect 150756 79908 150762 79960
rect 150814 79908 150820 79960
rect 151032 79908 151038 79960
rect 151090 79908 151096 79960
rect 151308 79908 151314 79960
rect 151366 79908 151372 79960
rect 151584 79908 151590 79960
rect 151642 79948 151648 79960
rect 151642 79920 151860 79948
rect 151642 79908 151648 79920
rect 147904 79840 147910 79892
rect 147962 79840 147968 79892
rect 148088 79840 148094 79892
rect 148146 79840 148152 79892
rect 147922 79688 147950 79840
rect 147922 79648 147956 79688
rect 147950 79636 147956 79648
rect 148008 79636 148014 79688
rect 148106 79608 148134 79840
rect 148382 79688 148410 79908
rect 148474 79744 148502 79908
rect 148916 79880 148922 79892
rect 148888 79840 148922 79880
rect 148974 79840 148980 79892
rect 149376 79880 149382 79892
rect 149348 79840 149382 79880
rect 149434 79840 149440 79892
rect 149468 79840 149474 79892
rect 149526 79840 149532 79892
rect 149560 79840 149566 79892
rect 149618 79840 149624 79892
rect 149836 79840 149842 79892
rect 149894 79840 149900 79892
rect 150112 79840 150118 79892
rect 150170 79880 150176 79892
rect 150170 79840 150204 79880
rect 150572 79840 150578 79892
rect 150630 79880 150636 79892
rect 150630 79840 150664 79880
rect 148474 79716 148824 79744
rect 148382 79648 148416 79688
rect 148410 79636 148416 79648
rect 148468 79636 148474 79688
rect 148796 79620 148824 79716
rect 148594 79608 148600 79620
rect 148106 79580 148600 79608
rect 148594 79568 148600 79580
rect 148652 79568 148658 79620
rect 148778 79568 148784 79620
rect 148836 79568 148842 79620
rect 148042 79540 148048 79552
rect 147692 79512 148048 79540
rect 147456 79500 147462 79512
rect 148042 79500 148048 79512
rect 148100 79500 148106 79552
rect 148134 79500 148140 79552
rect 148192 79540 148198 79552
rect 148888 79540 148916 79840
rect 149008 79772 149014 79824
rect 149066 79772 149072 79824
rect 149026 79688 149054 79772
rect 148962 79636 148968 79688
rect 149020 79648 149054 79688
rect 149020 79636 149026 79648
rect 148192 79512 148916 79540
rect 148192 79500 148198 79512
rect 145466 79472 145472 79484
rect 145300 79444 145472 79472
rect 145466 79432 145472 79444
rect 145524 79432 145530 79484
rect 145834 79432 145840 79484
rect 145892 79472 145898 79484
rect 149348 79472 149376 79840
rect 149486 79688 149514 79840
rect 149422 79636 149428 79688
rect 149480 79648 149514 79688
rect 149480 79636 149486 79648
rect 149578 79552 149606 79840
rect 149854 79552 149882 79840
rect 150176 79688 150204 79840
rect 150636 79756 150664 79840
rect 150774 79824 150802 79908
rect 150710 79772 150716 79824
rect 150768 79784 150802 79824
rect 151050 79824 151078 79908
rect 151050 79784 151084 79824
rect 150768 79772 150774 79784
rect 151078 79772 151084 79784
rect 151136 79772 151142 79824
rect 150618 79704 150624 79756
rect 150676 79704 150682 79756
rect 151326 79744 151354 79908
rect 151188 79716 151354 79744
rect 151188 79688 151216 79716
rect 150158 79636 150164 79688
rect 150216 79636 150222 79688
rect 151170 79636 151176 79688
rect 151228 79636 151234 79688
rect 151832 79620 151860 79920
rect 152136 79908 152142 79960
rect 152194 79908 152200 79960
rect 151952 79840 151958 79892
rect 152010 79880 152016 79892
rect 152010 79840 152044 79880
rect 152016 79688 152044 79840
rect 152154 79812 152182 79908
rect 152228 79840 152234 79892
rect 152286 79840 152292 79892
rect 152108 79784 152182 79812
rect 151998 79636 152004 79688
rect 152056 79636 152062 79688
rect 151814 79568 151820 79620
rect 151872 79568 151878 79620
rect 149578 79512 149612 79552
rect 149606 79500 149612 79512
rect 149664 79500 149670 79552
rect 149790 79500 149796 79552
rect 149848 79512 149882 79552
rect 150526 79540 150532 79552
rect 149946 79512 150532 79540
rect 149848 79500 149854 79512
rect 149422 79472 149428 79484
rect 145892 79444 149428 79472
rect 145892 79432 145898 79444
rect 149422 79432 149428 79444
rect 149480 79432 149486 79484
rect 149946 79404 149974 79512
rect 150526 79500 150532 79512
rect 150584 79500 150590 79552
rect 151538 79500 151544 79552
rect 151596 79540 151602 79552
rect 152108 79540 152136 79784
rect 152246 79756 152274 79840
rect 152182 79704 152188 79756
rect 152240 79716 152274 79756
rect 152240 79704 152246 79716
rect 151596 79512 152136 79540
rect 151596 79500 151602 79512
rect 145024 79376 149974 79404
rect 150268 79444 150480 79472
rect 109770 79296 109776 79348
rect 109828 79336 109834 79348
rect 132126 79336 132132 79348
rect 109828 79308 132132 79336
rect 109828 79296 109834 79308
rect 132126 79296 132132 79308
rect 132184 79296 132190 79348
rect 132218 79296 132224 79348
rect 132276 79336 132282 79348
rect 139578 79336 139584 79348
rect 132276 79308 139584 79336
rect 132276 79296 132282 79308
rect 139578 79296 139584 79308
rect 139636 79296 139642 79348
rect 139946 79296 139952 79348
rect 140004 79336 140010 79348
rect 140222 79336 140228 79348
rect 140004 79308 140228 79336
rect 140004 79296 140010 79308
rect 140222 79296 140228 79308
rect 140280 79296 140286 79348
rect 141234 79296 141240 79348
rect 141292 79336 141298 79348
rect 141418 79336 141424 79348
rect 141292 79308 141424 79336
rect 141292 79296 141298 79308
rect 141418 79296 141424 79308
rect 141476 79296 141482 79348
rect 143534 79296 143540 79348
rect 143592 79336 143598 79348
rect 144178 79336 144184 79348
rect 143592 79308 144184 79336
rect 143592 79296 143598 79308
rect 144178 79296 144184 79308
rect 144236 79296 144242 79348
rect 146202 79296 146208 79348
rect 146260 79336 146266 79348
rect 150268 79336 150296 79444
rect 150342 79364 150348 79416
rect 150400 79364 150406 79416
rect 146260 79308 150296 79336
rect 146260 79296 146266 79308
rect 119338 79228 119344 79280
rect 119396 79268 119402 79280
rect 147582 79268 147588 79280
rect 119396 79240 147588 79268
rect 119396 79228 119402 79240
rect 147582 79228 147588 79240
rect 147640 79268 147646 79280
rect 147858 79268 147864 79280
rect 147640 79240 147864 79268
rect 147640 79228 147646 79240
rect 147858 79228 147864 79240
rect 147916 79228 147922 79280
rect 149882 79228 149888 79280
rect 149940 79268 149946 79280
rect 150360 79268 150388 79364
rect 149940 79240 150388 79268
rect 150452 79268 150480 79444
rect 152090 79432 152096 79484
rect 152148 79472 152154 79484
rect 152338 79472 152366 79988
rect 152890 79960 152918 79988
rect 153442 79960 153470 80124
rect 161308 80084 161336 80260
rect 160756 80056 161336 80084
rect 153626 79988 154206 80016
rect 152412 79908 152418 79960
rect 152470 79908 152476 79960
rect 152688 79908 152694 79960
rect 152746 79908 152752 79960
rect 152780 79908 152786 79960
rect 152838 79908 152844 79960
rect 152872 79908 152878 79960
rect 152930 79908 152936 79960
rect 153240 79908 153246 79960
rect 153298 79908 153304 79960
rect 153424 79908 153430 79960
rect 153482 79908 153488 79960
rect 152430 79688 152458 79908
rect 152504 79772 152510 79824
rect 152562 79812 152568 79824
rect 152562 79772 152596 79812
rect 152430 79648 152464 79688
rect 152458 79636 152464 79648
rect 152516 79636 152522 79688
rect 152568 79540 152596 79772
rect 152706 79608 152734 79908
rect 152798 79688 152826 79908
rect 153148 79880 153154 79892
rect 152936 79852 153154 79880
rect 152936 79824 152964 79852
rect 153148 79840 153154 79852
rect 153206 79840 153212 79892
rect 152918 79772 152924 79824
rect 152976 79772 152982 79824
rect 153056 79772 153062 79824
rect 153114 79772 153120 79824
rect 153074 79688 153102 79772
rect 153258 79756 153286 79908
rect 153194 79704 153200 79756
rect 153252 79716 153286 79756
rect 153252 79704 153258 79716
rect 152798 79648 152832 79688
rect 152826 79636 152832 79648
rect 152884 79636 152890 79688
rect 153010 79636 153016 79688
rect 153068 79648 153102 79688
rect 153068 79636 153074 79648
rect 152706 79580 153516 79608
rect 152826 79540 152832 79552
rect 152568 79512 152832 79540
rect 152826 79500 152832 79512
rect 152884 79500 152890 79552
rect 152148 79444 152366 79472
rect 152148 79432 152154 79444
rect 153488 79268 153516 79580
rect 153626 79404 153654 79988
rect 154178 79960 154206 79988
rect 154822 79988 155218 80016
rect 154822 79960 154850 79988
rect 153792 79908 153798 79960
rect 153850 79908 153856 79960
rect 154068 79908 154074 79960
rect 154126 79908 154132 79960
rect 154160 79908 154166 79960
rect 154218 79908 154224 79960
rect 154436 79948 154442 79960
rect 154408 79908 154442 79948
rect 154494 79908 154500 79960
rect 154712 79908 154718 79960
rect 154770 79908 154776 79960
rect 154804 79908 154810 79960
rect 154862 79908 154868 79960
rect 154896 79908 154902 79960
rect 154954 79908 154960 79960
rect 153810 79880 153838 79908
rect 153810 79852 153884 79880
rect 153856 79688 153884 79852
rect 154086 79688 154114 79908
rect 154252 79840 154258 79892
rect 154310 79840 154316 79892
rect 154270 79688 154298 79840
rect 154408 79756 154436 79908
rect 154528 79840 154534 79892
rect 154586 79840 154592 79892
rect 154620 79840 154626 79892
rect 154678 79840 154684 79892
rect 154390 79704 154396 79756
rect 154448 79704 154454 79756
rect 154546 79688 154574 79840
rect 154638 79756 154666 79840
rect 154730 79824 154758 79908
rect 154730 79784 154764 79824
rect 154758 79772 154764 79784
rect 154816 79772 154822 79824
rect 154914 79756 154942 79908
rect 155080 79772 155086 79824
rect 155138 79772 155144 79824
rect 154638 79716 154672 79756
rect 154666 79704 154672 79716
rect 154724 79704 154730 79756
rect 154850 79704 154856 79756
rect 154908 79716 154942 79756
rect 154908 79704 154914 79716
rect 155098 79688 155126 79772
rect 153838 79636 153844 79688
rect 153896 79636 153902 79688
rect 153930 79636 153936 79688
rect 153988 79636 153994 79688
rect 154022 79636 154028 79688
rect 154080 79648 154114 79688
rect 154080 79636 154086 79648
rect 154206 79636 154212 79688
rect 154264 79648 154298 79688
rect 154264 79636 154270 79648
rect 154482 79636 154488 79688
rect 154540 79648 154574 79688
rect 154540 79636 154546 79648
rect 155034 79636 155040 79688
rect 155092 79648 155126 79688
rect 155092 79636 155098 79648
rect 153948 79608 153976 79636
rect 155190 79620 155218 79988
rect 157030 79988 158070 80016
rect 155264 79908 155270 79960
rect 155322 79908 155328 79960
rect 155448 79908 155454 79960
rect 155506 79908 155512 79960
rect 155540 79908 155546 79960
rect 155598 79908 155604 79960
rect 156184 79908 156190 79960
rect 156242 79908 156248 79960
rect 156368 79908 156374 79960
rect 156426 79908 156432 79960
rect 154942 79608 154948 79620
rect 153948 79580 154948 79608
rect 154942 79568 154948 79580
rect 155000 79568 155006 79620
rect 155126 79568 155132 79620
rect 155184 79580 155218 79620
rect 155184 79568 155190 79580
rect 155282 79472 155310 79908
rect 155466 79824 155494 79908
rect 155448 79772 155454 79824
rect 155506 79772 155512 79824
rect 155402 79568 155408 79620
rect 155460 79608 155466 79620
rect 155558 79608 155586 79908
rect 156000 79840 156006 79892
rect 156058 79840 156064 79892
rect 155460 79580 155586 79608
rect 156018 79620 156046 79840
rect 156018 79580 156052 79620
rect 155460 79568 155466 79580
rect 155558 79540 155586 79580
rect 156046 79568 156052 79580
rect 156104 79568 156110 79620
rect 155954 79540 155960 79552
rect 155558 79512 155960 79540
rect 155954 79500 155960 79512
rect 156012 79500 156018 79552
rect 156202 79540 156230 79908
rect 156386 79620 156414 79908
rect 156828 79772 156834 79824
rect 156886 79772 156892 79824
rect 156386 79580 156420 79620
rect 156414 79568 156420 79580
rect 156472 79568 156478 79620
rect 156690 79540 156696 79552
rect 156202 79512 156696 79540
rect 156690 79500 156696 79512
rect 156748 79500 156754 79552
rect 155678 79472 155684 79484
rect 155282 79444 155684 79472
rect 155678 79432 155684 79444
rect 155736 79432 155742 79484
rect 156846 79416 156874 79772
rect 157030 79620 157058 79988
rect 158042 79960 158070 79988
rect 159330 79988 159634 80016
rect 159330 79960 159358 79988
rect 157104 79908 157110 79960
rect 157162 79908 157168 79960
rect 157380 79908 157386 79960
rect 157438 79908 157444 79960
rect 157748 79908 157754 79960
rect 157806 79908 157812 79960
rect 158024 79908 158030 79960
rect 158082 79908 158088 79960
rect 158116 79908 158122 79960
rect 158174 79908 158180 79960
rect 158392 79908 158398 79960
rect 158450 79908 158456 79960
rect 158484 79908 158490 79960
rect 158542 79908 158548 79960
rect 158760 79908 158766 79960
rect 158818 79908 158824 79960
rect 159220 79908 159226 79960
rect 159278 79908 159284 79960
rect 159312 79908 159318 79960
rect 159370 79908 159376 79960
rect 159496 79908 159502 79960
rect 159554 79908 159560 79960
rect 157122 79688 157150 79908
rect 157196 79772 157202 79824
rect 157254 79812 157260 79824
rect 157254 79772 157288 79812
rect 157122 79648 157156 79688
rect 157150 79636 157156 79648
rect 157208 79636 157214 79688
rect 157260 79620 157288 79772
rect 157398 79620 157426 79908
rect 157766 79824 157794 79908
rect 158134 79824 158162 79908
rect 158410 79824 158438 79908
rect 157656 79772 157662 79824
rect 157714 79772 157720 79824
rect 157748 79772 157754 79824
rect 157806 79812 157812 79824
rect 157806 79784 157899 79812
rect 157806 79772 157812 79784
rect 158070 79772 158076 79824
rect 158128 79784 158162 79824
rect 158128 79772 158134 79784
rect 158392 79772 158398 79824
rect 158450 79772 158456 79824
rect 157030 79580 157064 79620
rect 157058 79568 157064 79580
rect 157116 79568 157122 79620
rect 157242 79568 157248 79620
rect 157300 79568 157306 79620
rect 157398 79580 157432 79620
rect 157426 79568 157432 79580
rect 157484 79568 157490 79620
rect 157674 79472 157702 79772
rect 157766 79552 157794 79772
rect 158502 79620 158530 79908
rect 158438 79568 158444 79620
rect 158496 79580 158530 79620
rect 158496 79568 158502 79580
rect 157766 79512 157800 79552
rect 157794 79500 157800 79512
rect 157852 79500 157858 79552
rect 158778 79540 158806 79908
rect 158944 79880 158950 79892
rect 158916 79840 158950 79880
rect 159002 79840 159008 79892
rect 159238 79880 159266 79908
rect 159100 79852 159266 79880
rect 158916 79756 158944 79840
rect 158898 79704 158904 79756
rect 158956 79704 158962 79756
rect 159100 79608 159128 79852
rect 159404 79840 159410 79892
rect 159462 79840 159468 79892
rect 159174 79772 159180 79824
rect 159232 79812 159238 79824
rect 159422 79812 159450 79840
rect 159232 79784 159450 79812
rect 159232 79772 159238 79784
rect 159514 79756 159542 79908
rect 159450 79704 159456 79756
rect 159508 79716 159542 79756
rect 159508 79704 159514 79716
rect 159358 79636 159364 79688
rect 159416 79676 159422 79688
rect 159606 79676 159634 79988
rect 159772 79908 159778 79960
rect 159830 79908 159836 79960
rect 160232 79908 160238 79960
rect 160290 79948 160296 79960
rect 160290 79908 160324 79948
rect 160416 79908 160422 79960
rect 160474 79908 160480 79960
rect 160600 79908 160606 79960
rect 160658 79908 160664 79960
rect 159790 79824 159818 79908
rect 159956 79880 159962 79892
rect 159726 79772 159732 79824
rect 159784 79784 159818 79824
rect 159928 79840 159962 79880
rect 160014 79840 160020 79892
rect 159784 79772 159790 79784
rect 159818 79704 159824 79756
rect 159876 79744 159882 79756
rect 159928 79744 159956 79840
rect 160296 79756 160324 79908
rect 159876 79716 159956 79744
rect 159876 79704 159882 79716
rect 160278 79704 160284 79756
rect 160336 79704 160342 79756
rect 159416 79648 159634 79676
rect 159416 79636 159422 79648
rect 160186 79636 160192 79688
rect 160244 79676 160250 79688
rect 160434 79676 160462 79908
rect 160618 79824 160646 79908
rect 160756 79892 160784 80056
rect 160876 79908 160882 79960
rect 160934 79908 160940 79960
rect 160968 79908 160974 79960
rect 161026 79908 161032 79960
rect 161060 79908 161066 79960
rect 161118 79908 161124 79960
rect 161152 79908 161158 79960
rect 161210 79908 161216 79960
rect 161428 79948 161434 79960
rect 161400 79908 161434 79948
rect 161486 79908 161492 79960
rect 161704 79908 161710 79960
rect 161762 79908 161768 79960
rect 161796 79908 161802 79960
rect 161854 79908 161860 79960
rect 162072 79948 162078 79960
rect 162044 79908 162078 79948
rect 162130 79908 162136 79960
rect 162256 79908 162262 79960
rect 162314 79908 162320 79960
rect 162624 79948 162630 79960
rect 162596 79908 162630 79948
rect 162682 79908 162688 79960
rect 162716 79908 162722 79960
rect 162774 79948 162780 79960
rect 162774 79908 162808 79948
rect 163176 79908 163182 79960
rect 163234 79908 163240 79960
rect 163360 79908 163366 79960
rect 163418 79908 163424 79960
rect 163544 79908 163550 79960
rect 163602 79908 163608 79960
rect 164096 79908 164102 79960
rect 164154 79908 164160 79960
rect 160692 79840 160698 79892
rect 160750 79840 160784 79892
rect 160600 79772 160606 79824
rect 160658 79772 160664 79824
rect 160244 79648 160462 79676
rect 160244 79636 160250 79648
rect 159266 79608 159272 79620
rect 159100 79580 159272 79608
rect 159266 79568 159272 79580
rect 159324 79568 159330 79620
rect 160554 79568 160560 79620
rect 160612 79608 160618 79620
rect 160756 79608 160784 79840
rect 160894 79824 160922 79908
rect 160876 79772 160882 79824
rect 160934 79772 160940 79824
rect 160986 79744 161014 79908
rect 160848 79716 161014 79744
rect 160848 79620 160876 79716
rect 161078 79676 161106 79908
rect 161170 79824 161198 79908
rect 161152 79772 161158 79824
rect 161210 79772 161216 79824
rect 161244 79772 161250 79824
rect 161302 79772 161308 79824
rect 161032 79648 161106 79676
rect 161262 79688 161290 79772
rect 161262 79648 161296 79688
rect 160612 79580 160784 79608
rect 160612 79568 160618 79580
rect 160830 79568 160836 79620
rect 160888 79568 160894 79620
rect 159542 79540 159548 79552
rect 158778 79512 159548 79540
rect 159542 79500 159548 79512
rect 159600 79500 159606 79552
rect 161032 79540 161060 79648
rect 161290 79636 161296 79648
rect 161348 79636 161354 79688
rect 161106 79568 161112 79620
rect 161164 79608 161170 79620
rect 161400 79608 161428 79908
rect 161722 79880 161750 79908
rect 161676 79852 161750 79880
rect 161676 79824 161704 79852
rect 161658 79772 161664 79824
rect 161716 79772 161722 79824
rect 161814 79756 161842 79908
rect 161888 79840 161894 79892
rect 161946 79840 161952 79892
rect 161750 79704 161756 79756
rect 161808 79716 161842 79756
rect 161808 79704 161814 79716
rect 161906 79620 161934 79840
rect 162044 79688 162072 79908
rect 162026 79636 162032 79688
rect 162084 79636 162090 79688
rect 161164 79580 161428 79608
rect 161164 79568 161170 79580
rect 161842 79568 161848 79620
rect 161900 79580 161934 79620
rect 161900 79568 161906 79580
rect 162274 79552 162302 79908
rect 162440 79812 162446 79824
rect 162412 79772 162446 79812
rect 162498 79772 162504 79824
rect 162412 79620 162440 79772
rect 162596 79620 162624 79908
rect 162670 79772 162676 79824
rect 162728 79772 162734 79824
rect 162394 79568 162400 79620
rect 162452 79568 162458 79620
rect 162578 79568 162584 79620
rect 162636 79568 162642 79620
rect 161198 79540 161204 79552
rect 161032 79512 161204 79540
rect 161198 79500 161204 79512
rect 161256 79500 161262 79552
rect 162274 79512 162308 79552
rect 162302 79500 162308 79512
rect 162360 79500 162366 79552
rect 162486 79500 162492 79552
rect 162544 79540 162550 79552
rect 162688 79540 162716 79772
rect 162544 79512 162716 79540
rect 162544 79500 162550 79512
rect 157978 79472 157984 79484
rect 157674 79444 157984 79472
rect 157978 79432 157984 79444
rect 158036 79432 158042 79484
rect 162780 79472 162808 79908
rect 163084 79880 163090 79892
rect 162872 79852 163090 79880
rect 162872 79688 162900 79852
rect 163084 79840 163090 79852
rect 163142 79840 163148 79892
rect 162992 79772 162998 79824
rect 163050 79772 163056 79824
rect 162854 79636 162860 79688
rect 162912 79636 162918 79688
rect 163010 79620 163038 79772
rect 163010 79580 163044 79620
rect 163038 79568 163044 79580
rect 163096 79568 163102 79620
rect 163194 79608 163222 79908
rect 163378 79824 163406 79908
rect 163314 79772 163320 79824
rect 163372 79784 163406 79824
rect 163562 79824 163590 79908
rect 163820 79880 163826 79892
rect 163792 79840 163826 79880
rect 163878 79840 163884 79892
rect 163562 79784 163596 79824
rect 163372 79772 163378 79784
rect 163590 79772 163596 79784
rect 163648 79772 163654 79824
rect 163792 79688 163820 79840
rect 163774 79636 163780 79688
rect 163832 79636 163838 79688
rect 163958 79608 163964 79620
rect 163194 79580 163964 79608
rect 163958 79568 163964 79580
rect 164016 79568 164022 79620
rect 162136 79444 162808 79472
rect 164114 79472 164142 79908
rect 164252 79688 164280 80328
rect 187142 80316 187148 80328
rect 187200 80356 187206 80368
rect 187200 80328 189074 80356
rect 187200 80316 187206 80328
rect 177758 80288 177764 80300
rect 166920 80260 177764 80288
rect 166920 80220 166948 80260
rect 177758 80248 177764 80260
rect 177816 80248 177822 80300
rect 178310 80220 178316 80232
rect 165126 80192 166948 80220
rect 167242 80192 178316 80220
rect 165126 79960 165154 80192
rect 167242 79960 167270 80192
rect 178310 80180 178316 80192
rect 178368 80180 178374 80232
rect 178126 80152 178132 80164
rect 173314 80124 178132 80152
rect 167978 80056 172284 80084
rect 167978 79960 168006 80056
rect 168070 79988 168696 80016
rect 168070 79960 168098 79988
rect 165108 79908 165114 79960
rect 165166 79908 165172 79960
rect 165200 79908 165206 79960
rect 165258 79948 165264 79960
rect 166304 79948 166310 79960
rect 165258 79908 165292 79948
rect 164464 79840 164470 79892
rect 164522 79840 164528 79892
rect 164556 79840 164562 79892
rect 164614 79880 164620 79892
rect 164614 79852 164740 79880
rect 164614 79840 164620 79852
rect 164482 79744 164510 79840
rect 164482 79716 164648 79744
rect 164620 79688 164648 79716
rect 164712 79688 164740 79852
rect 164832 79840 164838 79892
rect 164890 79880 164896 79892
rect 164890 79840 164924 79880
rect 165016 79840 165022 79892
rect 165074 79880 165080 79892
rect 165074 79852 165200 79880
rect 165074 79840 165080 79852
rect 164896 79688 164924 79840
rect 165172 79688 165200 79852
rect 164234 79636 164240 79688
rect 164292 79636 164298 79688
rect 164326 79636 164332 79688
rect 164384 79676 164390 79688
rect 164510 79676 164516 79688
rect 164384 79648 164516 79676
rect 164384 79636 164390 79648
rect 164510 79636 164516 79648
rect 164568 79636 164574 79688
rect 164602 79636 164608 79688
rect 164660 79636 164666 79688
rect 164694 79636 164700 79688
rect 164752 79636 164758 79688
rect 164878 79636 164884 79688
rect 164936 79636 164942 79688
rect 165154 79636 165160 79688
rect 165212 79636 165218 79688
rect 165062 79568 165068 79620
rect 165120 79608 165126 79620
rect 165264 79608 165292 79908
rect 165816 79920 166310 79948
rect 165384 79840 165390 79892
rect 165442 79840 165448 79892
rect 165120 79580 165292 79608
rect 165120 79568 165126 79580
rect 165402 79540 165430 79840
rect 165816 79688 165844 79920
rect 166304 79908 166310 79920
rect 166362 79908 166368 79960
rect 166672 79908 166678 79960
rect 166730 79908 166736 79960
rect 166764 79908 166770 79960
rect 166822 79908 166828 79960
rect 166948 79908 166954 79960
rect 167006 79908 167012 79960
rect 167132 79908 167138 79960
rect 167190 79908 167196 79960
rect 167224 79908 167230 79960
rect 167282 79908 167288 79960
rect 167316 79908 167322 79960
rect 167374 79908 167380 79960
rect 167592 79908 167598 79960
rect 167650 79908 167656 79960
rect 167684 79908 167690 79960
rect 167742 79908 167748 79960
rect 167960 79908 167966 79960
rect 168018 79908 168024 79960
rect 168052 79908 168058 79960
rect 168110 79908 168116 79960
rect 168144 79908 168150 79960
rect 168202 79948 168208 79960
rect 168512 79948 168518 79960
rect 168202 79920 168420 79948
rect 168202 79908 168208 79920
rect 166120 79880 166126 79892
rect 165908 79852 166126 79880
rect 165798 79636 165804 79688
rect 165856 79636 165862 79688
rect 165614 79568 165620 79620
rect 165672 79608 165678 79620
rect 165908 79608 165936 79852
rect 166120 79840 166126 79852
rect 166178 79840 166184 79892
rect 166028 79772 166034 79824
rect 166086 79772 166092 79824
rect 166212 79772 166218 79824
rect 166270 79772 166276 79824
rect 166488 79772 166494 79824
rect 166546 79772 166552 79824
rect 165672 79580 165936 79608
rect 165672 79568 165678 79580
rect 165890 79540 165896 79552
rect 165402 79512 165896 79540
rect 165890 79500 165896 79512
rect 165948 79500 165954 79552
rect 166046 79540 166074 79772
rect 166230 79620 166258 79772
rect 166506 79744 166534 79772
rect 166460 79716 166534 79744
rect 166460 79620 166488 79716
rect 166690 79688 166718 79908
rect 166626 79636 166632 79688
rect 166684 79648 166718 79688
rect 166782 79688 166810 79908
rect 166782 79648 166816 79688
rect 166684 79636 166690 79648
rect 166810 79636 166816 79648
rect 166868 79636 166874 79688
rect 166230 79580 166264 79620
rect 166258 79568 166264 79580
rect 166316 79568 166322 79620
rect 166442 79568 166448 79620
rect 166500 79568 166506 79620
rect 166810 79540 166816 79552
rect 166046 79512 166816 79540
rect 166810 79500 166816 79512
rect 166868 79500 166874 79552
rect 166442 79472 166448 79484
rect 164114 79444 166448 79472
rect 153838 79404 153844 79416
rect 153626 79376 153844 79404
rect 153838 79364 153844 79376
rect 153896 79404 153902 79416
rect 154390 79404 154396 79416
rect 153896 79376 154396 79404
rect 153896 79364 153902 79376
rect 154390 79364 154396 79376
rect 154448 79364 154454 79416
rect 155402 79364 155408 79416
rect 155460 79404 155466 79416
rect 155862 79404 155868 79416
rect 155460 79376 155868 79404
rect 155460 79364 155466 79376
rect 155862 79364 155868 79376
rect 155920 79364 155926 79416
rect 156846 79376 156880 79416
rect 156874 79364 156880 79376
rect 156932 79364 156938 79416
rect 157334 79364 157340 79416
rect 157392 79404 157398 79416
rect 157518 79404 157524 79416
rect 157392 79376 157524 79404
rect 157392 79364 157398 79376
rect 157518 79364 157524 79376
rect 157576 79364 157582 79416
rect 153654 79296 153660 79348
rect 153712 79336 153718 79348
rect 160278 79336 160284 79348
rect 153712 79308 160284 79336
rect 153712 79296 153718 79308
rect 160278 79296 160284 79308
rect 160336 79296 160342 79348
rect 162136 79280 162164 79444
rect 166442 79432 166448 79444
rect 166500 79432 166506 79484
rect 166966 79472 166994 79908
rect 167040 79840 167046 79892
rect 167098 79840 167104 79892
rect 167058 79540 167086 79840
rect 167150 79756 167178 79908
rect 167150 79716 167184 79756
rect 167178 79704 167184 79716
rect 167236 79704 167242 79756
rect 167334 79688 167362 79908
rect 167500 79840 167506 79892
rect 167558 79840 167564 79892
rect 167518 79744 167546 79840
rect 167472 79716 167546 79744
rect 167472 79688 167500 79716
rect 167610 79688 167638 79908
rect 167334 79648 167368 79688
rect 167362 79636 167368 79648
rect 167420 79636 167426 79688
rect 167454 79636 167460 79688
rect 167512 79636 167518 79688
rect 167546 79636 167552 79688
rect 167604 79648 167638 79688
rect 167604 79636 167610 79648
rect 167270 79568 167276 79620
rect 167328 79608 167334 79620
rect 167702 79608 167730 79908
rect 167978 79812 168006 79908
rect 168098 79812 168104 79824
rect 167978 79784 168104 79812
rect 168098 79772 168104 79784
rect 168156 79772 168162 79824
rect 167328 79580 167730 79608
rect 168392 79608 168420 79920
rect 168484 79908 168518 79948
rect 168570 79908 168576 79960
rect 168484 79824 168512 79908
rect 168466 79772 168472 79824
rect 168524 79772 168530 79824
rect 168558 79608 168564 79620
rect 168392 79580 168564 79608
rect 167328 79568 167334 79580
rect 168558 79568 168564 79580
rect 168616 79568 168622 79620
rect 168098 79540 168104 79552
rect 167058 79512 168104 79540
rect 168098 79500 168104 79512
rect 168156 79500 168162 79552
rect 167638 79472 167644 79484
rect 166966 79444 167644 79472
rect 167638 79432 167644 79444
rect 167696 79432 167702 79484
rect 167822 79432 167828 79484
rect 167880 79472 167886 79484
rect 168668 79472 168696 79988
rect 169082 79988 170076 80016
rect 169082 79960 169110 79988
rect 168788 79908 168794 79960
rect 168846 79908 168852 79960
rect 168972 79948 168978 79960
rect 168944 79908 168978 79948
rect 169030 79908 169036 79960
rect 169064 79908 169070 79960
rect 169122 79908 169128 79960
rect 169156 79908 169162 79960
rect 169214 79908 169220 79960
rect 169616 79908 169622 79960
rect 169674 79908 169680 79960
rect 167880 79444 168696 79472
rect 168806 79472 168834 79908
rect 168944 79688 168972 79908
rect 169174 79880 169202 79908
rect 169036 79852 169202 79880
rect 168926 79636 168932 79688
rect 168984 79636 168990 79688
rect 169036 79552 169064 79852
rect 169248 79840 169254 79892
rect 169306 79840 169312 79892
rect 169340 79840 169346 79892
rect 169398 79880 169404 79892
rect 169398 79852 169570 79880
rect 169398 79840 169404 79852
rect 169266 79620 169294 79840
rect 169432 79772 169438 79824
rect 169490 79772 169496 79824
rect 169450 79688 169478 79772
rect 169386 79636 169392 79688
rect 169444 79648 169478 79688
rect 169444 79636 169450 79648
rect 169542 79620 169570 79852
rect 169634 79756 169662 79908
rect 169892 79880 169898 79892
rect 169864 79840 169898 79880
rect 169950 79840 169956 79892
rect 169634 79716 169668 79756
rect 169662 79704 169668 79716
rect 169720 79704 169726 79756
rect 169864 79620 169892 79840
rect 170048 79620 170076 79988
rect 170260 79908 170266 79960
rect 170318 79908 170324 79960
rect 170812 79908 170818 79960
rect 170870 79908 170876 79960
rect 170996 79908 171002 79960
rect 171054 79948 171060 79960
rect 171054 79920 171180 79948
rect 171054 79908 171060 79920
rect 170278 79688 170306 79908
rect 170352 79840 170358 79892
rect 170410 79840 170416 79892
rect 170536 79840 170542 79892
rect 170594 79840 170600 79892
rect 170370 79756 170398 79840
rect 170370 79716 170404 79756
rect 170398 79704 170404 79716
rect 170456 79704 170462 79756
rect 170278 79648 170312 79688
rect 170306 79636 170312 79648
rect 170364 79636 170370 79688
rect 170554 79620 170582 79840
rect 170830 79824 170858 79908
rect 170766 79772 170772 79824
rect 170824 79784 170858 79824
rect 170824 79772 170830 79784
rect 170904 79772 170910 79824
rect 170962 79772 170968 79824
rect 170922 79744 170950 79772
rect 169202 79568 169208 79620
rect 169260 79580 169294 79620
rect 169260 79568 169266 79580
rect 169478 79568 169484 79620
rect 169536 79580 169570 79620
rect 169536 79568 169542 79580
rect 169846 79568 169852 79620
rect 169904 79568 169910 79620
rect 170030 79568 170036 79620
rect 170088 79568 170094 79620
rect 170490 79568 170496 79620
rect 170548 79580 170582 79620
rect 170784 79716 170950 79744
rect 170548 79568 170554 79580
rect 170784 79552 170812 79716
rect 171152 79620 171180 79920
rect 171272 79908 171278 79960
rect 171330 79908 171336 79960
rect 171640 79948 171646 79960
rect 171612 79908 171646 79948
rect 171698 79908 171704 79960
rect 171732 79908 171738 79960
rect 171790 79908 171796 79960
rect 171824 79908 171830 79960
rect 171882 79908 171888 79960
rect 171916 79908 171922 79960
rect 171974 79948 171980 79960
rect 172100 79948 172106 79960
rect 171974 79908 172008 79948
rect 171290 79812 171318 79908
rect 171456 79840 171462 79892
rect 171514 79880 171520 79892
rect 171514 79840 171548 79880
rect 171290 79784 171456 79812
rect 171428 79756 171456 79784
rect 171410 79704 171416 79756
rect 171468 79704 171474 79756
rect 171520 79688 171548 79840
rect 171502 79636 171508 79688
rect 171560 79636 171566 79688
rect 171134 79568 171140 79620
rect 171192 79568 171198 79620
rect 171612 79608 171640 79908
rect 171750 79824 171778 79908
rect 171842 79880 171870 79908
rect 171842 79852 171916 79880
rect 171686 79772 171692 79824
rect 171744 79784 171778 79824
rect 171744 79772 171750 79784
rect 171778 79704 171784 79756
rect 171836 79744 171842 79756
rect 171888 79744 171916 79852
rect 171980 79756 172008 79908
rect 172072 79908 172106 79948
rect 172158 79908 172164 79960
rect 172072 79756 172100 79908
rect 171836 79716 171916 79744
rect 171836 79704 171842 79716
rect 171778 79608 171784 79620
rect 171612 79580 171784 79608
rect 171778 79568 171784 79580
rect 171836 79568 171842 79620
rect 169018 79500 169024 79552
rect 169076 79500 169082 79552
rect 170766 79500 170772 79552
rect 170824 79500 170830 79552
rect 169294 79472 169300 79484
rect 168806 79444 169300 79472
rect 167880 79432 167886 79444
rect 169294 79432 169300 79444
rect 169352 79432 169358 79484
rect 171888 79472 171916 79716
rect 171962 79704 171968 79756
rect 172020 79704 172026 79756
rect 172054 79704 172060 79756
rect 172112 79704 172118 79756
rect 172256 79676 172284 80056
rect 173314 79960 173342 80124
rect 178126 80112 178132 80124
rect 178184 80112 178190 80164
rect 189046 80152 189074 80328
rect 252554 80152 252560 80164
rect 189046 80124 252560 80152
rect 252554 80112 252560 80124
rect 252612 80112 252618 80164
rect 177850 80084 177856 80096
rect 173590 80056 174630 80084
rect 173590 79960 173618 80056
rect 172376 79948 172382 79960
rect 172348 79908 172382 79948
rect 172434 79908 172440 79960
rect 172836 79948 172842 79960
rect 172808 79908 172842 79948
rect 172894 79908 172900 79960
rect 173020 79908 173026 79960
rect 173078 79908 173084 79960
rect 173112 79908 173118 79960
rect 173170 79948 173176 79960
rect 173170 79908 173204 79948
rect 173296 79908 173302 79960
rect 173354 79908 173360 79960
rect 173572 79908 173578 79960
rect 173630 79908 173636 79960
rect 173664 79908 173670 79960
rect 173722 79908 173728 79960
rect 173756 79908 173762 79960
rect 173814 79948 173820 79960
rect 173814 79908 173848 79948
rect 173940 79908 173946 79960
rect 173998 79948 174004 79960
rect 173998 79920 174216 79948
rect 173998 79908 174004 79920
rect 172348 79756 172376 79908
rect 172468 79840 172474 79892
rect 172526 79840 172532 79892
rect 172560 79840 172566 79892
rect 172618 79840 172624 79892
rect 172330 79704 172336 79756
rect 172388 79704 172394 79756
rect 172486 79744 172514 79840
rect 172578 79812 172606 79840
rect 172578 79784 172744 79812
rect 172486 79716 172560 79744
rect 172422 79676 172428 79688
rect 172256 79648 172428 79676
rect 172422 79636 172428 79648
rect 172480 79636 172486 79688
rect 172146 79568 172152 79620
rect 172204 79608 172210 79620
rect 172532 79608 172560 79716
rect 172204 79580 172560 79608
rect 172204 79568 172210 79580
rect 172716 79540 172744 79784
rect 172808 79620 172836 79908
rect 172928 79772 172934 79824
rect 172986 79772 172992 79824
rect 172946 79688 172974 79772
rect 172882 79636 172888 79688
rect 172940 79648 172974 79688
rect 172940 79636 172946 79648
rect 172790 79568 172796 79620
rect 172848 79568 172854 79620
rect 173038 79608 173066 79908
rect 173176 79688 173204 79908
rect 173682 79824 173710 79908
rect 173682 79784 173716 79824
rect 173710 79772 173716 79784
rect 173768 79772 173774 79824
rect 173158 79636 173164 79688
rect 173216 79636 173222 79688
rect 173250 79608 173256 79620
rect 173038 79580 173256 79608
rect 173250 79568 173256 79580
rect 173308 79568 173314 79620
rect 173820 79608 173848 79908
rect 174032 79880 174038 79892
rect 174004 79840 174038 79880
rect 174090 79840 174096 79892
rect 174004 79756 174032 79840
rect 173986 79704 173992 79756
rect 174044 79704 174050 79756
rect 173894 79636 173900 79688
rect 173952 79676 173958 79688
rect 173952 79648 174124 79676
rect 173952 79636 173958 79648
rect 173820 79580 174032 79608
rect 173342 79540 173348 79552
rect 172716 79512 173348 79540
rect 173342 79500 173348 79512
rect 173400 79500 173406 79552
rect 172882 79472 172888 79484
rect 171888 79444 172888 79472
rect 172882 79432 172888 79444
rect 172940 79432 172946 79484
rect 171594 79404 171600 79416
rect 162228 79376 171600 79404
rect 155862 79268 155868 79280
rect 150452 79240 153332 79268
rect 153488 79240 155868 79268
rect 149940 79228 149946 79240
rect 124122 79160 124128 79212
rect 124180 79200 124186 79212
rect 153304 79200 153332 79240
rect 155862 79228 155868 79240
rect 155920 79228 155926 79280
rect 162118 79228 162124 79280
rect 162176 79228 162182 79280
rect 162228 79200 162256 79376
rect 171594 79364 171600 79376
rect 171652 79364 171658 79416
rect 165154 79296 165160 79348
rect 165212 79336 165218 79348
rect 165522 79336 165528 79348
rect 165212 79308 165528 79336
rect 165212 79296 165218 79308
rect 165522 79296 165528 79308
rect 165580 79296 165586 79348
rect 173894 79336 173900 79348
rect 173268 79308 173900 79336
rect 173268 79268 173296 79308
rect 173894 79296 173900 79308
rect 173952 79296 173958 79348
rect 124180 79172 153240 79200
rect 153304 79172 162256 79200
rect 165540 79240 173296 79268
rect 124180 79160 124186 79172
rect 117958 79092 117964 79144
rect 118016 79132 118022 79144
rect 149054 79132 149060 79144
rect 118016 79104 149060 79132
rect 118016 79092 118022 79104
rect 149054 79092 149060 79104
rect 149112 79132 149118 79144
rect 149698 79132 149704 79144
rect 149112 79104 149704 79132
rect 149112 79092 149118 79104
rect 149698 79092 149704 79104
rect 149756 79092 149762 79144
rect 151078 79132 151084 79144
rect 150912 79104 151084 79132
rect 119062 79024 119068 79076
rect 119120 79064 119126 79076
rect 150912 79064 150940 79104
rect 151078 79092 151084 79104
rect 151136 79092 151142 79144
rect 153212 79132 153240 79172
rect 155770 79132 155776 79144
rect 153212 79104 155776 79132
rect 155770 79092 155776 79104
rect 155828 79092 155834 79144
rect 158806 79092 158812 79144
rect 158864 79132 158870 79144
rect 163498 79132 163504 79144
rect 158864 79104 163504 79132
rect 158864 79092 158870 79104
rect 163498 79092 163504 79104
rect 163556 79092 163562 79144
rect 119120 79036 150940 79064
rect 119120 79024 119126 79036
rect 150986 79024 150992 79076
rect 151044 79064 151050 79076
rect 165540 79064 165568 79240
rect 173434 79228 173440 79280
rect 173492 79268 173498 79280
rect 174004 79268 174032 79580
rect 174096 79404 174124 79648
rect 174188 79620 174216 79920
rect 174492 79908 174498 79960
rect 174550 79908 174556 79960
rect 174308 79840 174314 79892
rect 174366 79840 174372 79892
rect 174400 79840 174406 79892
rect 174458 79840 174464 79892
rect 174170 79568 174176 79620
rect 174228 79568 174234 79620
rect 174326 79608 174354 79840
rect 174418 79676 174446 79840
rect 174510 79824 174538 79908
rect 174492 79772 174498 79824
rect 174550 79772 174556 79824
rect 174602 79744 174630 80056
rect 175614 80056 177856 80084
rect 175614 80054 175642 80056
rect 175522 80026 175642 80054
rect 177850 80044 177856 80056
rect 177908 80044 177914 80096
rect 186498 80044 186504 80096
rect 186556 80084 186562 80096
rect 302234 80084 302240 80096
rect 186556 80056 302240 80084
rect 186556 80044 186562 80056
rect 302234 80044 302240 80056
rect 302292 80044 302298 80096
rect 175522 79960 175550 80026
rect 177942 80016 177948 80028
rect 175982 79988 177948 80016
rect 174676 79908 174682 79960
rect 174734 79948 174740 79960
rect 174734 79920 175136 79948
rect 174734 79908 174740 79920
rect 174952 79840 174958 79892
rect 175010 79840 175016 79892
rect 174970 79744 174998 79840
rect 175108 79812 175136 79920
rect 175504 79908 175510 79960
rect 175562 79908 175568 79960
rect 175688 79840 175694 79892
rect 175746 79840 175752 79892
rect 175872 79840 175878 79892
rect 175930 79880 175936 79892
rect 175982 79880 176010 79988
rect 177942 79976 177948 79988
rect 178000 79976 178006 80028
rect 178034 79976 178040 80028
rect 178092 80016 178098 80028
rect 178092 79988 179414 80016
rect 178092 79976 178098 79988
rect 176240 79908 176246 79960
rect 176298 79908 176304 79960
rect 176332 79908 176338 79960
rect 176390 79948 176396 79960
rect 178678 79948 178684 79960
rect 176390 79920 178684 79948
rect 176390 79908 176396 79920
rect 178678 79908 178684 79920
rect 178736 79908 178742 79960
rect 175930 79852 176010 79880
rect 175930 79840 175936 79852
rect 175458 79812 175464 79824
rect 175108 79784 175464 79812
rect 175458 79772 175464 79784
rect 175516 79772 175522 79824
rect 175706 79812 175734 79840
rect 176258 79824 176286 79908
rect 177068 79840 177074 79892
rect 177126 79880 177132 79892
rect 177758 79880 177764 79892
rect 177126 79852 177764 79880
rect 177126 79840 177132 79852
rect 177758 79840 177764 79852
rect 177816 79840 177822 79892
rect 175706 79784 175964 79812
rect 176258 79784 176292 79824
rect 175936 79756 175964 79784
rect 176286 79772 176292 79784
rect 176344 79772 176350 79824
rect 176516 79772 176522 79824
rect 176574 79772 176580 79824
rect 177252 79772 177258 79824
rect 177310 79812 177316 79824
rect 177850 79812 177856 79824
rect 177310 79784 177856 79812
rect 177310 79772 177316 79784
rect 177850 79772 177856 79784
rect 177908 79772 177914 79824
rect 179386 79812 179414 79988
rect 199470 79812 199476 79824
rect 179386 79784 199476 79812
rect 199470 79772 199476 79784
rect 199528 79772 199534 79824
rect 174602 79716 174906 79744
rect 174970 79716 175320 79744
rect 174538 79676 174544 79688
rect 174418 79648 174544 79676
rect 174538 79636 174544 79648
rect 174596 79636 174602 79688
rect 174446 79608 174452 79620
rect 174326 79580 174452 79608
rect 174446 79568 174452 79580
rect 174504 79568 174510 79620
rect 174878 79540 174906 79716
rect 175292 79620 175320 79716
rect 175918 79704 175924 79756
rect 175976 79704 175982 79756
rect 176534 79688 176562 79772
rect 197998 79744 198004 79756
rect 176470 79636 176476 79688
rect 176528 79648 176562 79688
rect 176626 79716 198004 79744
rect 176528 79636 176534 79648
rect 175274 79568 175280 79620
rect 175332 79568 175338 79620
rect 175642 79568 175648 79620
rect 175700 79608 175706 79620
rect 176626 79608 176654 79716
rect 197998 79704 198004 79716
rect 198056 79704 198062 79756
rect 175700 79580 176654 79608
rect 175700 79568 175706 79580
rect 178126 79568 178132 79620
rect 178184 79608 178190 79620
rect 197630 79608 197636 79620
rect 178184 79580 197636 79608
rect 178184 79568 178190 79580
rect 197630 79568 197636 79580
rect 197688 79568 197694 79620
rect 174878 79512 175136 79540
rect 174722 79432 174728 79484
rect 174780 79472 174786 79484
rect 174998 79472 175004 79484
rect 174780 79444 175004 79472
rect 174780 79432 174786 79444
rect 174998 79432 175004 79444
rect 175056 79432 175062 79484
rect 175108 79472 175136 79512
rect 178310 79500 178316 79552
rect 178368 79540 178374 79552
rect 193950 79540 193956 79552
rect 178368 79512 193956 79540
rect 178368 79500 178374 79512
rect 193950 79500 193956 79512
rect 194008 79540 194014 79552
rect 194502 79540 194508 79552
rect 194008 79512 194508 79540
rect 194008 79500 194014 79512
rect 194502 79500 194508 79512
rect 194560 79500 194566 79552
rect 176930 79472 176936 79484
rect 175108 79444 176936 79472
rect 176930 79432 176936 79444
rect 176988 79432 176994 79484
rect 178218 79472 178224 79484
rect 177040 79444 178224 79472
rect 177040 79404 177068 79444
rect 178218 79432 178224 79444
rect 178276 79472 178282 79484
rect 238754 79472 238760 79484
rect 178276 79444 238760 79472
rect 178276 79432 178282 79444
rect 238754 79432 238760 79444
rect 238812 79432 238818 79484
rect 174096 79376 177068 79404
rect 177390 79364 177396 79416
rect 177448 79404 177454 79416
rect 189902 79404 189908 79416
rect 177448 79376 189908 79404
rect 177448 79364 177454 79376
rect 189902 79364 189908 79376
rect 189960 79364 189966 79416
rect 175182 79296 175188 79348
rect 175240 79336 175246 79348
rect 178034 79336 178040 79348
rect 175240 79308 178040 79336
rect 175240 79296 175246 79308
rect 178034 79296 178040 79308
rect 178092 79296 178098 79348
rect 181898 79296 181904 79348
rect 181956 79336 181962 79348
rect 191282 79336 191288 79348
rect 181956 79308 191288 79336
rect 181956 79296 181962 79308
rect 191282 79296 191288 79308
rect 191340 79296 191346 79348
rect 194502 79296 194508 79348
rect 194560 79336 194566 79348
rect 448514 79336 448520 79348
rect 194560 79308 448520 79336
rect 194560 79296 194566 79308
rect 448514 79296 448520 79308
rect 448572 79296 448578 79348
rect 173492 79240 174032 79268
rect 173492 79228 173498 79240
rect 175826 79228 175832 79280
rect 175884 79268 175890 79280
rect 202322 79268 202328 79280
rect 175884 79240 202328 79268
rect 175884 79228 175890 79240
rect 202322 79228 202328 79240
rect 202380 79228 202386 79280
rect 173526 79160 173532 79212
rect 173584 79200 173590 79212
rect 203702 79200 203708 79212
rect 173584 79172 203708 79200
rect 173584 79160 173590 79172
rect 203702 79160 203708 79172
rect 203760 79160 203766 79212
rect 166166 79092 166172 79144
rect 166224 79132 166230 79144
rect 178402 79132 178408 79144
rect 166224 79104 178408 79132
rect 166224 79092 166230 79104
rect 178402 79092 178408 79104
rect 178460 79132 178466 79144
rect 178460 79104 179414 79132
rect 178460 79092 178466 79104
rect 151044 79036 165568 79064
rect 151044 79024 151050 79036
rect 171134 79024 171140 79076
rect 171192 79064 171198 79076
rect 173250 79064 173256 79076
rect 171192 79036 173256 79064
rect 171192 79024 171198 79036
rect 173250 79024 173256 79036
rect 173308 79024 173314 79076
rect 174538 79024 174544 79076
rect 174596 79064 174602 79076
rect 174814 79064 174820 79076
rect 174596 79036 174820 79064
rect 174596 79024 174602 79036
rect 174814 79024 174820 79036
rect 174872 79064 174878 79076
rect 175826 79064 175832 79076
rect 174872 79036 175832 79064
rect 174872 79024 174878 79036
rect 175826 79024 175832 79036
rect 175884 79024 175890 79076
rect 176746 79024 176752 79076
rect 176804 79064 176810 79076
rect 177206 79064 177212 79076
rect 176804 79036 177212 79064
rect 176804 79024 176810 79036
rect 177206 79024 177212 79036
rect 177264 79024 177270 79076
rect 179386 79064 179414 79104
rect 180150 79092 180156 79144
rect 180208 79132 180214 79144
rect 183738 79132 183744 79144
rect 180208 79104 183744 79132
rect 180208 79092 180214 79104
rect 183738 79092 183744 79104
rect 183796 79132 183802 79144
rect 285674 79132 285680 79144
rect 183796 79104 285680 79132
rect 183796 79092 183802 79104
rect 285674 79092 285680 79104
rect 285732 79092 285738 79144
rect 376754 79064 376760 79076
rect 179386 79036 376760 79064
rect 376754 79024 376760 79036
rect 376812 79024 376818 79076
rect 119246 78956 119252 79008
rect 119304 78996 119310 79008
rect 151538 78996 151544 79008
rect 119304 78968 151544 78996
rect 119304 78956 119310 78968
rect 151538 78956 151544 78968
rect 151596 78996 151602 79008
rect 153102 78996 153108 79008
rect 151596 78968 153108 78996
rect 151596 78956 151602 78968
rect 153102 78956 153108 78968
rect 153160 78956 153166 79008
rect 154666 78956 154672 79008
rect 154724 78996 154730 79008
rect 180150 78996 180156 79008
rect 154724 78968 180156 78996
rect 154724 78956 154730 78968
rect 180150 78956 180156 78968
rect 180208 78956 180214 79008
rect 198090 78956 198096 79008
rect 198148 78996 198154 79008
rect 483014 78996 483020 79008
rect 198148 78968 483020 78996
rect 198148 78956 198154 78968
rect 483014 78956 483020 78968
rect 483072 78956 483078 79008
rect 116486 78888 116492 78940
rect 116544 78928 116550 78940
rect 148134 78928 148140 78940
rect 116544 78900 148140 78928
rect 116544 78888 116550 78900
rect 148134 78888 148140 78900
rect 148192 78888 148198 78940
rect 157306 78900 167086 78928
rect 121086 78820 121092 78872
rect 121144 78860 121150 78872
rect 125594 78860 125600 78872
rect 121144 78832 125600 78860
rect 121144 78820 121150 78832
rect 125594 78820 125600 78832
rect 125652 78820 125658 78872
rect 129550 78820 129556 78872
rect 129608 78860 129614 78872
rect 142154 78860 142160 78872
rect 129608 78832 142160 78860
rect 129608 78820 129614 78832
rect 142154 78820 142160 78832
rect 142212 78820 142218 78872
rect 147950 78820 147956 78872
rect 148008 78860 148014 78872
rect 157306 78860 157334 78900
rect 148008 78832 157334 78860
rect 148008 78820 148014 78832
rect 161658 78820 161664 78872
rect 161716 78860 161722 78872
rect 166166 78860 166172 78872
rect 161716 78832 166172 78860
rect 161716 78820 161722 78832
rect 166166 78820 166172 78832
rect 166224 78820 166230 78872
rect 167058 78860 167086 78900
rect 171594 78888 171600 78940
rect 171652 78928 171658 78940
rect 178034 78928 178040 78940
rect 171652 78900 178040 78928
rect 171652 78888 171658 78900
rect 178034 78888 178040 78900
rect 178092 78928 178098 78940
rect 179322 78928 179328 78940
rect 178092 78900 179328 78928
rect 178092 78888 178098 78900
rect 179322 78888 179328 78900
rect 179380 78888 179386 78940
rect 195238 78888 195244 78940
rect 195296 78928 195302 78940
rect 500954 78928 500960 78940
rect 195296 78900 500960 78928
rect 195296 78888 195302 78900
rect 500954 78888 500960 78900
rect 501012 78888 501018 78940
rect 179966 78860 179972 78872
rect 167058 78832 179972 78860
rect 179966 78820 179972 78832
rect 180024 78820 180030 78872
rect 197998 78820 198004 78872
rect 198056 78860 198062 78872
rect 523126 78860 523132 78872
rect 198056 78832 523132 78860
rect 198056 78820 198062 78832
rect 523126 78820 523132 78832
rect 523184 78820 523190 78872
rect 130654 78752 130660 78804
rect 130712 78792 130718 78804
rect 144914 78792 144920 78804
rect 130712 78764 144920 78792
rect 130712 78752 130718 78764
rect 144914 78752 144920 78764
rect 144972 78752 144978 78804
rect 166258 78752 166264 78804
rect 166316 78792 166322 78804
rect 166994 78792 167000 78804
rect 166316 78764 167000 78792
rect 166316 78752 166322 78764
rect 166994 78752 167000 78764
rect 167052 78752 167058 78804
rect 176194 78752 176200 78804
rect 176252 78792 176258 78804
rect 178678 78792 178684 78804
rect 176252 78764 178684 78792
rect 176252 78752 176258 78764
rect 178678 78752 178684 78764
rect 178736 78752 178742 78804
rect 197630 78752 197636 78804
rect 197688 78792 197694 78804
rect 525794 78792 525800 78804
rect 197688 78764 525800 78792
rect 197688 78752 197694 78764
rect 525794 78752 525800 78764
rect 525852 78752 525858 78804
rect 142062 78724 142068 78736
rect 132374 78696 142068 78724
rect 132374 78668 132402 78696
rect 142062 78684 142068 78696
rect 142120 78684 142126 78736
rect 149514 78684 149520 78736
rect 149572 78724 149578 78736
rect 150158 78724 150164 78736
rect 149572 78696 150164 78724
rect 149572 78684 149578 78696
rect 150158 78684 150164 78696
rect 150216 78684 150222 78736
rect 160186 78684 160192 78736
rect 160244 78724 160250 78736
rect 195422 78724 195428 78736
rect 160244 78696 195428 78724
rect 160244 78684 160250 78696
rect 195422 78684 195428 78696
rect 195480 78684 195486 78736
rect 200758 78684 200764 78736
rect 200816 78724 200822 78736
rect 201402 78724 201408 78736
rect 200816 78696 201408 78724
rect 200816 78684 200822 78696
rect 201402 78684 201408 78696
rect 201460 78724 201466 78736
rect 536834 78724 536840 78736
rect 201460 78696 536840 78724
rect 201460 78684 201466 78696
rect 536834 78684 536840 78696
rect 536892 78684 536898 78736
rect 132310 78616 132316 78668
rect 132368 78628 132402 78668
rect 132368 78616 132374 78628
rect 135254 78616 135260 78668
rect 135312 78656 135318 78668
rect 135898 78656 135904 78668
rect 135312 78628 135904 78656
rect 135312 78616 135318 78628
rect 135898 78616 135904 78628
rect 135956 78616 135962 78668
rect 136726 78616 136732 78668
rect 136784 78656 136790 78668
rect 136910 78656 136916 78668
rect 136784 78628 136916 78656
rect 136784 78616 136790 78628
rect 136910 78616 136916 78628
rect 136968 78616 136974 78668
rect 137094 78616 137100 78668
rect 137152 78656 137158 78668
rect 137738 78656 137744 78668
rect 137152 78628 137744 78656
rect 137152 78616 137158 78628
rect 137738 78616 137744 78628
rect 137796 78616 137802 78668
rect 141234 78616 141240 78668
rect 141292 78656 141298 78668
rect 141510 78656 141516 78668
rect 141292 78628 141516 78656
rect 141292 78616 141298 78628
rect 141510 78616 141516 78628
rect 141568 78616 141574 78668
rect 142430 78656 142436 78668
rect 141620 78628 142436 78656
rect 102134 78548 102140 78600
rect 102192 78588 102198 78600
rect 102870 78588 102876 78600
rect 102192 78560 102876 78588
rect 102192 78548 102198 78560
rect 102870 78548 102876 78560
rect 102928 78588 102934 78600
rect 133874 78588 133880 78600
rect 102928 78560 133880 78588
rect 102928 78548 102934 78560
rect 133874 78548 133880 78560
rect 133932 78548 133938 78600
rect 137278 78548 137284 78600
rect 137336 78588 137342 78600
rect 137830 78588 137836 78600
rect 137336 78560 137836 78588
rect 137336 78548 137342 78560
rect 137830 78548 137836 78560
rect 137888 78588 137894 78600
rect 141620 78588 141648 78628
rect 142430 78616 142436 78628
rect 142488 78616 142494 78668
rect 143902 78616 143908 78668
rect 143960 78656 143966 78668
rect 150066 78656 150072 78668
rect 143960 78628 150072 78656
rect 143960 78616 143966 78628
rect 150066 78616 150072 78628
rect 150124 78616 150130 78668
rect 157978 78616 157984 78668
rect 158036 78656 158042 78668
rect 158438 78656 158444 78668
rect 158036 78628 158444 78656
rect 158036 78616 158042 78628
rect 158438 78616 158444 78628
rect 158496 78616 158502 78668
rect 162026 78616 162032 78668
rect 162084 78656 162090 78668
rect 162394 78656 162400 78668
rect 162084 78628 162400 78656
rect 162084 78616 162090 78628
rect 162394 78616 162400 78628
rect 162452 78616 162458 78668
rect 175182 78656 175188 78668
rect 167196 78628 175188 78656
rect 137888 78560 141648 78588
rect 137888 78548 137894 78560
rect 141970 78548 141976 78600
rect 142028 78588 142034 78600
rect 142706 78588 142712 78600
rect 142028 78560 142712 78588
rect 142028 78548 142034 78560
rect 142706 78548 142712 78560
rect 142764 78548 142770 78600
rect 162946 78548 162952 78600
rect 163004 78588 163010 78600
rect 163222 78588 163228 78600
rect 163004 78560 163228 78588
rect 163004 78548 163010 78560
rect 163222 78548 163228 78560
rect 163280 78548 163286 78600
rect 164418 78548 164424 78600
rect 164476 78588 164482 78600
rect 165522 78588 165528 78600
rect 164476 78560 165528 78588
rect 164476 78548 164482 78560
rect 165522 78548 165528 78560
rect 165580 78548 165586 78600
rect 75914 78480 75920 78532
rect 75972 78520 75978 78532
rect 106826 78520 106832 78532
rect 75972 78492 106832 78520
rect 75972 78480 75978 78492
rect 106826 78480 106832 78492
rect 106884 78520 106890 78532
rect 107194 78520 107200 78532
rect 106884 78492 107200 78520
rect 106884 78480 106890 78492
rect 107194 78480 107200 78492
rect 107252 78480 107258 78532
rect 137370 78480 137376 78532
rect 137428 78520 137434 78532
rect 137738 78520 137744 78532
rect 137428 78492 137744 78520
rect 137428 78480 137434 78492
rect 137738 78480 137744 78492
rect 137796 78480 137802 78532
rect 141510 78480 141516 78532
rect 141568 78520 141574 78532
rect 141694 78520 141700 78532
rect 141568 78492 141700 78520
rect 141568 78480 141574 78492
rect 141694 78480 141700 78492
rect 141752 78480 141758 78532
rect 157610 78480 157616 78532
rect 157668 78520 157674 78532
rect 161658 78520 161664 78532
rect 157668 78492 161664 78520
rect 157668 78480 157674 78492
rect 161658 78480 161664 78492
rect 161716 78480 161722 78532
rect 164234 78480 164240 78532
rect 164292 78520 164298 78532
rect 164878 78520 164884 78532
rect 164292 78492 164884 78520
rect 164292 78480 164298 78492
rect 164878 78480 164884 78492
rect 164936 78520 164942 78532
rect 167196 78520 167224 78628
rect 175182 78616 175188 78628
rect 175240 78616 175246 78668
rect 177022 78616 177028 78668
rect 177080 78656 177086 78668
rect 206278 78656 206284 78668
rect 177080 78628 206284 78656
rect 177080 78616 177086 78628
rect 206278 78616 206284 78628
rect 206336 78616 206342 78668
rect 174078 78548 174084 78600
rect 174136 78588 174142 78600
rect 178954 78588 178960 78600
rect 174136 78560 178960 78588
rect 174136 78548 174142 78560
rect 178954 78548 178960 78560
rect 179012 78548 179018 78600
rect 179322 78548 179328 78600
rect 179380 78588 179386 78600
rect 206462 78588 206468 78600
rect 179380 78560 206468 78588
rect 179380 78548 179386 78560
rect 206462 78548 206468 78560
rect 206520 78548 206526 78600
rect 164936 78492 167224 78520
rect 164936 78480 164942 78492
rect 168466 78480 168472 78532
rect 168524 78520 168530 78532
rect 193582 78520 193588 78532
rect 168524 78492 193588 78520
rect 168524 78480 168530 78492
rect 193582 78480 193588 78492
rect 193640 78520 193646 78532
rect 194502 78520 194508 78532
rect 193640 78492 194508 78520
rect 193640 78480 193646 78492
rect 194502 78480 194508 78492
rect 194560 78480 194566 78532
rect 107102 78452 107108 78464
rect 103486 78424 107108 78452
rect 60734 78276 60740 78328
rect 60792 78316 60798 78328
rect 103486 78316 103514 78424
rect 107102 78412 107108 78424
rect 107160 78452 107166 78464
rect 137186 78452 137192 78464
rect 107160 78424 137192 78452
rect 107160 78412 107166 78424
rect 137186 78412 137192 78424
rect 137244 78412 137250 78464
rect 144178 78412 144184 78464
rect 144236 78452 144242 78464
rect 152366 78452 152372 78464
rect 144236 78424 152372 78452
rect 144236 78412 144242 78424
rect 152366 78412 152372 78424
rect 152424 78412 152430 78464
rect 166258 78412 166264 78464
rect 166316 78452 166322 78464
rect 167638 78452 167644 78464
rect 166316 78424 167644 78452
rect 166316 78412 166322 78424
rect 167638 78412 167644 78424
rect 167696 78452 167702 78464
rect 177390 78452 177396 78464
rect 167696 78424 177396 78452
rect 167696 78412 167702 78424
rect 177390 78412 177396 78424
rect 177448 78412 177454 78464
rect 179966 78412 179972 78464
rect 180024 78452 180030 78464
rect 183462 78452 183468 78464
rect 180024 78424 183468 78452
rect 180024 78412 180030 78424
rect 183462 78412 183468 78424
rect 183520 78452 183526 78464
rect 206186 78452 206192 78464
rect 183520 78424 206192 78452
rect 183520 78412 183526 78424
rect 206186 78412 206192 78424
rect 206244 78412 206250 78464
rect 107010 78344 107016 78396
rect 107068 78384 107074 78396
rect 107194 78384 107200 78396
rect 107068 78356 107200 78384
rect 107068 78344 107074 78356
rect 107194 78344 107200 78356
rect 107252 78384 107258 78396
rect 135990 78384 135996 78396
rect 107252 78356 135996 78384
rect 107252 78344 107258 78356
rect 135990 78344 135996 78356
rect 136048 78344 136054 78396
rect 137554 78344 137560 78396
rect 137612 78384 137618 78396
rect 142614 78384 142620 78396
rect 137612 78356 142620 78384
rect 137612 78344 137618 78356
rect 142614 78344 142620 78356
rect 142672 78344 142678 78396
rect 148134 78344 148140 78396
rect 148192 78384 148198 78396
rect 148870 78384 148876 78396
rect 148192 78356 148876 78384
rect 148192 78344 148198 78356
rect 148870 78344 148876 78356
rect 148928 78344 148934 78396
rect 157426 78344 157432 78396
rect 157484 78384 157490 78396
rect 157702 78384 157708 78396
rect 157484 78356 157708 78384
rect 157484 78344 157490 78356
rect 157702 78344 157708 78356
rect 157760 78344 157766 78396
rect 163958 78344 163964 78396
rect 164016 78384 164022 78396
rect 166166 78384 166172 78396
rect 164016 78356 166172 78384
rect 164016 78344 164022 78356
rect 166166 78344 166172 78356
rect 166224 78344 166230 78396
rect 168282 78344 168288 78396
rect 168340 78384 168346 78396
rect 202230 78384 202236 78396
rect 168340 78356 202236 78384
rect 168340 78344 168346 78356
rect 202230 78344 202236 78356
rect 202288 78344 202294 78396
rect 135714 78316 135720 78328
rect 60792 78288 103514 78316
rect 113146 78288 135720 78316
rect 60792 78276 60798 78288
rect 57974 78208 57980 78260
rect 58032 78248 58038 78260
rect 108482 78248 108488 78260
rect 58032 78220 108488 78248
rect 58032 78208 58038 78220
rect 108482 78208 108488 78220
rect 108540 78248 108546 78260
rect 113146 78248 113174 78288
rect 135714 78276 135720 78288
rect 135772 78276 135778 78328
rect 138106 78276 138112 78328
rect 138164 78316 138170 78328
rect 138750 78316 138756 78328
rect 138164 78288 138756 78316
rect 138164 78276 138170 78288
rect 138750 78276 138756 78288
rect 138808 78276 138814 78328
rect 140130 78276 140136 78328
rect 140188 78316 140194 78328
rect 140498 78316 140504 78328
rect 140188 78288 140504 78316
rect 140188 78276 140194 78288
rect 140498 78276 140504 78288
rect 140556 78276 140562 78328
rect 146570 78276 146576 78328
rect 146628 78316 146634 78328
rect 171870 78316 171876 78328
rect 146628 78288 171876 78316
rect 146628 78276 146634 78288
rect 171870 78276 171876 78288
rect 171928 78276 171934 78328
rect 183002 78276 183008 78328
rect 183060 78316 183066 78328
rect 204806 78316 204812 78328
rect 183060 78288 204812 78316
rect 183060 78276 183066 78288
rect 204806 78276 204812 78288
rect 204864 78276 204870 78328
rect 108540 78220 113174 78248
rect 108540 78208 108546 78220
rect 122466 78208 122472 78260
rect 122524 78248 122530 78260
rect 148318 78248 148324 78260
rect 122524 78220 148324 78248
rect 122524 78208 122530 78220
rect 148318 78208 148324 78220
rect 148376 78208 148382 78260
rect 149330 78208 149336 78260
rect 149388 78248 149394 78260
rect 183554 78248 183560 78260
rect 149388 78220 183560 78248
rect 149388 78208 149394 78220
rect 183554 78208 183560 78220
rect 183612 78208 183618 78260
rect 46934 78140 46940 78192
rect 46992 78180 46998 78192
rect 107194 78180 107200 78192
rect 46992 78152 107200 78180
rect 46992 78140 46998 78152
rect 107194 78140 107200 78152
rect 107252 78140 107258 78192
rect 130930 78180 130936 78192
rect 113146 78152 130936 78180
rect 34514 78072 34520 78124
rect 34572 78112 34578 78124
rect 100754 78112 100760 78124
rect 34572 78084 100760 78112
rect 34572 78072 34578 78084
rect 100754 78072 100760 78084
rect 100812 78072 100818 78124
rect 108574 78112 108580 78124
rect 103486 78084 108580 78112
rect 20714 78004 20720 78056
rect 20772 78044 20778 78056
rect 102134 78044 102140 78056
rect 20772 78016 102140 78044
rect 20772 78004 20778 78016
rect 102134 78004 102140 78016
rect 102192 78004 102198 78056
rect 2774 77936 2780 77988
rect 2832 77976 2838 77988
rect 103486 77976 103514 78084
rect 108574 78072 108580 78084
rect 108632 78112 108638 78124
rect 113146 78112 113174 78152
rect 130930 78140 130936 78152
rect 130988 78140 130994 78192
rect 137646 78180 137652 78192
rect 132604 78152 137652 78180
rect 108632 78084 113174 78112
rect 108632 78072 108638 78084
rect 130838 78072 130844 78124
rect 130896 78112 130902 78124
rect 132604 78112 132632 78152
rect 137646 78140 137652 78152
rect 137704 78140 137710 78192
rect 139854 78140 139860 78192
rect 139912 78180 139918 78192
rect 140222 78180 140228 78192
rect 139912 78152 140228 78180
rect 139912 78140 139918 78152
rect 140222 78140 140228 78152
rect 140280 78140 140286 78192
rect 159818 78140 159824 78192
rect 159876 78180 159882 78192
rect 167270 78180 167276 78192
rect 159876 78152 167276 78180
rect 159876 78140 159882 78152
rect 167270 78140 167276 78152
rect 167328 78140 167334 78192
rect 170030 78140 170036 78192
rect 170088 78180 170094 78192
rect 170088 78152 171916 78180
rect 170088 78140 170094 78152
rect 130896 78084 132632 78112
rect 130896 78072 130902 78084
rect 132678 78072 132684 78124
rect 132736 78112 132742 78124
rect 142430 78112 142436 78124
rect 132736 78084 142436 78112
rect 132736 78072 132742 78084
rect 142430 78072 142436 78084
rect 142488 78072 142494 78124
rect 151998 78072 152004 78124
rect 152056 78112 152062 78124
rect 152550 78112 152556 78124
rect 152056 78084 152556 78112
rect 152056 78072 152062 78084
rect 152550 78072 152556 78084
rect 152608 78072 152614 78124
rect 156138 78072 156144 78124
rect 156196 78112 156202 78124
rect 163038 78112 163044 78124
rect 156196 78084 163044 78112
rect 156196 78072 156202 78084
rect 163038 78072 163044 78084
rect 163096 78112 163102 78124
rect 171888 78112 171916 78152
rect 172422 78140 172428 78192
rect 172480 78180 172486 78192
rect 255958 78180 255964 78192
rect 172480 78152 255964 78180
rect 172480 78140 172486 78152
rect 255958 78140 255964 78152
rect 256016 78140 256022 78192
rect 337378 78112 337384 78124
rect 163096 78084 171824 78112
rect 171888 78084 337384 78112
rect 163096 78072 163102 78084
rect 106918 78004 106924 78056
rect 106976 78044 106982 78056
rect 129918 78044 129924 78056
rect 106976 78016 129924 78044
rect 106976 78004 106982 78016
rect 129918 78004 129924 78016
rect 129976 78004 129982 78056
rect 130378 78004 130384 78056
rect 130436 78044 130442 78056
rect 150158 78044 150164 78056
rect 130436 78016 150164 78044
rect 130436 78004 130442 78016
rect 150158 78004 150164 78016
rect 150216 78004 150222 78056
rect 160094 78004 160100 78056
rect 160152 78044 160158 78056
rect 161106 78044 161112 78056
rect 160152 78016 161112 78044
rect 160152 78004 160158 78016
rect 161106 78004 161112 78016
rect 161164 78004 161170 78056
rect 171796 78044 171824 78084
rect 337378 78072 337384 78084
rect 337436 78072 337442 78124
rect 393314 78044 393320 78056
rect 171796 78016 393320 78044
rect 393314 78004 393320 78016
rect 393372 78004 393378 78056
rect 2832 77948 103514 77976
rect 2832 77936 2838 77948
rect 122834 77936 122840 77988
rect 122892 77976 122898 77988
rect 148410 77976 148416 77988
rect 122892 77948 148416 77976
rect 122892 77936 122898 77948
rect 148410 77936 148416 77948
rect 148468 77936 148474 77988
rect 148594 77936 148600 77988
rect 148652 77976 148658 77988
rect 148870 77976 148876 77988
rect 148652 77948 148876 77976
rect 148652 77936 148658 77948
rect 148870 77936 148876 77948
rect 148928 77936 148934 77988
rect 169662 77936 169668 77988
rect 169720 77976 169726 77988
rect 400858 77976 400864 77988
rect 169720 77948 400864 77976
rect 169720 77936 169726 77948
rect 400858 77936 400864 77948
rect 400916 77936 400922 77988
rect 130930 77868 130936 77920
rect 130988 77908 130994 77920
rect 132678 77908 132684 77920
rect 130988 77880 132684 77908
rect 130988 77868 130994 77880
rect 132678 77868 132684 77880
rect 132736 77868 132742 77920
rect 137830 77868 137836 77920
rect 137888 77908 137894 77920
rect 146754 77908 146760 77920
rect 137888 77880 146760 77908
rect 137888 77868 137894 77880
rect 146754 77868 146760 77880
rect 146812 77868 146818 77920
rect 166718 77868 166724 77920
rect 166776 77908 166782 77920
rect 182818 77908 182824 77920
rect 166776 77880 182824 77908
rect 166776 77868 166782 77880
rect 182818 77868 182824 77880
rect 182876 77868 182882 77920
rect 131206 77800 131212 77852
rect 131264 77840 131270 77852
rect 132126 77840 132132 77852
rect 131264 77812 132132 77840
rect 131264 77800 131270 77812
rect 132126 77800 132132 77812
rect 132184 77840 132190 77852
rect 141970 77840 141976 77852
rect 132184 77812 141976 77840
rect 132184 77800 132190 77812
rect 141970 77800 141976 77812
rect 142028 77800 142034 77852
rect 161934 77800 161940 77852
rect 161992 77840 161998 77852
rect 168650 77840 168656 77852
rect 161992 77812 168656 77840
rect 161992 77800 161998 77812
rect 168650 77800 168656 77812
rect 168708 77800 168714 77852
rect 171870 77800 171876 77852
rect 171928 77840 171934 77852
rect 180702 77840 180708 77852
rect 171928 77812 180708 77840
rect 171928 77800 171934 77812
rect 180702 77800 180708 77812
rect 180760 77840 180766 77852
rect 183002 77840 183008 77852
rect 180760 77812 183008 77840
rect 180760 77800 180766 77812
rect 183002 77800 183008 77812
rect 183060 77800 183066 77852
rect 100754 77732 100760 77784
rect 100812 77772 100818 77784
rect 101490 77772 101496 77784
rect 100812 77744 101496 77772
rect 100812 77732 100818 77744
rect 101490 77732 101496 77744
rect 101548 77772 101554 77784
rect 134978 77772 134984 77784
rect 101548 77744 134984 77772
rect 101548 77732 101554 77744
rect 134978 77732 134984 77744
rect 135036 77732 135042 77784
rect 146938 77732 146944 77784
rect 146996 77772 147002 77784
rect 147398 77772 147404 77784
rect 146996 77744 147404 77772
rect 146996 77732 147002 77744
rect 147398 77732 147404 77744
rect 147456 77732 147462 77784
rect 157058 77732 157064 77784
rect 157116 77772 157122 77784
rect 157426 77772 157432 77784
rect 157116 77744 157432 77772
rect 157116 77732 157122 77744
rect 157426 77732 157432 77744
rect 157484 77732 157490 77784
rect 165798 77732 165804 77784
rect 165856 77772 165862 77784
rect 181622 77772 181628 77784
rect 165856 77744 181628 77772
rect 165856 77732 165862 77744
rect 181622 77732 181628 77744
rect 181680 77732 181686 77784
rect 133966 77664 133972 77716
rect 134024 77704 134030 77716
rect 140038 77704 140044 77716
rect 134024 77676 140044 77704
rect 134024 77664 134030 77676
rect 140038 77664 140044 77676
rect 140096 77664 140102 77716
rect 142706 77664 142712 77716
rect 142764 77704 142770 77716
rect 143258 77704 143264 77716
rect 142764 77676 143264 77704
rect 142764 77664 142770 77676
rect 143258 77664 143264 77676
rect 143316 77664 143322 77716
rect 165430 77664 165436 77716
rect 165488 77704 165494 77716
rect 181898 77704 181904 77716
rect 165488 77676 181904 77704
rect 165488 77664 165494 77676
rect 181898 77664 181904 77676
rect 181956 77664 181962 77716
rect 106826 77596 106832 77648
rect 106884 77636 106890 77648
rect 136726 77636 136732 77648
rect 106884 77608 136732 77636
rect 106884 77596 106890 77608
rect 136726 77596 136732 77608
rect 136784 77596 136790 77648
rect 147766 77596 147772 77648
rect 147824 77636 147830 77648
rect 148502 77636 148508 77648
rect 147824 77608 148508 77636
rect 147824 77596 147830 77608
rect 148502 77596 148508 77608
rect 148560 77596 148566 77648
rect 166442 77596 166448 77648
rect 166500 77636 166506 77648
rect 178770 77636 178776 77648
rect 166500 77608 178776 77636
rect 166500 77596 166506 77608
rect 178770 77596 178776 77608
rect 178828 77596 178834 77648
rect 131666 77528 131672 77580
rect 131724 77568 131730 77580
rect 142246 77568 142252 77580
rect 131724 77540 142252 77568
rect 131724 77528 131730 77540
rect 142246 77528 142252 77540
rect 142304 77528 142310 77580
rect 143074 77528 143080 77580
rect 143132 77568 143138 77580
rect 143258 77568 143264 77580
rect 143132 77540 143264 77568
rect 143132 77528 143138 77540
rect 143258 77528 143264 77540
rect 143316 77528 143322 77580
rect 143442 77528 143448 77580
rect 143500 77568 143506 77580
rect 144178 77568 144184 77580
rect 143500 77540 144184 77568
rect 143500 77528 143506 77540
rect 144178 77528 144184 77540
rect 144236 77528 144242 77580
rect 148318 77528 148324 77580
rect 148376 77568 148382 77580
rect 148594 77568 148600 77580
rect 148376 77540 148600 77568
rect 148376 77528 148382 77540
rect 148594 77528 148600 77540
rect 148652 77528 148658 77580
rect 146754 77460 146760 77512
rect 146812 77500 146818 77512
rect 147306 77500 147312 77512
rect 146812 77472 147312 77500
rect 146812 77460 146818 77472
rect 147306 77460 147312 77472
rect 147364 77460 147370 77512
rect 165522 77460 165528 77512
rect 165580 77500 165586 77512
rect 180334 77500 180340 77512
rect 165580 77472 180340 77500
rect 165580 77460 165586 77472
rect 180334 77460 180340 77472
rect 180392 77460 180398 77512
rect 134334 77392 134340 77444
rect 134392 77432 134398 77444
rect 134794 77432 134800 77444
rect 134392 77404 134800 77432
rect 134392 77392 134398 77404
rect 134794 77392 134800 77404
rect 134852 77392 134858 77444
rect 140774 77392 140780 77444
rect 140832 77432 140838 77444
rect 141234 77432 141240 77444
rect 140832 77404 141240 77432
rect 140832 77392 140838 77404
rect 141234 77392 141240 77404
rect 141292 77392 141298 77444
rect 134794 77256 134800 77308
rect 134852 77296 134858 77308
rect 136910 77296 136916 77308
rect 134852 77268 136916 77296
rect 134852 77256 134858 77268
rect 136910 77256 136916 77268
rect 136968 77256 136974 77308
rect 140498 77256 140504 77308
rect 140556 77296 140562 77308
rect 142982 77296 142988 77308
rect 140556 77268 142988 77296
rect 140556 77256 140562 77268
rect 142982 77256 142988 77268
rect 143040 77296 143046 77308
rect 143626 77296 143632 77308
rect 143040 77268 143632 77296
rect 143040 77256 143046 77268
rect 143626 77256 143632 77268
rect 143684 77256 143690 77308
rect 143718 77256 143724 77308
rect 143776 77296 143782 77308
rect 143902 77296 143908 77308
rect 143776 77268 143908 77296
rect 143776 77256 143782 77268
rect 143902 77256 143908 77268
rect 143960 77256 143966 77308
rect 145006 77256 145012 77308
rect 145064 77296 145070 77308
rect 146110 77296 146116 77308
rect 145064 77268 146116 77296
rect 145064 77256 145070 77268
rect 146110 77256 146116 77268
rect 146168 77256 146174 77308
rect 151814 77296 151820 77308
rect 151372 77268 151820 77296
rect 126974 77188 126980 77240
rect 127032 77228 127038 77240
rect 127618 77228 127624 77240
rect 127032 77200 127624 77228
rect 127032 77188 127038 77200
rect 127618 77188 127624 77200
rect 127676 77228 127682 77240
rect 129642 77228 129648 77240
rect 127676 77200 129648 77228
rect 127676 77188 127682 77200
rect 129642 77188 129648 77200
rect 129700 77188 129706 77240
rect 136634 77188 136640 77240
rect 136692 77228 136698 77240
rect 137186 77228 137192 77240
rect 136692 77200 137192 77228
rect 136692 77188 136698 77200
rect 137186 77188 137192 77200
rect 137244 77188 137250 77240
rect 151262 77188 151268 77240
rect 151320 77228 151326 77240
rect 151372 77228 151400 77268
rect 151814 77256 151820 77268
rect 151872 77256 151878 77308
rect 162302 77256 162308 77308
rect 162360 77296 162366 77308
rect 163590 77296 163596 77308
rect 162360 77268 163596 77296
rect 162360 77256 162366 77268
rect 163590 77256 163596 77268
rect 163648 77256 163654 77308
rect 170858 77256 170864 77308
rect 170916 77296 170922 77308
rect 171134 77296 171140 77308
rect 170916 77268 171140 77296
rect 170916 77256 170922 77268
rect 171134 77256 171140 77268
rect 171192 77256 171198 77308
rect 177022 77256 177028 77308
rect 177080 77296 177086 77308
rect 177666 77296 177672 77308
rect 177080 77268 177672 77296
rect 177080 77256 177086 77268
rect 177666 77256 177672 77268
rect 177724 77256 177730 77308
rect 194502 77256 194508 77308
rect 194560 77296 194566 77308
rect 269758 77296 269764 77308
rect 194560 77268 269764 77296
rect 194560 77256 194566 77268
rect 269758 77256 269764 77268
rect 269816 77256 269822 77308
rect 196710 77228 196716 77240
rect 151320 77200 151400 77228
rect 162320 77200 196716 77228
rect 151320 77188 151326 77200
rect 162320 77172 162348 77200
rect 196710 77188 196716 77200
rect 196768 77188 196774 77240
rect 119706 77120 119712 77172
rect 119764 77160 119770 77172
rect 153470 77160 153476 77172
rect 119764 77132 153476 77160
rect 119764 77120 119770 77132
rect 153470 77120 153476 77132
rect 153528 77120 153534 77172
rect 162302 77120 162308 77172
rect 162360 77120 162366 77172
rect 169754 77120 169760 77172
rect 169812 77160 169818 77172
rect 203150 77160 203156 77172
rect 169812 77132 203156 77160
rect 169812 77120 169818 77132
rect 203150 77120 203156 77132
rect 203208 77120 203214 77172
rect 115658 77052 115664 77104
rect 115716 77092 115722 77104
rect 115716 77064 138014 77092
rect 115716 77052 115722 77064
rect 104066 77024 104072 77036
rect 103486 76996 104072 77024
rect 66254 76644 66260 76696
rect 66312 76684 66318 76696
rect 103486 76684 103514 76996
rect 104066 76984 104072 76996
rect 104124 77024 104130 77036
rect 137462 77024 137468 77036
rect 104124 76996 137468 77024
rect 104124 76984 104130 76996
rect 137462 76984 137468 76996
rect 137520 76984 137526 77036
rect 137986 77024 138014 77064
rect 155402 77052 155408 77104
rect 155460 77092 155466 77104
rect 187418 77092 187424 77104
rect 155460 77064 187424 77092
rect 155460 77052 155466 77064
rect 187418 77052 187424 77064
rect 187476 77092 187482 77104
rect 188798 77092 188804 77104
rect 187476 77064 188804 77092
rect 187476 77052 187482 77064
rect 188798 77052 188804 77064
rect 188856 77052 188862 77104
rect 148226 77024 148232 77036
rect 137986 76996 148232 77024
rect 148226 76984 148232 76996
rect 148284 76984 148290 77036
rect 171594 76984 171600 77036
rect 171652 77024 171658 77036
rect 191466 77024 191472 77036
rect 171652 76996 191472 77024
rect 171652 76984 171658 76996
rect 191466 76984 191472 76996
rect 191524 77024 191530 77036
rect 191742 77024 191748 77036
rect 191524 76996 191748 77024
rect 191524 76984 191530 76996
rect 191742 76984 191748 76996
rect 191800 76984 191806 77036
rect 117222 76916 117228 76968
rect 117280 76956 117286 76968
rect 148778 76956 148784 76968
rect 117280 76928 148784 76956
rect 117280 76916 117286 76928
rect 148778 76916 148784 76928
rect 148836 76916 148842 76968
rect 154850 76916 154856 76968
rect 154908 76956 154914 76968
rect 184474 76956 184480 76968
rect 154908 76928 184480 76956
rect 154908 76916 154914 76928
rect 184474 76916 184480 76928
rect 184532 76916 184538 76968
rect 120534 76848 120540 76900
rect 120592 76888 120598 76900
rect 120592 76860 142844 76888
rect 120592 76848 120598 76860
rect 115750 76780 115756 76832
rect 115808 76820 115814 76832
rect 115808 76792 138060 76820
rect 115808 76780 115814 76792
rect 108298 76752 108304 76764
rect 66312 76656 103514 76684
rect 106292 76724 108304 76752
rect 66312 76644 66318 76656
rect 59354 76576 59360 76628
rect 59412 76616 59418 76628
rect 106292 76616 106320 76724
rect 108298 76712 108304 76724
rect 108356 76752 108362 76764
rect 108356 76724 131804 76752
rect 108356 76712 108362 76724
rect 106366 76644 106372 76696
rect 106424 76684 106430 76696
rect 131666 76684 131672 76696
rect 106424 76656 131672 76684
rect 106424 76644 106430 76656
rect 131666 76644 131672 76656
rect 131724 76644 131730 76696
rect 59412 76588 106320 76616
rect 131776 76616 131804 76724
rect 138032 76684 138060 76792
rect 142816 76752 142844 76860
rect 151078 76848 151084 76900
rect 151136 76888 151142 76900
rect 151136 76860 157334 76888
rect 151136 76848 151142 76860
rect 156966 76780 156972 76832
rect 157024 76820 157030 76832
rect 157150 76820 157156 76832
rect 157024 76792 157156 76820
rect 157024 76780 157030 76792
rect 157150 76780 157156 76792
rect 157208 76780 157214 76832
rect 157306 76820 157334 76860
rect 172514 76848 172520 76900
rect 172572 76888 172578 76900
rect 173526 76888 173532 76900
rect 172572 76860 173532 76888
rect 172572 76848 172578 76860
rect 173526 76848 173532 76860
rect 173584 76848 173590 76900
rect 184198 76848 184204 76900
rect 184256 76888 184262 76900
rect 200850 76888 200856 76900
rect 184256 76860 200856 76888
rect 184256 76848 184262 76860
rect 200850 76848 200856 76860
rect 200908 76848 200914 76900
rect 224218 76820 224224 76832
rect 157306 76792 224224 76820
rect 224218 76780 224224 76792
rect 224276 76780 224282 76832
rect 151262 76752 151268 76764
rect 142816 76724 151268 76752
rect 151262 76712 151268 76724
rect 151320 76752 151326 76764
rect 247034 76752 247040 76764
rect 151320 76724 247040 76752
rect 151320 76712 151326 76724
rect 247034 76712 247040 76724
rect 247092 76712 247098 76764
rect 146018 76684 146024 76696
rect 138032 76656 146024 76684
rect 146018 76644 146024 76656
rect 146076 76684 146082 76696
rect 151078 76684 151084 76696
rect 146076 76656 151084 76684
rect 146076 76644 146082 76656
rect 151078 76644 151084 76656
rect 151136 76644 151142 76696
rect 153102 76644 153108 76696
rect 153160 76684 153166 76696
rect 253934 76684 253940 76696
rect 153160 76656 253940 76684
rect 153160 76644 153166 76656
rect 253934 76644 253940 76656
rect 253992 76644 253998 76696
rect 134794 76616 134800 76628
rect 131776 76588 134800 76616
rect 59412 76576 59418 76588
rect 134794 76576 134800 76588
rect 134852 76576 134858 76628
rect 150710 76576 150716 76628
rect 150768 76616 150774 76628
rect 150894 76616 150900 76628
rect 150768 76588 150900 76616
rect 150768 76576 150774 76588
rect 150894 76576 150900 76588
rect 150952 76576 150958 76628
rect 181346 76616 181352 76628
rect 158686 76588 181352 76616
rect 52454 76508 52460 76560
rect 52512 76548 52518 76560
rect 135990 76548 135996 76560
rect 52512 76520 135996 76548
rect 52512 76508 52518 76520
rect 135990 76508 135996 76520
rect 136048 76508 136054 76560
rect 150066 76508 150072 76560
rect 150124 76548 150130 76560
rect 158686 76548 158714 76588
rect 181346 76576 181352 76588
rect 181404 76576 181410 76628
rect 191742 76576 191748 76628
rect 191800 76616 191806 76628
rect 353294 76616 353300 76628
rect 191800 76588 353300 76616
rect 191800 76576 191806 76588
rect 353294 76576 353300 76588
rect 353352 76576 353358 76628
rect 150124 76520 158714 76548
rect 150124 76508 150130 76520
rect 162578 76508 162584 76560
rect 162636 76548 162642 76560
rect 389174 76548 389180 76560
rect 162636 76520 389180 76548
rect 162636 76508 162642 76520
rect 389174 76508 389180 76520
rect 389232 76508 389238 76560
rect 123018 76440 123024 76492
rect 123076 76480 123082 76492
rect 141602 76480 141608 76492
rect 123076 76452 141608 76480
rect 123076 76440 123082 76452
rect 141602 76440 141608 76452
rect 141660 76440 141666 76492
rect 114370 76372 114376 76424
rect 114428 76412 114434 76424
rect 141050 76412 141056 76424
rect 114428 76384 141056 76412
rect 114428 76372 114434 76384
rect 141050 76372 141056 76384
rect 141108 76372 141114 76424
rect 177206 76372 177212 76424
rect 177264 76412 177270 76424
rect 207106 76412 207112 76424
rect 177264 76384 207112 76412
rect 177264 76372 177270 76384
rect 207106 76372 207112 76384
rect 207164 76372 207170 76424
rect 115474 76304 115480 76356
rect 115532 76344 115538 76356
rect 149790 76344 149796 76356
rect 115532 76316 149796 76344
rect 115532 76304 115538 76316
rect 149790 76304 149796 76316
rect 149848 76304 149854 76356
rect 169754 76304 169760 76356
rect 169812 76344 169818 76356
rect 170582 76344 170588 76356
rect 169812 76316 170588 76344
rect 169812 76304 169818 76316
rect 170582 76304 170588 76316
rect 170640 76304 170646 76356
rect 173342 76304 173348 76356
rect 173400 76344 173406 76356
rect 184198 76344 184204 76356
rect 173400 76316 184204 76344
rect 173400 76304 173406 76316
rect 184198 76304 184204 76316
rect 184256 76304 184262 76356
rect 131666 76236 131672 76288
rect 131724 76276 131730 76288
rect 139578 76276 139584 76288
rect 131724 76248 139584 76276
rect 131724 76236 131730 76248
rect 139578 76236 139584 76248
rect 139636 76236 139642 76288
rect 164418 76236 164424 76288
rect 164476 76276 164482 76288
rect 165430 76276 165436 76288
rect 164476 76248 165436 76276
rect 164476 76236 164482 76248
rect 165430 76236 165436 76248
rect 165488 76236 165494 76288
rect 173434 76236 173440 76288
rect 173492 76276 173498 76288
rect 173710 76276 173716 76288
rect 173492 76248 173716 76276
rect 173492 76236 173498 76248
rect 173710 76236 173716 76248
rect 173768 76236 173774 76288
rect 129642 76168 129648 76220
rect 129700 76208 129706 76220
rect 141786 76208 141792 76220
rect 129700 76180 141792 76208
rect 129700 76168 129706 76180
rect 141786 76168 141792 76180
rect 141844 76168 141850 76220
rect 143350 76168 143356 76220
rect 143408 76208 143414 76220
rect 144730 76208 144736 76220
rect 143408 76180 144736 76208
rect 143408 76168 143414 76180
rect 144730 76168 144736 76180
rect 144788 76168 144794 76220
rect 165246 76100 165252 76152
rect 165304 76140 165310 76152
rect 165430 76140 165436 76152
rect 165304 76112 165436 76140
rect 165304 76100 165310 76112
rect 165430 76100 165436 76112
rect 165488 76100 165494 76152
rect 145374 76032 145380 76084
rect 145432 76072 145438 76084
rect 146018 76072 146024 76084
rect 145432 76044 146024 76072
rect 145432 76032 145438 76044
rect 146018 76032 146024 76044
rect 146076 76032 146082 76084
rect 173066 75964 173072 76016
rect 173124 76004 173130 76016
rect 173802 76004 173808 76016
rect 173124 75976 173808 76004
rect 173124 75964 173130 75976
rect 173802 75964 173808 75976
rect 173860 75964 173866 76016
rect 174354 75964 174360 76016
rect 174412 76004 174418 76016
rect 175182 76004 175188 76016
rect 174412 75976 175188 76004
rect 174412 75964 174418 75976
rect 175182 75964 175188 75976
rect 175240 75964 175246 76016
rect 184474 75964 184480 76016
rect 184532 76004 184538 76016
rect 289814 76004 289820 76016
rect 184532 75976 289820 76004
rect 184532 75964 184538 75976
rect 289814 75964 289820 75976
rect 289872 75964 289878 76016
rect 111794 75896 111800 75948
rect 111852 75936 111858 75948
rect 113634 75936 113640 75948
rect 111852 75908 113640 75936
rect 111852 75896 111858 75908
rect 113634 75896 113640 75908
rect 113692 75936 113698 75948
rect 114370 75936 114376 75948
rect 113692 75908 114376 75936
rect 113692 75896 113698 75908
rect 114370 75896 114376 75908
rect 114428 75896 114434 75948
rect 134518 75896 134524 75948
rect 134576 75936 134582 75948
rect 134702 75936 134708 75948
rect 134576 75908 134708 75936
rect 134576 75896 134582 75908
rect 134702 75896 134708 75908
rect 134760 75896 134766 75948
rect 173894 75896 173900 75948
rect 173952 75936 173958 75948
rect 174538 75936 174544 75948
rect 173952 75908 174544 75936
rect 173952 75896 173958 75908
rect 174538 75896 174544 75908
rect 174596 75896 174602 75948
rect 177206 75896 177212 75948
rect 177264 75936 177270 75948
rect 177666 75936 177672 75948
rect 177264 75908 177672 75936
rect 177264 75896 177270 75908
rect 177666 75896 177672 75908
rect 177724 75896 177730 75948
rect 188798 75896 188804 75948
rect 188856 75936 188862 75948
rect 296714 75936 296720 75948
rect 188856 75908 296720 75936
rect 188856 75896 188862 75908
rect 296714 75896 296720 75908
rect 296772 75896 296778 75948
rect 118234 75828 118240 75880
rect 118292 75868 118298 75880
rect 145098 75868 145104 75880
rect 118292 75840 145104 75868
rect 118292 75828 118298 75840
rect 145098 75828 145104 75840
rect 145156 75868 145162 75880
rect 148318 75868 148324 75880
rect 145156 75840 148324 75868
rect 145156 75828 145162 75840
rect 148318 75828 148324 75840
rect 148376 75828 148382 75880
rect 168834 75828 168840 75880
rect 168892 75868 168898 75880
rect 169570 75868 169576 75880
rect 168892 75840 169576 75868
rect 168892 75828 168898 75840
rect 169570 75828 169576 75840
rect 169628 75828 169634 75880
rect 105538 75760 105544 75812
rect 105596 75800 105602 75812
rect 139486 75800 139492 75812
rect 105596 75772 139492 75800
rect 105596 75760 105602 75772
rect 139486 75760 139492 75772
rect 139544 75760 139550 75812
rect 161382 75760 161388 75812
rect 161440 75800 161446 75812
rect 195514 75800 195520 75812
rect 161440 75772 195520 75800
rect 161440 75760 161446 75772
rect 195514 75760 195520 75772
rect 195572 75760 195578 75812
rect 113726 75692 113732 75744
rect 113784 75732 113790 75744
rect 146662 75732 146668 75744
rect 113784 75704 146668 75732
rect 113784 75692 113790 75704
rect 146662 75692 146668 75704
rect 146720 75692 146726 75744
rect 156322 75692 156328 75744
rect 156380 75732 156386 75744
rect 156690 75732 156696 75744
rect 156380 75704 156696 75732
rect 156380 75692 156386 75704
rect 156690 75692 156696 75704
rect 156748 75732 156754 75744
rect 190638 75732 190644 75744
rect 156748 75704 190644 75732
rect 156748 75692 156754 75704
rect 190638 75692 190644 75704
rect 190696 75692 190702 75744
rect 113082 75624 113088 75676
rect 113140 75664 113146 75676
rect 145650 75664 145656 75676
rect 113140 75636 145656 75664
rect 113140 75624 113146 75636
rect 145650 75624 145656 75636
rect 145708 75624 145714 75676
rect 146478 75624 146484 75676
rect 146536 75664 146542 75676
rect 180794 75664 180800 75676
rect 146536 75636 180800 75664
rect 146536 75624 146542 75636
rect 180794 75624 180800 75636
rect 180852 75624 180858 75676
rect 115906 75568 120120 75596
rect 114094 75488 114100 75540
rect 114152 75528 114158 75540
rect 115906 75528 115934 75568
rect 114152 75500 115934 75528
rect 120092 75528 120120 75568
rect 120718 75556 120724 75608
rect 120776 75596 120782 75608
rect 135438 75596 135444 75608
rect 120776 75568 135444 75596
rect 120776 75556 120782 75568
rect 135438 75556 135444 75568
rect 135496 75556 135502 75608
rect 148042 75556 148048 75608
rect 148100 75596 148106 75608
rect 181530 75596 181536 75608
rect 148100 75568 181536 75596
rect 148100 75556 148106 75568
rect 181530 75556 181536 75568
rect 181588 75556 181594 75608
rect 120092 75500 133000 75528
rect 114152 75488 114158 75500
rect 104250 75420 104256 75472
rect 104308 75460 104314 75472
rect 120718 75460 120724 75472
rect 104308 75432 120724 75460
rect 104308 75420 104314 75432
rect 120718 75420 120724 75432
rect 120776 75420 120782 75472
rect 132972 75460 133000 75500
rect 133202 75500 138014 75528
rect 133202 75460 133230 75500
rect 132972 75432 133230 75460
rect 134058 75420 134064 75472
rect 134116 75460 134122 75472
rect 134518 75460 134524 75472
rect 134116 75432 134524 75460
rect 134116 75420 134122 75432
rect 134518 75420 134524 75432
rect 134576 75420 134582 75472
rect 137986 75460 138014 75500
rect 147674 75488 147680 75540
rect 147732 75528 147738 75540
rect 198734 75528 198740 75540
rect 147732 75500 198740 75528
rect 147732 75488 147738 75500
rect 198734 75488 198740 75500
rect 198792 75488 198798 75540
rect 147122 75460 147128 75472
rect 137986 75432 147128 75460
rect 147122 75420 147128 75432
rect 147180 75460 147186 75472
rect 187694 75460 187700 75472
rect 147180 75432 187700 75460
rect 147180 75420 147186 75432
rect 187694 75420 187700 75432
rect 187752 75420 187758 75472
rect 114462 75352 114468 75404
rect 114520 75392 114526 75404
rect 145466 75392 145472 75404
rect 114520 75364 145472 75392
rect 114520 75352 114526 75364
rect 145466 75352 145472 75364
rect 145524 75352 145530 75404
rect 148870 75352 148876 75404
rect 148928 75392 148934 75404
rect 201494 75392 201500 75404
rect 148928 75364 201500 75392
rect 148928 75352 148934 75364
rect 201494 75352 201500 75364
rect 201552 75352 201558 75404
rect 96614 75284 96620 75336
rect 96672 75324 96678 75336
rect 108758 75324 108764 75336
rect 96672 75296 108764 75324
rect 96672 75284 96678 75296
rect 108758 75284 108764 75296
rect 108816 75324 108822 75336
rect 140222 75324 140228 75336
rect 108816 75296 140228 75324
rect 108816 75284 108822 75296
rect 140222 75284 140228 75296
rect 140280 75284 140286 75336
rect 173250 75284 173256 75336
rect 173308 75324 173314 75336
rect 453298 75324 453304 75336
rect 173308 75296 453304 75324
rect 173308 75284 173314 75296
rect 453298 75284 453304 75296
rect 453356 75284 453362 75336
rect 81434 75216 81440 75268
rect 81492 75256 81498 75268
rect 138750 75256 138756 75268
rect 81492 75228 138756 75256
rect 81492 75216 81498 75228
rect 138750 75216 138756 75228
rect 138808 75216 138814 75268
rect 149422 75216 149428 75268
rect 149480 75256 149486 75268
rect 150066 75256 150072 75268
rect 149480 75228 150072 75256
rect 149480 75216 149486 75228
rect 150066 75216 150072 75228
rect 150124 75216 150130 75268
rect 163038 75216 163044 75268
rect 163096 75256 163102 75268
rect 163682 75256 163688 75268
rect 163096 75228 163688 75256
rect 163096 75216 163102 75228
rect 163682 75216 163688 75228
rect 163740 75216 163746 75268
rect 172882 75216 172888 75268
rect 172940 75256 172946 75268
rect 506474 75256 506480 75268
rect 172940 75228 506480 75256
rect 172940 75216 172946 75228
rect 506474 75216 506480 75228
rect 506532 75216 506538 75268
rect 27614 75148 27620 75200
rect 27672 75188 27678 75200
rect 100110 75188 100116 75200
rect 27672 75160 100116 75188
rect 27672 75148 27678 75160
rect 100110 75148 100116 75160
rect 100168 75188 100174 75200
rect 141418 75188 141424 75200
rect 100168 75160 103514 75188
rect 100168 75148 100174 75160
rect 103486 75052 103514 75160
rect 115124 75160 141424 75188
rect 115124 75132 115152 75160
rect 141418 75148 141424 75160
rect 141476 75148 141482 75200
rect 163130 75148 163136 75200
rect 163188 75188 163194 75200
rect 164050 75188 164056 75200
rect 163188 75160 164056 75188
rect 163188 75148 163194 75160
rect 164050 75148 164056 75160
rect 164108 75148 164114 75200
rect 172330 75148 172336 75200
rect 172388 75188 172394 75200
rect 511258 75188 511264 75200
rect 172388 75160 511264 75188
rect 172388 75148 172394 75160
rect 511258 75148 511264 75160
rect 511316 75148 511322 75200
rect 114554 75080 114560 75132
rect 114612 75120 114618 75132
rect 115106 75120 115112 75132
rect 114612 75092 115112 75120
rect 114612 75080 114618 75092
rect 115106 75080 115112 75092
rect 115164 75080 115170 75132
rect 121270 75080 121276 75132
rect 121328 75120 121334 75132
rect 147214 75120 147220 75132
rect 121328 75092 147220 75120
rect 121328 75080 121334 75092
rect 147214 75080 147220 75092
rect 147272 75080 147278 75132
rect 167822 75080 167828 75132
rect 167880 75120 167886 75132
rect 192662 75120 192668 75132
rect 167880 75092 192668 75120
rect 167880 75080 167886 75092
rect 192662 75080 192668 75092
rect 192720 75080 192726 75132
rect 132402 75052 132408 75064
rect 103486 75024 132408 75052
rect 132402 75012 132408 75024
rect 132460 75012 132466 75064
rect 114002 74944 114008 74996
rect 114060 74984 114066 74996
rect 146478 74984 146484 74996
rect 114060 74956 146484 74984
rect 114060 74944 114066 74956
rect 146478 74944 146484 74956
rect 146536 74944 146542 74996
rect 155862 74944 155868 74996
rect 155920 74984 155926 74996
rect 156782 74984 156788 74996
rect 155920 74956 156788 74984
rect 155920 74944 155926 74956
rect 156782 74944 156788 74956
rect 156840 74984 156846 74996
rect 190730 74984 190736 74996
rect 156840 74956 190736 74984
rect 156840 74944 156846 74956
rect 190730 74944 190736 74956
rect 190788 74944 190794 74996
rect 173986 74876 173992 74928
rect 174044 74916 174050 74928
rect 174906 74916 174912 74928
rect 174044 74888 174912 74916
rect 174044 74876 174050 74888
rect 174906 74876 174912 74888
rect 174964 74876 174970 74928
rect 145650 74808 145656 74860
rect 145708 74848 145714 74860
rect 145926 74848 145932 74860
rect 145708 74820 145932 74848
rect 145708 74808 145714 74820
rect 145926 74808 145932 74820
rect 145984 74808 145990 74860
rect 173986 74740 173992 74792
rect 174044 74780 174050 74792
rect 174262 74780 174268 74792
rect 174044 74752 174268 74780
rect 174044 74740 174050 74752
rect 174262 74740 174268 74752
rect 174320 74740 174326 74792
rect 165062 74604 165068 74656
rect 165120 74644 165126 74656
rect 178862 74644 178868 74656
rect 165120 74616 178868 74644
rect 165120 74604 165126 74616
rect 178862 74604 178868 74616
rect 178920 74604 178926 74656
rect 121362 74468 121368 74520
rect 121420 74508 121426 74520
rect 131114 74508 131120 74520
rect 121420 74480 131120 74508
rect 121420 74468 121426 74480
rect 131114 74468 131120 74480
rect 131172 74508 131178 74520
rect 132310 74508 132316 74520
rect 131172 74480 132316 74508
rect 131172 74468 131178 74480
rect 132310 74468 132316 74480
rect 132368 74468 132374 74520
rect 143902 74468 143908 74520
rect 143960 74508 143966 74520
rect 144454 74508 144460 74520
rect 143960 74480 144460 74508
rect 143960 74468 143966 74480
rect 144454 74468 144460 74480
rect 144512 74468 144518 74520
rect 145558 74468 145564 74520
rect 145616 74508 145622 74520
rect 145834 74508 145840 74520
rect 145616 74480 145840 74508
rect 145616 74468 145622 74480
rect 145834 74468 145840 74480
rect 145892 74468 145898 74520
rect 154022 74468 154028 74520
rect 154080 74508 154086 74520
rect 154206 74508 154212 74520
rect 154080 74480 154212 74508
rect 154080 74468 154086 74480
rect 154206 74468 154212 74480
rect 154264 74468 154270 74520
rect 157886 74468 157892 74520
rect 157944 74508 157950 74520
rect 158162 74508 158168 74520
rect 157944 74480 158168 74508
rect 157944 74468 157950 74480
rect 158162 74468 158168 74480
rect 158220 74508 158226 74520
rect 192294 74508 192300 74520
rect 158220 74480 192300 74508
rect 158220 74468 158226 74480
rect 192294 74468 192300 74480
rect 192352 74468 192358 74520
rect 110138 74400 110144 74452
rect 110196 74440 110202 74452
rect 144638 74440 144644 74452
rect 110196 74412 144644 74440
rect 110196 74400 110202 74412
rect 144638 74400 144644 74412
rect 144696 74400 144702 74452
rect 161198 74400 161204 74452
rect 161256 74440 161262 74452
rect 164878 74440 164884 74452
rect 161256 74412 164884 74440
rect 161256 74400 161262 74412
rect 164878 74400 164884 74412
rect 164936 74400 164942 74452
rect 166994 74400 167000 74452
rect 167052 74440 167058 74452
rect 200574 74440 200580 74452
rect 167052 74412 200580 74440
rect 167052 74400 167058 74412
rect 200574 74400 200580 74412
rect 200632 74400 200638 74452
rect 115566 74332 115572 74384
rect 115624 74372 115630 74384
rect 115624 74344 147674 74372
rect 115624 74332 115630 74344
rect 112714 74264 112720 74316
rect 112772 74304 112778 74316
rect 146110 74304 146116 74316
rect 112772 74276 146116 74304
rect 112772 74264 112778 74276
rect 146110 74264 146116 74276
rect 146168 74264 146174 74316
rect 111150 74196 111156 74248
rect 111208 74236 111214 74248
rect 143166 74236 143172 74248
rect 111208 74208 143172 74236
rect 111208 74196 111214 74208
rect 143166 74196 143172 74208
rect 143224 74196 143230 74248
rect 147646 74236 147674 74344
rect 153378 74332 153384 74384
rect 153436 74372 153442 74384
rect 154206 74372 154212 74384
rect 153436 74344 154212 74372
rect 153436 74332 153442 74344
rect 154206 74332 154212 74344
rect 154264 74372 154270 74384
rect 188522 74372 188528 74384
rect 154264 74344 188528 74372
rect 154264 74332 154270 74344
rect 188522 74332 188528 74344
rect 188580 74332 188586 74384
rect 160738 74264 160744 74316
rect 160796 74304 160802 74316
rect 161290 74304 161296 74316
rect 160796 74276 161296 74304
rect 160796 74264 160802 74276
rect 161290 74264 161296 74276
rect 161348 74264 161354 74316
rect 171318 74264 171324 74316
rect 171376 74304 171382 74316
rect 172146 74304 172152 74316
rect 171376 74276 172152 74304
rect 171376 74264 171382 74276
rect 172146 74264 172152 74276
rect 172204 74264 172210 74316
rect 175366 74264 175372 74316
rect 175424 74304 175430 74316
rect 176194 74304 176200 74316
rect 175424 74276 176200 74304
rect 175424 74264 175430 74276
rect 176194 74264 176200 74276
rect 176252 74304 176258 74316
rect 205910 74304 205916 74316
rect 176252 74276 205916 74304
rect 176252 74264 176258 74276
rect 205910 74264 205916 74276
rect 205968 74264 205974 74316
rect 149974 74236 149980 74248
rect 147646 74208 149980 74236
rect 149974 74196 149980 74208
rect 150032 74236 150038 74248
rect 203702 74236 203708 74248
rect 150032 74208 203708 74236
rect 150032 74196 150038 74208
rect 203702 74196 203708 74208
rect 203760 74196 203766 74248
rect 104342 74128 104348 74180
rect 104400 74168 104406 74180
rect 134242 74168 134248 74180
rect 104400 74140 134248 74168
rect 104400 74128 104406 74140
rect 134242 74128 134248 74140
rect 134300 74168 134306 74180
rect 135162 74168 135168 74180
rect 134300 74140 135168 74168
rect 134300 74128 134306 74140
rect 135162 74128 135168 74140
rect 135220 74128 135226 74180
rect 136910 74128 136916 74180
rect 136968 74168 136974 74180
rect 137922 74168 137928 74180
rect 136968 74140 137928 74168
rect 136968 74128 136974 74140
rect 137922 74128 137928 74140
rect 137980 74128 137986 74180
rect 152734 74128 152740 74180
rect 152792 74168 152798 74180
rect 262214 74168 262220 74180
rect 152792 74140 262220 74168
rect 152792 74128 152798 74140
rect 262214 74128 262220 74140
rect 262272 74128 262278 74180
rect 116670 74060 116676 74112
rect 116728 74100 116734 74112
rect 145834 74100 145840 74112
rect 116728 74072 145840 74100
rect 116728 74060 116734 74072
rect 145834 74060 145840 74072
rect 145892 74060 145898 74112
rect 154482 74060 154488 74112
rect 154540 74100 154546 74112
rect 284294 74100 284300 74112
rect 154540 74072 284300 74100
rect 154540 74060 154546 74072
rect 284294 74060 284300 74072
rect 284352 74060 284358 74112
rect 118050 73992 118056 74044
rect 118108 74032 118114 74044
rect 143994 74032 144000 74044
rect 118108 74004 144000 74032
rect 118108 73992 118114 74004
rect 143994 73992 144000 74004
rect 144052 73992 144058 74044
rect 144270 73992 144276 74044
rect 144328 74032 144334 74044
rect 144638 74032 144644 74044
rect 144328 74004 144644 74032
rect 144328 73992 144334 74004
rect 144638 73992 144644 74004
rect 144696 73992 144702 74044
rect 155954 73992 155960 74044
rect 156012 74032 156018 74044
rect 297358 74032 297364 74044
rect 156012 74004 297364 74032
rect 156012 73992 156018 74004
rect 297358 73992 297364 74004
rect 297416 73992 297422 74044
rect 119614 73924 119620 73976
rect 119672 73964 119678 73976
rect 119672 73936 142982 73964
rect 119672 73924 119678 73936
rect 99374 73856 99380 73908
rect 99432 73896 99438 73908
rect 140314 73896 140320 73908
rect 99432 73868 140320 73896
rect 99432 73856 99438 73868
rect 140314 73856 140320 73868
rect 140372 73856 140378 73908
rect 142954 73896 142982 73936
rect 144086 73924 144092 73976
rect 144144 73964 144150 73976
rect 149698 73964 149704 73976
rect 144144 73936 149704 73964
rect 144144 73924 144150 73936
rect 149698 73924 149704 73936
rect 149756 73924 149762 73976
rect 159174 73924 159180 73976
rect 159232 73964 159238 73976
rect 347774 73964 347780 73976
rect 159232 73936 347780 73964
rect 159232 73924 159238 73936
rect 347774 73924 347780 73936
rect 347832 73924 347838 73976
rect 145190 73896 145196 73908
rect 142954 73868 145196 73896
rect 145190 73856 145196 73868
rect 145248 73856 145254 73908
rect 153470 73856 153476 73908
rect 153528 73896 153534 73908
rect 269114 73896 269120 73908
rect 153528 73868 269120 73896
rect 153528 73856 153534 73868
rect 269114 73856 269120 73868
rect 269172 73856 269178 73908
rect 269758 73856 269764 73908
rect 269816 73896 269822 73908
rect 465166 73896 465172 73908
rect 269816 73868 465172 73896
rect 269816 73856 269822 73868
rect 465166 73856 465172 73868
rect 465224 73856 465230 73908
rect 78674 73788 78680 73840
rect 78732 73828 78738 73840
rect 138290 73828 138296 73840
rect 78732 73800 138296 73828
rect 78732 73788 78738 73800
rect 138290 73788 138296 73800
rect 138348 73788 138354 73840
rect 151722 73788 151728 73840
rect 151780 73828 151786 73840
rect 248414 73828 248420 73840
rect 151780 73800 248420 73828
rect 151780 73788 151786 73800
rect 248414 73788 248420 73800
rect 248472 73788 248478 73840
rect 255958 73788 255964 73840
rect 256016 73828 256022 73840
rect 456794 73828 456800 73840
rect 256016 73800 456800 73828
rect 256016 73788 256022 73800
rect 456794 73788 456800 73800
rect 456852 73788 456858 73840
rect 119522 73720 119528 73772
rect 119580 73760 119586 73772
rect 144454 73760 144460 73772
rect 119580 73732 144460 73760
rect 119580 73720 119586 73732
rect 144454 73720 144460 73732
rect 144512 73720 144518 73772
rect 153194 73720 153200 73772
rect 153252 73760 153258 73772
rect 154298 73760 154304 73772
rect 153252 73732 154304 73760
rect 153252 73720 153258 73732
rect 154298 73720 154304 73732
rect 154356 73720 154362 73772
rect 171318 73720 171324 73772
rect 171376 73760 171382 73772
rect 171686 73760 171692 73772
rect 171376 73732 171692 73760
rect 171376 73720 171382 73732
rect 171686 73720 171692 73732
rect 171744 73720 171750 73772
rect 175550 73720 175556 73772
rect 175608 73760 175614 73772
rect 176470 73760 176476 73772
rect 175608 73732 176476 73760
rect 175608 73720 175614 73732
rect 176470 73720 176476 73732
rect 176528 73760 176534 73772
rect 206002 73760 206008 73772
rect 176528 73732 206008 73760
rect 176528 73720 176534 73732
rect 206002 73720 206008 73732
rect 206060 73720 206066 73772
rect 124858 73652 124864 73704
rect 124916 73692 124922 73704
rect 125594 73692 125600 73704
rect 124916 73664 125600 73692
rect 124916 73652 124922 73664
rect 125594 73652 125600 73664
rect 125652 73652 125658 73704
rect 132678 73652 132684 73704
rect 132736 73692 132742 73704
rect 133690 73692 133696 73704
rect 132736 73664 133696 73692
rect 132736 73652 132742 73664
rect 133690 73652 133696 73664
rect 133748 73652 133754 73704
rect 172146 73652 172152 73704
rect 172204 73692 172210 73704
rect 194962 73692 194968 73704
rect 172204 73664 194968 73692
rect 172204 73652 172210 73664
rect 194962 73652 194968 73664
rect 195020 73652 195026 73704
rect 114738 73584 114744 73636
rect 114796 73624 114802 73636
rect 149146 73624 149152 73636
rect 114796 73596 149152 73624
rect 114796 73584 114802 73596
rect 149146 73584 149152 73596
rect 149204 73624 149210 73636
rect 149974 73624 149980 73636
rect 149204 73596 149980 73624
rect 149204 73584 149210 73596
rect 149974 73584 149980 73596
rect 150032 73584 150038 73636
rect 168466 73584 168472 73636
rect 168524 73624 168530 73636
rect 169202 73624 169208 73636
rect 168524 73596 169208 73624
rect 168524 73584 168530 73596
rect 169202 73584 169208 73596
rect 169260 73584 169266 73636
rect 166350 73516 166356 73568
rect 166408 73556 166414 73568
rect 183738 73556 183744 73568
rect 166408 73528 183744 73556
rect 166408 73516 166414 73528
rect 183738 73516 183744 73528
rect 183796 73516 183802 73568
rect 145190 73448 145196 73500
rect 145248 73488 145254 73500
rect 145650 73488 145656 73500
rect 145248 73460 145656 73488
rect 145248 73448 145254 73460
rect 145650 73448 145656 73460
rect 145708 73448 145714 73500
rect 164326 73176 164332 73228
rect 164384 73216 164390 73228
rect 164970 73216 164976 73228
rect 164384 73188 164976 73216
rect 164384 73176 164390 73188
rect 164970 73176 164976 73188
rect 165028 73176 165034 73228
rect 118602 73108 118608 73160
rect 118660 73148 118666 73160
rect 152274 73148 152280 73160
rect 118660 73120 152280 73148
rect 118660 73108 118666 73120
rect 152274 73108 152280 73120
rect 152332 73108 152338 73160
rect 163314 73108 163320 73160
rect 163372 73148 163378 73160
rect 163682 73148 163688 73160
rect 163372 73120 163688 73148
rect 163372 73108 163378 73120
rect 163682 73108 163688 73120
rect 163740 73108 163746 73160
rect 167178 73108 167184 73160
rect 167236 73148 167242 73160
rect 208486 73148 208492 73160
rect 167236 73120 208492 73148
rect 167236 73108 167242 73120
rect 208486 73108 208492 73120
rect 208544 73148 208550 73160
rect 208544 73120 209774 73148
rect 208544 73108 208550 73120
rect 109862 73040 109868 73092
rect 109920 73080 109926 73092
rect 143902 73080 143908 73092
rect 109920 73052 143908 73080
rect 109920 73040 109926 73052
rect 143902 73040 143908 73052
rect 143960 73080 143966 73092
rect 147030 73080 147036 73092
rect 143960 73052 147036 73080
rect 143960 73040 143966 73052
rect 147030 73040 147036 73052
rect 147088 73040 147094 73092
rect 168098 73040 168104 73092
rect 168156 73080 168162 73092
rect 202138 73080 202144 73092
rect 168156 73052 202144 73080
rect 168156 73040 168162 73052
rect 202138 73040 202144 73052
rect 202196 73040 202202 73092
rect 102134 72972 102140 73024
rect 102192 73012 102198 73024
rect 102778 73012 102784 73024
rect 102192 72984 102784 73012
rect 102192 72972 102198 72984
rect 102778 72972 102784 72984
rect 102836 73012 102842 73024
rect 135530 73012 135536 73024
rect 102836 72984 135536 73012
rect 102836 72972 102842 72984
rect 135530 72972 135536 72984
rect 135588 72972 135594 73024
rect 155218 72972 155224 73024
rect 155276 73012 155282 73024
rect 155402 73012 155408 73024
rect 155276 72984 155408 73012
rect 155276 72972 155282 72984
rect 155402 72972 155408 72984
rect 155460 73012 155466 73024
rect 189994 73012 190000 73024
rect 155460 72984 190000 73012
rect 155460 72972 155466 72984
rect 189994 72972 190000 72984
rect 190052 72972 190058 73024
rect 105722 72904 105728 72956
rect 105780 72944 105786 72956
rect 139302 72944 139308 72956
rect 105780 72916 139308 72944
rect 105780 72904 105786 72916
rect 139302 72904 139308 72916
rect 139360 72904 139366 72956
rect 163682 72904 163688 72956
rect 163740 72944 163746 72956
rect 198182 72944 198188 72956
rect 163740 72916 198188 72944
rect 163740 72904 163746 72916
rect 198182 72904 198188 72916
rect 198240 72904 198246 72956
rect 108666 72836 108672 72888
rect 108724 72876 108730 72888
rect 140590 72876 140596 72888
rect 108724 72848 140596 72876
rect 108724 72836 108730 72848
rect 140590 72836 140596 72848
rect 140648 72836 140654 72888
rect 159634 72836 159640 72888
rect 159692 72876 159698 72888
rect 189810 72876 189816 72888
rect 159692 72848 189816 72876
rect 159692 72836 159698 72848
rect 189810 72836 189816 72848
rect 189868 72836 189874 72888
rect 111242 72768 111248 72820
rect 111300 72808 111306 72820
rect 142798 72808 142804 72820
rect 111300 72780 142804 72808
rect 111300 72768 111306 72780
rect 142798 72768 142804 72780
rect 142856 72768 142862 72820
rect 146662 72768 146668 72820
rect 146720 72808 146726 72820
rect 180334 72808 180340 72820
rect 146720 72780 180340 72808
rect 146720 72768 146726 72780
rect 180334 72768 180340 72780
rect 180392 72768 180398 72820
rect 181990 72768 181996 72820
rect 182048 72808 182054 72820
rect 204254 72808 204260 72820
rect 182048 72780 204260 72808
rect 182048 72768 182054 72780
rect 204254 72768 204260 72780
rect 204312 72768 204318 72820
rect 209746 72808 209774 73120
rect 327718 73108 327724 73160
rect 327776 73148 327782 73160
rect 579982 73148 579988 73160
rect 327776 73120 579988 73148
rect 327776 73108 327782 73120
rect 579982 73108 579988 73120
rect 580040 73108 580046 73160
rect 220078 72808 220084 72820
rect 209746 72780 220084 72808
rect 220078 72768 220084 72780
rect 220136 72768 220142 72820
rect 111426 72700 111432 72752
rect 111484 72740 111490 72752
rect 143074 72740 143080 72752
rect 111484 72712 143080 72740
rect 111484 72700 111490 72712
rect 143074 72700 143080 72712
rect 143132 72700 143138 72752
rect 156598 72700 156604 72752
rect 156656 72740 156662 72752
rect 311158 72740 311164 72752
rect 156656 72712 311164 72740
rect 156656 72700 156662 72712
rect 311158 72700 311164 72712
rect 311216 72700 311222 72752
rect 85574 72632 85580 72684
rect 85632 72672 85638 72684
rect 105722 72672 105728 72684
rect 85632 72644 105728 72672
rect 85632 72632 85638 72644
rect 105722 72632 105728 72644
rect 105780 72632 105786 72684
rect 119798 72632 119804 72684
rect 119856 72672 119862 72684
rect 144362 72672 144368 72684
rect 119856 72644 144368 72672
rect 119856 72632 119862 72644
rect 144362 72632 144368 72644
rect 144420 72632 144426 72684
rect 157242 72632 157248 72684
rect 157300 72672 157306 72684
rect 318794 72672 318800 72684
rect 157300 72644 318800 72672
rect 157300 72632 157306 72644
rect 318794 72632 318800 72644
rect 318852 72632 318858 72684
rect 43438 72564 43444 72616
rect 43496 72604 43502 72616
rect 102134 72604 102140 72616
rect 43496 72576 102140 72604
rect 43496 72564 43502 72576
rect 102134 72564 102140 72576
rect 102192 72564 102198 72616
rect 122098 72564 122104 72616
rect 122156 72604 122162 72616
rect 123018 72604 123024 72616
rect 122156 72576 123024 72604
rect 122156 72564 122162 72576
rect 123018 72564 123024 72576
rect 123076 72564 123082 72616
rect 124214 72564 124220 72616
rect 124272 72604 124278 72616
rect 140774 72604 140780 72616
rect 124272 72576 140780 72604
rect 124272 72564 124278 72576
rect 140774 72564 140780 72576
rect 140832 72564 140838 72616
rect 157794 72564 157800 72616
rect 157852 72604 157858 72616
rect 324958 72604 324964 72616
rect 157852 72576 324964 72604
rect 157852 72564 157858 72576
rect 324958 72564 324964 72576
rect 325016 72564 325022 72616
rect 67634 72496 67640 72548
rect 67692 72536 67698 72548
rect 137738 72536 137744 72548
rect 67692 72508 137744 72536
rect 67692 72496 67698 72508
rect 137738 72496 137744 72508
rect 137796 72496 137802 72548
rect 158254 72496 158260 72548
rect 158312 72536 158318 72548
rect 332594 72536 332600 72548
rect 158312 72508 332600 72536
rect 158312 72496 158318 72508
rect 332594 72496 332600 72508
rect 332652 72496 332658 72548
rect 14458 72428 14464 72480
rect 14516 72468 14522 72480
rect 14516 72440 103514 72468
rect 14516 72428 14522 72440
rect 103486 72400 103514 72440
rect 111610 72428 111616 72480
rect 111668 72468 111674 72480
rect 130010 72468 130016 72480
rect 111668 72440 130016 72468
rect 111668 72428 111674 72440
rect 130010 72428 130016 72440
rect 130068 72468 130074 72480
rect 131022 72468 131028 72480
rect 130068 72440 131028 72468
rect 130068 72428 130074 72440
rect 131022 72428 131028 72440
rect 131080 72428 131086 72480
rect 132494 72428 132500 72480
rect 132552 72468 132558 72480
rect 133506 72468 133512 72480
rect 132552 72440 133512 72468
rect 132552 72428 132558 72440
rect 133506 72428 133512 72440
rect 133564 72428 133570 72480
rect 167086 72428 167092 72480
rect 167144 72468 167150 72480
rect 168374 72468 168380 72480
rect 167144 72440 168380 72468
rect 167144 72428 167150 72440
rect 168374 72428 168380 72440
rect 168432 72428 168438 72480
rect 168650 72428 168656 72480
rect 168708 72468 168714 72480
rect 375374 72468 375380 72480
rect 168708 72440 375380 72468
rect 168708 72428 168714 72440
rect 375374 72428 375380 72440
rect 375432 72428 375438 72480
rect 104526 72400 104532 72412
rect 103486 72372 104532 72400
rect 104526 72360 104532 72372
rect 104584 72400 104590 72412
rect 129090 72400 129096 72412
rect 104584 72372 129096 72400
rect 104584 72360 104590 72372
rect 129090 72360 129096 72372
rect 129148 72360 129154 72412
rect 161658 72360 161664 72412
rect 161716 72400 161722 72412
rect 179690 72400 179696 72412
rect 161716 72372 179696 72400
rect 161716 72360 161722 72372
rect 179690 72360 179696 72372
rect 179748 72400 179754 72412
rect 180610 72400 180616 72412
rect 179748 72372 180616 72400
rect 179748 72360 179754 72372
rect 180610 72360 180616 72372
rect 180668 72360 180674 72412
rect 171502 72292 171508 72344
rect 171560 72332 171566 72344
rect 172238 72332 172244 72344
rect 171560 72304 172244 72332
rect 171560 72292 171566 72304
rect 172238 72292 172244 72304
rect 172296 72292 172302 72344
rect 178402 72292 178408 72344
rect 178460 72332 178466 72344
rect 181990 72332 181996 72344
rect 178460 72304 181996 72332
rect 178460 72292 178466 72304
rect 181990 72292 181996 72304
rect 182048 72292 182054 72344
rect 156414 72224 156420 72276
rect 156472 72264 156478 72276
rect 181254 72264 181260 72276
rect 156472 72236 181260 72264
rect 156472 72224 156478 72236
rect 181254 72224 181260 72236
rect 181312 72224 181318 72276
rect 152274 72088 152280 72140
rect 152332 72128 152338 72140
rect 152734 72128 152740 72140
rect 152332 72100 152740 72128
rect 152332 72088 152338 72100
rect 152734 72088 152740 72100
rect 152792 72088 152798 72140
rect 160186 72020 160192 72072
rect 160244 72060 160250 72072
rect 160554 72060 160560 72072
rect 160244 72032 160560 72060
rect 160244 72020 160250 72032
rect 160554 72020 160560 72032
rect 160612 72020 160618 72072
rect 181254 71816 181260 71868
rect 181312 71856 181318 71868
rect 304258 71856 304264 71868
rect 181312 71828 304264 71856
rect 181312 71816 181318 71828
rect 304258 71816 304264 71828
rect 304316 71816 304322 71868
rect 107654 71748 107660 71800
rect 107712 71788 107718 71800
rect 108666 71788 108672 71800
rect 107712 71760 108672 71788
rect 107712 71748 107718 71760
rect 108666 71748 108672 71760
rect 108724 71748 108730 71800
rect 161768 71760 162716 71788
rect 118326 71680 118332 71732
rect 118384 71720 118390 71732
rect 151906 71720 151912 71732
rect 118384 71692 151912 71720
rect 118384 71680 118390 71692
rect 151906 71680 151912 71692
rect 151964 71720 151970 71732
rect 152642 71720 152648 71732
rect 151964 71692 152648 71720
rect 151964 71680 151970 71692
rect 152642 71680 152648 71692
rect 152700 71680 152706 71732
rect 157702 71680 157708 71732
rect 157760 71720 157766 71732
rect 158070 71720 158076 71732
rect 157760 71692 158076 71720
rect 157760 71680 157766 71692
rect 158070 71680 158076 71692
rect 158128 71680 158134 71732
rect 158346 71680 158352 71732
rect 158404 71720 158410 71732
rect 158622 71720 158628 71732
rect 158404 71692 158628 71720
rect 158404 71680 158410 71692
rect 158622 71680 158628 71692
rect 158680 71680 158686 71732
rect 159082 71680 159088 71732
rect 159140 71720 159146 71732
rect 159910 71720 159916 71732
rect 159140 71692 159916 71720
rect 159140 71680 159146 71692
rect 159910 71680 159916 71692
rect 159968 71680 159974 71732
rect 161768 71720 161796 71760
rect 161676 71692 161796 71720
rect 3510 71612 3516 71664
rect 3568 71652 3574 71664
rect 8938 71652 8944 71664
rect 3568 71624 8944 71652
rect 3568 71612 3574 71624
rect 8938 71612 8944 71624
rect 8996 71612 9002 71664
rect 116302 71612 116308 71664
rect 116360 71652 116366 71664
rect 151170 71652 151176 71664
rect 116360 71624 151176 71652
rect 116360 71612 116366 71624
rect 151170 71612 151176 71624
rect 151228 71612 151234 71664
rect 159542 71612 159548 71664
rect 159600 71652 159606 71664
rect 161676 71652 161704 71692
rect 159600 71624 161704 71652
rect 159600 71612 159606 71624
rect 161750 71612 161756 71664
rect 161808 71652 161814 71664
rect 162578 71652 162584 71664
rect 161808 71624 162584 71652
rect 161808 71612 161814 71624
rect 162578 71612 162584 71624
rect 162636 71612 162642 71664
rect 162688 71652 162716 71760
rect 180610 71748 180616 71800
rect 180668 71788 180674 71800
rect 322934 71788 322940 71800
rect 180668 71760 322940 71788
rect 180668 71748 180674 71760
rect 322934 71748 322940 71760
rect 322992 71748 322998 71800
rect 183554 71680 183560 71732
rect 183612 71720 183618 71732
rect 204714 71720 204720 71732
rect 183612 71692 204720 71720
rect 183612 71680 183618 71692
rect 204714 71680 204720 71692
rect 204772 71680 204778 71732
rect 194318 71652 194324 71664
rect 162688 71624 194324 71652
rect 194318 71612 194324 71624
rect 194376 71612 194382 71664
rect 121178 71544 121184 71596
rect 121236 71584 121242 71596
rect 152458 71584 152464 71596
rect 121236 71556 152464 71584
rect 121236 71544 121242 71556
rect 152458 71544 152464 71556
rect 152516 71544 152522 71596
rect 161106 71544 161112 71596
rect 161164 71584 161170 71596
rect 195146 71584 195152 71596
rect 161164 71556 195152 71584
rect 161164 71544 161170 71556
rect 195146 71544 195152 71556
rect 195204 71544 195210 71596
rect 102134 71476 102140 71528
rect 102192 71516 102198 71528
rect 102962 71516 102968 71528
rect 102192 71488 102968 71516
rect 102192 71476 102198 71488
rect 102962 71476 102968 71488
rect 103020 71516 103026 71528
rect 134702 71516 134708 71528
rect 103020 71488 134708 71516
rect 103020 71476 103026 71488
rect 134702 71476 134708 71488
rect 134760 71476 134766 71528
rect 135438 71476 135444 71528
rect 135496 71516 135502 71528
rect 136542 71516 136548 71528
rect 135496 71488 136548 71516
rect 135496 71476 135502 71488
rect 136542 71476 136548 71488
rect 136600 71476 136606 71528
rect 141418 71476 141424 71528
rect 141476 71516 141482 71528
rect 142798 71516 142804 71528
rect 141476 71488 142804 71516
rect 141476 71476 141482 71488
rect 142798 71476 142804 71488
rect 142856 71476 142862 71528
rect 160370 71476 160376 71528
rect 160428 71516 160434 71528
rect 162118 71516 162124 71528
rect 160428 71488 162124 71516
rect 160428 71476 160434 71488
rect 162118 71476 162124 71488
rect 162176 71476 162182 71528
rect 162578 71476 162584 71528
rect 162636 71516 162642 71528
rect 196802 71516 196808 71528
rect 162636 71488 196808 71516
rect 162636 71476 162642 71488
rect 196802 71476 196808 71488
rect 196860 71476 196866 71528
rect 112162 71408 112168 71460
rect 112220 71448 112226 71460
rect 142430 71448 142436 71460
rect 112220 71420 142436 71448
rect 112220 71408 112226 71420
rect 142430 71408 142436 71420
rect 142488 71448 142494 71460
rect 143258 71448 143264 71460
rect 142488 71420 143264 71448
rect 142488 71408 142494 71420
rect 143258 71408 143264 71420
rect 143316 71408 143322 71460
rect 159910 71408 159916 71460
rect 159968 71448 159974 71460
rect 193858 71448 193864 71460
rect 159968 71420 193864 71448
rect 159968 71408 159974 71420
rect 193858 71408 193864 71420
rect 193916 71408 193922 71460
rect 105630 71340 105636 71392
rect 105688 71380 105694 71392
rect 135438 71380 135444 71392
rect 105688 71352 135444 71380
rect 105688 71340 105694 71352
rect 135438 71340 135444 71352
rect 135496 71340 135502 71392
rect 142798 71340 142804 71392
rect 142856 71380 142862 71392
rect 143166 71380 143172 71392
rect 142856 71352 143172 71380
rect 142856 71340 142862 71352
rect 143166 71340 143172 71352
rect 143224 71340 143230 71392
rect 161566 71340 161572 71392
rect 161624 71380 161630 71392
rect 196894 71380 196900 71392
rect 161624 71352 196900 71380
rect 161624 71340 161630 71352
rect 196894 71340 196900 71352
rect 196952 71340 196958 71392
rect 107470 71272 107476 71324
rect 107528 71312 107534 71324
rect 135714 71312 135720 71324
rect 107528 71284 135720 71312
rect 107528 71272 107534 71284
rect 135714 71272 135720 71284
rect 135772 71272 135778 71324
rect 142154 71312 142160 71324
rect 137986 71284 142160 71312
rect 102778 71204 102784 71256
rect 102836 71244 102842 71256
rect 106734 71244 106740 71256
rect 102836 71216 106740 71244
rect 102836 71204 102842 71216
rect 106734 71204 106740 71216
rect 106792 71204 106798 71256
rect 53834 71136 53840 71188
rect 53892 71176 53898 71188
rect 107488 71176 107516 71272
rect 113542 71204 113548 71256
rect 113600 71244 113606 71256
rect 137986 71244 138014 71284
rect 142154 71272 142160 71284
rect 142212 71312 142218 71324
rect 143442 71312 143448 71324
rect 142212 71284 143448 71312
rect 142212 71272 142218 71284
rect 143442 71272 143448 71284
rect 143500 71272 143506 71324
rect 172422 71272 172428 71324
rect 172480 71312 172486 71324
rect 200390 71312 200396 71324
rect 172480 71284 200396 71312
rect 172480 71272 172486 71284
rect 200390 71272 200396 71284
rect 200448 71272 200454 71324
rect 113600 71216 138014 71244
rect 113600 71204 113606 71216
rect 158990 71204 158996 71256
rect 159048 71244 159054 71256
rect 193490 71244 193496 71256
rect 159048 71216 193496 71244
rect 159048 71204 159054 71216
rect 193490 71204 193496 71216
rect 193548 71244 193554 71256
rect 193548 71216 200114 71244
rect 193548 71204 193554 71216
rect 53892 71148 107516 71176
rect 53892 71136 53898 71148
rect 112530 71136 112536 71188
rect 112588 71176 112594 71188
rect 138014 71176 138020 71188
rect 112588 71148 138020 71176
rect 112588 71136 112594 71148
rect 138014 71136 138020 71148
rect 138072 71176 138078 71188
rect 139118 71176 139124 71188
rect 138072 71148 139124 71176
rect 138072 71136 138078 71148
rect 139118 71136 139124 71148
rect 139176 71136 139182 71188
rect 142982 71136 142988 71188
rect 143040 71176 143046 71188
rect 143442 71176 143448 71188
rect 143040 71148 143448 71176
rect 143040 71136 143046 71148
rect 143442 71136 143448 71148
rect 143500 71136 143506 71188
rect 158622 71136 158628 71188
rect 158680 71176 158686 71188
rect 191190 71176 191196 71188
rect 158680 71148 191196 71176
rect 158680 71136 158686 71148
rect 191190 71136 191196 71148
rect 191248 71136 191254 71188
rect 31018 71068 31024 71120
rect 31076 71108 31082 71120
rect 102134 71108 102140 71120
rect 31076 71080 102140 71108
rect 31076 71068 31082 71080
rect 102134 71068 102140 71080
rect 102192 71068 102198 71120
rect 116210 71068 116216 71120
rect 116268 71108 116274 71120
rect 128354 71108 128360 71120
rect 116268 71080 128360 71108
rect 116268 71068 116274 71080
rect 128354 71068 128360 71080
rect 128412 71108 128418 71120
rect 129550 71108 129556 71120
rect 128412 71080 129556 71108
rect 128412 71068 128418 71080
rect 129550 71068 129556 71080
rect 129608 71068 129614 71120
rect 158438 71068 158444 71120
rect 158496 71108 158502 71120
rect 191098 71108 191104 71120
rect 158496 71080 191104 71108
rect 158496 71068 158502 71080
rect 191098 71068 191104 71080
rect 191156 71068 191162 71120
rect 200086 71108 200114 71216
rect 204714 71136 204720 71188
rect 204772 71176 204778 71188
rect 217318 71176 217324 71188
rect 204772 71148 217324 71176
rect 204772 71136 204778 71148
rect 217318 71136 217324 71148
rect 217376 71136 217382 71188
rect 335998 71108 336004 71120
rect 200086 71080 336004 71108
rect 335998 71068 336004 71080
rect 336056 71068 336062 71120
rect 31754 71000 31760 71052
rect 31812 71040 31818 71052
rect 133414 71040 133420 71052
rect 31812 71012 133420 71040
rect 31812 71000 31818 71012
rect 133414 71000 133420 71012
rect 133472 71000 133478 71052
rect 160830 71000 160836 71052
rect 160888 71040 160894 71052
rect 192570 71040 192576 71052
rect 160888 71012 192576 71040
rect 160888 71000 160894 71012
rect 192570 71000 192576 71012
rect 192628 71040 192634 71052
rect 367094 71040 367100 71052
rect 192628 71012 367100 71040
rect 192628 71000 192634 71012
rect 367094 71000 367100 71012
rect 367152 71000 367158 71052
rect 174906 70932 174912 70984
rect 174964 70972 174970 70984
rect 204346 70972 204352 70984
rect 174964 70944 204352 70972
rect 174964 70932 174970 70944
rect 204346 70932 204352 70944
rect 204404 70932 204410 70984
rect 162578 70864 162584 70916
rect 162636 70904 162642 70916
rect 186406 70904 186412 70916
rect 162636 70876 186412 70904
rect 162636 70864 162642 70876
rect 186406 70864 186412 70876
rect 186464 70864 186470 70916
rect 158070 70796 158076 70848
rect 158128 70836 158134 70848
rect 192754 70836 192760 70848
rect 158128 70808 192760 70836
rect 158128 70796 158134 70808
rect 192754 70796 192760 70808
rect 192812 70796 192818 70848
rect 159634 70456 159640 70508
rect 159692 70496 159698 70508
rect 160002 70496 160008 70508
rect 159692 70468 160008 70496
rect 159692 70456 159698 70468
rect 160002 70456 160008 70468
rect 160060 70456 160066 70508
rect 168374 70388 168380 70440
rect 168432 70428 168438 70440
rect 169110 70428 169116 70440
rect 168432 70400 169116 70428
rect 168432 70388 168438 70400
rect 169110 70388 169116 70400
rect 169168 70388 169174 70440
rect 192110 70388 192116 70440
rect 192168 70428 192174 70440
rect 192294 70428 192300 70440
rect 192168 70400 192300 70428
rect 192168 70388 192174 70400
rect 192294 70388 192300 70400
rect 192352 70388 192358 70440
rect 100294 70320 100300 70372
rect 100352 70360 100358 70372
rect 134150 70360 134156 70372
rect 100352 70332 134156 70360
rect 100352 70320 100358 70332
rect 134150 70320 134156 70332
rect 134208 70320 134214 70372
rect 166718 70320 166724 70372
rect 166776 70360 166782 70372
rect 200666 70360 200672 70372
rect 166776 70332 200672 70360
rect 166776 70320 166782 70332
rect 200666 70320 200672 70332
rect 200724 70320 200730 70372
rect 102134 70252 102140 70304
rect 102192 70292 102198 70304
rect 103054 70292 103060 70304
rect 102192 70264 103060 70292
rect 102192 70252 102198 70264
rect 103054 70252 103060 70264
rect 103112 70292 103118 70304
rect 137002 70292 137008 70304
rect 103112 70264 137008 70292
rect 103112 70252 103118 70264
rect 137002 70252 137008 70264
rect 137060 70252 137066 70304
rect 165246 70252 165252 70304
rect 165304 70292 165310 70304
rect 199378 70292 199384 70304
rect 165304 70264 199384 70292
rect 165304 70252 165310 70264
rect 199378 70252 199384 70264
rect 199436 70252 199442 70304
rect 105906 70184 105912 70236
rect 105964 70224 105970 70236
rect 139578 70224 139584 70236
rect 105964 70196 139584 70224
rect 105964 70184 105970 70196
rect 139578 70184 139584 70196
rect 139636 70184 139642 70236
rect 165706 70184 165712 70236
rect 165764 70224 165770 70236
rect 166350 70224 166356 70236
rect 165764 70196 166356 70224
rect 165764 70184 165770 70196
rect 166350 70184 166356 70196
rect 166408 70224 166414 70236
rect 200482 70224 200488 70236
rect 166408 70196 200488 70224
rect 166408 70184 166414 70196
rect 200482 70184 200488 70196
rect 200540 70184 200546 70236
rect 100386 70116 100392 70168
rect 100444 70156 100450 70168
rect 132494 70156 132500 70168
rect 100444 70128 132500 70156
rect 100444 70116 100450 70128
rect 132494 70116 132500 70128
rect 132552 70116 132558 70168
rect 165522 70116 165528 70168
rect 165580 70156 165586 70168
rect 199746 70156 199752 70168
rect 165580 70128 199752 70156
rect 165580 70116 165586 70128
rect 199746 70116 199752 70128
rect 199804 70116 199810 70168
rect 102226 70048 102232 70100
rect 102284 70088 102290 70100
rect 103238 70088 103244 70100
rect 102284 70060 103244 70088
rect 102284 70048 102290 70060
rect 103238 70048 103244 70060
rect 103296 70088 103302 70100
rect 133598 70088 133604 70100
rect 103296 70060 133604 70088
rect 103296 70048 103302 70060
rect 133598 70048 133604 70060
rect 133656 70048 133662 70100
rect 164050 70048 164056 70100
rect 164108 70088 164114 70100
rect 197722 70088 197728 70100
rect 164108 70060 197728 70088
rect 164108 70048 164114 70060
rect 197722 70048 197728 70060
rect 197780 70048 197786 70100
rect 116762 69980 116768 70032
rect 116820 70020 116826 70032
rect 138198 70020 138204 70032
rect 116820 69992 138204 70020
rect 116820 69980 116826 69992
rect 138198 69980 138204 69992
rect 138256 69980 138262 70032
rect 164602 69980 164608 70032
rect 164660 70020 164666 70032
rect 199010 70020 199016 70032
rect 164660 69992 199016 70020
rect 164660 69980 164666 69992
rect 199010 69980 199016 69992
rect 199068 69980 199074 70032
rect 164510 69912 164516 69964
rect 164568 69952 164574 69964
rect 165246 69952 165252 69964
rect 164568 69924 165252 69952
rect 164568 69912 164574 69924
rect 165246 69912 165252 69924
rect 165304 69912 165310 69964
rect 196526 69952 196532 69964
rect 166092 69924 196532 69952
rect 62114 69844 62120 69896
rect 62172 69884 62178 69896
rect 102134 69884 102140 69896
rect 62172 69856 102140 69884
rect 62172 69844 62178 69856
rect 102134 69844 102140 69856
rect 102192 69844 102198 69896
rect 103514 69844 103520 69896
rect 103572 69884 103578 69896
rect 105906 69884 105912 69896
rect 103572 69856 105912 69884
rect 103572 69844 103578 69856
rect 105906 69844 105912 69856
rect 105964 69844 105970 69896
rect 163130 69844 163136 69896
rect 163188 69884 163194 69896
rect 163958 69884 163964 69896
rect 163188 69856 163964 69884
rect 163188 69844 163194 69856
rect 163958 69844 163964 69856
rect 164016 69884 164022 69896
rect 164016 69856 164648 69884
rect 164016 69844 164022 69856
rect 85666 69776 85672 69828
rect 85724 69816 85730 69828
rect 138106 69816 138112 69828
rect 85724 69788 138112 69816
rect 85724 69776 85730 69788
rect 138106 69776 138112 69788
rect 138164 69776 138170 69828
rect 163222 69776 163228 69828
rect 163280 69816 163286 69828
rect 164050 69816 164056 69828
rect 163280 69788 164056 69816
rect 163280 69776 163286 69788
rect 164050 69776 164056 69788
rect 164108 69776 164114 69828
rect 164620 69816 164648 69856
rect 164694 69844 164700 69896
rect 164752 69884 164758 69896
rect 165522 69884 165528 69896
rect 164752 69856 165528 69884
rect 164752 69844 164758 69856
rect 165522 69844 165528 69856
rect 165580 69844 165586 69896
rect 166092 69816 166120 69924
rect 196526 69912 196532 69924
rect 196584 69912 196590 69964
rect 168926 69844 168932 69896
rect 168984 69884 168990 69896
rect 169386 69884 169392 69896
rect 168984 69856 169392 69884
rect 168984 69844 168990 69856
rect 169386 69844 169392 69856
rect 169444 69844 169450 69896
rect 171042 69844 171048 69896
rect 171100 69884 171106 69896
rect 199102 69884 199108 69896
rect 171100 69856 199108 69884
rect 171100 69844 171106 69856
rect 199102 69844 199108 69856
rect 199160 69844 199166 69896
rect 164620 69788 166120 69816
rect 167270 69776 167276 69828
rect 167328 69816 167334 69828
rect 354674 69816 354680 69828
rect 167328 69788 354680 69816
rect 167328 69776 167334 69788
rect 354674 69776 354680 69788
rect 354732 69776 354738 69828
rect 18598 69708 18604 69760
rect 18656 69748 18662 69760
rect 102226 69748 102232 69760
rect 18656 69720 102232 69748
rect 18656 69708 18662 69720
rect 102226 69708 102232 69720
rect 102284 69708 102290 69760
rect 147122 69708 147128 69760
rect 147180 69748 147186 69760
rect 185578 69748 185584 69760
rect 147180 69720 185584 69748
rect 147180 69708 147186 69720
rect 185578 69708 185584 69720
rect 185636 69708 185642 69760
rect 199010 69708 199016 69760
rect 199068 69748 199074 69760
rect 199286 69748 199292 69760
rect 199068 69720 199292 69748
rect 199068 69708 199074 69720
rect 199286 69708 199292 69720
rect 199344 69748 199350 69760
rect 412634 69748 412640 69760
rect 199344 69720 412640 69748
rect 199344 69708 199350 69720
rect 412634 69708 412640 69720
rect 412692 69708 412698 69760
rect 45554 69640 45560 69692
rect 45612 69680 45618 69692
rect 135254 69680 135260 69692
rect 45612 69652 135260 69680
rect 45612 69640 45618 69652
rect 135254 69640 135260 69652
rect 135312 69640 135318 69692
rect 148226 69640 148232 69692
rect 148284 69680 148290 69692
rect 148284 69652 191880 69680
rect 148284 69640 148290 69652
rect 143994 69572 144000 69624
rect 144052 69612 144058 69624
rect 147122 69612 147128 69624
rect 144052 69584 147128 69612
rect 144052 69572 144058 69584
rect 147122 69572 147128 69584
rect 147180 69572 147186 69624
rect 168742 69572 168748 69624
rect 168800 69612 168806 69624
rect 169478 69612 169484 69624
rect 168800 69584 169484 69612
rect 168800 69572 168806 69584
rect 169478 69572 169484 69584
rect 169536 69572 169542 69624
rect 176930 69572 176936 69624
rect 176988 69612 176994 69624
rect 191852 69612 191880 69652
rect 191926 69640 191932 69692
rect 191984 69680 191990 69692
rect 192110 69680 192116 69692
rect 191984 69652 192116 69680
rect 191984 69640 191990 69652
rect 192110 69640 192116 69652
rect 192168 69640 192174 69692
rect 199102 69640 199108 69692
rect 199160 69680 199166 69692
rect 199654 69680 199660 69692
rect 199160 69652 199660 69680
rect 199160 69640 199166 69652
rect 199654 69640 199660 69652
rect 199712 69680 199718 69692
rect 498194 69680 498200 69692
rect 199712 69652 498200 69680
rect 199712 69640 199718 69652
rect 498194 69640 498200 69652
rect 498252 69640 498258 69692
rect 196618 69612 196624 69624
rect 176988 69584 180794 69612
rect 191852 69584 196624 69612
rect 176988 69572 176994 69584
rect 146386 69504 146392 69556
rect 146444 69544 146450 69556
rect 179414 69544 179420 69556
rect 146444 69516 179420 69544
rect 146444 69504 146450 69516
rect 179414 69504 179420 69516
rect 179472 69504 179478 69556
rect 180766 69544 180794 69584
rect 196618 69572 196624 69584
rect 196676 69572 196682 69624
rect 195146 69544 195152 69556
rect 180766 69516 195152 69544
rect 195146 69504 195152 69516
rect 195204 69504 195210 69556
rect 153746 69368 153752 69420
rect 153804 69408 153810 69420
rect 181162 69408 181168 69420
rect 153804 69380 181168 69408
rect 153804 69368 153810 69380
rect 181162 69368 181168 69380
rect 181220 69368 181226 69420
rect 195146 69028 195152 69080
rect 195204 69068 195210 69080
rect 529934 69068 529940 69080
rect 195204 69040 529940 69068
rect 195204 69028 195210 69040
rect 529934 69028 529940 69040
rect 529992 69028 529998 69080
rect 116118 68960 116124 69012
rect 116176 69000 116182 69012
rect 116176 68972 144408 69000
rect 116176 68960 116182 68972
rect 118510 68892 118516 68944
rect 118568 68932 118574 68944
rect 118568 68904 144316 68932
rect 118568 68892 118574 68904
rect 105998 68824 106004 68876
rect 106056 68864 106062 68876
rect 138658 68864 138664 68876
rect 106056 68836 138664 68864
rect 106056 68824 106062 68836
rect 138658 68824 138664 68836
rect 138716 68824 138722 68876
rect 140774 68824 140780 68876
rect 140832 68864 140838 68876
rect 142154 68864 142160 68876
rect 140832 68836 142160 68864
rect 140832 68824 140838 68836
rect 142154 68824 142160 68836
rect 142212 68824 142218 68876
rect 110230 68756 110236 68808
rect 110288 68796 110294 68808
rect 142246 68796 142252 68808
rect 110288 68768 142252 68796
rect 110288 68756 110294 68768
rect 142246 68756 142252 68768
rect 142304 68796 142310 68808
rect 142706 68796 142712 68808
rect 142304 68768 142712 68796
rect 142304 68756 142310 68768
rect 142706 68756 142712 68768
rect 142764 68756 142770 68808
rect 144288 68796 144316 68904
rect 144380 68864 144408 68972
rect 144454 68960 144460 69012
rect 144512 69000 144518 69012
rect 146294 69000 146300 69012
rect 144512 68972 146300 69000
rect 144512 68960 144518 68972
rect 146294 68960 146300 68972
rect 146352 68960 146358 69012
rect 150618 68960 150624 69012
rect 150676 69000 150682 69012
rect 151170 69000 151176 69012
rect 150676 68972 151176 69000
rect 150676 68960 150682 68972
rect 151170 68960 151176 68972
rect 151228 68960 151234 69012
rect 167362 68960 167368 69012
rect 167420 69000 167426 69012
rect 168006 69000 168012 69012
rect 167420 68972 168012 69000
rect 167420 68960 167426 68972
rect 168006 68960 168012 68972
rect 168064 69000 168070 69012
rect 201954 69000 201960 69012
rect 168064 68972 201960 69000
rect 168064 68960 168070 68972
rect 201954 68960 201960 68972
rect 202012 68960 202018 69012
rect 152550 68932 152556 68944
rect 151786 68904 152556 68932
rect 150618 68864 150624 68876
rect 144380 68836 150624 68864
rect 150618 68824 150624 68836
rect 150676 68824 150682 68876
rect 151786 68796 151814 68904
rect 152550 68892 152556 68904
rect 152608 68892 152614 68944
rect 161750 68892 161756 68944
rect 161808 68932 161814 68944
rect 162486 68932 162492 68944
rect 161808 68904 162492 68932
rect 161808 68892 161814 68904
rect 162486 68892 162492 68904
rect 162544 68892 162550 68944
rect 168834 68892 168840 68944
rect 168892 68932 168898 68944
rect 169570 68932 169576 68944
rect 168892 68904 169576 68932
rect 168892 68892 168898 68904
rect 169570 68892 169576 68904
rect 169628 68932 169634 68944
rect 203610 68932 203616 68944
rect 169628 68904 203616 68932
rect 169628 68892 169634 68904
rect 203610 68892 203616 68904
rect 203668 68892 203674 68944
rect 161566 68824 161572 68876
rect 161624 68864 161630 68876
rect 162394 68864 162400 68876
rect 161624 68836 162400 68864
rect 161624 68824 161630 68836
rect 162394 68824 162400 68836
rect 162452 68824 162458 68876
rect 169478 68824 169484 68876
rect 169536 68864 169542 68876
rect 203426 68864 203432 68876
rect 169536 68836 203432 68864
rect 169536 68824 169542 68836
rect 203426 68824 203432 68836
rect 203484 68824 203490 68876
rect 144288 68768 151814 68796
rect 169386 68756 169392 68808
rect 169444 68796 169450 68808
rect 203518 68796 203524 68808
rect 169444 68768 203524 68796
rect 169444 68756 169450 68768
rect 203518 68756 203524 68768
rect 203576 68756 203582 68808
rect 104434 68688 104440 68740
rect 104492 68728 104498 68740
rect 104618 68728 104624 68740
rect 104492 68700 104624 68728
rect 104492 68688 104498 68700
rect 104618 68688 104624 68700
rect 104676 68728 104682 68740
rect 135714 68728 135720 68740
rect 104676 68700 135720 68728
rect 104676 68688 104682 68700
rect 135714 68688 135720 68700
rect 135772 68688 135778 68740
rect 183830 68688 183836 68740
rect 183888 68728 183894 68740
rect 203058 68728 203064 68740
rect 183888 68700 203064 68728
rect 183888 68688 183894 68700
rect 203058 68688 203064 68700
rect 203116 68728 203122 68740
rect 204162 68728 204168 68740
rect 203116 68700 204168 68728
rect 203116 68688 203122 68700
rect 204162 68688 204168 68700
rect 204220 68688 204226 68740
rect 114278 68620 114284 68672
rect 114336 68660 114342 68672
rect 142338 68660 142344 68672
rect 114336 68632 142344 68660
rect 114336 68620 114342 68632
rect 142338 68620 142344 68632
rect 142396 68660 142402 68672
rect 142890 68660 142896 68672
rect 142396 68632 142896 68660
rect 142396 68620 142402 68632
rect 142890 68620 142896 68632
rect 142948 68620 142954 68672
rect 163038 68620 163044 68672
rect 163096 68660 163102 68672
rect 188246 68660 188252 68672
rect 163096 68632 188252 68660
rect 163096 68620 163102 68632
rect 188246 68620 188252 68632
rect 188304 68620 188310 68672
rect 111150 68552 111156 68604
rect 111208 68592 111214 68604
rect 112254 68592 112260 68604
rect 111208 68564 112260 68592
rect 111208 68552 111214 68564
rect 112254 68552 112260 68564
rect 112312 68552 112318 68604
rect 180702 68552 180708 68604
rect 180760 68592 180766 68604
rect 182174 68592 182180 68604
rect 180760 68564 182180 68592
rect 180760 68552 180766 68564
rect 182174 68552 182180 68564
rect 182232 68552 182238 68604
rect 201402 68592 201408 68604
rect 190426 68564 201408 68592
rect 176746 68484 176752 68536
rect 176804 68524 176810 68536
rect 190426 68524 190454 68564
rect 201402 68552 201408 68564
rect 201460 68552 201466 68604
rect 176804 68496 190454 68524
rect 176804 68484 176810 68496
rect 120074 68416 120080 68468
rect 120132 68456 120138 68468
rect 141602 68456 141608 68468
rect 120132 68428 141608 68456
rect 120132 68416 120138 68428
rect 141602 68416 141608 68428
rect 141660 68416 141666 68468
rect 89714 68348 89720 68400
rect 89772 68388 89778 68400
rect 105998 68388 106004 68400
rect 89772 68360 106004 68388
rect 89772 68348 89778 68360
rect 105998 68348 106004 68360
rect 106056 68348 106062 68400
rect 117314 68348 117320 68400
rect 117372 68388 117378 68400
rect 141142 68388 141148 68400
rect 117372 68360 141148 68388
rect 117372 68348 117378 68360
rect 141142 68348 141148 68360
rect 141200 68348 141206 68400
rect 48314 68280 48320 68332
rect 48372 68320 48378 68332
rect 104618 68320 104624 68332
rect 48372 68292 104624 68320
rect 48372 68280 48378 68292
rect 104618 68280 104624 68292
rect 104676 68280 104682 68332
rect 113174 68280 113180 68332
rect 113232 68320 113238 68332
rect 140958 68320 140964 68332
rect 113232 68292 140964 68320
rect 113232 68280 113238 68292
rect 140958 68280 140964 68292
rect 141016 68280 141022 68332
rect 204162 68280 204168 68332
rect 204220 68320 204226 68332
rect 464338 68320 464344 68332
rect 204220 68292 464344 68320
rect 204220 68280 204226 68292
rect 464338 68280 464344 68292
rect 464396 68280 464402 68332
rect 188246 67668 188252 67720
rect 188304 67708 188310 67720
rect 402974 67708 402980 67720
rect 188304 67680 402980 67708
rect 188304 67668 188310 67680
rect 402974 67668 402980 67680
rect 403032 67668 403038 67720
rect 201402 67600 201408 67652
rect 201460 67640 201466 67652
rect 552658 67640 552664 67652
rect 201460 67612 552664 67640
rect 201460 67600 201466 67612
rect 552658 67600 552664 67612
rect 552716 67600 552722 67652
rect 105998 67532 106004 67584
rect 106056 67572 106062 67584
rect 137094 67572 137100 67584
rect 106056 67544 137100 67572
rect 106056 67532 106062 67544
rect 137094 67532 137100 67544
rect 137152 67532 137158 67584
rect 146018 67532 146024 67584
rect 146076 67572 146082 67584
rect 148410 67572 148416 67584
rect 146076 67544 148416 67572
rect 146076 67532 146082 67544
rect 148410 67532 148416 67544
rect 148468 67532 148474 67584
rect 155126 67532 155132 67584
rect 155184 67572 155190 67584
rect 189166 67572 189172 67584
rect 155184 67544 189172 67572
rect 155184 67532 155190 67544
rect 189166 67532 189172 67544
rect 189224 67532 189230 67584
rect 104526 67464 104532 67516
rect 104584 67504 104590 67516
rect 134794 67504 134800 67516
rect 104584 67476 134800 67504
rect 104584 67464 104590 67476
rect 134794 67464 134800 67476
rect 134852 67464 134858 67516
rect 72418 66920 72424 66972
rect 72476 66960 72482 66972
rect 105998 66960 106004 66972
rect 72476 66932 106004 66960
rect 72476 66920 72482 66932
rect 105998 66920 106004 66932
rect 106056 66920 106062 66972
rect 35158 66852 35164 66904
rect 35216 66892 35222 66904
rect 104526 66892 104532 66904
rect 35216 66864 104532 66892
rect 35216 66852 35222 66864
rect 104526 66852 104532 66864
rect 104584 66852 104590 66904
rect 189166 66852 189172 66904
rect 189224 66892 189230 66904
rect 295334 66892 295340 66904
rect 189224 66864 295340 66892
rect 189224 66852 189230 66864
rect 295334 66852 295340 66864
rect 295392 66852 295398 66904
rect 102134 66172 102140 66224
rect 102192 66212 102198 66224
rect 103146 66212 103152 66224
rect 102192 66184 103152 66212
rect 102192 66172 102198 66184
rect 103146 66172 103152 66184
rect 103204 66212 103210 66224
rect 137186 66212 137192 66224
rect 103204 66184 137192 66212
rect 103204 66172 103210 66184
rect 137186 66172 137192 66184
rect 137244 66172 137250 66224
rect 157334 66172 157340 66224
rect 157392 66212 157398 66224
rect 192294 66212 192300 66224
rect 157392 66184 192300 66212
rect 157392 66172 157398 66184
rect 192294 66172 192300 66184
rect 192352 66212 192358 66224
rect 193122 66212 193128 66224
rect 192352 66184 193128 66212
rect 192352 66172 192358 66184
rect 193122 66172 193128 66184
rect 193180 66172 193186 66224
rect 159358 66104 159364 66156
rect 159416 66144 159422 66156
rect 188062 66144 188068 66156
rect 159416 66116 188068 66144
rect 159416 66104 159422 66116
rect 188062 66104 188068 66116
rect 188120 66104 188126 66156
rect 177114 66036 177120 66088
rect 177172 66076 177178 66088
rect 197538 66076 197544 66088
rect 177172 66048 197544 66076
rect 177172 66036 177178 66048
rect 197538 66036 197544 66048
rect 197596 66036 197602 66088
rect 148778 65560 148784 65612
rect 148836 65600 148842 65612
rect 207014 65600 207020 65612
rect 148836 65572 207020 65600
rect 148836 65560 148842 65572
rect 207014 65560 207020 65572
rect 207072 65560 207078 65612
rect 58618 65492 58624 65544
rect 58676 65532 58682 65544
rect 102134 65532 102140 65544
rect 58676 65504 102140 65532
rect 58676 65492 58682 65504
rect 102134 65492 102140 65504
rect 102192 65492 102198 65544
rect 193122 65492 193128 65544
rect 193180 65532 193186 65544
rect 324314 65532 324320 65544
rect 193180 65504 324320 65532
rect 193180 65492 193186 65504
rect 324314 65492 324320 65504
rect 324372 65492 324378 65544
rect 188614 64948 188620 65000
rect 188672 64988 188678 65000
rect 346394 64988 346400 65000
rect 188672 64960 346400 64988
rect 188672 64948 188678 64960
rect 346394 64948 346400 64960
rect 346452 64948 346458 65000
rect 197538 64880 197544 64932
rect 197596 64920 197602 64932
rect 574738 64920 574744 64932
rect 197596 64892 574744 64920
rect 197596 64880 197602 64892
rect 574738 64880 574744 64892
rect 574796 64880 574802 64932
rect 102134 64812 102140 64864
rect 102192 64852 102198 64864
rect 106090 64852 106096 64864
rect 102192 64824 106096 64852
rect 102192 64812 102198 64824
rect 106090 64812 106096 64824
rect 106148 64852 106154 64864
rect 139854 64852 139860 64864
rect 106148 64824 139860 64852
rect 106148 64812 106154 64824
rect 139854 64812 139860 64824
rect 139912 64812 139918 64864
rect 160462 64812 160468 64864
rect 160520 64852 160526 64864
rect 194870 64852 194876 64864
rect 160520 64824 194876 64852
rect 160520 64812 160526 64824
rect 194870 64812 194876 64824
rect 194928 64812 194934 64864
rect 108942 64744 108948 64796
rect 109000 64784 109006 64796
rect 138474 64784 138480 64796
rect 109000 64756 138480 64784
rect 109000 64744 109006 64756
rect 138474 64744 138480 64756
rect 138532 64744 138538 64796
rect 169018 64744 169024 64796
rect 169076 64784 169082 64796
rect 202966 64784 202972 64796
rect 169076 64756 202972 64784
rect 169076 64744 169082 64756
rect 202966 64744 202972 64756
rect 203024 64744 203030 64796
rect 149790 64268 149796 64320
rect 149848 64308 149854 64320
rect 224954 64308 224960 64320
rect 149848 64280 224960 64308
rect 149848 64268 149854 64280
rect 224954 64268 224960 64280
rect 225012 64268 225018 64320
rect 84838 64200 84844 64252
rect 84896 64240 84902 64252
rect 108942 64240 108948 64252
rect 84896 64212 108948 64240
rect 84896 64200 84902 64212
rect 108942 64200 108948 64212
rect 109000 64200 109006 64252
rect 194870 64200 194876 64252
rect 194928 64240 194934 64252
rect 358814 64240 358820 64252
rect 194928 64212 358820 64240
rect 194928 64200 194934 64212
rect 358814 64200 358820 64212
rect 358872 64200 358878 64252
rect 35894 64132 35900 64184
rect 35952 64172 35958 64184
rect 134334 64172 134340 64184
rect 35952 64144 134340 64172
rect 35952 64132 35958 64144
rect 134334 64132 134340 64144
rect 134392 64132 134398 64184
rect 147306 64132 147312 64184
rect 147364 64172 147370 64184
rect 183554 64172 183560 64184
rect 147364 64144 183560 64172
rect 147364 64132 147370 64144
rect 183554 64132 183560 64144
rect 183612 64132 183618 64184
rect 202966 64132 202972 64184
rect 203024 64172 203030 64184
rect 472618 64172 472624 64184
rect 203024 64144 472624 64172
rect 203024 64132 203030 64144
rect 472618 64132 472624 64144
rect 472676 64132 472682 64184
rect 140038 63520 140044 63572
rect 140096 63560 140102 63572
rect 142982 63560 142988 63572
rect 140096 63532 142988 63560
rect 140096 63520 140102 63532
rect 142982 63520 142988 63532
rect 143040 63520 143046 63572
rect 146110 63520 146116 63572
rect 146168 63560 146174 63572
rect 147214 63560 147220 63572
rect 146168 63532 147220 63560
rect 146168 63520 146174 63532
rect 147214 63520 147220 63532
rect 147272 63520 147278 63572
rect 104710 63452 104716 63504
rect 104768 63492 104774 63504
rect 132770 63492 132776 63504
rect 104768 63464 132776 63492
rect 104768 63452 104774 63464
rect 132770 63452 132776 63464
rect 132828 63452 132834 63504
rect 159450 63452 159456 63504
rect 159508 63492 159514 63504
rect 193398 63492 193404 63504
rect 159508 63464 193404 63492
rect 159508 63452 159514 63464
rect 193398 63452 193404 63464
rect 193456 63452 193462 63504
rect 144362 63044 144368 63096
rect 144420 63084 144426 63096
rect 149790 63084 149796 63096
rect 144420 63056 149796 63084
rect 144420 63044 144426 63056
rect 149790 63044 149796 63056
rect 149848 63044 149854 63096
rect 150250 62840 150256 62892
rect 150308 62880 150314 62892
rect 227714 62880 227720 62892
rect 150308 62852 227720 62880
rect 150308 62840 150314 62852
rect 227714 62840 227720 62852
rect 227772 62840 227778 62892
rect 10318 62772 10324 62824
rect 10376 62812 10382 62824
rect 104710 62812 104716 62824
rect 10376 62784 104716 62812
rect 10376 62772 10382 62784
rect 104710 62772 104716 62784
rect 104768 62772 104774 62824
rect 147398 62772 147404 62824
rect 147456 62812 147462 62824
rect 190454 62812 190460 62824
rect 147456 62784 190460 62812
rect 147456 62772 147462 62784
rect 190454 62772 190460 62784
rect 190512 62772 190518 62824
rect 193398 62772 193404 62824
rect 193456 62812 193462 62824
rect 349154 62812 349160 62824
rect 193456 62784 349160 62812
rect 193456 62772 193462 62784
rect 349154 62772 349160 62784
rect 349212 62772 349218 62824
rect 139394 62296 139400 62348
rect 139452 62336 139458 62348
rect 142798 62336 142804 62348
rect 139452 62308 142804 62336
rect 139452 62296 139458 62308
rect 142798 62296 142804 62308
rect 142856 62296 142862 62348
rect 102226 62024 102232 62076
rect 102284 62064 102290 62076
rect 103422 62064 103428 62076
rect 102284 62036 103428 62064
rect 102284 62024 102290 62036
rect 103422 62024 103428 62036
rect 103480 62064 103486 62076
rect 134426 62064 134432 62076
rect 103480 62036 134432 62064
rect 103480 62024 103486 62036
rect 134426 62024 134432 62036
rect 134484 62024 134490 62076
rect 26234 61412 26240 61464
rect 26292 61452 26298 61464
rect 102226 61452 102232 61464
rect 26292 61424 102232 61452
rect 26292 61412 26298 61424
rect 102226 61412 102232 61424
rect 102284 61412 102290 61464
rect 44818 61344 44824 61396
rect 44876 61384 44882 61396
rect 135622 61384 135628 61396
rect 44876 61356 135628 61384
rect 44876 61344 44882 61356
rect 135622 61344 135628 61356
rect 135680 61344 135686 61396
rect 154758 61208 154764 61260
rect 154816 61248 154822 61260
rect 155218 61248 155224 61260
rect 154816 61220 155224 61248
rect 154816 61208 154822 61220
rect 155218 61208 155224 61220
rect 155276 61208 155282 61260
rect 99466 60664 99472 60716
rect 99524 60704 99530 60716
rect 100570 60704 100576 60716
rect 99524 60676 100576 60704
rect 99524 60664 99530 60676
rect 100570 60664 100576 60676
rect 100628 60704 100634 60716
rect 132678 60704 132684 60716
rect 100628 60676 132684 60704
rect 100628 60664 100634 60676
rect 132678 60664 132684 60676
rect 132736 60664 132742 60716
rect 166166 60664 166172 60716
rect 166224 60704 166230 60716
rect 197446 60704 197452 60716
rect 166224 60676 197452 60704
rect 166224 60664 166230 60676
rect 197446 60664 197452 60676
rect 197504 60704 197510 60716
rect 197814 60704 197820 60716
rect 197504 60676 197820 60704
rect 197504 60664 197510 60676
rect 197814 60664 197820 60676
rect 197872 60664 197878 60716
rect 162946 60596 162952 60648
rect 163004 60636 163010 60648
rect 189350 60636 189356 60648
rect 163004 60608 189356 60636
rect 163004 60596 163010 60608
rect 189350 60596 189356 60608
rect 189408 60596 189414 60648
rect 151906 60120 151912 60172
rect 151964 60160 151970 60172
rect 263594 60160 263600 60172
rect 151964 60132 263600 60160
rect 151964 60120 151970 60132
rect 263594 60120 263600 60132
rect 263652 60120 263658 60172
rect 197446 60052 197452 60104
rect 197504 60092 197510 60104
rect 396074 60092 396080 60104
rect 197504 60064 396080 60092
rect 197504 60052 197510 60064
rect 396074 60052 396080 60064
rect 396132 60052 396138 60104
rect 22738 59984 22744 60036
rect 22796 60024 22802 60036
rect 99466 60024 99472 60036
rect 22796 59996 99472 60024
rect 22796 59984 22802 59996
rect 99466 59984 99472 59996
rect 99524 59984 99530 60036
rect 145926 59984 145932 60036
rect 145984 60024 145990 60036
rect 147306 60024 147312 60036
rect 145984 59996 147312 60024
rect 145984 59984 145990 59996
rect 147306 59984 147312 59996
rect 147364 59984 147370 60036
rect 189350 59984 189356 60036
rect 189408 60024 189414 60036
rect 398834 60024 398840 60036
rect 189408 59996 398840 60024
rect 189408 59984 189414 59996
rect 398834 59984 398840 59996
rect 398892 59984 398898 60036
rect 110414 59848 110420 59900
rect 110472 59888 110478 59900
rect 115014 59888 115020 59900
rect 110472 59860 115020 59888
rect 110472 59848 110478 59860
rect 115014 59848 115020 59860
rect 115072 59848 115078 59900
rect 3510 59304 3516 59356
rect 3568 59344 3574 59356
rect 111058 59344 111064 59356
rect 3568 59316 111064 59344
rect 3568 59304 3574 59316
rect 111058 59304 111064 59316
rect 111116 59304 111122 59356
rect 146386 58760 146392 58812
rect 146444 58800 146450 58812
rect 186314 58800 186320 58812
rect 146444 58772 186320 58800
rect 146444 58760 146450 58772
rect 186314 58760 186320 58772
rect 186372 58760 186378 58812
rect 154022 58692 154028 58744
rect 154080 58732 154086 58744
rect 281534 58732 281540 58744
rect 154080 58704 281540 58732
rect 154080 58692 154086 58704
rect 281534 58692 281540 58704
rect 281592 58692 281598 58744
rect 60826 58624 60832 58676
rect 60884 58664 60890 58676
rect 137370 58664 137376 58676
rect 60884 58636 137376 58664
rect 60884 58624 60890 58636
rect 137370 58624 137376 58636
rect 137428 58624 137434 58676
rect 144270 58624 144276 58676
rect 144328 58664 144334 58676
rect 156598 58664 156604 58676
rect 144328 58636 156604 58664
rect 144328 58624 144334 58636
rect 156598 58624 156604 58636
rect 156656 58624 156662 58676
rect 169294 58624 169300 58676
rect 169352 58664 169358 58676
rect 467834 58664 467840 58676
rect 169352 58636 467840 58664
rect 169352 58624 169358 58636
rect 467834 58624 467840 58636
rect 467892 58624 467898 58676
rect 100754 57876 100760 57928
rect 100812 57916 100818 57928
rect 101674 57916 101680 57928
rect 100812 57888 101680 57916
rect 100812 57876 100818 57888
rect 101674 57876 101680 57888
rect 101732 57916 101738 57928
rect 134518 57916 134524 57928
rect 101732 57888 134524 57916
rect 101732 57876 101738 57888
rect 134518 57876 134524 57888
rect 134576 57876 134582 57928
rect 168466 57876 168472 57928
rect 168524 57916 168530 57928
rect 203334 57916 203340 57928
rect 168524 57888 203340 57916
rect 168524 57876 168530 57888
rect 203334 57876 203340 57888
rect 203392 57916 203398 57928
rect 204162 57916 204168 57928
rect 203392 57888 204168 57916
rect 203392 57876 203398 57888
rect 204162 57876 204168 57888
rect 204220 57876 204226 57928
rect 159266 57808 159272 57860
rect 159324 57848 159330 57860
rect 194134 57848 194140 57860
rect 159324 57820 194140 57848
rect 159324 57808 159330 57820
rect 194134 57808 194140 57820
rect 194192 57848 194198 57860
rect 194502 57848 194508 57860
rect 194192 57820 194508 57848
rect 194192 57808 194198 57820
rect 194502 57808 194508 57820
rect 194560 57808 194566 57860
rect 149974 57400 149980 57452
rect 150032 57440 150038 57452
rect 215294 57440 215300 57452
rect 150032 57412 215300 57440
rect 150032 57400 150038 57412
rect 215294 57400 215300 57412
rect 215352 57400 215358 57452
rect 151998 57332 152004 57384
rect 152056 57372 152062 57384
rect 255314 57372 255320 57384
rect 152056 57344 255320 57372
rect 152056 57332 152062 57344
rect 255314 57332 255320 57344
rect 255372 57332 255378 57384
rect 194502 57264 194508 57316
rect 194560 57304 194566 57316
rect 345014 57304 345020 57316
rect 194560 57276 345020 57304
rect 194560 57264 194566 57276
rect 345014 57264 345020 57276
rect 345072 57264 345078 57316
rect 22094 57196 22100 57248
rect 22152 57236 22158 57248
rect 100754 57236 100760 57248
rect 22152 57208 100760 57236
rect 22152 57196 22158 57208
rect 100754 57196 100760 57208
rect 100812 57196 100818 57248
rect 204162 57196 204168 57248
rect 204220 57236 204226 57248
rect 473446 57236 473452 57248
rect 204220 57208 473452 57236
rect 204220 57196 204226 57208
rect 473446 57196 473452 57208
rect 473504 57196 473510 57248
rect 99466 56516 99472 56568
rect 99524 56556 99530 56568
rect 100662 56556 100668 56568
rect 99524 56528 100668 56556
rect 99524 56516 99530 56528
rect 100662 56516 100668 56528
rect 100720 56556 100726 56568
rect 132954 56556 132960 56568
rect 100720 56528 132960 56556
rect 100720 56516 100726 56528
rect 132954 56516 132960 56528
rect 133012 56516 133018 56568
rect 162854 56516 162860 56568
rect 162912 56556 162918 56568
rect 197630 56556 197636 56568
rect 162912 56528 197636 56556
rect 162912 56516 162918 56528
rect 197630 56516 197636 56528
rect 197688 56516 197694 56568
rect 88334 55904 88340 55956
rect 88392 55944 88398 55956
rect 138750 55944 138756 55956
rect 88392 55916 138756 55944
rect 88392 55904 88398 55916
rect 138750 55904 138756 55916
rect 138808 55904 138814 55956
rect 12434 55836 12440 55888
rect 12492 55876 12498 55888
rect 99466 55876 99472 55888
rect 12492 55848 99472 55876
rect 12492 55836 12498 55848
rect 99466 55836 99472 55848
rect 99524 55836 99530 55888
rect 197630 55836 197636 55888
rect 197688 55876 197694 55888
rect 394694 55876 394700 55888
rect 197688 55848 394700 55876
rect 197688 55836 197694 55848
rect 394694 55836 394700 55848
rect 394752 55836 394758 55888
rect 113818 55156 113824 55208
rect 113876 55196 113882 55208
rect 140130 55196 140136 55208
rect 113876 55168 140136 55196
rect 113876 55156 113882 55168
rect 140130 55156 140136 55168
rect 140188 55156 140194 55208
rect 168374 55156 168380 55208
rect 168432 55196 168438 55208
rect 202874 55196 202880 55208
rect 168432 55168 202880 55196
rect 168432 55156 168438 55168
rect 202874 55156 202880 55168
rect 202932 55156 202938 55208
rect 202874 54476 202880 54528
rect 202932 54516 202938 54528
rect 468478 54516 468484 54528
rect 202932 54488 468484 54516
rect 202932 54476 202938 54488
rect 468478 54476 468484 54488
rect 468536 54476 468542 54528
rect 468570 54476 468576 54528
rect 468628 54516 468634 54528
rect 581086 54516 581092 54528
rect 468628 54488 581092 54516
rect 468628 54476 468634 54488
rect 581086 54476 581092 54488
rect 581144 54476 581150 54528
rect 138658 53796 138664 53848
rect 138716 53836 138722 53848
rect 142430 53836 142436 53848
rect 138716 53808 142436 53836
rect 138716 53796 138722 53808
rect 142430 53796 142436 53808
rect 142488 53796 142494 53848
rect 100478 53728 100484 53780
rect 100536 53768 100542 53780
rect 132862 53768 132868 53780
rect 100536 53740 132868 53768
rect 100536 53728 100542 53740
rect 132862 53728 132868 53740
rect 132920 53728 132926 53780
rect 143626 53388 143632 53440
rect 143684 53428 143690 53440
rect 147674 53428 147680 53440
rect 143684 53400 147680 53428
rect 143684 53388 143690 53400
rect 147674 53388 147680 53400
rect 147732 53388 147738 53440
rect 147858 53184 147864 53236
rect 147916 53224 147922 53236
rect 197446 53224 197452 53236
rect 147916 53196 197452 53224
rect 147916 53184 147922 53196
rect 197446 53184 197452 53196
rect 197504 53184 197510 53236
rect 95234 53116 95240 53168
rect 95292 53156 95298 53168
rect 139762 53156 139768 53168
rect 95292 53128 139768 53156
rect 95292 53116 95298 53128
rect 139762 53116 139768 53128
rect 139820 53116 139826 53168
rect 151538 53116 151544 53168
rect 151596 53156 151602 53168
rect 237374 53156 237380 53168
rect 151596 53128 237380 53156
rect 151596 53116 151602 53128
rect 237374 53116 237380 53128
rect 237432 53116 237438 53168
rect 9674 53048 9680 53100
rect 9732 53088 9738 53100
rect 100478 53088 100484 53100
rect 9732 53060 100484 53088
rect 9732 53048 9738 53060
rect 100478 53048 100484 53060
rect 100536 53048 100542 53100
rect 176010 53048 176016 53100
rect 176068 53088 176074 53100
rect 556154 53088 556160 53100
rect 176068 53060 556160 53088
rect 176068 53048 176074 53060
rect 556154 53048 556160 53060
rect 556212 53048 556218 53100
rect 148134 51756 148140 51808
rect 148192 51796 148198 51808
rect 211154 51796 211160 51808
rect 148192 51768 211160 51796
rect 148192 51756 148198 51768
rect 211154 51756 211160 51768
rect 211212 51756 211218 51808
rect 93946 51688 93952 51740
rect 94004 51728 94010 51740
rect 105538 51728 105544 51740
rect 94004 51700 105544 51728
rect 94004 51688 94010 51700
rect 105538 51688 105544 51700
rect 105596 51688 105602 51740
rect 145834 51688 145840 51740
rect 145892 51728 145898 51740
rect 168466 51728 168472 51740
rect 145892 51700 168472 51728
rect 145892 51688 145898 51700
rect 168466 51688 168472 51700
rect 168524 51688 168530 51740
rect 177482 51688 177488 51740
rect 177540 51728 177546 51740
rect 578234 51728 578240 51740
rect 177540 51700 578240 51728
rect 177540 51688 177546 51700
rect 578234 51688 578240 51700
rect 578292 51688 578298 51740
rect 100754 51008 100760 51060
rect 100812 51048 100818 51060
rect 101858 51048 101864 51060
rect 100812 51020 101864 51048
rect 100812 51008 100818 51020
rect 101858 51008 101864 51020
rect 101916 51048 101922 51060
rect 134610 51048 134616 51060
rect 101916 51020 134616 51048
rect 101916 51008 101922 51020
rect 134610 51008 134616 51020
rect 134668 51008 134674 51060
rect 147582 50396 147588 50448
rect 147640 50436 147646 50448
rect 191834 50436 191840 50448
rect 147640 50408 191840 50436
rect 147640 50396 147646 50408
rect 191834 50396 191840 50408
rect 191892 50396 191898 50448
rect 30374 50328 30380 50380
rect 30432 50368 30438 50380
rect 100754 50368 100760 50380
rect 30432 50340 100760 50368
rect 30432 50328 30438 50340
rect 100754 50328 100760 50340
rect 100812 50328 100818 50380
rect 164970 50328 164976 50380
rect 165028 50368 165034 50380
rect 368474 50368 368480 50380
rect 165028 50340 368480 50368
rect 165028 50328 165034 50340
rect 368474 50328 368480 50340
rect 368532 50328 368538 50380
rect 148686 49240 148692 49292
rect 148744 49280 148750 49292
rect 201586 49280 201592 49292
rect 148744 49252 201592 49280
rect 148744 49240 148750 49252
rect 201586 49240 201592 49252
rect 201644 49240 201650 49292
rect 150066 49036 150072 49088
rect 150124 49076 150130 49088
rect 218146 49076 218152 49088
rect 150124 49048 218152 49076
rect 150124 49036 150130 49048
rect 218146 49036 218152 49048
rect 218204 49036 218210 49088
rect 171410 48968 171416 49020
rect 171468 49008 171474 49020
rect 499574 49008 499580 49020
rect 171468 48980 499580 49008
rect 171468 48968 171474 48980
rect 499574 48968 499580 48980
rect 499632 48968 499638 49020
rect 152734 47676 152740 47728
rect 152792 47716 152798 47728
rect 256694 47716 256700 47728
rect 152792 47688 256700 47716
rect 152792 47676 152798 47688
rect 256694 47676 256700 47688
rect 256752 47676 256758 47728
rect 166258 47608 166264 47660
rect 166316 47648 166322 47660
rect 444374 47648 444380 47660
rect 166316 47620 444380 47648
rect 166316 47608 166322 47620
rect 444374 47608 444380 47620
rect 444432 47608 444438 47660
rect 174722 47540 174728 47592
rect 174780 47580 174786 47592
rect 542354 47580 542360 47592
rect 174780 47552 542360 47580
rect 174780 47540 174786 47552
rect 542354 47540 542360 47552
rect 542412 47540 542418 47592
rect 148594 46248 148600 46300
rect 148652 46288 148658 46300
rect 204254 46288 204260 46300
rect 148652 46260 204260 46288
rect 148652 46248 148658 46260
rect 204254 46248 204260 46260
rect 204312 46248 204318 46300
rect 144914 46180 144920 46232
rect 144972 46220 144978 46232
rect 166994 46220 167000 46232
rect 144972 46192 167000 46220
rect 144972 46180 144978 46192
rect 166994 46180 167000 46192
rect 167052 46180 167058 46232
rect 167914 46180 167920 46232
rect 167972 46220 167978 46232
rect 449894 46220 449900 46232
rect 167972 46192 449900 46220
rect 167972 46180 167978 46192
rect 449894 46180 449900 46192
rect 449952 46180 449958 46232
rect 135254 45568 135260 45620
rect 135312 45608 135318 45620
rect 142338 45608 142344 45620
rect 135312 45580 142344 45608
rect 135312 45568 135318 45580
rect 142338 45568 142344 45580
rect 142396 45568 142402 45620
rect 167822 44956 167828 45008
rect 167880 44996 167886 45008
rect 458174 44996 458180 45008
rect 167880 44968 458180 44996
rect 167880 44956 167886 44968
rect 458174 44956 458180 44968
rect 458232 44956 458238 45008
rect 175274 44888 175280 44940
rect 175332 44928 175338 44940
rect 560294 44928 560300 44940
rect 175332 44900 560300 44928
rect 175332 44888 175338 44900
rect 560294 44888 560300 44900
rect 560352 44888 560358 44940
rect 177574 44820 177580 44872
rect 177632 44860 177638 44872
rect 571978 44860 571984 44872
rect 177632 44832 571984 44860
rect 177632 44820 177638 44832
rect 571978 44820 571984 44832
rect 572036 44820 572042 44872
rect 149146 43596 149152 43648
rect 149204 43636 149210 43648
rect 216674 43636 216680 43648
rect 149204 43608 216680 43636
rect 149204 43596 149210 43608
rect 216674 43596 216680 43608
rect 216732 43596 216738 43648
rect 162118 43528 162124 43580
rect 162176 43568 162182 43580
rect 361574 43568 361580 43580
rect 162176 43540 361580 43568
rect 162176 43528 162182 43540
rect 361574 43528 361580 43540
rect 361632 43528 361638 43580
rect 164418 43460 164424 43512
rect 164476 43500 164482 43512
rect 426434 43500 426440 43512
rect 164476 43472 426440 43500
rect 164476 43460 164482 43472
rect 426434 43460 426440 43472
rect 426492 43460 426498 43512
rect 63494 43392 63500 43444
rect 63552 43432 63558 43444
rect 136634 43432 136640 43444
rect 63552 43404 136640 43432
rect 63552 43392 63558 43404
rect 136634 43392 136640 43404
rect 136692 43392 136698 43444
rect 172238 43392 172244 43444
rect 172296 43432 172302 43444
rect 502334 43432 502340 43444
rect 172296 43404 502340 43432
rect 172296 43392 172302 43404
rect 502334 43392 502340 43404
rect 502392 43392 502398 43444
rect 150526 42304 150532 42356
rect 150584 42344 150590 42356
rect 233234 42344 233240 42356
rect 150584 42316 233240 42344
rect 150584 42304 150590 42316
rect 233234 42304 233240 42316
rect 233292 42304 233298 42356
rect 155402 42236 155408 42288
rect 155460 42276 155466 42288
rect 292666 42276 292672 42288
rect 155460 42248 292672 42276
rect 155460 42236 155466 42248
rect 292666 42236 292672 42248
rect 292724 42236 292730 42288
rect 158162 42168 158168 42220
rect 158220 42208 158226 42220
rect 328454 42208 328460 42220
rect 158220 42180 328460 42208
rect 158220 42168 158226 42180
rect 328454 42168 328460 42180
rect 328512 42168 328518 42220
rect 172146 42100 172152 42152
rect 172204 42140 172210 42152
rect 498286 42140 498292 42152
rect 172204 42112 498292 42140
rect 172204 42100 172210 42112
rect 498286 42100 498292 42112
rect 498344 42100 498350 42152
rect 70394 42032 70400 42084
rect 70452 42072 70458 42084
rect 136910 42072 136916 42084
rect 70452 42044 136916 42072
rect 70452 42032 70458 42044
rect 136910 42032 136916 42044
rect 136968 42032 136974 42084
rect 174814 42032 174820 42084
rect 174872 42072 174878 42084
rect 538858 42072 538864 42084
rect 174872 42044 538864 42072
rect 174872 42032 174878 42044
rect 538858 42032 538864 42044
rect 538916 42032 538922 42084
rect 155494 40944 155500 40996
rect 155552 40984 155558 40996
rect 300854 40984 300860 40996
rect 155552 40956 300860 40984
rect 155552 40944 155558 40956
rect 300854 40944 300860 40956
rect 300912 40944 300918 40996
rect 156690 40876 156696 40928
rect 156748 40916 156754 40928
rect 309134 40916 309140 40928
rect 156748 40888 309140 40916
rect 156748 40876 156754 40888
rect 309134 40876 309140 40888
rect 309192 40876 309198 40928
rect 166350 40808 166356 40860
rect 166408 40848 166414 40860
rect 427814 40848 427820 40860
rect 166408 40820 427820 40848
rect 166408 40808 166414 40820
rect 427814 40808 427820 40820
rect 427872 40808 427878 40860
rect 167086 40740 167092 40792
rect 167144 40780 167150 40792
rect 462314 40780 462320 40792
rect 167144 40752 462320 40780
rect 167144 40740 167150 40752
rect 462314 40740 462320 40752
rect 462372 40740 462378 40792
rect 74534 40672 74540 40724
rect 74592 40712 74598 40724
rect 138198 40712 138204 40724
rect 74592 40684 138204 40712
rect 74592 40672 74598 40684
rect 138198 40672 138204 40684
rect 138256 40672 138262 40724
rect 173526 40672 173532 40724
rect 173584 40712 173590 40724
rect 516134 40712 516140 40724
rect 173584 40684 516140 40712
rect 173584 40672 173590 40684
rect 516134 40672 516140 40684
rect 516192 40672 516198 40724
rect 152642 39584 152648 39636
rect 152700 39624 152706 39636
rect 251174 39624 251180 39636
rect 152700 39596 251180 39624
rect 152700 39584 152706 39596
rect 251174 39584 251180 39596
rect 251232 39584 251238 39636
rect 163498 39516 163504 39568
rect 163556 39556 163562 39568
rect 340966 39556 340972 39568
rect 163556 39528 340972 39556
rect 163556 39516 163562 39528
rect 340966 39516 340972 39528
rect 341024 39516 341030 39568
rect 169386 39448 169392 39500
rect 169444 39488 169450 39500
rect 470594 39488 470600 39500
rect 169444 39460 470600 39488
rect 169444 39448 169450 39460
rect 470594 39448 470600 39460
rect 470652 39448 470658 39500
rect 170582 39380 170588 39432
rect 170640 39420 170646 39432
rect 481634 39420 481640 39432
rect 170640 39392 481640 39420
rect 170640 39380 170646 39392
rect 481634 39380 481640 39392
rect 481692 39380 481698 39432
rect 77386 39312 77392 39364
rect 77444 39352 77450 39364
rect 138290 39352 138296 39364
rect 77444 39324 138296 39352
rect 77444 39312 77450 39324
rect 138290 39312 138296 39324
rect 138348 39312 138354 39364
rect 174078 39312 174084 39364
rect 174136 39352 174142 39364
rect 534074 39352 534080 39364
rect 174136 39324 534080 39352
rect 174136 39312 174142 39324
rect 534074 39312 534080 39324
rect 534132 39312 534138 39364
rect 154206 38156 154212 38208
rect 154264 38196 154270 38208
rect 267826 38196 267832 38208
rect 154264 38168 267832 38196
rect 154264 38156 154270 38168
rect 267826 38156 267832 38168
rect 267884 38156 267890 38208
rect 161198 38088 161204 38140
rect 161256 38128 161262 38140
rect 372614 38128 372620 38140
rect 161256 38100 372620 38128
rect 161256 38088 161262 38100
rect 372614 38088 372620 38100
rect 372672 38088 372678 38140
rect 170674 38020 170680 38072
rect 170732 38060 170738 38072
rect 488534 38060 488540 38072
rect 170732 38032 488540 38060
rect 170732 38020 170738 38032
rect 488534 38020 488540 38032
rect 488592 38020 488598 38072
rect 173618 37952 173624 38004
rect 173676 37992 173682 38004
rect 528554 37992 528560 38004
rect 173676 37964 528560 37992
rect 173676 37952 173682 37964
rect 528554 37952 528560 37964
rect 528612 37952 528618 38004
rect 13814 37884 13820 37936
rect 13872 37924 13878 37936
rect 132494 37924 132500 37936
rect 13872 37896 132500 37924
rect 13872 37884 13878 37896
rect 132494 37884 132500 37896
rect 132552 37884 132558 37936
rect 176194 37884 176200 37936
rect 176252 37924 176258 37936
rect 552014 37924 552020 37936
rect 176252 37896 552020 37924
rect 176252 37884 176258 37896
rect 552014 37884 552020 37896
rect 552072 37884 552078 37936
rect 147766 36864 147772 36916
rect 147824 36904 147830 36916
rect 208394 36904 208400 36916
rect 147824 36876 208400 36904
rect 147824 36864 147830 36876
rect 208394 36864 208400 36876
rect 208452 36864 208458 36916
rect 149054 36796 149060 36848
rect 149112 36836 149118 36848
rect 222194 36836 222200 36848
rect 149112 36808 222200 36836
rect 149112 36796 149118 36808
rect 222194 36796 222200 36808
rect 222252 36796 222258 36848
rect 156782 36728 156788 36780
rect 156840 36768 156846 36780
rect 303614 36768 303620 36780
rect 156840 36740 303620 36768
rect 156840 36728 156846 36740
rect 303614 36728 303620 36740
rect 303672 36728 303678 36780
rect 165614 36660 165620 36712
rect 165672 36700 165678 36712
rect 440326 36700 440332 36712
rect 165672 36672 440332 36700
rect 165672 36660 165678 36672
rect 440326 36660 440332 36672
rect 440384 36660 440390 36712
rect 175826 36592 175832 36644
rect 175884 36632 175890 36644
rect 558914 36632 558920 36644
rect 175884 36604 558920 36632
rect 175884 36592 175890 36604
rect 558914 36592 558920 36604
rect 558972 36592 558978 36644
rect 104158 36524 104164 36576
rect 104216 36564 104222 36576
rect 140406 36564 140412 36576
rect 104216 36536 140412 36564
rect 104216 36524 104222 36536
rect 140406 36524 140412 36536
rect 140464 36524 140470 36576
rect 177666 36524 177672 36576
rect 177724 36564 177730 36576
rect 571334 36564 571340 36576
rect 177724 36536 571340 36564
rect 177724 36524 177730 36536
rect 571334 36524 571340 36536
rect 571392 36524 571398 36576
rect 153286 35436 153292 35488
rect 153344 35476 153350 35488
rect 276014 35476 276020 35488
rect 153344 35448 276020 35476
rect 153344 35436 153350 35448
rect 276014 35436 276020 35448
rect 276072 35436 276078 35488
rect 158070 35368 158076 35420
rect 158128 35408 158134 35420
rect 321554 35408 321560 35420
rect 158128 35380 321560 35408
rect 158128 35368 158134 35380
rect 321554 35368 321560 35380
rect 321612 35368 321618 35420
rect 165154 35300 165160 35352
rect 165212 35340 165218 35352
rect 418154 35340 418160 35352
rect 165212 35312 418160 35340
rect 165212 35300 165218 35312
rect 418154 35300 418160 35312
rect 418212 35300 418218 35352
rect 170766 35232 170772 35284
rect 170824 35272 170830 35284
rect 491294 35272 491300 35284
rect 170824 35244 491300 35272
rect 170824 35232 170830 35244
rect 491294 35232 491300 35244
rect 491352 35232 491358 35284
rect 38654 35164 38660 35216
rect 38712 35204 38718 35216
rect 136358 35204 136364 35216
rect 38712 35176 136364 35204
rect 38712 35164 38718 35176
rect 136358 35164 136364 35176
rect 136416 35164 136422 35216
rect 145650 35164 145656 35216
rect 145708 35204 145714 35216
rect 165614 35204 165620 35216
rect 145708 35176 165620 35204
rect 145708 35164 145714 35176
rect 165614 35164 165620 35176
rect 165672 35164 165678 35216
rect 177758 35164 177764 35216
rect 177816 35204 177822 35216
rect 576854 35204 576860 35216
rect 177816 35176 576860 35204
rect 177816 35164 177822 35176
rect 576854 35164 576860 35176
rect 576912 35164 576918 35216
rect 155586 34008 155592 34060
rect 155644 34048 155650 34060
rect 299566 34048 299572 34060
rect 155644 34020 299572 34048
rect 155644 34008 155650 34020
rect 299566 34008 299572 34020
rect 299624 34008 299630 34060
rect 162302 33940 162308 33992
rect 162360 33980 162366 33992
rect 385034 33980 385040 33992
rect 162360 33952 385040 33980
rect 162360 33940 162366 33952
rect 385034 33940 385040 33952
rect 385092 33940 385098 33992
rect 169662 33872 169668 33924
rect 169720 33912 169726 33924
rect 474734 33912 474740 33924
rect 169720 33884 474740 33912
rect 169720 33872 169726 33884
rect 474734 33872 474740 33884
rect 474792 33872 474798 33924
rect 170858 33804 170864 33856
rect 170916 33844 170922 33856
rect 490006 33844 490012 33856
rect 170916 33816 490012 33844
rect 170916 33804 170922 33816
rect 490006 33804 490012 33816
rect 490064 33804 490070 33856
rect 175918 33736 175924 33788
rect 175976 33776 175982 33788
rect 563698 33776 563704 33788
rect 175976 33748 563704 33776
rect 175976 33736 175982 33748
rect 563698 33736 563704 33748
rect 563756 33736 563762 33788
rect 148502 32648 148508 32700
rect 148560 32688 148566 32700
rect 205634 32688 205640 32700
rect 148560 32660 205640 32688
rect 148560 32648 148566 32660
rect 205634 32648 205640 32660
rect 205692 32648 205698 32700
rect 150894 32580 150900 32632
rect 150952 32620 150958 32632
rect 235994 32620 236000 32632
rect 150952 32592 236000 32620
rect 150952 32580 150958 32592
rect 235994 32580 236000 32592
rect 236052 32580 236058 32632
rect 161106 32512 161112 32564
rect 161164 32552 161170 32564
rect 357434 32552 357440 32564
rect 161164 32524 357440 32552
rect 161164 32512 161170 32524
rect 357434 32512 357440 32524
rect 357492 32512 357498 32564
rect 173710 32444 173716 32496
rect 173768 32484 173774 32496
rect 531406 32484 531412 32496
rect 173768 32456 531412 32484
rect 173768 32444 173774 32456
rect 531406 32444 531412 32456
rect 531464 32444 531470 32496
rect 176654 32376 176660 32428
rect 176712 32416 176718 32428
rect 582374 32416 582380 32428
rect 176712 32388 582380 32416
rect 176712 32376 176718 32388
rect 582374 32376 582380 32388
rect 582432 32376 582438 32428
rect 156874 31220 156880 31272
rect 156932 31260 156938 31272
rect 317414 31260 317420 31272
rect 156932 31232 317420 31260
rect 156932 31220 156938 31232
rect 317414 31220 317420 31232
rect 317472 31220 317478 31272
rect 164326 31152 164332 31204
rect 164384 31192 164390 31204
rect 420914 31192 420920 31204
rect 164384 31164 420920 31192
rect 164384 31152 164390 31164
rect 420914 31152 420920 31164
rect 420972 31152 420978 31204
rect 169478 31084 169484 31136
rect 169536 31124 169542 31136
rect 466454 31124 466460 31136
rect 169536 31096 466460 31124
rect 169536 31084 169542 31096
rect 466454 31084 466460 31096
rect 466512 31084 466518 31136
rect 177298 31016 177304 31068
rect 177356 31056 177362 31068
rect 554774 31056 554780 31068
rect 177356 31028 554780 31056
rect 177356 31016 177362 31028
rect 554774 31016 554780 31028
rect 554832 31016 554838 31068
rect 151262 29860 151268 29912
rect 151320 29900 151326 29912
rect 242986 29900 242992 29912
rect 151320 29872 242992 29900
rect 151320 29860 151326 29872
rect 242986 29860 242992 29872
rect 243044 29860 243050 29912
rect 157978 29792 157984 29844
rect 158036 29832 158042 29844
rect 332686 29832 332692 29844
rect 158036 29804 332692 29832
rect 158036 29792 158042 29804
rect 332686 29792 332692 29804
rect 332744 29792 332750 29844
rect 161290 29724 161296 29776
rect 161348 29764 161354 29776
rect 365806 29764 365812 29776
rect 161348 29736 365812 29764
rect 161348 29724 161354 29736
rect 365806 29724 365812 29736
rect 365864 29724 365870 29776
rect 166442 29656 166448 29708
rect 166500 29696 166506 29708
rect 441614 29696 441620 29708
rect 166500 29668 441620 29696
rect 166500 29656 166506 29668
rect 441614 29656 441620 29668
rect 441672 29656 441678 29708
rect 171318 29588 171324 29640
rect 171376 29628 171382 29640
rect 506566 29628 506572 29640
rect 171376 29600 506572 29628
rect 171376 29588 171382 29600
rect 506566 29588 506572 29600
rect 506624 29588 506630 29640
rect 159726 28432 159732 28484
rect 159784 28472 159790 28484
rect 339494 28472 339500 28484
rect 159784 28444 339500 28472
rect 159784 28432 159790 28444
rect 339494 28432 339500 28444
rect 339552 28432 339558 28484
rect 163866 28364 163872 28416
rect 163924 28404 163930 28416
rect 397454 28404 397460 28416
rect 163924 28376 397460 28404
rect 163924 28364 163930 28376
rect 397454 28364 397460 28376
rect 397512 28364 397518 28416
rect 169570 28296 169576 28348
rect 169628 28336 169634 28348
rect 477494 28336 477500 28348
rect 169628 28308 477500 28336
rect 169628 28296 169634 28308
rect 477494 28296 477500 28308
rect 477552 28296 477558 28348
rect 52546 28228 52552 28280
rect 52604 28268 52610 28280
rect 135438 28268 135444 28280
rect 52604 28240 135444 28268
rect 52604 28228 52610 28240
rect 135438 28228 135444 28240
rect 135496 28228 135502 28280
rect 171226 28228 171232 28280
rect 171284 28268 171290 28280
rect 509234 28268 509240 28280
rect 171284 28240 509240 28268
rect 171284 28228 171290 28240
rect 509234 28228 509240 28240
rect 509292 28228 509298 28280
rect 153194 27140 153200 27192
rect 153252 27180 153258 27192
rect 282914 27180 282920 27192
rect 153252 27152 282920 27180
rect 153252 27140 153258 27152
rect 282914 27140 282920 27152
rect 282972 27140 282978 27192
rect 162394 27072 162400 27124
rect 162452 27112 162458 27124
rect 374086 27112 374092 27124
rect 162452 27084 374092 27112
rect 162452 27072 162458 27084
rect 374086 27072 374092 27084
rect 374144 27072 374150 27124
rect 165338 27004 165344 27056
rect 165396 27044 165402 27056
rect 425054 27044 425060 27056
rect 165396 27016 425060 27044
rect 165396 27004 165402 27016
rect 425054 27004 425060 27016
rect 425112 27004 425118 27056
rect 171870 26936 171876 26988
rect 171928 26976 171934 26988
rect 513374 26976 513380 26988
rect 171928 26948 513380 26976
rect 171928 26936 171934 26948
rect 513374 26936 513380 26948
rect 513432 26936 513438 26988
rect 35986 26868 35992 26920
rect 36044 26908 36050 26920
rect 134242 26908 134248 26920
rect 36044 26880 134248 26908
rect 36044 26868 36050 26880
rect 134242 26868 134248 26880
rect 134300 26868 134306 26920
rect 174906 26868 174912 26920
rect 174964 26908 174970 26920
rect 535454 26908 535460 26920
rect 174964 26880 535460 26908
rect 174964 26868 174970 26880
rect 535454 26868 535460 26880
rect 535512 26868 535518 26920
rect 156966 25780 156972 25832
rect 157024 25820 157030 25832
rect 310514 25820 310520 25832
rect 157024 25792 310520 25820
rect 157024 25780 157030 25792
rect 310514 25780 310520 25792
rect 310572 25780 310578 25832
rect 163774 25712 163780 25764
rect 163832 25752 163838 25764
rect 391934 25752 391940 25764
rect 163832 25724 391940 25752
rect 163832 25712 163838 25724
rect 391934 25712 391940 25724
rect 391992 25712 391998 25764
rect 181622 25644 181628 25696
rect 181680 25684 181686 25696
rect 436094 25684 436100 25696
rect 181680 25656 436100 25684
rect 181680 25644 181686 25656
rect 436094 25644 436100 25656
rect 436152 25644 436158 25696
rect 172606 25576 172612 25628
rect 172664 25616 172670 25628
rect 520274 25616 520280 25628
rect 172664 25588 520280 25616
rect 172664 25576 172670 25588
rect 520274 25576 520280 25588
rect 520332 25576 520338 25628
rect 145742 25508 145748 25560
rect 145800 25548 145806 25560
rect 171778 25548 171784 25560
rect 145800 25520 171784 25548
rect 145800 25508 145806 25520
rect 171778 25508 171784 25520
rect 171836 25508 171842 25560
rect 174998 25508 175004 25560
rect 175056 25548 175062 25560
rect 546494 25548 546500 25560
rect 175056 25520 546500 25548
rect 175056 25508 175062 25520
rect 546494 25508 546500 25520
rect 546552 25508 546558 25560
rect 157058 24352 157064 24404
rect 157116 24392 157122 24404
rect 314654 24392 314660 24404
rect 157116 24364 314660 24392
rect 157116 24352 157122 24364
rect 314654 24352 314660 24364
rect 314712 24352 314718 24404
rect 165246 24284 165252 24336
rect 165304 24324 165310 24336
rect 409874 24324 409880 24336
rect 165304 24296 409880 24324
rect 165304 24284 165310 24296
rect 409874 24284 409880 24296
rect 409932 24284 409938 24336
rect 182818 24216 182824 24268
rect 182876 24256 182882 24268
rect 442994 24256 443000 24268
rect 182876 24228 443000 24256
rect 182876 24216 182882 24228
rect 442994 24216 443000 24228
rect 443052 24216 443058 24268
rect 172514 24148 172520 24200
rect 172572 24188 172578 24200
rect 527174 24188 527180 24200
rect 172572 24160 527180 24188
rect 172572 24148 172578 24160
rect 527174 24148 527180 24160
rect 527232 24148 527238 24200
rect 40034 24080 40040 24132
rect 40092 24120 40098 24132
rect 135346 24120 135352 24132
rect 40092 24092 135352 24120
rect 40092 24080 40098 24092
rect 135346 24080 135352 24092
rect 135404 24080 135410 24132
rect 145558 24080 145564 24132
rect 145616 24120 145622 24132
rect 164878 24120 164884 24132
rect 145616 24092 164884 24120
rect 145616 24080 145622 24092
rect 164878 24080 164884 24092
rect 164936 24080 164942 24132
rect 176286 24080 176292 24132
rect 176344 24120 176350 24132
rect 564526 24120 564532 24132
rect 176344 24092 564532 24120
rect 176344 24080 176350 24092
rect 564526 24080 564532 24092
rect 564584 24080 564590 24132
rect 144178 23468 144184 23520
rect 144236 23508 144242 23520
rect 144914 23508 144920 23520
rect 144236 23480 144920 23508
rect 144236 23468 144242 23480
rect 144914 23468 144920 23480
rect 144972 23468 144978 23520
rect 150158 22992 150164 23044
rect 150216 23032 150222 23044
rect 219434 23032 219440 23044
rect 150216 23004 219440 23032
rect 150216 22992 150222 23004
rect 219434 22992 219440 23004
rect 219492 22992 219498 23044
rect 157150 22924 157156 22976
rect 157208 22964 157214 22976
rect 316126 22964 316132 22976
rect 157208 22936 316132 22964
rect 157208 22924 157214 22936
rect 316126 22924 316132 22936
rect 316184 22924 316190 22976
rect 164234 22856 164240 22908
rect 164292 22896 164298 22908
rect 416774 22896 416780 22908
rect 164292 22868 416780 22896
rect 164292 22856 164298 22868
rect 416774 22856 416780 22868
rect 416832 22856 416838 22908
rect 168190 22788 168196 22840
rect 168248 22828 168254 22840
rect 460934 22828 460940 22840
rect 168248 22800 460940 22828
rect 168248 22788 168254 22800
rect 460934 22788 460940 22800
rect 460992 22788 460998 22840
rect 173986 22720 173992 22772
rect 174044 22760 174050 22772
rect 538214 22760 538220 22772
rect 174044 22732 538220 22760
rect 174044 22720 174050 22732
rect 538214 22720 538220 22732
rect 538272 22720 538278 22772
rect 157426 21632 157432 21684
rect 157484 21672 157490 21684
rect 329834 21672 329840 21684
rect 157484 21644 329840 21672
rect 157484 21632 157490 21644
rect 329834 21632 329840 21644
rect 329892 21632 329898 21684
rect 157518 21564 157524 21616
rect 157576 21604 157582 21616
rect 336734 21604 336740 21616
rect 157576 21576 336740 21604
rect 157576 21564 157582 21576
rect 336734 21564 336740 21576
rect 336792 21564 336798 21616
rect 337378 21564 337384 21616
rect 337436 21604 337442 21616
rect 471974 21604 471980 21616
rect 337436 21576 471980 21604
rect 337436 21564 337442 21576
rect 471974 21564 471980 21576
rect 472032 21564 472038 21616
rect 158714 21496 158720 21548
rect 158772 21536 158778 21548
rect 343634 21536 343640 21548
rect 158772 21508 343640 21536
rect 158772 21496 158778 21508
rect 343634 21496 343640 21508
rect 343692 21496 343698 21548
rect 159818 21428 159824 21480
rect 159876 21468 159882 21480
rect 350534 21468 350540 21480
rect 159876 21440 350540 21468
rect 159876 21428 159882 21440
rect 350534 21428 350540 21440
rect 350592 21428 350598 21480
rect 178862 21360 178868 21412
rect 178920 21400 178926 21412
rect 422294 21400 422300 21412
rect 178920 21372 422300 21400
rect 178920 21360 178926 21372
rect 422294 21360 422300 21372
rect 422352 21360 422358 21412
rect 286318 20612 286324 20664
rect 286376 20652 286382 20664
rect 579982 20652 579988 20664
rect 286376 20624 579988 20652
rect 286376 20612 286382 20624
rect 579982 20612 579988 20624
rect 580040 20612 580046 20664
rect 154390 20204 154396 20256
rect 154448 20244 154454 20256
rect 280154 20244 280160 20256
rect 154448 20216 280160 20244
rect 154448 20204 154454 20216
rect 280154 20204 280160 20216
rect 280212 20204 280218 20256
rect 155218 20136 155224 20188
rect 155276 20176 155282 20188
rect 287054 20176 287060 20188
rect 155276 20148 287060 20176
rect 155276 20136 155282 20148
rect 287054 20136 287060 20148
rect 287112 20136 287118 20188
rect 155678 20068 155684 20120
rect 155736 20108 155742 20120
rect 293954 20108 293960 20120
rect 155736 20080 293960 20108
rect 155736 20068 155742 20080
rect 293954 20068 293960 20080
rect 294012 20068 294018 20120
rect 161934 20000 161940 20052
rect 161992 20040 161998 20052
rect 379514 20040 379520 20052
rect 161992 20012 379520 20040
rect 161992 20000 161998 20012
rect 379514 20000 379520 20012
rect 379572 20000 379578 20052
rect 155770 19932 155776 19984
rect 155828 19972 155834 19984
rect 291194 19972 291200 19984
rect 155828 19944 291200 19972
rect 155828 19932 155834 19944
rect 291194 19932 291200 19944
rect 291252 19932 291258 19984
rect 291838 19932 291844 19984
rect 291896 19972 291902 19984
rect 518894 19972 518900 19984
rect 291896 19944 518900 19972
rect 291896 19932 291902 19944
rect 518894 19932 518900 19944
rect 518952 19932 518958 19984
rect 153010 18844 153016 18896
rect 153068 18884 153074 18896
rect 266354 18884 266360 18896
rect 153068 18856 266360 18884
rect 153068 18844 153074 18856
rect 266354 18844 266360 18856
rect 266412 18844 266418 18896
rect 160278 18776 160284 18828
rect 160336 18816 160342 18828
rect 357526 18816 357532 18828
rect 160336 18788 357532 18816
rect 160336 18776 160342 18788
rect 357526 18776 357532 18788
rect 357584 18776 357590 18828
rect 166810 18708 166816 18760
rect 166868 18748 166874 18760
rect 431954 18748 431960 18760
rect 166868 18720 431960 18748
rect 166868 18708 166874 18720
rect 431954 18708 431960 18720
rect 432012 18708 432018 18760
rect 176378 18640 176384 18692
rect 176436 18680 176442 18692
rect 567194 18680 567200 18692
rect 176436 18652 567200 18680
rect 176436 18640 176442 18652
rect 567194 18640 567200 18652
rect 567252 18640 567258 18692
rect 177942 18572 177948 18624
rect 178000 18612 178006 18624
rect 574094 18612 574100 18624
rect 178000 18584 574100 18612
rect 178000 18572 178006 18584
rect 574094 18572 574100 18584
rect 574152 18572 574158 18624
rect 151170 17484 151176 17536
rect 151228 17524 151234 17536
rect 234706 17524 234712 17536
rect 151228 17496 234712 17524
rect 151228 17484 151234 17496
rect 234706 17484 234712 17496
rect 234764 17484 234770 17536
rect 180426 17416 180432 17468
rect 180484 17456 180490 17468
rect 415486 17456 415492 17468
rect 180484 17428 415492 17456
rect 180484 17416 180490 17428
rect 415486 17416 415492 17428
rect 415544 17416 415550 17468
rect 168098 17348 168104 17400
rect 168156 17388 168162 17400
rect 445754 17388 445760 17400
rect 168156 17360 445760 17388
rect 168156 17348 168162 17360
rect 445754 17348 445760 17360
rect 445812 17348 445818 17400
rect 168006 17280 168012 17332
rect 168064 17320 168070 17332
rect 448606 17320 448612 17332
rect 168064 17292 448612 17320
rect 168064 17280 168070 17292
rect 448606 17280 448612 17292
rect 448664 17280 448670 17332
rect 171962 17212 171968 17264
rect 172020 17252 172026 17264
rect 503714 17252 503720 17264
rect 172020 17224 503720 17252
rect 172020 17212 172026 17224
rect 503714 17212 503720 17224
rect 503772 17212 503778 17264
rect 152826 16056 152832 16108
rect 152884 16096 152890 16108
rect 259546 16096 259552 16108
rect 152884 16068 259552 16096
rect 152884 16056 152890 16068
rect 259546 16056 259552 16068
rect 259604 16056 259610 16108
rect 160094 15988 160100 16040
rect 160152 16028 160158 16040
rect 361114 16028 361120 16040
rect 160152 16000 361120 16028
rect 160152 15988 160158 16000
rect 361114 15988 361120 16000
rect 361172 15988 361178 16040
rect 160186 15920 160192 15972
rect 160244 15960 160250 15972
rect 364610 15960 364616 15972
rect 160244 15932 364616 15960
rect 160244 15920 160250 15932
rect 364610 15920 364616 15932
rect 364668 15920 364674 15972
rect 400858 15920 400864 15972
rect 400916 15960 400922 15972
rect 478874 15960 478880 15972
rect 400916 15932 478880 15960
rect 400916 15920 400922 15932
rect 478874 15920 478880 15932
rect 478932 15920 478938 15972
rect 166626 15852 166632 15904
rect 166684 15892 166690 15904
rect 432046 15892 432052 15904
rect 166684 15864 432052 15892
rect 166684 15852 166690 15864
rect 432046 15852 432052 15864
rect 432104 15852 432110 15904
rect 153930 14696 153936 14748
rect 153988 14736 153994 14748
rect 276106 14736 276112 14748
rect 153988 14708 276112 14736
rect 153988 14696 153994 14708
rect 276106 14696 276112 14708
rect 276164 14696 276170 14748
rect 158530 14628 158536 14680
rect 158588 14668 158594 14680
rect 324406 14668 324412 14680
rect 158588 14640 324412 14668
rect 158588 14628 158594 14640
rect 324406 14628 324412 14640
rect 324464 14628 324470 14680
rect 178770 14560 178776 14612
rect 178828 14600 178834 14612
rect 407206 14600 407212 14612
rect 178828 14572 407212 14600
rect 178828 14560 178834 14572
rect 407206 14560 407212 14572
rect 407264 14560 407270 14612
rect 163958 14492 163964 14544
rect 164016 14532 164022 14544
rect 407114 14532 407120 14544
rect 164016 14504 407120 14532
rect 164016 14492 164022 14504
rect 407114 14492 407120 14504
rect 407172 14492 407178 14544
rect 172054 14424 172060 14476
rect 172112 14464 172118 14476
rect 511258 14464 511264 14476
rect 172112 14436 511264 14464
rect 172112 14424 172118 14436
rect 511258 14424 511264 14436
rect 511316 14424 511322 14476
rect 152458 13268 152464 13320
rect 152516 13308 152522 13320
rect 258258 13308 258264 13320
rect 152516 13280 258264 13308
rect 152516 13268 152522 13280
rect 258258 13268 258264 13280
rect 258316 13268 258322 13320
rect 156506 13200 156512 13252
rect 156564 13240 156570 13252
rect 307938 13240 307944 13252
rect 156564 13212 307944 13240
rect 156564 13200 156570 13212
rect 307938 13200 307944 13212
rect 307996 13200 308002 13252
rect 164050 13132 164056 13184
rect 164108 13172 164114 13184
rect 398926 13172 398932 13184
rect 164108 13144 398932 13172
rect 164108 13132 164114 13144
rect 398926 13132 398932 13144
rect 398984 13132 398990 13184
rect 170950 13064 170956 13116
rect 171008 13104 171014 13116
rect 493042 13104 493048 13116
rect 171008 13076 493048 13104
rect 171008 13064 171014 13076
rect 493042 13064 493048 13076
rect 493100 13064 493106 13116
rect 152550 11908 152556 11960
rect 152608 11948 152614 11960
rect 252370 11948 252376 11960
rect 152608 11920 252376 11948
rect 152608 11908 152614 11920
rect 252370 11908 252376 11920
rect 252428 11908 252434 11960
rect 160002 11840 160008 11892
rect 160060 11880 160066 11892
rect 349246 11880 349252 11892
rect 160060 11852 349252 11880
rect 160060 11840 160066 11852
rect 349246 11840 349252 11852
rect 349304 11840 349310 11892
rect 166718 11772 166724 11824
rect 166776 11812 166782 11824
rect 439130 11812 439136 11824
rect 166776 11784 439136 11812
rect 166776 11772 166782 11784
rect 439130 11772 439136 11784
rect 439188 11772 439194 11824
rect 175090 11704 175096 11756
rect 175148 11744 175154 11756
rect 548610 11744 548616 11756
rect 175148 11716 548616 11744
rect 175148 11704 175154 11716
rect 548610 11704 548616 11716
rect 548668 11704 548674 11756
rect 201494 11636 201500 11688
rect 201552 11676 201558 11688
rect 202690 11676 202696 11688
rect 201552 11648 202696 11676
rect 201552 11636 201558 11648
rect 202690 11636 202696 11648
rect 202748 11636 202754 11688
rect 234614 11636 234620 11688
rect 234672 11676 234678 11688
rect 235810 11676 235816 11688
rect 234672 11648 235816 11676
rect 234672 11636 234678 11648
rect 235810 11636 235816 11648
rect 235868 11636 235874 11688
rect 259454 11636 259460 11688
rect 259512 11676 259518 11688
rect 260650 11676 260656 11688
rect 259512 11648 260656 11676
rect 259512 11636 259518 11648
rect 260650 11636 260656 11648
rect 260708 11636 260714 11688
rect 151630 10548 151636 10600
rect 151688 10588 151694 10600
rect 245194 10588 245200 10600
rect 151688 10560 245200 10588
rect 151688 10548 151694 10560
rect 245194 10548 245200 10560
rect 245252 10548 245258 10600
rect 159910 10480 159916 10532
rect 159968 10520 159974 10532
rect 342898 10520 342904 10532
rect 159968 10492 342904 10520
rect 159968 10480 159974 10492
rect 342898 10480 342904 10492
rect 342956 10480 342962 10532
rect 162670 10412 162676 10464
rect 162728 10452 162734 10464
rect 386690 10452 386696 10464
rect 162728 10424 386696 10452
rect 162728 10412 162734 10424
rect 386690 10412 386696 10424
rect 386748 10412 386754 10464
rect 166902 10344 166908 10396
rect 166960 10384 166966 10396
rect 435082 10384 435088 10396
rect 166960 10356 435088 10384
rect 166960 10344 166966 10356
rect 435082 10344 435088 10356
rect 435140 10344 435146 10396
rect 176562 10276 176568 10328
rect 176620 10316 176626 10328
rect 563054 10316 563060 10328
rect 176620 10288 563060 10316
rect 176620 10276 176626 10288
rect 563054 10276 563060 10288
rect 563112 10276 563118 10328
rect 150802 9188 150808 9240
rect 150860 9228 150866 9240
rect 241698 9228 241704 9240
rect 150860 9200 241704 9228
rect 150860 9188 150866 9200
rect 241698 9188 241704 9200
rect 241756 9188 241762 9240
rect 161382 9120 161388 9172
rect 161440 9160 161446 9172
rect 371694 9160 371700 9172
rect 161440 9132 371700 9160
rect 161440 9120 161446 9132
rect 371694 9120 371700 9132
rect 371752 9120 371758 9172
rect 164142 9052 164148 9104
rect 164200 9092 164206 9104
rect 404814 9092 404820 9104
rect 164200 9064 404820 9092
rect 164200 9052 164206 9064
rect 404814 9052 404820 9064
rect 404872 9052 404878 9104
rect 168282 8984 168288 9036
rect 168340 9024 168346 9036
rect 456886 9024 456892 9036
rect 168340 8996 456892 9024
rect 168340 8984 168346 8996
rect 456886 8984 456892 8996
rect 456944 8984 456950 9036
rect 176470 8916 176476 8968
rect 176528 8956 176534 8968
rect 556154 8956 556160 8968
rect 176528 8928 556160 8956
rect 176528 8916 176534 8928
rect 556154 8916 556160 8928
rect 556212 8916 556218 8968
rect 150342 7828 150348 7880
rect 150400 7868 150406 7880
rect 227530 7868 227536 7880
rect 150400 7840 227536 7868
rect 150400 7828 150406 7840
rect 227530 7828 227536 7840
rect 227588 7828 227594 7880
rect 162486 7760 162492 7812
rect 162544 7800 162550 7812
rect 378870 7800 378876 7812
rect 162544 7772 378876 7800
rect 162544 7760 162550 7772
rect 378870 7760 378876 7772
rect 378928 7760 378934 7812
rect 162026 7692 162032 7744
rect 162084 7732 162090 7744
rect 390646 7732 390652 7744
rect 162084 7704 390652 7732
rect 162084 7692 162090 7704
rect 390646 7692 390652 7704
rect 390704 7692 390710 7744
rect 169754 7624 169760 7676
rect 169812 7664 169818 7676
rect 482830 7664 482836 7676
rect 169812 7636 482836 7664
rect 169812 7624 169818 7636
rect 482830 7624 482836 7636
rect 482888 7624 482894 7676
rect 24210 7556 24216 7608
rect 24268 7596 24274 7608
rect 134150 7596 134156 7608
rect 24268 7568 134156 7596
rect 24268 7556 24274 7568
rect 134150 7556 134156 7568
rect 134208 7556 134214 7608
rect 173894 7556 173900 7608
rect 173952 7596 173958 7608
rect 545482 7596 545488 7608
rect 173952 7568 545488 7596
rect 173952 7556 173958 7568
rect 545482 7556 545488 7568
rect 545540 7556 545546 7608
rect 576118 6808 576124 6860
rect 576176 6848 576182 6860
rect 580166 6848 580172 6860
rect 576176 6820 580172 6848
rect 576176 6808 576182 6820
rect 580166 6808 580172 6820
rect 580224 6808 580230 6860
rect 153838 6400 153844 6452
rect 153896 6440 153902 6452
rect 272426 6440 272432 6452
rect 153896 6412 272432 6440
rect 153896 6400 153902 6412
rect 272426 6400 272432 6412
rect 272484 6400 272490 6452
rect 158622 6332 158628 6384
rect 158680 6372 158686 6384
rect 336274 6372 336280 6384
rect 158680 6344 336280 6372
rect 158680 6332 158686 6344
rect 336274 6332 336280 6344
rect 336332 6332 336338 6384
rect 165430 6264 165436 6316
rect 165488 6304 165494 6316
rect 411898 6304 411904 6316
rect 165488 6276 411904 6304
rect 165488 6264 165494 6276
rect 411898 6264 411904 6276
rect 411956 6264 411962 6316
rect 165522 6196 165528 6248
rect 165580 6236 165586 6248
rect 414290 6236 414296 6248
rect 165580 6208 414296 6236
rect 165580 6196 165586 6208
rect 414290 6196 414296 6208
rect 414348 6196 414354 6248
rect 87966 6128 87972 6180
rect 88024 6168 88030 6180
rect 138014 6168 138020 6180
rect 88024 6140 138020 6168
rect 88024 6128 88030 6140
rect 138014 6128 138020 6140
rect 138072 6128 138078 6180
rect 143534 6128 143540 6180
rect 143592 6168 143598 6180
rect 155402 6168 155408 6180
rect 143592 6140 155408 6168
rect 143592 6128 143598 6140
rect 155402 6128 155408 6140
rect 155460 6128 155466 6180
rect 173802 6128 173808 6180
rect 173860 6168 173866 6180
rect 525426 6168 525432 6180
rect 173860 6140 525432 6168
rect 173860 6128 173866 6140
rect 525426 6128 525432 6140
rect 525484 6128 525490 6180
rect 154114 5040 154120 5092
rect 154172 5080 154178 5092
rect 273622 5080 273628 5092
rect 154172 5052 273628 5080
rect 154172 5040 154178 5052
rect 273622 5040 273628 5052
rect 273680 5040 273686 5092
rect 162578 4972 162584 5024
rect 162636 5012 162642 5024
rect 382366 5012 382372 5024
rect 162636 4984 382372 5012
rect 162636 4972 162642 4984
rect 382366 4972 382372 4984
rect 382424 4972 382430 5024
rect 180150 4904 180156 4956
rect 180208 4944 180214 4956
rect 429654 4944 429660 4956
rect 180208 4916 429660 4944
rect 180208 4904 180214 4916
rect 429654 4904 429660 4916
rect 429712 4904 429718 4956
rect 138842 4836 138848 4888
rect 138900 4876 138906 4888
rect 142246 4876 142252 4888
rect 138900 4848 142252 4876
rect 138900 4836 138906 4848
rect 142246 4836 142252 4848
rect 142304 4836 142310 4888
rect 170306 4836 170312 4888
rect 170364 4876 170370 4888
rect 486418 4876 486424 4888
rect 170364 4848 486424 4876
rect 170364 4836 170370 4848
rect 486418 4836 486424 4848
rect 486476 4836 486482 4888
rect 175182 4768 175188 4820
rect 175240 4808 175246 4820
rect 541986 4808 541992 4820
rect 175240 4780 541992 4808
rect 175240 4768 175246 4780
rect 541986 4768 541992 4780
rect 542044 4768 542050 4820
rect 566 4088 572 4140
rect 624 4128 630 4140
rect 7558 4128 7564 4140
rect 624 4100 7564 4128
rect 624 4088 630 4100
rect 7558 4088 7564 4100
rect 7616 4088 7622 4140
rect 73798 4088 73804 4140
rect 73856 4128 73862 4140
rect 75178 4128 75184 4140
rect 73856 4100 75184 4128
rect 73856 4088 73862 4100
rect 75178 4088 75184 4100
rect 75236 4088 75242 4140
rect 103330 4088 103336 4140
rect 103388 4128 103394 4140
rect 104158 4128 104164 4140
rect 103388 4100 104164 4128
rect 103388 4088 103394 4100
rect 104158 4088 104164 4100
rect 104216 4088 104222 4140
rect 146938 4088 146944 4140
rect 146996 4128 147002 4140
rect 147398 4128 147404 4140
rect 146996 4100 147404 4128
rect 146996 4088 147002 4100
rect 147398 4088 147404 4100
rect 147456 4088 147462 4140
rect 149698 4088 149704 4140
rect 149756 4128 149762 4140
rect 151814 4128 151820 4140
rect 149756 4100 151820 4128
rect 149756 4088 149762 4100
rect 151814 4088 151820 4100
rect 151872 4088 151878 4140
rect 196618 4088 196624 4140
rect 196676 4128 196682 4140
rect 203886 4128 203892 4140
rect 196676 4100 203892 4128
rect 196676 4088 196682 4100
rect 203886 4088 203892 4100
rect 203944 4088 203950 4140
rect 304258 4088 304264 4140
rect 304316 4128 304322 4140
rect 309042 4128 309048 4140
rect 304316 4100 309048 4128
rect 304316 4088 304322 4100
rect 309042 4088 309048 4100
rect 309100 4088 309106 4140
rect 450538 4088 450544 4140
rect 450596 4128 450602 4140
rect 450998 4128 451004 4140
rect 450596 4100 451004 4128
rect 450596 4088 450602 4100
rect 450998 4088 451004 4100
rect 451056 4088 451062 4140
rect 6454 4020 6460 4072
rect 6512 4060 6518 4072
rect 7650 4060 7656 4072
rect 6512 4032 7656 4060
rect 6512 4020 6518 4032
rect 7650 4020 7656 4032
rect 7708 4020 7714 4072
rect 180334 4020 180340 4072
rect 180392 4060 180398 4072
rect 186130 4060 186136 4072
rect 180392 4032 186136 4060
rect 180392 4020 180398 4032
rect 186130 4020 186136 4032
rect 186188 4020 186194 4072
rect 189810 4020 189816 4072
rect 189868 4060 189874 4072
rect 193214 4060 193220 4072
rect 189868 4032 193220 4060
rect 189868 4020 189874 4032
rect 193214 4020 193220 4032
rect 193272 4020 193278 4072
rect 193858 4020 193864 4072
rect 193916 4060 193922 4072
rect 196802 4060 196808 4072
rect 193916 4032 196808 4060
rect 193916 4020 193922 4032
rect 196802 4020 196808 4032
rect 196860 4020 196866 4072
rect 203702 4020 203708 4072
rect 203760 4060 203766 4072
rect 223942 4060 223948 4072
rect 203760 4032 223948 4060
rect 203760 4020 203766 4032
rect 223942 4020 223948 4032
rect 224000 4020 224006 4072
rect 224218 4020 224224 4072
rect 224276 4060 224282 4072
rect 240502 4060 240508 4072
rect 224276 4032 240508 4060
rect 224276 4020 224282 4032
rect 240502 4020 240508 4032
rect 240560 4020 240566 4072
rect 164878 3952 164884 4004
rect 164936 3992 164942 4004
rect 168374 3992 168380 4004
rect 164936 3964 168380 3992
rect 164936 3952 164942 3964
rect 168374 3952 168380 3964
rect 168432 3952 168438 4004
rect 181438 3952 181444 4004
rect 181496 3992 181502 4004
rect 226334 3992 226340 4004
rect 181496 3964 226340 3992
rect 181496 3952 181502 3964
rect 226334 3952 226340 3964
rect 226392 3952 226398 4004
rect 276014 3952 276020 4004
rect 276072 3992 276078 4004
rect 276750 3992 276756 4004
rect 276072 3964 276756 3992
rect 276072 3952 276078 3964
rect 276750 3952 276756 3964
rect 276808 3952 276814 4004
rect 299566 3952 299572 4004
rect 299624 3992 299630 4004
rect 300762 3992 300768 4004
rect 299624 3964 300768 3992
rect 299624 3952 299630 3964
rect 300762 3952 300768 3964
rect 300820 3952 300826 4004
rect 147122 3884 147128 3936
rect 147180 3924 147186 3936
rect 150618 3924 150624 3936
rect 147180 3896 150624 3924
rect 147180 3884 147186 3896
rect 150618 3884 150624 3896
rect 150676 3884 150682 3936
rect 155862 3884 155868 3936
rect 155920 3924 155926 3936
rect 306742 3924 306748 3936
rect 155920 3896 306748 3924
rect 155920 3884 155926 3896
rect 306742 3884 306748 3896
rect 306800 3884 306806 3936
rect 311158 3884 311164 3936
rect 311216 3924 311222 3936
rect 312630 3924 312636 3936
rect 311216 3896 312636 3924
rect 311216 3884 311222 3896
rect 312630 3884 312636 3896
rect 312688 3884 312694 3936
rect 44266 3816 44272 3868
rect 44324 3856 44330 3868
rect 46198 3856 46204 3868
rect 44324 3828 46204 3856
rect 44324 3816 44330 3828
rect 46198 3816 46204 3828
rect 46256 3816 46262 3868
rect 69106 3816 69112 3868
rect 69164 3856 69170 3868
rect 69164 3828 74534 3856
rect 69164 3816 69170 3828
rect 65518 3748 65524 3800
rect 65576 3788 65582 3800
rect 65576 3760 72648 3788
rect 65576 3748 65582 3760
rect 19426 3612 19432 3664
rect 19484 3652 19490 3664
rect 21358 3652 21364 3664
rect 19484 3624 21364 3652
rect 19484 3612 19490 3624
rect 21358 3612 21364 3624
rect 21416 3612 21422 3664
rect 43070 3612 43076 3664
rect 43128 3652 43134 3664
rect 44818 3652 44824 3664
rect 43128 3624 44824 3652
rect 43128 3612 43134 3624
rect 44818 3612 44824 3624
rect 44876 3612 44882 3664
rect 51350 3612 51356 3664
rect 51408 3652 51414 3664
rect 54478 3652 54484 3664
rect 51408 3624 54484 3652
rect 51408 3612 51414 3624
rect 54478 3612 54484 3624
rect 54536 3612 54542 3664
rect 70302 3612 70308 3664
rect 70360 3652 70366 3664
rect 72418 3652 72424 3664
rect 70360 3624 72424 3652
rect 70360 3612 70366 3624
rect 72418 3612 72424 3624
rect 72476 3612 72482 3664
rect 72620 3652 72648 3760
rect 74506 3720 74534 3828
rect 122282 3816 122288 3868
rect 122340 3856 122346 3868
rect 127618 3856 127624 3868
rect 122340 3828 127624 3856
rect 122340 3816 122346 3828
rect 127618 3816 127624 3828
rect 127676 3816 127682 3868
rect 147214 3816 147220 3868
rect 147272 3856 147278 3868
rect 163682 3856 163688 3868
rect 147272 3828 163688 3856
rect 147272 3816 147278 3828
rect 163682 3816 163688 3828
rect 163740 3816 163746 3868
rect 178678 3816 178684 3868
rect 178736 3856 178742 3868
rect 401318 3856 401324 3868
rect 178736 3828 401324 3856
rect 178736 3816 178742 3828
rect 401318 3816 401324 3828
rect 401376 3816 401382 3868
rect 111610 3748 111616 3800
rect 111668 3788 111674 3800
rect 131758 3788 131764 3800
rect 111668 3760 131764 3788
rect 111668 3748 111674 3760
rect 131758 3748 131764 3760
rect 131816 3748 131822 3800
rect 148318 3748 148324 3800
rect 148376 3788 148382 3800
rect 164878 3788 164884 3800
rect 148376 3760 164884 3788
rect 148376 3748 148382 3760
rect 164878 3748 164884 3760
rect 164936 3748 164942 3800
rect 170398 3748 170404 3800
rect 170456 3788 170462 3800
rect 174262 3788 174268 3800
rect 170456 3760 174268 3788
rect 170456 3748 170462 3760
rect 174262 3748 174268 3760
rect 174320 3748 174326 3800
rect 183462 3748 183468 3800
rect 183520 3788 183526 3800
rect 200298 3788 200304 3800
rect 183520 3760 200304 3788
rect 183520 3748 183526 3760
rect 200298 3748 200304 3760
rect 200356 3748 200362 3800
rect 200758 3748 200764 3800
rect 200816 3788 200822 3800
rect 210970 3788 210976 3800
rect 200816 3760 210976 3788
rect 200816 3748 200822 3760
rect 210970 3748 210976 3760
rect 211028 3748 211034 3800
rect 220078 3748 220084 3800
rect 220136 3788 220142 3800
rect 447410 3788 447416 3800
rect 220136 3760 447416 3788
rect 220136 3748 220142 3760
rect 447410 3748 447416 3760
rect 447468 3748 447474 3800
rect 453390 3748 453396 3800
rect 453448 3788 453454 3800
rect 497090 3788 497096 3800
rect 453448 3760 497096 3788
rect 453448 3748 453454 3760
rect 497090 3748 497096 3760
rect 497148 3748 497154 3800
rect 129826 3720 129832 3732
rect 74506 3692 129832 3720
rect 129826 3680 129832 3692
rect 129884 3680 129890 3732
rect 131022 3680 131028 3732
rect 131080 3720 131086 3732
rect 143534 3720 143540 3732
rect 131080 3692 143540 3720
rect 131080 3680 131086 3692
rect 143534 3680 143540 3692
rect 143592 3680 143598 3732
rect 148410 3680 148416 3732
rect 148468 3720 148474 3732
rect 170766 3720 170772 3732
rect 148468 3692 170772 3720
rect 148468 3680 148474 3692
rect 170766 3680 170772 3692
rect 170824 3680 170830 3732
rect 179230 3680 179236 3732
rect 179288 3720 179294 3732
rect 179288 3692 180196 3720
rect 179288 3680 179294 3692
rect 137278 3652 137284 3664
rect 72620 3624 137284 3652
rect 137278 3612 137284 3624
rect 137336 3612 137342 3664
rect 147030 3612 147036 3664
rect 147088 3652 147094 3664
rect 149514 3652 149520 3664
rect 147088 3624 149520 3652
rect 147088 3612 147094 3624
rect 149514 3612 149520 3624
rect 149572 3612 149578 3664
rect 171962 3652 171968 3664
rect 149624 3624 171968 3652
rect 7650 3544 7656 3596
rect 7708 3584 7714 3596
rect 129918 3584 129924 3596
rect 7708 3556 129924 3584
rect 7708 3544 7714 3556
rect 129918 3544 129924 3556
rect 129976 3544 129982 3596
rect 130930 3544 130936 3596
rect 130988 3584 130994 3596
rect 130988 3556 142154 3584
rect 130988 3544 130994 3556
rect 4062 3476 4068 3528
rect 4120 3516 4126 3528
rect 4798 3516 4804 3528
rect 4120 3488 4804 3516
rect 4120 3476 4126 3488
rect 4798 3476 4804 3488
rect 4856 3476 4862 3528
rect 5258 3476 5264 3528
rect 5316 3516 5322 3528
rect 5316 3488 126928 3516
rect 5316 3476 5322 3488
rect 8754 3408 8760 3460
rect 8812 3448 8818 3460
rect 10318 3448 10324 3460
rect 8812 3420 10324 3448
rect 8812 3408 8818 3420
rect 10318 3408 10324 3420
rect 10376 3408 10382 3460
rect 17034 3408 17040 3460
rect 17092 3448 17098 3460
rect 18598 3448 18604 3460
rect 17092 3420 18604 3448
rect 17092 3408 17098 3420
rect 18598 3408 18604 3420
rect 18656 3408 18662 3460
rect 20622 3408 20628 3460
rect 20680 3448 20686 3460
rect 20680 3420 126836 3448
rect 20680 3408 20686 3420
rect 27614 3340 27620 3392
rect 27672 3380 27678 3392
rect 28534 3380 28540 3392
rect 27672 3352 28540 3380
rect 27672 3340 27678 3352
rect 28534 3340 28540 3352
rect 28592 3340 28598 3392
rect 33594 3340 33600 3392
rect 33652 3380 33658 3392
rect 35158 3380 35164 3392
rect 33652 3352 35164 3380
rect 33652 3340 33658 3352
rect 35158 3340 35164 3352
rect 35216 3340 35222 3392
rect 41874 3340 41880 3392
rect 41932 3380 41938 3392
rect 43438 3380 43444 3392
rect 41932 3352 43444 3380
rect 41932 3340 41938 3352
rect 43438 3340 43444 3352
rect 43496 3340 43502 3392
rect 52454 3340 52460 3392
rect 52512 3380 52518 3392
rect 53374 3380 53380 3392
rect 52512 3352 53380 3380
rect 52512 3340 52518 3352
rect 53374 3340 53380 3352
rect 53432 3340 53438 3392
rect 60734 3340 60740 3392
rect 60792 3380 60798 3392
rect 61654 3380 61660 3392
rect 60792 3352 61660 3380
rect 60792 3340 60798 3352
rect 61654 3340 61660 3352
rect 61712 3340 61718 3392
rect 85574 3340 85580 3392
rect 85632 3380 85638 3392
rect 86494 3380 86500 3392
rect 85632 3352 86500 3380
rect 85632 3340 85638 3352
rect 86494 3340 86500 3352
rect 86552 3340 86558 3392
rect 91554 3340 91560 3392
rect 91612 3380 91618 3392
rect 93118 3380 93124 3392
rect 91612 3352 93124 3380
rect 91612 3340 91618 3352
rect 93118 3340 93124 3352
rect 93176 3340 93182 3392
rect 93854 3340 93860 3392
rect 93912 3380 93918 3392
rect 94774 3380 94780 3392
rect 93912 3352 94780 3380
rect 93912 3340 93918 3352
rect 94774 3340 94780 3352
rect 94832 3340 94838 3392
rect 101030 3340 101036 3392
rect 101088 3380 101094 3392
rect 102778 3380 102784 3392
rect 101088 3352 102784 3380
rect 101088 3340 101094 3352
rect 102778 3340 102784 3352
rect 102836 3340 102842 3392
rect 109310 3340 109316 3392
rect 109368 3380 109374 3392
rect 111150 3380 111156 3392
rect 109368 3352 111156 3380
rect 109368 3340 109374 3352
rect 111150 3340 111156 3352
rect 111208 3340 111214 3392
rect 119890 3340 119896 3392
rect 119948 3380 119954 3392
rect 120718 3380 120724 3392
rect 119948 3352 120724 3380
rect 119948 3340 119954 3352
rect 120718 3340 120724 3352
rect 120776 3340 120782 3392
rect 15930 3272 15936 3324
rect 15988 3312 15994 3324
rect 17218 3312 17224 3324
rect 15988 3284 17224 3312
rect 15988 3272 15994 3284
rect 17218 3272 17224 3284
rect 17276 3272 17282 3324
rect 83274 3272 83280 3324
rect 83332 3312 83338 3324
rect 84838 3312 84844 3324
rect 83332 3284 84844 3312
rect 83332 3272 83338 3284
rect 84838 3272 84844 3284
rect 84896 3272 84902 3324
rect 123478 3272 123484 3324
rect 123536 3312 123542 3324
rect 124858 3312 124864 3324
rect 123536 3284 124864 3312
rect 123536 3272 123542 3284
rect 124858 3272 124864 3284
rect 124916 3272 124922 3324
rect 126808 3312 126836 3420
rect 126900 3380 126928 3488
rect 126974 3476 126980 3528
rect 127032 3516 127038 3528
rect 128354 3516 128360 3528
rect 127032 3488 128360 3516
rect 127032 3476 127038 3488
rect 128354 3476 128360 3488
rect 128412 3476 128418 3528
rect 129366 3476 129372 3528
rect 129424 3516 129430 3528
rect 130010 3516 130016 3528
rect 129424 3488 130016 3516
rect 129424 3476 129430 3488
rect 130010 3476 130016 3488
rect 130068 3476 130074 3528
rect 137646 3476 137652 3528
rect 137704 3516 137710 3528
rect 138658 3516 138664 3528
rect 137704 3488 138664 3516
rect 137704 3476 137710 3488
rect 138658 3476 138664 3488
rect 138716 3476 138722 3528
rect 128170 3408 128176 3460
rect 128228 3448 128234 3460
rect 130378 3448 130384 3460
rect 128228 3420 130384 3448
rect 128228 3408 128234 3420
rect 130378 3408 130384 3420
rect 130436 3408 130442 3460
rect 131850 3380 131856 3392
rect 126900 3352 131856 3380
rect 131850 3340 131856 3352
rect 131908 3340 131914 3392
rect 142126 3380 142154 3556
rect 147306 3544 147312 3596
rect 147364 3584 147370 3596
rect 149624 3584 149652 3624
rect 171962 3612 171968 3624
rect 172020 3612 172026 3664
rect 180168 3652 180196 3692
rect 180242 3680 180248 3732
rect 180300 3720 180306 3732
rect 454494 3720 454500 3732
rect 180300 3692 454500 3720
rect 180300 3680 180306 3692
rect 454494 3680 454500 3692
rect 454552 3680 454558 3732
rect 180168 3624 180794 3652
rect 162486 3584 162492 3596
rect 147364 3556 149652 3584
rect 149808 3556 162492 3584
rect 147364 3544 147370 3556
rect 143442 3476 143448 3528
rect 143500 3516 143506 3528
rect 144730 3516 144736 3528
rect 143500 3488 144736 3516
rect 143500 3476 143506 3488
rect 144730 3476 144736 3488
rect 144788 3476 144794 3528
rect 149808 3380 149836 3556
rect 162486 3544 162492 3556
rect 162544 3544 162550 3596
rect 171870 3544 171876 3596
rect 171928 3584 171934 3596
rect 177850 3584 177856 3596
rect 171928 3556 177856 3584
rect 171928 3544 171934 3556
rect 177850 3544 177856 3556
rect 177908 3544 177914 3596
rect 180766 3584 180794 3624
rect 182082 3612 182088 3664
rect 182140 3652 182146 3664
rect 480530 3652 480536 3664
rect 182140 3624 480536 3652
rect 182140 3612 182146 3624
rect 480530 3612 480536 3624
rect 480588 3612 480594 3664
rect 486510 3612 486516 3664
rect 486568 3652 486574 3664
rect 518342 3652 518348 3664
rect 486568 3624 518348 3652
rect 486568 3612 486574 3624
rect 518342 3612 518348 3624
rect 518400 3612 518406 3664
rect 487614 3584 487620 3596
rect 180766 3556 487620 3584
rect 487614 3544 487620 3556
rect 487672 3544 487678 3596
rect 489914 3544 489920 3596
rect 489972 3584 489978 3596
rect 490742 3584 490748 3596
rect 489972 3556 490748 3584
rect 489972 3544 489978 3556
rect 490742 3544 490748 3556
rect 490800 3544 490806 3596
rect 504358 3544 504364 3596
rect 504416 3584 504422 3596
rect 505370 3584 505376 3596
rect 504416 3556 505376 3584
rect 504416 3544 504422 3556
rect 505370 3544 505376 3556
rect 505428 3544 505434 3596
rect 506474 3544 506480 3596
rect 506532 3584 506538 3596
rect 507302 3584 507308 3596
rect 506532 3556 507308 3584
rect 506532 3544 506538 3556
rect 507302 3544 507308 3556
rect 507360 3544 507366 3596
rect 520918 3544 520924 3596
rect 520976 3584 520982 3596
rect 524230 3584 524236 3596
rect 520976 3556 524236 3584
rect 520976 3544 520982 3556
rect 524230 3544 524236 3556
rect 524288 3544 524294 3596
rect 525058 3544 525064 3596
rect 525116 3584 525122 3596
rect 533706 3584 533712 3596
rect 525116 3556 533712 3584
rect 525116 3544 525122 3556
rect 533706 3544 533712 3556
rect 533764 3544 533770 3596
rect 572714 3584 572720 3596
rect 567166 3556 572720 3584
rect 151078 3476 151084 3528
rect 151136 3516 151142 3528
rect 151136 3488 171732 3516
rect 151136 3476 151142 3488
rect 171704 3448 171732 3488
rect 171778 3476 171784 3528
rect 171836 3516 171842 3528
rect 173158 3516 173164 3528
rect 171836 3488 173164 3516
rect 171836 3476 171842 3488
rect 173158 3476 173164 3488
rect 173216 3476 173222 3528
rect 179322 3476 179328 3528
rect 179380 3516 179386 3528
rect 531314 3516 531320 3528
rect 179380 3488 531320 3516
rect 179380 3476 179386 3488
rect 531314 3476 531320 3488
rect 531372 3476 531378 3528
rect 538858 3476 538864 3528
rect 538916 3516 538922 3528
rect 539594 3516 539600 3528
rect 538916 3488 539600 3516
rect 538916 3476 538922 3488
rect 539594 3476 539600 3488
rect 539652 3476 539658 3528
rect 545758 3476 545764 3528
rect 545816 3516 545822 3528
rect 551462 3516 551468 3528
rect 545816 3488 551468 3516
rect 545816 3476 545822 3488
rect 551462 3476 551468 3488
rect 551520 3476 551526 3528
rect 552750 3476 552756 3528
rect 552808 3516 552814 3528
rect 567166 3516 567194 3556
rect 572714 3544 572720 3556
rect 572772 3544 572778 3596
rect 574738 3544 574744 3596
rect 574796 3584 574802 3596
rect 576302 3584 576308 3596
rect 574796 3556 576308 3584
rect 574796 3544 574802 3556
rect 576302 3544 576308 3556
rect 576360 3544 576366 3596
rect 552808 3488 567194 3516
rect 552808 3476 552814 3488
rect 567838 3476 567844 3528
rect 567896 3516 567902 3528
rect 569126 3516 569132 3528
rect 567896 3488 569132 3516
rect 567896 3476 567902 3488
rect 569126 3476 569132 3488
rect 569184 3476 569190 3528
rect 175458 3448 175464 3460
rect 142126 3352 149836 3380
rect 151786 3420 161474 3448
rect 171704 3420 175464 3448
rect 131942 3312 131948 3324
rect 126808 3284 131948 3312
rect 131942 3272 131948 3284
rect 132000 3272 132006 3324
rect 132954 3272 132960 3324
rect 133012 3312 133018 3324
rect 141418 3312 141424 3324
rect 133012 3284 141424 3312
rect 133012 3272 133018 3284
rect 141418 3272 141424 3284
rect 141476 3272 141482 3324
rect 147398 3272 147404 3324
rect 147456 3312 147462 3324
rect 151786 3312 151814 3420
rect 156598 3340 156604 3392
rect 156656 3380 156662 3392
rect 157794 3380 157800 3392
rect 156656 3352 157800 3380
rect 156656 3340 156662 3352
rect 157794 3340 157800 3352
rect 157852 3340 157858 3392
rect 161446 3380 161474 3420
rect 175458 3408 175464 3420
rect 175516 3408 175522 3460
rect 580994 3448 581000 3460
rect 180766 3420 581000 3448
rect 176654 3380 176660 3392
rect 161446 3352 176660 3380
rect 176654 3340 176660 3352
rect 176712 3340 176718 3392
rect 180334 3340 180340 3392
rect 180392 3380 180398 3392
rect 180766 3380 180794 3420
rect 580994 3408 581000 3420
rect 581052 3408 581058 3460
rect 180392 3352 180794 3380
rect 180392 3340 180398 3352
rect 185578 3340 185584 3392
rect 185636 3380 185642 3392
rect 189718 3380 189724 3392
rect 185636 3352 189724 3380
rect 185636 3340 185642 3352
rect 189718 3340 189724 3352
rect 189776 3340 189782 3392
rect 217318 3340 217324 3392
rect 217376 3380 217382 3392
rect 218054 3380 218060 3392
rect 217376 3352 218060 3380
rect 217376 3340 217382 3352
rect 218054 3340 218060 3352
rect 218112 3340 218118 3392
rect 229738 3340 229744 3392
rect 229796 3380 229802 3392
rect 231026 3380 231032 3392
rect 229796 3352 231032 3380
rect 229796 3340 229802 3352
rect 231026 3340 231032 3352
rect 231084 3340 231090 3392
rect 324406 3340 324412 3392
rect 324464 3380 324470 3392
rect 325602 3380 325608 3392
rect 324464 3352 325608 3380
rect 324464 3340 324470 3352
rect 325602 3340 325608 3352
rect 325660 3340 325666 3392
rect 332594 3340 332600 3392
rect 332652 3380 332658 3392
rect 333882 3380 333888 3392
rect 332652 3352 333888 3380
rect 332652 3340 332658 3352
rect 333882 3340 333888 3352
rect 333940 3340 333946 3392
rect 349246 3340 349252 3392
rect 349304 3380 349310 3392
rect 350442 3380 350448 3392
rect 349304 3352 350448 3380
rect 349304 3340 349310 3352
rect 350442 3340 350448 3352
rect 350500 3340 350506 3392
rect 357526 3340 357532 3392
rect 357584 3380 357590 3392
rect 358722 3380 358728 3392
rect 357584 3352 358728 3380
rect 357584 3340 357590 3352
rect 358722 3340 358728 3352
rect 358780 3340 358786 3392
rect 364978 3340 364984 3392
rect 365036 3380 365042 3392
rect 367002 3380 367008 3392
rect 365036 3352 367008 3380
rect 365036 3340 365042 3352
rect 367002 3340 367008 3352
rect 367060 3340 367066 3392
rect 374086 3340 374092 3392
rect 374144 3380 374150 3392
rect 375282 3380 375288 3392
rect 374144 3352 375288 3380
rect 374144 3340 374150 3352
rect 375282 3340 375288 3352
rect 375340 3340 375346 3392
rect 382274 3340 382280 3392
rect 382332 3380 382338 3392
rect 383562 3380 383568 3392
rect 382332 3352 383568 3380
rect 382332 3340 382338 3352
rect 383562 3340 383568 3352
rect 383620 3340 383626 3392
rect 390554 3340 390560 3392
rect 390612 3380 390618 3392
rect 391842 3380 391848 3392
rect 390612 3352 391848 3380
rect 390612 3340 390618 3352
rect 391842 3340 391848 3352
rect 391900 3340 391906 3392
rect 398926 3340 398932 3392
rect 398984 3380 398990 3392
rect 400122 3380 400128 3392
rect 398984 3352 400128 3380
rect 398984 3340 398990 3352
rect 400122 3340 400128 3352
rect 400180 3340 400186 3392
rect 400950 3340 400956 3392
rect 401008 3380 401014 3392
rect 402514 3380 402520 3392
rect 401008 3352 402520 3380
rect 401008 3340 401014 3352
rect 402514 3340 402520 3352
rect 402572 3340 402578 3392
rect 407206 3340 407212 3392
rect 407264 3380 407270 3392
rect 408402 3380 408408 3392
rect 407264 3352 408408 3380
rect 407264 3340 407270 3352
rect 408402 3340 408408 3352
rect 408460 3340 408466 3392
rect 414658 3340 414664 3392
rect 414716 3380 414722 3392
rect 416682 3380 416688 3392
rect 414716 3352 416688 3380
rect 414716 3340 414722 3352
rect 416682 3340 416688 3352
rect 416740 3340 416746 3392
rect 418798 3340 418804 3392
rect 418856 3380 418862 3392
rect 420178 3380 420184 3392
rect 418856 3352 420184 3380
rect 418856 3340 418862 3352
rect 420178 3340 420184 3352
rect 420236 3340 420242 3392
rect 423674 3340 423680 3392
rect 423732 3380 423738 3392
rect 424962 3380 424968 3392
rect 423732 3352 424968 3380
rect 423732 3340 423738 3352
rect 424962 3340 424968 3352
rect 425020 3340 425026 3392
rect 432598 3340 432604 3392
rect 432656 3380 432662 3392
rect 434438 3380 434444 3392
rect 432656 3352 434444 3380
rect 432656 3340 432662 3352
rect 434438 3340 434444 3352
rect 434496 3340 434502 3392
rect 440234 3340 440240 3392
rect 440292 3380 440298 3392
rect 441522 3380 441528 3392
rect 440292 3352 441528 3380
rect 440292 3340 440298 3352
rect 441522 3340 441528 3352
rect 441580 3340 441586 3392
rect 448606 3340 448612 3392
rect 448664 3380 448670 3392
rect 449802 3380 449808 3392
rect 448664 3352 449808 3380
rect 448664 3340 448670 3352
rect 449802 3340 449808 3352
rect 449860 3340 449866 3392
rect 456794 3340 456800 3392
rect 456852 3380 456858 3392
rect 458082 3380 458088 3392
rect 456852 3352 458088 3380
rect 456852 3340 456858 3352
rect 458082 3340 458088 3352
rect 458140 3340 458146 3392
rect 464338 3340 464344 3392
rect 464396 3380 464402 3392
rect 466270 3380 466276 3392
rect 464396 3352 466276 3380
rect 464396 3340 464402 3352
rect 466270 3340 466276 3352
rect 466328 3340 466334 3392
rect 468478 3340 468484 3392
rect 468536 3380 468542 3392
rect 469858 3380 469864 3392
rect 468536 3352 469864 3380
rect 468536 3340 468542 3352
rect 469858 3340 469864 3352
rect 469916 3340 469922 3392
rect 472618 3340 472624 3392
rect 472676 3380 472682 3392
rect 473446 3380 473452 3392
rect 472676 3352 473452 3380
rect 472676 3340 472682 3352
rect 473446 3340 473452 3352
rect 473504 3340 473510 3392
rect 147456 3284 151814 3312
rect 147456 3272 147462 3284
rect 315298 3272 315304 3324
rect 315356 3312 315362 3324
rect 317322 3312 317328 3324
rect 315356 3284 317328 3312
rect 315356 3272 315362 3284
rect 317322 3272 317328 3284
rect 317380 3272 317386 3324
rect 431954 3272 431960 3324
rect 432012 3312 432018 3324
rect 433242 3312 433248 3324
rect 432012 3284 433248 3312
rect 432012 3272 432018 3284
rect 433242 3272 433248 3284
rect 433300 3272 433306 3324
rect 1670 3204 1676 3256
rect 1728 3244 1734 3256
rect 8938 3244 8944 3256
rect 1728 3216 8944 3244
rect 1728 3204 1734 3216
rect 8938 3204 8944 3216
rect 8996 3204 9002 3256
rect 136450 3204 136456 3256
rect 136508 3244 136514 3256
rect 140038 3244 140044 3256
rect 136508 3216 140044 3244
rect 136508 3204 136514 3216
rect 140038 3204 140044 3216
rect 140096 3204 140102 3256
rect 18230 3136 18236 3188
rect 18288 3176 18294 3188
rect 22738 3176 22744 3188
rect 18288 3148 22744 3176
rect 18288 3136 18294 3148
rect 22738 3136 22744 3148
rect 22796 3136 22802 3188
rect 30098 3136 30104 3188
rect 30156 3176 30162 3188
rect 31018 3176 31024 3188
rect 30156 3148 31024 3176
rect 30156 3136 30162 3148
rect 31018 3136 31024 3148
rect 31076 3136 31082 3188
rect 38378 3136 38384 3188
rect 38436 3176 38442 3188
rect 39298 3176 39304 3188
rect 38436 3148 39304 3176
rect 38436 3136 38442 3148
rect 39298 3136 39304 3148
rect 39356 3136 39362 3188
rect 125870 3136 125876 3188
rect 125928 3176 125934 3188
rect 131114 3176 131120 3188
rect 125928 3148 131120 3176
rect 125928 3136 125934 3148
rect 131114 3136 131120 3148
rect 131172 3136 131178 3188
rect 181530 3136 181536 3188
rect 181588 3176 181594 3188
rect 184934 3176 184940 3188
rect 181588 3148 184940 3176
rect 181588 3136 181594 3148
rect 184934 3136 184940 3148
rect 184992 3136 184998 3188
rect 324958 3136 324964 3188
rect 325016 3176 325022 3188
rect 326798 3176 326804 3188
rect 325016 3148 326804 3176
rect 325016 3136 325022 3148
rect 326798 3136 326804 3148
rect 326856 3136 326862 3188
rect 335998 3136 336004 3188
rect 336056 3176 336062 3188
rect 342162 3176 342168 3188
rect 336056 3148 342168 3176
rect 336056 3136 336062 3148
rect 342162 3136 342168 3148
rect 342220 3136 342226 3188
rect 382918 3136 382924 3188
rect 382976 3176 382982 3188
rect 384758 3176 384764 3188
rect 382976 3148 384764 3176
rect 382976 3136 382982 3148
rect 384758 3136 384764 3148
rect 384816 3136 384822 3188
rect 450998 3136 451004 3188
rect 451056 3176 451062 3188
rect 452102 3176 452108 3188
rect 451056 3148 452108 3176
rect 451056 3136 451062 3148
rect 452102 3136 452108 3148
rect 452160 3136 452166 3188
rect 511350 3136 511356 3188
rect 511408 3176 511414 3188
rect 514754 3176 514760 3188
rect 511408 3148 514760 3176
rect 511408 3136 511414 3148
rect 514754 3136 514760 3148
rect 514812 3136 514818 3188
rect 56042 3000 56048 3052
rect 56100 3040 56106 3052
rect 58618 3040 58624 3052
rect 56100 3012 58624 3040
rect 56100 3000 56106 3012
rect 58618 3000 58624 3012
rect 58676 3000 58682 3052
rect 118786 3000 118792 3052
rect 118844 3040 118850 3052
rect 122098 3040 122104 3052
rect 118844 3012 122104 3040
rect 118844 3000 118850 3012
rect 122098 3000 122104 3012
rect 122156 3000 122162 3052
rect 297358 3000 297364 3052
rect 297416 3040 297422 3052
rect 298462 3040 298468 3052
rect 297416 3012 298468 3040
rect 297416 3000 297422 3012
rect 298462 3000 298468 3012
rect 298520 3000 298526 3052
rect 514018 3000 514024 3052
rect 514076 3040 514082 3052
rect 515950 3040 515956 3052
rect 514076 3012 515956 3040
rect 514076 3000 514082 3012
rect 515950 3000 515956 3012
rect 516008 3000 516014 3052
rect 563698 3000 563704 3052
rect 563756 3040 563762 3052
rect 565630 3040 565636 3052
rect 563756 3012 565636 3040
rect 563756 3000 563762 3012
rect 565630 3000 565636 3012
rect 565688 3000 565694 3052
rect 571978 3000 571984 3052
rect 572036 3040 572042 3052
rect 573910 3040 573916 3052
rect 572036 3012 573916 3040
rect 572036 3000 572042 3012
rect 573910 3000 573916 3012
rect 573968 3000 573974 3052
rect 12342 2932 12348 2984
rect 12400 2972 12406 2984
rect 14458 2972 14464 2984
rect 12400 2944 14464 2972
rect 12400 2932 12406 2944
rect 14458 2932 14464 2944
rect 14516 2932 14522 2984
rect 149790 2864 149796 2916
rect 149848 2904 149854 2916
rect 154206 2904 154212 2916
rect 149848 2876 154212 2904
rect 149848 2864 149854 2876
rect 154206 2864 154212 2876
rect 154264 2864 154270 2916
rect 454678 2864 454684 2916
rect 454736 2904 454742 2916
rect 455690 2904 455696 2916
rect 454736 2876 455696 2904
rect 454736 2864 454742 2876
rect 455690 2864 455696 2876
rect 455748 2864 455754 2916
<< via1 >>
rect 157340 700680 157392 700732
rect 202788 700680 202840 700732
rect 89168 700612 89220 700664
rect 160744 700612 160796 700664
rect 72976 700544 73028 700596
rect 160100 700544 160152 700596
rect 157248 700476 157300 700528
rect 283840 700476 283892 700528
rect 8116 700408 8168 700460
rect 162124 700408 162176 700460
rect 153200 700340 153252 700392
rect 332508 700340 332560 700392
rect 525064 700340 525116 700392
rect 559656 700340 559708 700392
rect 149704 700272 149756 700324
rect 543464 700272 543516 700324
rect 24308 699660 24360 699712
rect 25504 699660 25556 699712
rect 105452 699660 105504 699712
rect 106924 699660 106976 699712
rect 137836 699660 137888 699712
rect 140044 699660 140096 699712
rect 265624 699660 265676 699712
rect 267648 699660 267700 699712
rect 396724 699660 396776 699712
rect 397460 699660 397512 699712
rect 428464 699660 428516 699712
rect 429844 699660 429896 699712
rect 146576 696940 146628 696992
rect 580172 696940 580224 696992
rect 148324 683136 148376 683188
rect 580172 683136 580224 683188
rect 3332 670760 3384 670812
rect 164884 670760 164936 670812
rect 146944 670692 146996 670744
rect 580172 670692 580224 670744
rect 3516 658112 3568 658164
rect 7564 658112 7616 658164
rect 144920 643084 144972 643136
rect 580172 643084 580224 643136
rect 3516 632068 3568 632120
rect 164240 632068 164292 632120
rect 147036 630640 147088 630692
rect 580172 630640 580224 630692
rect 3516 618264 3568 618316
rect 166264 618264 166316 618316
rect 145564 616836 145616 616888
rect 580172 616836 580224 616888
rect 3516 605820 3568 605872
rect 166356 605820 166408 605872
rect 157616 605072 157668 605124
rect 169760 605072 169812 605124
rect 143724 590656 143776 590708
rect 579804 590656 579856 590708
rect 3332 579640 3384 579692
rect 165620 579640 165672 579692
rect 143816 576852 143868 576904
rect 580172 576852 580224 576904
rect 3240 565836 3292 565888
rect 167644 565836 167696 565888
rect 144184 563048 144236 563100
rect 579804 563048 579856 563100
rect 3332 553392 3384 553444
rect 167736 553392 167788 553444
rect 142160 536800 142212 536852
rect 580172 536800 580224 536852
rect 2780 527144 2832 527196
rect 4804 527144 4856 527196
rect 142252 524424 142304 524476
rect 580172 524424 580224 524476
rect 3516 514768 3568 514820
rect 10324 514768 10376 514820
rect 180064 510620 180116 510672
rect 580172 510620 580224 510672
rect 3056 500964 3108 501016
rect 152464 500964 152516 501016
rect 181444 484372 181496 484424
rect 580172 484372 580224 484424
rect 3056 474716 3108 474768
rect 169760 474716 169812 474768
rect 192484 470568 192536 470620
rect 579988 470568 580040 470620
rect 3516 462340 3568 462392
rect 171784 462340 171836 462392
rect 178684 456764 178736 456816
rect 580172 456764 580224 456816
rect 3148 448536 3200 448588
rect 170404 448536 170456 448588
rect 138020 430584 138072 430636
rect 580172 430584 580224 430636
rect 3516 422288 3568 422340
rect 171140 422288 171192 422340
rect 140136 418140 140188 418192
rect 580172 418140 580224 418192
rect 2872 409844 2924 409896
rect 13084 409844 13136 409896
rect 138664 404336 138716 404388
rect 580172 404336 580224 404388
rect 3516 397468 3568 397520
rect 171876 397468 171928 397520
rect 185584 378156 185636 378208
rect 580172 378156 580224 378208
rect 3516 371288 3568 371340
rect 8944 371288 8996 371340
rect 3148 357416 3200 357468
rect 174544 357416 174596 357468
rect 140228 351908 140280 351960
rect 580172 351908 580224 351960
rect 3332 345040 3384 345092
rect 173900 345040 173952 345092
rect 135536 324300 135588 324352
rect 580172 324300 580224 324352
rect 3332 318792 3384 318844
rect 173992 318792 174044 318844
rect 135904 311856 135956 311908
rect 579988 311856 580040 311908
rect 3516 304988 3568 305040
rect 175924 304988 175976 305040
rect 135996 298120 136048 298172
rect 580172 298120 580224 298172
rect 3516 292544 3568 292596
rect 176016 292544 176068 292596
rect 13084 286288 13136 286340
rect 173164 286288 173216 286340
rect 25504 284928 25556 284980
rect 163504 284928 163556 284980
rect 141424 283568 141476 283620
rect 192484 283568 192536 283620
rect 137284 282140 137336 282192
rect 185584 282140 185636 282192
rect 186412 280780 186464 280832
rect 396724 280780 396776 280832
rect 151820 280168 151872 280220
rect 186412 280168 186464 280220
rect 151084 279420 151136 279472
rect 462320 279420 462372 279472
rect 149244 277992 149296 278044
rect 527180 277992 527232 278044
rect 40040 276632 40092 276684
rect 161480 276632 161532 276684
rect 10324 275272 10376 275324
rect 169116 275272 169168 275324
rect 186688 275272 186740 275324
rect 364340 275272 364392 275324
rect 153384 274660 153436 274712
rect 186504 274660 186556 274712
rect 186688 274660 186740 274712
rect 7564 273912 7616 273964
rect 163596 273912 163648 273964
rect 187700 273912 187752 273964
rect 234620 273912 234672 273964
rect 155960 273232 156012 273284
rect 187700 273232 187752 273284
rect 152464 272484 152516 272536
rect 169024 272484 169076 272536
rect 134524 271872 134576 271924
rect 580172 271872 580224 271924
rect 140044 271124 140096 271176
rect 158720 271124 158772 271176
rect 8944 269832 8996 269884
rect 172520 269832 172572 269884
rect 149152 269764 149204 269816
rect 494060 269764 494112 269816
rect 106924 268404 106976 268456
rect 160192 268404 160244 268456
rect 147680 268336 147732 268388
rect 525064 268336 525116 268388
rect 141056 266976 141108 267028
rect 181444 266976 181496 267028
rect 3056 266364 3108 266416
rect 176660 266364 176712 266416
rect 171692 265752 171744 265804
rect 176108 265752 176160 265804
rect 141608 265684 141660 265736
rect 180064 265684 180116 265736
rect 3424 265616 3476 265668
rect 163504 265616 163556 265668
rect 176016 265616 176068 265668
rect 192300 265616 192352 265668
rect 175924 265548 175976 265600
rect 196440 265548 196492 265600
rect 171968 265480 172020 265532
rect 193864 265480 193916 265532
rect 173164 265412 173216 265464
rect 196256 265412 196308 265464
rect 174544 265344 174596 265396
rect 197728 265344 197780 265396
rect 169116 265276 169168 265328
rect 169576 265276 169628 265328
rect 193588 265276 193640 265328
rect 175832 265208 175884 265260
rect 176016 265208 176068 265260
rect 176108 265208 176160 265260
rect 197636 265208 197688 265260
rect 164884 265140 164936 265192
rect 195152 265140 195204 265192
rect 153292 265072 153344 265124
rect 158812 265072 158864 265124
rect 160744 265072 160796 265124
rect 161296 265072 161348 265124
rect 193220 265072 193272 265124
rect 190460 265004 190512 265056
rect 114284 264936 114336 264988
rect 135904 264936 135956 264988
rect 156328 264936 156380 264988
rect 157248 264936 157300 264988
rect 158812 264936 158864 264988
rect 159640 264936 159692 264988
rect 193772 264936 193824 264988
rect 119160 264392 119212 264444
rect 145564 264392 145616 264444
rect 139768 264324 139820 264376
rect 118148 264256 118200 264308
rect 137192 264256 137244 264308
rect 178684 264256 178736 264308
rect 4804 264188 4856 264240
rect 168380 264188 168432 264240
rect 188252 264188 188304 264240
rect 299480 264188 299532 264240
rect 117136 264120 117188 264172
rect 133972 264120 134024 264172
rect 134524 264120 134576 264172
rect 119804 264052 119856 264104
rect 138664 264052 138716 264104
rect 117044 263984 117096 264036
rect 135352 263984 135404 264036
rect 135996 263984 136048 264036
rect 137100 263984 137152 264036
rect 141056 263984 141108 264036
rect 119620 263916 119672 263968
rect 141608 263916 141660 263968
rect 114192 263848 114244 263900
rect 137284 263848 137336 263900
rect 121000 263780 121052 263832
rect 143632 263780 143684 263832
rect 144184 263780 144236 263832
rect 118332 263712 118384 263764
rect 137100 263712 137152 263764
rect 137192 263712 137244 263764
rect 140228 263712 140280 263764
rect 176660 263712 176712 263764
rect 190920 263712 190972 263764
rect 121092 263644 121144 263696
rect 139768 263644 139820 263696
rect 140320 263644 140372 263696
rect 168380 263644 168432 263696
rect 189264 263644 189316 263696
rect 120908 263576 120960 263628
rect 149152 263576 149204 263628
rect 149980 263576 150032 263628
rect 155224 263576 155276 263628
rect 188252 263576 188304 263628
rect 138296 263508 138348 263560
rect 580264 263508 580316 263560
rect 151820 263440 151872 263492
rect 152188 263440 152240 263492
rect 187976 263440 188028 263492
rect 347780 263440 347832 263492
rect 146392 263168 146444 263220
rect 147036 263168 147088 263220
rect 112444 263032 112496 263084
rect 131212 263032 131264 263084
rect 133696 263032 133748 263084
rect 580356 263032 580408 263084
rect 115204 262964 115256 263016
rect 132592 262964 132644 263016
rect 133788 262964 133840 263016
rect 3424 262896 3476 262948
rect 178776 262896 178828 262948
rect 180432 262896 180484 262948
rect 187148 262896 187200 262948
rect 118056 262828 118108 262880
rect 133144 262828 133196 262880
rect 178132 262828 178184 262880
rect 189632 262828 189684 262880
rect 191748 262828 191800 262880
rect 218060 262828 218112 262880
rect 111064 262760 111116 262812
rect 129740 262760 129792 262812
rect 133788 262760 133840 262812
rect 580448 262760 580500 262812
rect 116952 262692 117004 262744
rect 128452 262692 128504 262744
rect 170404 262692 170456 262744
rect 192484 262692 192536 262744
rect 117964 262624 118016 262676
rect 146392 262624 146444 262676
rect 169024 262624 169076 262676
rect 193680 262624 193732 262676
rect 120632 262556 120684 262608
rect 150440 262556 150492 262608
rect 158352 262556 158404 262608
rect 190828 262556 190880 262608
rect 191748 262556 191800 262608
rect 119436 262488 119488 262540
rect 149704 262488 149756 262540
rect 155040 262488 155092 262540
rect 187976 262488 188028 262540
rect 3516 262420 3568 262472
rect 177764 262420 177816 262472
rect 180616 262420 180668 262472
rect 192208 262420 192260 262472
rect 117872 262352 117924 262404
rect 130108 262352 130160 262404
rect 183192 262352 183244 262404
rect 196532 262352 196584 262404
rect 119528 262284 119580 262336
rect 125140 262284 125192 262336
rect 121184 262216 121236 262268
rect 126980 262216 127032 262268
rect 182088 262216 182140 262268
rect 187056 262216 187108 262268
rect 181536 261332 181588 261384
rect 192668 261332 192720 261384
rect 133144 261264 133196 261316
rect 133696 261264 133748 261316
rect 472624 261264 472676 261316
rect 4804 261196 4856 261248
rect 178132 261196 178184 261248
rect 116768 261128 116820 261180
rect 131120 261128 131172 261180
rect 178684 261128 178736 261180
rect 192576 261196 192628 261248
rect 112352 261060 112404 261112
rect 135168 261060 135220 261112
rect 187792 261060 187844 261112
rect 120540 260992 120592 261044
rect 178684 260992 178736 261044
rect 178776 260992 178828 261044
rect 179512 260992 179564 261044
rect 196624 260992 196676 261044
rect 177764 260924 177816 260976
rect 196716 260924 196768 260976
rect 113824 260856 113876 260908
rect 130660 260856 130712 260908
rect 184848 260856 184900 260908
rect 196348 260856 196400 260908
rect 175188 260448 175240 260500
rect 189540 260448 189592 260500
rect 157340 260380 157392 260432
rect 191104 260380 191156 260432
rect 7564 260312 7616 260364
rect 177028 260312 177080 260364
rect 182640 260312 182692 260364
rect 192392 260312 192444 260364
rect 131120 260244 131172 260296
rect 132040 260244 132092 260296
rect 471244 260244 471296 260296
rect 146576 260176 146628 260228
rect 147542 260176 147594 260228
rect 147680 260176 147732 260228
rect 148646 260176 148698 260228
rect 153200 260176 153252 260228
rect 154166 260176 154218 260228
rect 157616 260176 157668 260228
rect 158582 260176 158634 260228
rect 165620 260176 165672 260228
rect 166862 260176 166914 260228
rect 170174 260176 170226 260228
rect 189448 260176 189500 260228
rect 171140 260108 171192 260160
rect 171830 260108 171882 260160
rect 172520 260108 172572 260160
rect 173486 260108 173538 260160
rect 173992 260108 174044 260160
rect 175142 260108 175194 260160
rect 123484 260040 123536 260092
rect 116584 259972 116636 260024
rect 113916 259904 113968 259956
rect 127348 259904 127400 259956
rect 115388 259836 115440 259888
rect 123484 259836 123536 259888
rect 116676 259768 116728 259820
rect 124220 259768 124272 259820
rect 186964 260108 187016 260160
rect 184940 259972 184992 260024
rect 189816 259972 189868 260024
rect 187884 259904 187936 259956
rect 135536 259836 135588 259888
rect 167000 259836 167052 259888
rect 186688 259836 186740 259888
rect 142160 259768 142212 259820
rect 160560 259768 160612 259820
rect 186780 259768 186832 259820
rect 118240 259700 118292 259752
rect 146576 259700 146628 259752
rect 158720 259700 158772 259752
rect 188068 259700 188120 259752
rect 119344 259632 119396 259684
rect 147680 259632 147732 259684
rect 159456 259632 159508 259684
rect 191012 259632 191064 259684
rect 119252 259564 119304 259616
rect 153200 259564 153252 259616
rect 174360 259564 174412 259616
rect 184940 259564 184992 259616
rect 115296 259496 115348 259548
rect 124588 259496 124640 259548
rect 177672 259496 177724 259548
rect 189908 259564 189960 259616
rect 185308 259496 185360 259548
rect 187240 259496 187292 259548
rect 115112 259428 115164 259480
rect 129004 259428 129056 259480
rect 184296 259428 184348 259480
rect 195060 259428 195112 259480
rect 120816 259360 120868 259412
rect 123484 259360 123536 259412
rect 187792 259360 187844 259412
rect 580172 259360 580224 259412
rect 183652 259292 183704 259344
rect 188252 259292 188304 259344
rect 187792 259224 187844 259276
rect 188344 259224 188396 259276
rect 472624 245556 472676 245608
rect 580172 245556 580224 245608
rect 3516 241068 3568 241120
rect 7564 241068 7616 241120
rect 2780 215228 2832 215280
rect 4804 215228 4856 215280
rect 471244 206932 471296 206984
rect 579804 206932 579856 206984
rect 106924 199860 106976 199912
rect 131304 199860 131356 199912
rect 132040 199860 132092 199912
rect 132546 199860 132598 199912
rect 134110 199860 134162 199912
rect 134294 199860 134346 199912
rect 135030 199860 135082 199912
rect 131948 199792 132000 199844
rect 132822 199792 132874 199844
rect 133834 199792 133886 199844
rect 133650 199724 133702 199776
rect 133742 199724 133794 199776
rect 131672 199656 131724 199708
rect 104440 199452 104492 199504
rect 133420 199588 133472 199640
rect 133788 199588 133840 199640
rect 134018 199792 134070 199844
rect 134064 199656 134116 199708
rect 133880 199520 133932 199572
rect 133604 199452 133656 199504
rect 134846 199724 134898 199776
rect 135214 199860 135266 199912
rect 135490 199860 135542 199912
rect 135582 199860 135634 199912
rect 135674 199860 135726 199912
rect 135950 199860 136002 199912
rect 136410 199860 136462 199912
rect 136502 199860 136554 199912
rect 136870 199860 136922 199912
rect 136962 199860 137014 199912
rect 137054 199860 137106 199912
rect 137238 199860 137290 199912
rect 135398 199792 135450 199844
rect 135260 199724 135312 199776
rect 135076 199588 135128 199640
rect 135260 199588 135312 199640
rect 135444 199656 135496 199708
rect 135536 199656 135588 199708
rect 135766 199792 135818 199844
rect 135812 199656 135864 199708
rect 136134 199792 136186 199844
rect 136226 199792 136278 199844
rect 136318 199792 136370 199844
rect 135720 199588 135772 199640
rect 135996 199588 136048 199640
rect 136088 199588 136140 199640
rect 135904 199520 135956 199572
rect 136180 199520 136232 199572
rect 134340 199452 134392 199504
rect 136778 199792 136830 199844
rect 136548 199724 136600 199776
rect 136456 199656 136508 199708
rect 136916 199724 136968 199776
rect 137100 199656 137152 199708
rect 137606 199860 137658 199912
rect 137790 199860 137842 199912
rect 137974 199860 138026 199912
rect 138250 199860 138302 199912
rect 138342 199860 138394 199912
rect 138710 199860 138762 199912
rect 139262 199860 139314 199912
rect 137330 199724 137382 199776
rect 136732 199588 136784 199640
rect 137008 199588 137060 199640
rect 137284 199588 137336 199640
rect 137928 199656 137980 199708
rect 138020 199656 138072 199708
rect 138296 199588 138348 199640
rect 138388 199520 138440 199572
rect 139630 199860 139682 199912
rect 139906 199860 139958 199912
rect 140826 199860 140878 199912
rect 141102 199860 141154 199912
rect 141562 199860 141614 199912
rect 141654 199860 141706 199912
rect 141838 199860 141890 199912
rect 139584 199724 139636 199776
rect 140780 199724 140832 199776
rect 139216 199588 139268 199640
rect 139860 199588 139912 199640
rect 136456 199452 136508 199504
rect 136640 199452 136692 199504
rect 137468 199452 137520 199504
rect 138020 199452 138072 199504
rect 140044 199452 140096 199504
rect 141608 199656 141660 199708
rect 141700 199588 141752 199640
rect 140688 199520 140740 199572
rect 136364 199384 136416 199436
rect 140412 199384 140464 199436
rect 140872 199452 140924 199504
rect 141792 199452 141844 199504
rect 142206 199860 142258 199912
rect 142390 199860 142442 199912
rect 142758 199860 142810 199912
rect 142712 199724 142764 199776
rect 142436 199656 142488 199708
rect 142252 199588 142304 199640
rect 143126 199860 143178 199912
rect 143218 199860 143270 199912
rect 143402 199860 143454 199912
rect 143494 199860 143546 199912
rect 143678 199860 143730 199912
rect 144046 199860 144098 199912
rect 144230 199860 144282 199912
rect 144322 199860 144374 199912
rect 144874 199860 144926 199912
rect 143172 199724 143224 199776
rect 143356 199588 143408 199640
rect 143632 199588 143684 199640
rect 143448 199520 143500 199572
rect 144276 199656 144328 199708
rect 144184 199588 144236 199640
rect 144828 199588 144880 199640
rect 145426 199860 145478 199912
rect 145518 199860 145570 199912
rect 145794 199860 145846 199912
rect 145978 199860 146030 199912
rect 145242 199792 145294 199844
rect 145334 199792 145386 199844
rect 145288 199656 145340 199708
rect 145380 199656 145432 199708
rect 145748 199724 145800 199776
rect 145564 199588 145616 199640
rect 144552 199520 144604 199572
rect 144000 199452 144052 199504
rect 112996 199316 113048 199368
rect 115756 199248 115808 199300
rect 140044 199248 140096 199300
rect 147358 199860 147410 199912
rect 147542 199860 147594 199912
rect 148094 199860 148146 199912
rect 148278 199860 148330 199912
rect 148140 199724 148192 199776
rect 147680 199588 147732 199640
rect 148232 199520 148284 199572
rect 148646 199860 148698 199912
rect 148738 199860 148790 199912
rect 148830 199860 148882 199912
rect 148922 199860 148974 199912
rect 149106 199860 149158 199912
rect 149198 199860 149250 199912
rect 149382 199860 149434 199912
rect 149658 199860 149710 199912
rect 148692 199724 148744 199776
rect 148784 199724 148836 199776
rect 149060 199724 149112 199776
rect 149152 199724 149204 199776
rect 149244 199724 149296 199776
rect 148876 199656 148928 199708
rect 149336 199656 149388 199708
rect 149842 199656 149894 199708
rect 149520 199588 149572 199640
rect 150026 199860 150078 199912
rect 150118 199860 150170 199912
rect 150762 199860 150814 199912
rect 151222 199860 151274 199912
rect 151406 199860 151458 199912
rect 151590 199860 151642 199912
rect 151682 199860 151734 199912
rect 151958 199860 152010 199912
rect 152050 199860 152102 199912
rect 152418 199860 152470 199912
rect 152602 199860 152654 199912
rect 152970 199860 153022 199912
rect 153246 199860 153298 199912
rect 150394 199724 150446 199776
rect 150072 199656 150124 199708
rect 151176 199724 151228 199776
rect 150348 199588 150400 199640
rect 150808 199588 150860 199640
rect 151636 199656 151688 199708
rect 151084 199588 151136 199640
rect 151452 199520 151504 199572
rect 151544 199520 151596 199572
rect 147496 199452 147548 199504
rect 149888 199452 149940 199504
rect 152464 199588 152516 199640
rect 152188 199452 152240 199504
rect 152832 199520 152884 199572
rect 153338 199792 153390 199844
rect 153200 199452 153252 199504
rect 153292 199452 153344 199504
rect 153522 199860 153574 199912
rect 153614 199860 153666 199912
rect 153982 199860 154034 199912
rect 154074 199860 154126 199912
rect 154166 199860 154218 199912
rect 154258 199860 154310 199912
rect 154534 199860 154586 199912
rect 154626 199860 154678 199912
rect 154902 199860 154954 199912
rect 155086 199860 155138 199912
rect 155178 199860 155230 199912
rect 155270 199860 155322 199912
rect 153568 199724 153620 199776
rect 154120 199724 154172 199776
rect 154212 199724 154264 199776
rect 154028 199656 154080 199708
rect 154488 199724 154540 199776
rect 154580 199724 154632 199776
rect 153660 199588 153712 199640
rect 154304 199588 154356 199640
rect 155132 199724 155184 199776
rect 155224 199724 155276 199776
rect 155040 199588 155092 199640
rect 155546 199860 155598 199912
rect 156190 199860 156242 199912
rect 156282 199860 156334 199912
rect 156374 199860 156426 199912
rect 156742 199860 156794 199912
rect 157018 199860 157070 199912
rect 157110 199860 157162 199912
rect 157386 199860 157438 199912
rect 157570 199860 157622 199912
rect 157662 199860 157714 199912
rect 157754 199860 157806 199912
rect 157938 199860 157990 199912
rect 158398 199860 158450 199912
rect 158766 199860 158818 199912
rect 158950 199860 159002 199912
rect 159410 199860 159462 199912
rect 159502 199860 159554 199912
rect 160330 199860 160382 199912
rect 160422 199860 160474 199912
rect 160606 199860 160658 199912
rect 156236 199724 156288 199776
rect 156328 199724 156380 199776
rect 156420 199656 156472 199708
rect 157064 199724 157116 199776
rect 157156 199656 157208 199708
rect 156696 199588 156748 199640
rect 155408 199520 155460 199572
rect 155592 199520 155644 199572
rect 153384 199384 153436 199436
rect 157708 199656 157760 199708
rect 158352 199724 158404 199776
rect 157892 199588 157944 199640
rect 158904 199588 158956 199640
rect 158260 199520 158312 199572
rect 158812 199520 158864 199572
rect 159180 199520 159232 199572
rect 160238 199792 160290 199844
rect 159456 199724 159508 199776
rect 160192 199656 160244 199708
rect 160284 199588 160336 199640
rect 160468 199588 160520 199640
rect 157708 199452 157760 199504
rect 158536 199316 158588 199368
rect 161894 199860 161946 199912
rect 161986 199860 162038 199912
rect 162170 199860 162222 199912
rect 162262 199860 162314 199912
rect 162354 199860 162406 199912
rect 162446 199860 162498 199912
rect 162538 199860 162590 199912
rect 162814 199860 162866 199912
rect 160974 199792 161026 199844
rect 161526 199792 161578 199844
rect 161158 199724 161210 199776
rect 161250 199724 161302 199776
rect 160928 199656 160980 199708
rect 160836 199520 160888 199572
rect 161940 199724 161992 199776
rect 162216 199656 162268 199708
rect 162308 199656 162360 199708
rect 163090 199792 163142 199844
rect 163182 199792 163234 199844
rect 162584 199724 162636 199776
rect 162906 199724 162958 199776
rect 162492 199656 162544 199708
rect 162124 199588 162176 199640
rect 163136 199656 163188 199708
rect 163044 199588 163096 199640
rect 163366 199860 163418 199912
rect 163550 199860 163602 199912
rect 163642 199860 163694 199912
rect 163412 199656 163464 199708
rect 163826 199792 163878 199844
rect 163688 199724 163740 199776
rect 163504 199588 163556 199640
rect 161296 199520 161348 199572
rect 161480 199520 161532 199572
rect 162952 199520 163004 199572
rect 163320 199520 163372 199572
rect 163596 199520 163648 199572
rect 164010 199860 164062 199912
rect 164102 199860 164154 199912
rect 164194 199860 164246 199912
rect 164286 199860 164338 199912
rect 164378 199860 164430 199912
rect 164470 199860 164522 199912
rect 164056 199656 164108 199708
rect 164148 199656 164200 199708
rect 164562 199792 164614 199844
rect 164424 199656 164476 199708
rect 164516 199656 164568 199708
rect 164240 199588 164292 199640
rect 164838 199860 164890 199912
rect 164930 199860 164982 199912
rect 165022 199860 165074 199912
rect 165114 199860 165166 199912
rect 165482 199860 165534 199912
rect 165850 199860 165902 199912
rect 166034 199860 166086 199912
rect 166126 199860 166178 199912
rect 166218 199860 166270 199912
rect 166310 199860 166362 199912
rect 166494 199860 166546 199912
rect 166862 199860 166914 199912
rect 167230 199860 167282 199912
rect 167414 199860 167466 199912
rect 167506 199860 167558 199912
rect 167598 199860 167650 199912
rect 164792 199724 164844 199776
rect 164884 199656 164936 199708
rect 164976 199656 165028 199708
rect 165068 199656 165120 199708
rect 165666 199792 165718 199844
rect 165482 199588 165534 199640
rect 165712 199588 165764 199640
rect 164700 199520 164752 199572
rect 166080 199656 166132 199708
rect 166172 199656 166224 199708
rect 165988 199588 166040 199640
rect 166356 199588 166408 199640
rect 166678 199792 166730 199844
rect 166770 199792 166822 199844
rect 167138 199792 167190 199844
rect 166908 199724 166960 199776
rect 166816 199656 166868 199708
rect 166724 199588 166776 199640
rect 167276 199588 167328 199640
rect 166264 199520 166316 199572
rect 166540 199520 166592 199572
rect 167184 199520 167236 199572
rect 163872 199452 163924 199504
rect 165436 199384 165488 199436
rect 166264 199316 166316 199368
rect 167460 199520 167512 199572
rect 167966 199860 168018 199912
rect 168334 199860 168386 199912
rect 168518 199860 168570 199912
rect 168702 199860 168754 199912
rect 168978 199860 169030 199912
rect 169070 199860 169122 199912
rect 169162 199860 169214 199912
rect 169346 199860 169398 199912
rect 169438 199860 169490 199912
rect 168150 199792 168202 199844
rect 168288 199656 168340 199708
rect 168196 199588 168248 199640
rect 168748 199588 168800 199640
rect 168472 199520 168524 199572
rect 168932 199656 168984 199708
rect 169208 199588 169260 199640
rect 169300 199588 169352 199640
rect 169990 199860 170042 199912
rect 170082 199860 170134 199912
rect 170174 199860 170226 199912
rect 170266 199860 170318 199912
rect 170450 199860 170502 199912
rect 169806 199792 169858 199844
rect 169668 199588 169720 199640
rect 169116 199520 169168 199572
rect 169392 199520 169444 199572
rect 170036 199656 170088 199708
rect 170128 199588 170180 199640
rect 170220 199588 170272 199640
rect 169944 199520 169996 199572
rect 170726 199860 170778 199912
rect 170818 199860 170870 199912
rect 170910 199860 170962 199912
rect 171094 199860 171146 199912
rect 171278 199860 171330 199912
rect 171370 199860 171422 199912
rect 171462 199860 171514 199912
rect 171646 199860 171698 199912
rect 171738 199860 171790 199912
rect 171830 199860 171882 199912
rect 171922 199860 171974 199912
rect 172014 199860 172066 199912
rect 172198 199860 172250 199912
rect 172382 199860 172434 199912
rect 172566 199860 172618 199912
rect 172658 199860 172710 199912
rect 172750 199860 172802 199912
rect 172934 199860 172986 199912
rect 173026 199860 173078 199912
rect 173118 199860 173170 199912
rect 170772 199724 170824 199776
rect 170588 199588 170640 199640
rect 170680 199520 170732 199572
rect 167920 199384 167972 199436
rect 167644 199316 167696 199368
rect 151360 199248 151412 199300
rect 162400 199248 162452 199300
rect 167552 199248 167604 199300
rect 170036 199452 170088 199504
rect 171048 199724 171100 199776
rect 171600 199724 171652 199776
rect 171324 199656 171376 199708
rect 171416 199656 171468 199708
rect 171876 199656 171928 199708
rect 171968 199656 172020 199708
rect 171232 199588 171284 199640
rect 171692 199588 171744 199640
rect 171784 199520 171836 199572
rect 172612 199656 172664 199708
rect 172704 199656 172756 199708
rect 172152 199588 172204 199640
rect 172244 199588 172296 199640
rect 173302 199860 173354 199912
rect 173578 199860 173630 199912
rect 173670 199860 173722 199912
rect 173854 199860 173906 199912
rect 173946 199860 173998 199912
rect 174406 199860 174458 199912
rect 174590 199860 174642 199912
rect 174774 199860 174826 199912
rect 175142 199860 175194 199912
rect 175234 199860 175286 199912
rect 173072 199724 173124 199776
rect 173164 199724 173216 199776
rect 172888 199588 172940 199640
rect 172980 199520 173032 199572
rect 172888 199452 172940 199504
rect 173348 199588 173400 199640
rect 169760 199384 169812 199436
rect 171508 199384 171560 199436
rect 173164 199384 173216 199436
rect 173624 199724 173676 199776
rect 173900 199656 173952 199708
rect 174268 199588 174320 199640
rect 175188 199724 175240 199776
rect 174912 199588 174964 199640
rect 175280 199588 175332 199640
rect 174636 199452 174688 199504
rect 174544 199384 174596 199436
rect 175786 199860 175838 199912
rect 176062 199860 176114 199912
rect 176154 199860 176206 199912
rect 176246 199860 176298 199912
rect 176430 199860 176482 199912
rect 176706 199860 176758 199912
rect 176798 199860 176850 199912
rect 176982 199860 177034 199912
rect 177166 199860 177218 199912
rect 177350 199860 177402 199912
rect 177626 199860 177678 199912
rect 177764 199860 177816 199912
rect 175694 199792 175746 199844
rect 175740 199656 175792 199708
rect 176016 199656 176068 199708
rect 176292 199724 176344 199776
rect 176200 199656 176252 199708
rect 176384 199656 176436 199708
rect 176844 199724 176896 199776
rect 177856 199792 177908 199844
rect 187240 199724 187292 199776
rect 176936 199656 176988 199708
rect 179052 199588 179104 199640
rect 175648 199520 175700 199572
rect 201500 199452 201552 199504
rect 175556 199384 175608 199436
rect 178960 199384 179012 199436
rect 187148 199384 187200 199436
rect 174084 199316 174136 199368
rect 183192 199316 183244 199368
rect 195612 199248 195664 199300
rect 118424 199180 118476 199232
rect 148692 199180 148744 199232
rect 173808 199180 173860 199232
rect 208584 199180 208636 199232
rect 117228 199112 117280 199164
rect 114468 199044 114520 199096
rect 141332 199112 141384 199164
rect 143908 199112 143960 199164
rect 158628 199112 158680 199164
rect 180248 199112 180300 199164
rect 180800 199112 180852 199164
rect 187056 199112 187108 199164
rect 111616 198976 111668 199028
rect 148416 199044 148468 199096
rect 113088 198908 113140 198960
rect 144828 198976 144880 199028
rect 169944 198976 169996 199028
rect 174084 198976 174136 199028
rect 174728 198976 174780 199028
rect 202420 198976 202472 199028
rect 136364 198840 136416 198892
rect 136640 198840 136692 198892
rect 137836 198840 137888 198892
rect 138940 198840 138992 198892
rect 142436 198908 142488 198960
rect 150716 198908 150768 198960
rect 173808 198908 173860 198960
rect 142620 198840 142672 198892
rect 167184 198840 167236 198892
rect 208492 198840 208544 198892
rect 126244 198772 126296 198824
rect 145564 198772 145616 198824
rect 153200 198772 153252 198824
rect 208400 198772 208452 198824
rect 182824 198704 182876 198756
rect 188252 198704 188304 198756
rect 155132 198568 155184 198620
rect 174820 198568 174872 198620
rect 132316 198500 132368 198552
rect 150808 198500 150860 198552
rect 122748 198228 122800 198280
rect 149152 198228 149204 198280
rect 162860 198160 162912 198212
rect 163320 198160 163372 198212
rect 167920 198160 167972 198212
rect 169668 198160 169720 198212
rect 198004 198160 198056 198212
rect 167644 198092 167696 198144
rect 171048 198092 171100 198144
rect 199660 198092 199712 198144
rect 132040 198024 132092 198076
rect 132500 198024 132552 198076
rect 136088 198024 136140 198076
rect 136272 198024 136324 198076
rect 173440 198024 173492 198076
rect 198832 198024 198884 198076
rect 131948 197956 132000 198008
rect 132868 197956 132920 198008
rect 183192 197956 183244 198008
rect 203156 197956 203208 198008
rect 129648 197888 129700 197940
rect 150072 197888 150124 197940
rect 133972 197752 134024 197804
rect 134432 197752 134484 197804
rect 163228 197752 163280 197804
rect 163596 197752 163648 197804
rect 115664 197616 115716 197668
rect 142344 197616 142396 197668
rect 155316 197548 155368 197600
rect 173440 197548 173492 197600
rect 134524 197480 134576 197532
rect 134892 197480 134944 197532
rect 163044 197276 163096 197328
rect 197544 197276 197596 197328
rect 154488 197208 154540 197260
rect 187056 197208 187108 197260
rect 156696 197140 156748 197192
rect 190552 197140 190604 197192
rect 162216 197072 162268 197124
rect 196072 197072 196124 197124
rect 118240 197004 118292 197056
rect 145196 197004 145248 197056
rect 166264 197004 166316 197056
rect 194692 197004 194744 197056
rect 157984 196936 158036 196988
rect 191932 196936 191984 196988
rect 111432 196868 111484 196920
rect 142896 196868 142948 196920
rect 163688 196868 163740 196920
rect 197452 196868 197504 196920
rect 110144 196800 110196 196852
rect 144644 196800 144696 196852
rect 160284 196800 160336 196852
rect 194876 196800 194928 196852
rect 105912 196732 105964 196784
rect 131028 196732 131080 196784
rect 159456 196732 159508 196784
rect 193404 196732 193456 196784
rect 115480 196664 115532 196716
rect 149520 196664 149572 196716
rect 161940 196664 161992 196716
rect 196164 196664 196216 196716
rect 112628 196596 112680 196648
rect 147588 196596 147640 196648
rect 157708 196596 157760 196648
rect 192116 196596 192168 196648
rect 158904 196528 158956 196580
rect 193496 196528 193548 196580
rect 154764 196460 154816 196512
rect 189724 196460 189776 196512
rect 169944 196052 169996 196104
rect 183100 196052 183152 196104
rect 167000 195916 167052 195968
rect 182916 195916 182968 195968
rect 119896 195848 119948 195900
rect 150348 195848 150400 195900
rect 156236 195848 156288 195900
rect 190736 195848 190788 195900
rect 159640 195780 159692 195832
rect 180156 195780 180208 195832
rect 111248 195712 111300 195764
rect 120356 195712 120408 195764
rect 159272 195712 159324 195764
rect 194140 195712 194192 195764
rect 111156 195644 111208 195696
rect 143172 195644 143224 195696
rect 110236 195576 110288 195628
rect 142252 195576 142304 195628
rect 157340 195576 157392 195628
rect 180064 195644 180116 195696
rect 106004 195508 106056 195560
rect 138664 195508 138716 195560
rect 161572 195508 161624 195560
rect 194600 195508 194652 195560
rect 105728 195440 105780 195492
rect 139124 195440 139176 195492
rect 160100 195440 160152 195492
rect 193312 195440 193364 195492
rect 109776 195372 109828 195424
rect 142528 195372 142580 195424
rect 160376 195372 160428 195424
rect 190644 195372 190696 195424
rect 106832 195304 106884 195356
rect 137836 195304 137888 195356
rect 158352 195304 158404 195356
rect 191840 195304 191892 195356
rect 105544 195236 105596 195288
rect 139584 195236 139636 195288
rect 158076 195236 158128 195288
rect 192024 195236 192076 195288
rect 173440 194964 173492 195016
rect 189172 194964 189224 195016
rect 153476 194896 153528 194948
rect 188252 194896 188304 194948
rect 174820 194828 174872 194880
rect 189080 194828 189132 194880
rect 128268 194692 128320 194744
rect 138756 194692 138808 194744
rect 127900 194488 127952 194540
rect 153292 194488 153344 194540
rect 100668 194352 100720 194404
rect 104440 194352 104492 194404
rect 115848 194284 115900 194336
rect 148232 194284 148284 194336
rect 112812 194216 112864 194268
rect 145840 194216 145892 194268
rect 114100 194148 114152 194200
rect 146944 194148 146996 194200
rect 174176 194148 174228 194200
rect 200764 194148 200816 194200
rect 112720 194080 112772 194132
rect 145012 194080 145064 194132
rect 114008 194012 114060 194064
rect 146392 194012 146444 194064
rect 174360 194012 174412 194064
rect 174728 194012 174780 194064
rect 177120 194012 177172 194064
rect 207020 194012 207072 194064
rect 102048 193944 102100 193996
rect 135260 193944 135312 193996
rect 169944 193944 169996 193996
rect 202880 193944 202932 193996
rect 118516 193876 118568 193928
rect 151544 193876 151596 193928
rect 167828 193876 167880 193928
rect 202512 193876 202564 193928
rect 106096 193808 106148 193860
rect 140228 193808 140280 193860
rect 166724 193808 166776 193860
rect 200120 193808 200172 193860
rect 108948 193672 109000 193724
rect 128268 193672 128320 193724
rect 131948 193672 132000 193724
rect 154672 193672 154724 193724
rect 130476 193604 130528 193656
rect 150624 193604 150676 193656
rect 162584 193264 162636 193316
rect 183468 193264 183520 193316
rect 164700 193196 164752 193248
rect 184112 193196 184164 193248
rect 156144 193128 156196 193180
rect 181536 193128 181588 193180
rect 188436 193128 188488 193180
rect 580172 193128 580224 193180
rect 171968 193060 172020 193112
rect 205640 193060 205692 193112
rect 164976 192992 165028 193044
rect 194784 192992 194836 193044
rect 110972 192924 111024 192976
rect 140688 192924 140740 192976
rect 173992 192924 174044 192976
rect 204352 192924 204404 192976
rect 108672 192856 108724 192908
rect 138664 192856 138716 192908
rect 176844 192856 176896 192908
rect 207112 192856 207164 192908
rect 168748 192788 168800 192840
rect 180340 192788 180392 192840
rect 183100 192788 183152 192840
rect 203064 192788 203116 192840
rect 167460 192720 167512 192772
rect 201776 192720 201828 192772
rect 103336 192652 103388 192704
rect 135812 192652 135864 192704
rect 169208 192652 169260 192704
rect 202972 192652 203024 192704
rect 104072 192584 104124 192636
rect 137652 192584 137704 192636
rect 103060 192516 103112 192568
rect 138020 192516 138072 192568
rect 164148 192516 164200 192568
rect 197360 192516 197412 192568
rect 103152 192448 103204 192500
rect 137468 192448 137520 192500
rect 153384 192448 153436 192500
rect 162216 192448 162268 192500
rect 174084 192448 174136 192500
rect 174912 192448 174964 192500
rect 183468 192448 183520 192500
rect 195980 192448 196032 192500
rect 116860 192380 116912 192432
rect 144552 192380 144604 192432
rect 173992 192380 174044 192432
rect 175004 192380 175056 192432
rect 184112 192380 184164 192432
rect 199108 192380 199160 192432
rect 110328 192312 110380 192364
rect 138020 192312 138072 192364
rect 125048 192244 125100 192296
rect 141700 192244 141752 192296
rect 166080 192244 166132 192296
rect 200212 192312 200264 192364
rect 168288 192176 168340 192228
rect 185584 192244 185636 192296
rect 166448 192040 166500 192092
rect 183008 192040 183060 192092
rect 161388 191632 161440 191684
rect 183100 191632 183152 191684
rect 122104 191360 122156 191412
rect 139860 191360 139912 191412
rect 111340 191292 111392 191344
rect 143080 191292 143132 191344
rect 101956 191224 102008 191276
rect 134340 191224 134392 191276
rect 109868 191156 109920 191208
rect 141332 191224 141384 191276
rect 109684 191088 109736 191140
rect 144184 191088 144236 191140
rect 131764 190952 131816 191004
rect 138940 190952 138992 191004
rect 123576 190884 123628 190936
rect 145288 190884 145340 190936
rect 127716 190680 127768 190732
rect 144000 190680 144052 190732
rect 168104 190680 168156 190732
rect 178868 190680 178920 190732
rect 110052 190408 110104 190460
rect 141424 190408 141476 190460
rect 110880 190340 110932 190392
rect 141884 190340 141936 190392
rect 107568 190272 107620 190324
rect 139952 190272 140004 190324
rect 106188 190204 106240 190256
rect 138296 190204 138348 190256
rect 100576 190136 100628 190188
rect 133788 190136 133840 190188
rect 101864 190068 101916 190120
rect 134800 190068 134852 190120
rect 111524 190000 111576 190052
rect 139400 190000 139452 190052
rect 101588 189932 101640 189984
rect 104808 189932 104860 189984
rect 101772 189864 101824 189916
rect 133972 189864 134024 189916
rect 101680 189796 101732 189848
rect 133604 189796 133656 189848
rect 104808 189728 104860 189780
rect 138848 189728 138900 189780
rect 107384 189660 107436 189712
rect 138572 189660 138624 189712
rect 108856 189592 108908 189644
rect 138940 189592 138992 189644
rect 112536 189524 112588 189576
rect 120172 189524 120224 189576
rect 165620 189048 165672 189100
rect 178776 189048 178828 189100
rect 3424 188980 3476 189032
rect 120540 188980 120592 189032
rect 131856 188912 131908 188964
rect 140780 188912 140832 188964
rect 126336 188844 126388 188896
rect 146024 188844 146076 188896
rect 127624 187960 127676 188012
rect 143724 187960 143776 188012
rect 130384 187416 130436 187468
rect 142804 187416 142856 187468
rect 163964 187280 164016 187332
rect 181444 187280 181496 187332
rect 102784 186940 102836 186992
rect 135536 186940 135588 186992
rect 163412 186940 163464 186992
rect 178684 186940 178736 186992
rect 124128 186872 124180 186924
rect 148324 186872 148376 186924
rect 171324 186668 171376 186720
rect 195244 186668 195296 186720
rect 160008 186600 160060 186652
rect 171232 186600 171284 186652
rect 171600 186600 171652 186652
rect 199016 186600 199068 186652
rect 172888 186464 172940 186516
rect 199200 186464 199252 186516
rect 154856 186396 154908 186448
rect 155500 186396 155552 186448
rect 174268 186396 174320 186448
rect 198740 186396 198792 186448
rect 172796 186328 172848 186380
rect 205732 186328 205784 186380
rect 136548 186260 136600 186312
rect 137192 186260 137244 186312
rect 158904 186260 158956 186312
rect 159548 186260 159600 186312
rect 161572 186260 161624 186312
rect 162032 186260 162084 186312
rect 169852 186260 169904 186312
rect 170864 186260 170916 186312
rect 171048 186260 171100 186312
rect 171508 186260 171560 186312
rect 176844 186260 176896 186312
rect 177212 186260 177264 186312
rect 107292 186192 107344 186244
rect 136456 186192 136508 186244
rect 148968 186192 149020 186244
rect 157800 186192 157852 186244
rect 176752 186192 176804 186244
rect 177488 186192 177540 186244
rect 148324 186124 148376 186176
rect 148784 186124 148836 186176
rect 176660 186124 176712 186176
rect 177764 186124 177816 186176
rect 154488 185784 154540 185836
rect 158812 185784 158864 185836
rect 103428 185716 103480 185768
rect 134248 185716 134300 185768
rect 105820 185648 105872 185700
rect 137284 185648 137336 185700
rect 153936 185648 153988 185700
rect 154396 185648 154448 185700
rect 155500 185648 155552 185700
rect 155776 185648 155828 185700
rect 158812 185648 158864 185700
rect 159824 185648 159876 185700
rect 164148 185648 164200 185700
rect 167276 185648 167328 185700
rect 174636 185648 174688 185700
rect 201684 185648 201736 185700
rect 104624 185580 104676 185632
rect 134524 185580 134576 185632
rect 141148 185580 141200 185632
rect 141516 185580 141568 185632
rect 149612 185580 149664 185632
rect 150164 185580 150216 185632
rect 151912 185580 151964 185632
rect 152464 185580 152516 185632
rect 153384 185580 153436 185632
rect 154120 185580 154172 185632
rect 154764 185580 154816 185632
rect 155684 185580 155736 185632
rect 156144 185580 156196 185632
rect 157064 185580 157116 185632
rect 157524 185580 157576 185632
rect 158444 185580 158496 185632
rect 160100 185580 160152 185632
rect 160928 185580 160980 185632
rect 161388 185580 161440 185632
rect 168380 185580 168432 185632
rect 169760 185580 169812 185632
rect 170312 185580 170364 185632
rect 172612 185580 172664 185632
rect 173256 185580 173308 185632
rect 175280 185580 175332 185632
rect 175832 185580 175884 185632
rect 104348 185512 104400 185564
rect 135168 185512 135220 185564
rect 142436 185512 142488 185564
rect 142712 185512 142764 185564
rect 156788 185512 156840 185564
rect 157248 185512 157300 185564
rect 167276 185512 167328 185564
rect 167644 185512 167696 185564
rect 121368 185308 121420 185360
rect 142160 185308 142212 185360
rect 108580 185172 108632 185224
rect 132500 185172 132552 185224
rect 127808 185104 127860 185156
rect 144276 185104 144328 185156
rect 108396 184968 108448 185020
rect 137744 184968 137796 185020
rect 160284 184968 160336 185020
rect 160652 184968 160704 185020
rect 150624 184560 150676 184612
rect 150992 184560 151044 184612
rect 107016 184356 107068 184408
rect 136088 184356 136140 184408
rect 126888 184288 126940 184340
rect 144920 184288 144972 184340
rect 150808 184288 150860 184340
rect 151268 184288 151320 184340
rect 102876 184152 102928 184204
rect 134064 184152 134116 184204
rect 146760 184152 146812 184204
rect 148048 184152 148100 184204
rect 172428 184016 172480 184068
rect 196808 184016 196860 184068
rect 121276 183744 121328 183796
rect 139124 183744 139176 183796
rect 164424 183268 164476 183320
rect 165344 183268 165396 183320
rect 175464 183064 175516 183116
rect 176200 183064 176252 183116
rect 150348 182996 150400 183048
rect 156328 182996 156380 183048
rect 164240 182860 164292 182912
rect 164608 182860 164660 182912
rect 164240 182724 164292 182776
rect 165068 182724 165120 182776
rect 147588 182656 147640 182708
rect 155224 182656 155276 182708
rect 104532 182520 104584 182572
rect 133328 182520 133380 182572
rect 108488 182112 108540 182164
rect 136824 182112 136876 182164
rect 149520 181976 149572 182028
rect 149980 181976 150032 182028
rect 172520 181976 172572 182028
rect 173624 181976 173676 182028
rect 104164 181568 104216 181620
rect 132592 181568 132644 181620
rect 132592 181432 132644 181484
rect 133052 181432 133104 181484
rect 160192 181432 160244 181484
rect 161296 181432 161348 181484
rect 150532 181160 150584 181212
rect 151636 181160 151688 181212
rect 146852 180480 146904 180532
rect 147404 180480 147456 180532
rect 129004 180344 129056 180396
rect 140872 180344 140924 180396
rect 152004 179936 152056 179988
rect 152648 179936 152700 179988
rect 161664 179936 161716 179988
rect 162308 179936 162360 179988
rect 157432 179800 157484 179852
rect 157892 179800 157944 179852
rect 161296 179120 161348 179172
rect 162124 179120 162176 179172
rect 163136 179120 163188 179172
rect 163780 179120 163832 179172
rect 135628 178984 135680 179036
rect 136180 178984 136232 179036
rect 145564 178984 145616 179036
rect 149060 178984 149112 179036
rect 149704 178712 149756 178764
rect 153568 178712 153620 178764
rect 108212 178440 108264 178492
rect 137928 178440 137980 178492
rect 142436 178440 142488 178492
rect 143264 178440 143316 178492
rect 171232 178236 171284 178288
rect 172336 178236 172388 178288
rect 175648 178032 175700 178084
rect 176384 178032 176436 178084
rect 188436 178032 188488 178084
rect 580172 178032 580224 178084
rect 146944 177148 146996 177200
rect 147772 177148 147824 177200
rect 102968 176944 103020 176996
rect 134616 176944 134668 176996
rect 167092 176944 167144 176996
rect 168196 176944 168248 176996
rect 104716 176400 104768 176452
rect 132960 176400 133012 176452
rect 145196 175856 145248 175908
rect 146300 175856 146352 175908
rect 164332 175720 164384 175772
rect 164792 175720 164844 175772
rect 158996 175176 159048 175228
rect 159364 175176 159416 175228
rect 171324 175176 171376 175228
rect 171784 175176 171836 175228
rect 107108 174224 107160 174276
rect 136272 174224 136324 174276
rect 132684 174088 132736 174140
rect 133512 174088 133564 174140
rect 137008 173544 137060 173596
rect 137376 173544 137428 173596
rect 117872 166268 117924 166320
rect 580172 166268 580224 166320
rect 165804 155660 165856 155712
rect 200396 155660 200448 155712
rect 167276 155592 167328 155644
rect 201868 155592 201920 155644
rect 167368 155524 167420 155576
rect 201960 155524 202012 155576
rect 165896 155456 165948 155508
rect 200580 155456 200632 155508
rect 168656 155388 168708 155440
rect 203340 155388 203392 155440
rect 168564 155320 168616 155372
rect 203524 155320 203576 155372
rect 168472 155252 168524 155304
rect 203432 155252 203484 155304
rect 167184 155184 167236 155236
rect 202144 155184 202196 155236
rect 160376 153144 160428 153196
rect 185676 153144 185728 153196
rect 159088 153076 159140 153128
rect 184388 153076 184440 153128
rect 160284 153008 160336 153060
rect 185768 153008 185820 153060
rect 158996 152940 159048 152992
rect 184480 152940 184532 152992
rect 158904 152872 158956 152924
rect 185860 152872 185912 152924
rect 163228 152804 163280 152856
rect 198188 152804 198240 152856
rect 164516 152736 164568 152788
rect 199752 152736 199804 152788
rect 164608 152668 164660 152720
rect 199384 152668 199436 152720
rect 149336 152600 149388 152652
rect 204720 152600 204772 152652
rect 146484 152532 146536 152584
rect 204812 152532 204864 152584
rect 147864 152464 147916 152516
rect 206192 152464 206244 152516
rect 160468 152396 160520 152448
rect 184572 152396 184624 152448
rect 161756 152328 161808 152380
rect 184664 152328 184716 152380
rect 161664 152260 161716 152312
rect 184204 152260 184256 152312
rect 161388 151036 161440 151088
rect 203248 151036 203300 151088
rect 179052 150356 179104 150408
rect 205824 150356 205876 150408
rect 176844 150288 176896 150340
rect 204904 150288 204956 150340
rect 174084 150220 174136 150272
rect 202328 150220 202380 150272
rect 175648 150152 175700 150204
rect 204444 150152 204496 150204
rect 176936 150084 176988 150136
rect 206284 150084 206336 150136
rect 175556 150016 175608 150068
rect 205916 150016 205968 150068
rect 175464 149948 175516 150000
rect 206100 149948 206152 150000
rect 175372 149880 175424 149932
rect 206008 149880 206060 149932
rect 172888 149812 172940 149864
rect 203708 149812 203760 149864
rect 175280 149744 175332 149796
rect 206376 149744 206428 149796
rect 148968 149676 149020 149728
rect 184756 149676 184808 149728
rect 173072 149608 173124 149660
rect 186964 149608 187016 149660
rect 182088 149540 182140 149592
rect 192668 149540 192720 149592
rect 3424 149064 3476 149116
rect 180892 149064 180944 149116
rect 182088 149064 182140 149116
rect 122380 148996 122432 149048
rect 152188 148996 152240 149048
rect 162952 148996 163004 149048
rect 185308 148996 185360 149048
rect 112168 148928 112220 148980
rect 142988 148928 143040 148980
rect 161572 148928 161624 148980
rect 186320 148928 186372 148980
rect 108120 148860 108172 148912
rect 139860 148860 139912 148912
rect 164424 148860 164476 148912
rect 197912 148860 197964 148912
rect 100208 148792 100260 148844
rect 132868 148792 132920 148844
rect 163044 148792 163096 148844
rect 197820 148792 197872 148844
rect 100392 148724 100444 148776
rect 132684 148724 132736 148776
rect 161480 148724 161532 148776
rect 196900 148724 196952 148776
rect 117688 148656 117740 148708
rect 150716 148656 150768 148708
rect 167092 148656 167144 148708
rect 202052 148656 202104 148708
rect 102692 148588 102744 148640
rect 135628 148588 135680 148640
rect 166816 148588 166868 148640
rect 200672 148588 200724 148640
rect 103980 148520 104032 148572
rect 137192 148520 137244 148572
rect 164332 148520 164384 148572
rect 199476 148520 199528 148572
rect 100300 148452 100352 148504
rect 134248 148452 134300 148504
rect 167920 148452 167972 148504
rect 202236 148452 202288 148504
rect 116308 148384 116360 148436
rect 150808 148384 150860 148436
rect 169208 148384 169260 148436
rect 203616 148384 203668 148436
rect 100116 148316 100168 148368
rect 134340 148316 134392 148368
rect 164240 148316 164292 148368
rect 199568 148316 199620 148368
rect 123944 148248 123996 148300
rect 152096 148248 152148 148300
rect 185032 148248 185084 148300
rect 199292 148248 199344 148300
rect 113548 148180 113600 148232
rect 142436 148180 142488 148232
rect 180156 148180 180208 148232
rect 192852 148180 192904 148232
rect 122196 148112 122248 148164
rect 149704 148112 149756 148164
rect 179328 147568 179380 147620
rect 196716 147568 196768 147620
rect 171508 147500 171560 147552
rect 194968 147500 195020 147552
rect 171232 147432 171284 147484
rect 195336 147432 195388 147484
rect 171324 147364 171376 147416
rect 196992 147364 197044 147416
rect 169944 147296 169996 147348
rect 197084 147296 197136 147348
rect 171416 147228 171468 147280
rect 198096 147228 198148 147280
rect 172796 147160 172848 147212
rect 200948 147160 201000 147212
rect 172704 147092 172756 147144
rect 200856 147092 200908 147144
rect 164148 147024 164200 147076
rect 193956 147024 194008 147076
rect 111064 146956 111116 147008
rect 130200 146956 130252 147008
rect 172612 146956 172664 147008
rect 204536 146956 204588 147008
rect 113456 146888 113508 146940
rect 142712 146888 142764 146940
rect 170036 146888 170088 146940
rect 204628 146888 204680 146940
rect 178592 146820 178644 146872
rect 196440 146820 196492 146872
rect 130200 146276 130252 146328
rect 580356 146276 580408 146328
rect 3516 146208 3568 146260
rect 179052 146208 179104 146260
rect 179788 146208 179840 146260
rect 192300 146208 192352 146260
rect 113824 146140 113876 146192
rect 130752 146140 130804 146192
rect 183468 146140 183520 146192
rect 196532 146140 196584 146192
rect 114284 146072 114336 146124
rect 132408 146072 132460 146124
rect 178040 146072 178092 146124
rect 192576 146072 192628 146124
rect 112352 146004 112404 146056
rect 131028 146004 131080 146056
rect 131764 146004 131816 146056
rect 132224 146004 132276 146056
rect 179604 146004 179656 146056
rect 196624 146004 196676 146056
rect 117964 145936 118016 145988
rect 146300 145936 146352 145988
rect 162216 145936 162268 145988
rect 188528 145936 188580 145988
rect 119068 145868 119120 145920
rect 150624 145868 150676 145920
rect 160192 145868 160244 145920
rect 195520 145868 195572 145920
rect 117964 145800 118016 145852
rect 149244 145800 149296 145852
rect 158536 145800 158588 145852
rect 192760 145800 192812 145852
rect 114836 145732 114888 145784
rect 149520 145732 149572 145784
rect 157432 145732 157484 145784
rect 192300 145732 192352 145784
rect 114928 145664 114980 145716
rect 149612 145664 149664 145716
rect 154488 145664 154540 145716
rect 194324 145664 194376 145716
rect 114744 145596 114796 145648
rect 145564 145596 145616 145648
rect 147588 145596 147640 145648
rect 190000 145596 190052 145648
rect 112352 145528 112404 145580
rect 142528 145528 142580 145580
rect 145196 145528 145248 145580
rect 206468 145528 206520 145580
rect 115204 145460 115256 145512
rect 130568 145460 130620 145512
rect 178132 145460 178184 145512
rect 189632 145460 189684 145512
rect 115112 145392 115164 145444
rect 129556 145392 129608 145444
rect 179512 145392 179564 145444
rect 190920 145392 190972 145444
rect 179420 145324 179472 145376
rect 189908 145324 189960 145376
rect 116124 144848 116176 144900
rect 130476 144848 130528 144900
rect 180064 144848 180116 144900
rect 191380 144848 191432 144900
rect 114284 144780 114336 144832
rect 130384 144780 130436 144832
rect 174360 144780 174412 144832
rect 189816 144780 189868 144832
rect 113640 144712 113692 144764
rect 129004 144712 129056 144764
rect 171048 144712 171100 144764
rect 192484 144712 192536 144764
rect 114192 144644 114244 144696
rect 137284 144644 137336 144696
rect 172428 144644 172480 144696
rect 193864 144644 193916 144696
rect 116584 144576 116636 144628
rect 142252 144576 142304 144628
rect 162492 144576 162544 144628
rect 191012 144576 191064 144628
rect 120540 144508 120592 144560
rect 150532 144508 150584 144560
rect 158352 144508 158404 144560
rect 190828 144508 190880 144560
rect 119436 144440 119488 144492
rect 149428 144440 149480 144492
rect 157800 144440 157852 144492
rect 191104 144440 191156 144492
rect 119252 144372 119304 144424
rect 154028 144372 154080 144424
rect 156696 144372 156748 144424
rect 190460 144372 190512 144424
rect 120632 144304 120684 144356
rect 151268 144304 151320 144356
rect 153108 144304 153160 144356
rect 186596 144304 186648 144356
rect 113732 144236 113784 144288
rect 148048 144236 148100 144288
rect 159916 144236 159968 144288
rect 193772 144236 193824 144288
rect 112444 144168 112496 144220
rect 131488 144168 131540 144220
rect 188436 144168 188488 144220
rect 129556 143488 129608 143540
rect 580264 143488 580316 143540
rect 177672 143420 177724 143472
rect 179420 143420 179472 143472
rect 181536 143420 181588 143472
rect 189632 143420 189684 143472
rect 117872 143352 117924 143404
rect 130108 143352 130160 143404
rect 116768 143284 116820 143336
rect 132040 143352 132092 143404
rect 176568 143352 176620 143404
rect 178592 143352 178644 143404
rect 185584 143352 185636 143404
rect 188344 143352 188396 143404
rect 131856 143284 131908 143336
rect 138020 143284 138072 143336
rect 176016 143284 176068 143336
rect 179788 143284 179840 143336
rect 184296 143284 184348 143336
rect 195060 143284 195112 143336
rect 118056 143216 118108 143268
rect 133420 143216 133472 143268
rect 184664 143216 184716 143268
rect 196808 143216 196860 143268
rect 119804 143148 119856 143200
rect 138388 143148 138440 143200
rect 175188 143148 175240 143200
rect 189540 143148 189592 143200
rect 117044 143080 117096 143132
rect 135260 143080 135312 143132
rect 168840 143080 168892 143132
rect 189264 143080 189316 143132
rect 121092 143012 121144 143064
rect 140044 143012 140096 143064
rect 166908 143012 166960 143064
rect 186688 143012 186740 143064
rect 118148 142944 118200 142996
rect 136732 142944 136784 142996
rect 165528 142944 165580 142996
rect 187976 142944 188028 142996
rect 119620 142876 119672 142928
rect 141700 142876 141752 142928
rect 160560 142876 160612 142928
rect 186780 142876 186832 142928
rect 121000 142808 121052 142860
rect 143540 142808 143592 142860
rect 155040 142808 155092 142860
rect 157708 142808 157760 142860
rect 158628 142808 158680 142860
rect 188068 142808 188120 142860
rect 132408 142740 132460 142792
rect 136180 142740 136232 142792
rect 177120 142740 177172 142792
rect 179512 142740 179564 142792
rect 119712 142672 119764 142724
rect 127900 142672 127952 142724
rect 131028 142672 131080 142724
rect 134524 142672 134576 142724
rect 179052 142672 179104 142724
rect 179788 142672 179840 142724
rect 177948 142604 178000 142656
rect 179328 142604 179380 142656
rect 130568 142468 130620 142520
rect 132500 142468 132552 142520
rect 3424 142264 3476 142316
rect 185584 142264 185636 142316
rect 125600 142196 125652 142248
rect 126520 142196 126572 142248
rect 188160 142196 188212 142248
rect 116676 142128 116728 142180
rect 124220 142128 124272 142180
rect 118332 142060 118384 142112
rect 140780 142128 140832 142180
rect 155868 142128 155920 142180
rect 157340 142128 157392 142180
rect 159456 142128 159508 142180
rect 162492 142128 162544 142180
rect 184388 142060 184440 142112
rect 193864 142060 193916 142112
rect 121184 141992 121236 142044
rect 127072 141992 127124 142044
rect 182272 141992 182324 142044
rect 192392 141992 192444 142044
rect 120816 141924 120868 141976
rect 123760 141924 123812 141976
rect 183100 141924 183152 141976
rect 194232 141924 194284 141976
rect 119528 141856 119580 141908
rect 125140 141856 125192 141908
rect 184572 141856 184624 141908
rect 195152 141856 195204 141908
rect 115296 141788 115348 141840
rect 124588 141788 124640 141840
rect 180156 141788 180208 141840
rect 192208 141788 192260 141840
rect 116952 141720 117004 141772
rect 129004 141720 129056 141772
rect 184848 141720 184900 141772
rect 196348 141720 196400 141772
rect 113916 141652 113968 141704
rect 126980 141652 127032 141704
rect 172152 141652 172204 141704
rect 187884 141652 187936 141704
rect 117136 141584 117188 141636
rect 133972 141584 134024 141636
rect 170496 141584 170548 141636
rect 189448 141584 189500 141636
rect 112260 141516 112312 141568
rect 131672 141516 131724 141568
rect 174728 141516 174780 141568
rect 197728 141516 197780 141568
rect 115388 141448 115440 141500
rect 135628 141448 135680 141500
rect 169392 141448 169444 141500
rect 193680 141448 193732 141500
rect 121184 141380 121236 141432
rect 151912 141380 151964 141432
rect 160744 141380 160796 141432
rect 189356 141380 189408 141432
rect 118700 141108 118752 141160
rect 180156 141108 180208 141160
rect 180616 141108 180668 141160
rect 111064 141040 111116 141092
rect 184848 141040 184900 141092
rect 8944 140972 8996 141024
rect 182824 140972 182876 141024
rect 127072 140904 127124 140956
rect 549904 140904 549956 140956
rect 129004 140836 129056 140888
rect 580540 140836 580592 140888
rect 126980 140768 127032 140820
rect 127624 140768 127676 140820
rect 580448 140768 580500 140820
rect 119804 140700 119856 140752
rect 127808 140700 127860 140752
rect 169760 140700 169812 140752
rect 193680 140700 193732 140752
rect 119528 140632 119580 140684
rect 127532 140632 127584 140684
rect 178040 140632 178092 140684
rect 178684 140632 178736 140684
rect 120816 140564 120868 140616
rect 127716 140564 127768 140616
rect 172520 140564 172572 140616
rect 193220 140632 193272 140684
rect 185676 140564 185728 140616
rect 116676 140428 116728 140480
rect 126244 140496 126296 140548
rect 181444 140496 181496 140548
rect 116584 140360 116636 140412
rect 126336 140360 126388 140412
rect 178776 140360 178828 140412
rect 189356 140360 189408 140412
rect 195428 140428 195480 140480
rect 120908 140292 120960 140344
rect 148140 140292 148192 140344
rect 185860 140292 185912 140344
rect 189816 140292 189868 140344
rect 192208 140292 192260 140344
rect 119344 140224 119396 140276
rect 146944 140224 146996 140276
rect 178868 140224 178920 140276
rect 191288 140224 191340 140276
rect 117780 140156 117832 140208
rect 146852 140156 146904 140208
rect 183100 140156 183152 140208
rect 189908 140156 189960 140208
rect 116400 140088 116452 140140
rect 146760 140088 146812 140140
rect 179236 140088 179288 140140
rect 192668 140088 192720 140140
rect 116492 140020 116544 140072
rect 148232 140020 148284 140072
rect 160100 140020 160152 140072
rect 192576 140020 192628 140072
rect 119620 139952 119672 140004
rect 123576 139952 123628 140004
rect 184204 139952 184256 140004
rect 196716 139952 196768 140004
rect 168288 139816 168340 139868
rect 178592 139816 178644 139868
rect 173256 139748 173308 139800
rect 196256 139748 196308 139800
rect 121000 139680 121052 139732
rect 125048 139680 125100 139732
rect 169760 139680 169812 139732
rect 193588 139680 193640 139732
rect 118332 139612 118384 139664
rect 123944 139612 123996 139664
rect 171600 139612 171652 139664
rect 197636 139612 197688 139664
rect 126152 139544 126204 139596
rect 179880 139544 179932 139596
rect 125048 139476 125100 139528
rect 180432 139476 180484 139528
rect 113916 139408 113968 139460
rect 122104 139408 122156 139460
rect 124036 139408 124088 139460
rect 182088 139408 182140 139460
rect 121920 139340 121972 139392
rect 123668 139340 123720 139392
rect 155132 139340 155184 139392
rect 155500 139340 155552 139392
rect 185768 139340 185820 139392
rect 186412 139340 186464 139392
rect 188160 138660 188212 138712
rect 580264 138660 580316 138712
rect 3516 137912 3568 137964
rect 118700 137912 118752 137964
rect 118056 136280 118108 136332
rect 120816 136280 120868 136332
rect 3148 111732 3200 111784
rect 31024 111732 31076 111784
rect 549904 86912 549956 86964
rect 580172 86912 580224 86964
rect 108396 80928 108448 80980
rect 123484 80928 123536 80980
rect 120908 80860 120960 80912
rect 108212 80792 108264 80844
rect 124036 80792 124088 80844
rect 116400 80724 116452 80776
rect 71780 80656 71832 80708
rect 108212 80656 108264 80708
rect 117688 80656 117740 80708
rect 123484 80656 123536 80708
rect 129832 80656 129884 80708
rect 115020 80180 115072 80232
rect 132040 80112 132092 80164
rect 129832 80044 129884 80096
rect 130844 80044 130896 80096
rect 106832 79840 106884 79892
rect 131948 79908 132000 79960
rect 132730 79908 132782 79960
rect 132822 79908 132874 79960
rect 133006 79908 133058 79960
rect 124036 79840 124088 79892
rect 114836 79772 114888 79824
rect 129924 79840 129976 79892
rect 132914 79840 132966 79892
rect 109684 79704 109736 79756
rect 123484 79704 123536 79756
rect 132316 79704 132368 79756
rect 117872 79636 117924 79688
rect 130752 79636 130804 79688
rect 132224 79636 132276 79688
rect 132776 79704 132828 79756
rect 133190 79908 133242 79960
rect 133282 79908 133334 79960
rect 133374 79908 133426 79960
rect 133466 79908 133518 79960
rect 133328 79704 133380 79756
rect 133650 79908 133702 79960
rect 133742 79908 133794 79960
rect 133834 79840 133886 79892
rect 133696 79772 133748 79824
rect 133788 79704 133840 79756
rect 133236 79636 133288 79688
rect 133512 79636 133564 79688
rect 133604 79636 133656 79688
rect 110880 79568 110932 79620
rect 121092 79568 121144 79620
rect 106740 79500 106792 79552
rect 123024 79568 123076 79620
rect 129096 79568 129148 79620
rect 134386 79908 134438 79960
rect 135398 79908 135450 79960
rect 135858 79908 135910 79960
rect 134294 79840 134346 79892
rect 134110 79772 134162 79824
rect 134570 79840 134622 79892
rect 134432 79772 134484 79824
rect 134340 79704 134392 79756
rect 134064 79568 134116 79620
rect 110972 79432 111024 79484
rect 126980 79500 127032 79552
rect 131672 79500 131724 79552
rect 132408 79500 132460 79552
rect 135122 79840 135174 79892
rect 135214 79840 135266 79892
rect 135306 79840 135358 79892
rect 135030 79772 135082 79824
rect 135168 79704 135220 79756
rect 135076 79568 135128 79620
rect 134800 79500 134852 79552
rect 134984 79500 135036 79552
rect 135674 79840 135726 79892
rect 135950 79840 136002 79892
rect 135812 79772 135864 79824
rect 135904 79704 135956 79756
rect 135628 79568 135680 79620
rect 135720 79568 135772 79620
rect 136778 79908 136830 79960
rect 136870 79908 136922 79960
rect 136318 79840 136370 79892
rect 137238 79908 137290 79960
rect 137422 79908 137474 79960
rect 137606 79908 137658 79960
rect 137054 79840 137106 79892
rect 137146 79772 137198 79824
rect 137008 79704 137060 79756
rect 136916 79636 136968 79688
rect 136272 79568 136324 79620
rect 136180 79500 136232 79552
rect 137376 79636 137428 79688
rect 137974 79908 138026 79960
rect 138342 79908 138394 79960
rect 138802 79908 138854 79960
rect 138894 79908 138946 79960
rect 139262 79908 139314 79960
rect 138434 79840 138486 79892
rect 138158 79772 138210 79824
rect 138020 79636 138072 79688
rect 137284 79568 137336 79620
rect 137836 79568 137888 79620
rect 138388 79636 138440 79688
rect 138480 79568 138532 79620
rect 139170 79840 139222 79892
rect 139354 79840 139406 79892
rect 138940 79772 138992 79824
rect 139032 79636 139084 79688
rect 139124 79568 139176 79620
rect 137560 79500 137612 79552
rect 138204 79500 138256 79552
rect 139216 79500 139268 79552
rect 140182 79908 140234 79960
rect 140734 79908 140786 79960
rect 140826 79908 140878 79960
rect 140918 79908 140970 79960
rect 141838 79908 141890 79960
rect 141930 79908 141982 79960
rect 142114 79908 142166 79960
rect 142298 79908 142350 79960
rect 142390 79908 142442 79960
rect 142758 79908 142810 79960
rect 140458 79840 140510 79892
rect 139814 79772 139866 79824
rect 139768 79636 139820 79688
rect 139676 79568 139728 79620
rect 140596 79568 140648 79620
rect 141194 79840 141246 79892
rect 142022 79840 142074 79892
rect 140872 79636 140924 79688
rect 140964 79636 141016 79688
rect 141470 79772 141522 79824
rect 141838 79772 141890 79824
rect 141930 79772 141982 79824
rect 142206 79840 142258 79892
rect 142114 79772 142166 79824
rect 142298 79772 142350 79824
rect 142160 79636 142212 79688
rect 142344 79636 142396 79688
rect 141148 79568 141200 79620
rect 141516 79568 141568 79620
rect 142666 79840 142718 79892
rect 142942 79840 142994 79892
rect 143126 79840 143178 79892
rect 142620 79636 142672 79688
rect 142988 79636 143040 79688
rect 142804 79568 142856 79620
rect 143264 79568 143316 79620
rect 139584 79500 139636 79552
rect 143494 79908 143546 79960
rect 143586 79908 143638 79960
rect 143770 79908 143822 79960
rect 144322 79908 144374 79960
rect 144598 79908 144650 79960
rect 144690 79908 144742 79960
rect 144782 79908 144834 79960
rect 144138 79840 144190 79892
rect 144092 79568 144144 79620
rect 144276 79568 144328 79620
rect 144736 79704 144788 79756
rect 144828 79636 144880 79688
rect 144644 79568 144696 79620
rect 143632 79500 143684 79552
rect 143724 79500 143776 79552
rect 109960 79364 110012 79416
rect 123484 79364 123536 79416
rect 143540 79432 143592 79484
rect 132316 79364 132368 79416
rect 143908 79364 143960 79416
rect 145702 79908 145754 79960
rect 146346 79908 146398 79960
rect 146438 79908 146490 79960
rect 146714 79908 146766 79960
rect 146806 79908 146858 79960
rect 145150 79840 145202 79892
rect 145426 79840 145478 79892
rect 145610 79840 145662 79892
rect 145104 79500 145156 79552
rect 145794 79840 145846 79892
rect 146162 79840 146214 79892
rect 146254 79840 146306 79892
rect 145978 79772 146030 79824
rect 145656 79636 145708 79688
rect 145748 79636 145800 79688
rect 146024 79636 146076 79688
rect 146116 79636 146168 79688
rect 146208 79568 146260 79620
rect 146484 79568 146536 79620
rect 145380 79500 145432 79552
rect 146668 79500 146720 79552
rect 147174 79908 147226 79960
rect 147266 79840 147318 79892
rect 147542 79840 147594 79892
rect 147128 79568 147180 79620
rect 147496 79568 147548 79620
rect 146944 79500 146996 79552
rect 147404 79500 147456 79552
rect 188160 81200 188212 81252
rect 186412 80860 186464 80912
rect 199568 80860 199620 80912
rect 188160 80792 188212 80844
rect 208584 80792 208636 80844
rect 234620 80792 234672 80844
rect 188252 80724 188304 80776
rect 270500 80724 270552 80776
rect 177856 80656 177908 80708
rect 183652 80656 183704 80708
rect 183836 80656 183888 80708
rect 189724 80656 189776 80708
rect 288440 80656 288492 80708
rect 177764 80588 177816 80640
rect 186412 80452 186464 80504
rect 194048 80384 194100 80436
rect 148370 79908 148422 79960
rect 148462 79908 148514 79960
rect 148554 79908 148606 79960
rect 150670 79908 150722 79960
rect 150762 79908 150814 79960
rect 151038 79908 151090 79960
rect 151314 79908 151366 79960
rect 151590 79908 151642 79960
rect 147910 79840 147962 79892
rect 148094 79840 148146 79892
rect 147956 79636 148008 79688
rect 148922 79840 148974 79892
rect 149382 79840 149434 79892
rect 149474 79840 149526 79892
rect 149566 79840 149618 79892
rect 149842 79840 149894 79892
rect 150118 79840 150170 79892
rect 150578 79840 150630 79892
rect 148416 79636 148468 79688
rect 148600 79568 148652 79620
rect 148784 79568 148836 79620
rect 148048 79500 148100 79552
rect 148140 79500 148192 79552
rect 149014 79772 149066 79824
rect 148968 79636 149020 79688
rect 145472 79432 145524 79484
rect 145840 79432 145892 79484
rect 149428 79636 149480 79688
rect 150716 79772 150768 79824
rect 151084 79772 151136 79824
rect 150624 79704 150676 79756
rect 150164 79636 150216 79688
rect 151176 79636 151228 79688
rect 152142 79908 152194 79960
rect 151958 79840 152010 79892
rect 152234 79840 152286 79892
rect 152004 79636 152056 79688
rect 151820 79568 151872 79620
rect 149612 79500 149664 79552
rect 149796 79500 149848 79552
rect 149428 79432 149480 79484
rect 150532 79500 150584 79552
rect 151544 79500 151596 79552
rect 152188 79704 152240 79756
rect 109776 79296 109828 79348
rect 132132 79296 132184 79348
rect 132224 79296 132276 79348
rect 139584 79296 139636 79348
rect 139952 79296 140004 79348
rect 140228 79296 140280 79348
rect 141240 79296 141292 79348
rect 141424 79296 141476 79348
rect 143540 79296 143592 79348
rect 144184 79296 144236 79348
rect 146208 79296 146260 79348
rect 150348 79364 150400 79416
rect 119344 79228 119396 79280
rect 147588 79228 147640 79280
rect 147864 79228 147916 79280
rect 149888 79228 149940 79280
rect 152096 79432 152148 79484
rect 152418 79908 152470 79960
rect 152694 79908 152746 79960
rect 152786 79908 152838 79960
rect 152878 79908 152930 79960
rect 153246 79908 153298 79960
rect 153430 79908 153482 79960
rect 152510 79772 152562 79824
rect 152464 79636 152516 79688
rect 153154 79840 153206 79892
rect 152924 79772 152976 79824
rect 153062 79772 153114 79824
rect 153200 79704 153252 79756
rect 152832 79636 152884 79688
rect 153016 79636 153068 79688
rect 152832 79500 152884 79552
rect 153798 79908 153850 79960
rect 154074 79908 154126 79960
rect 154166 79908 154218 79960
rect 154442 79908 154494 79960
rect 154718 79908 154770 79960
rect 154810 79908 154862 79960
rect 154902 79908 154954 79960
rect 154258 79840 154310 79892
rect 154534 79840 154586 79892
rect 154626 79840 154678 79892
rect 154396 79704 154448 79756
rect 154764 79772 154816 79824
rect 155086 79772 155138 79824
rect 154672 79704 154724 79756
rect 154856 79704 154908 79756
rect 153844 79636 153896 79688
rect 153936 79636 153988 79688
rect 154028 79636 154080 79688
rect 154212 79636 154264 79688
rect 154488 79636 154540 79688
rect 155040 79636 155092 79688
rect 155270 79908 155322 79960
rect 155454 79908 155506 79960
rect 155546 79908 155598 79960
rect 156190 79908 156242 79960
rect 156374 79908 156426 79960
rect 154948 79568 155000 79620
rect 155132 79568 155184 79620
rect 155454 79772 155506 79824
rect 155408 79568 155460 79620
rect 156006 79840 156058 79892
rect 156052 79568 156104 79620
rect 155960 79500 156012 79552
rect 156834 79772 156886 79824
rect 156420 79568 156472 79620
rect 156696 79500 156748 79552
rect 155684 79432 155736 79484
rect 157110 79908 157162 79960
rect 157386 79908 157438 79960
rect 157754 79908 157806 79960
rect 158030 79908 158082 79960
rect 158122 79908 158174 79960
rect 158398 79908 158450 79960
rect 158490 79908 158542 79960
rect 158766 79908 158818 79960
rect 159226 79908 159278 79960
rect 159318 79908 159370 79960
rect 159502 79908 159554 79960
rect 157202 79772 157254 79824
rect 157156 79636 157208 79688
rect 157662 79772 157714 79824
rect 157754 79772 157806 79824
rect 158076 79772 158128 79824
rect 158398 79772 158450 79824
rect 157064 79568 157116 79620
rect 157248 79568 157300 79620
rect 157432 79568 157484 79620
rect 158444 79568 158496 79620
rect 157800 79500 157852 79552
rect 158950 79840 159002 79892
rect 158904 79704 158956 79756
rect 159410 79840 159462 79892
rect 159180 79772 159232 79824
rect 159456 79704 159508 79756
rect 159364 79636 159416 79688
rect 159778 79908 159830 79960
rect 160238 79908 160290 79960
rect 160422 79908 160474 79960
rect 160606 79908 160658 79960
rect 159732 79772 159784 79824
rect 159962 79840 160014 79892
rect 159824 79704 159876 79756
rect 160284 79704 160336 79756
rect 160192 79636 160244 79688
rect 160882 79908 160934 79960
rect 160974 79908 161026 79960
rect 161066 79908 161118 79960
rect 161158 79908 161210 79960
rect 161434 79908 161486 79960
rect 161710 79908 161762 79960
rect 161802 79908 161854 79960
rect 162078 79908 162130 79960
rect 162262 79908 162314 79960
rect 162630 79908 162682 79960
rect 162722 79908 162774 79960
rect 163182 79908 163234 79960
rect 163366 79908 163418 79960
rect 163550 79908 163602 79960
rect 164102 79908 164154 79960
rect 160698 79840 160750 79892
rect 160606 79772 160658 79824
rect 159272 79568 159324 79620
rect 160560 79568 160612 79620
rect 160882 79772 160934 79824
rect 161158 79772 161210 79824
rect 161250 79772 161302 79824
rect 160836 79568 160888 79620
rect 159548 79500 159600 79552
rect 161296 79636 161348 79688
rect 161112 79568 161164 79620
rect 161664 79772 161716 79824
rect 161894 79840 161946 79892
rect 161756 79704 161808 79756
rect 162032 79636 162084 79688
rect 161848 79568 161900 79620
rect 162446 79772 162498 79824
rect 162676 79772 162728 79824
rect 162400 79568 162452 79620
rect 162584 79568 162636 79620
rect 161204 79500 161256 79552
rect 162308 79500 162360 79552
rect 162492 79500 162544 79552
rect 157984 79432 158036 79484
rect 163090 79840 163142 79892
rect 162998 79772 163050 79824
rect 162860 79636 162912 79688
rect 163044 79568 163096 79620
rect 163320 79772 163372 79824
rect 163826 79840 163878 79892
rect 163596 79772 163648 79824
rect 163780 79636 163832 79688
rect 163964 79568 164016 79620
rect 187148 80316 187200 80368
rect 177764 80248 177816 80300
rect 178316 80180 178368 80232
rect 165114 79908 165166 79960
rect 165206 79908 165258 79960
rect 164470 79840 164522 79892
rect 164562 79840 164614 79892
rect 164838 79840 164890 79892
rect 165022 79840 165074 79892
rect 164240 79636 164292 79688
rect 164332 79636 164384 79688
rect 164516 79636 164568 79688
rect 164608 79636 164660 79688
rect 164700 79636 164752 79688
rect 164884 79636 164936 79688
rect 165160 79636 165212 79688
rect 165068 79568 165120 79620
rect 165390 79840 165442 79892
rect 166310 79908 166362 79960
rect 166678 79908 166730 79960
rect 166770 79908 166822 79960
rect 166954 79908 167006 79960
rect 167138 79908 167190 79960
rect 167230 79908 167282 79960
rect 167322 79908 167374 79960
rect 167598 79908 167650 79960
rect 167690 79908 167742 79960
rect 167966 79908 168018 79960
rect 168058 79908 168110 79960
rect 168150 79908 168202 79960
rect 165804 79636 165856 79688
rect 165620 79568 165672 79620
rect 166126 79840 166178 79892
rect 166034 79772 166086 79824
rect 166218 79772 166270 79824
rect 166494 79772 166546 79824
rect 165896 79500 165948 79552
rect 166632 79636 166684 79688
rect 166816 79636 166868 79688
rect 166264 79568 166316 79620
rect 166448 79568 166500 79620
rect 166816 79500 166868 79552
rect 153844 79364 153896 79416
rect 154396 79364 154448 79416
rect 155408 79364 155460 79416
rect 155868 79364 155920 79416
rect 156880 79364 156932 79416
rect 157340 79364 157392 79416
rect 157524 79364 157576 79416
rect 153660 79296 153712 79348
rect 160284 79296 160336 79348
rect 166448 79432 166500 79484
rect 167046 79840 167098 79892
rect 167184 79704 167236 79756
rect 167506 79840 167558 79892
rect 167368 79636 167420 79688
rect 167460 79636 167512 79688
rect 167552 79636 167604 79688
rect 167276 79568 167328 79620
rect 168104 79772 168156 79824
rect 168518 79908 168570 79960
rect 168472 79772 168524 79824
rect 168564 79568 168616 79620
rect 168104 79500 168156 79552
rect 167644 79432 167696 79484
rect 167828 79432 167880 79484
rect 168794 79908 168846 79960
rect 168978 79908 169030 79960
rect 169070 79908 169122 79960
rect 169162 79908 169214 79960
rect 169622 79908 169674 79960
rect 168932 79636 168984 79688
rect 169254 79840 169306 79892
rect 169346 79840 169398 79892
rect 169438 79772 169490 79824
rect 169392 79636 169444 79688
rect 169898 79840 169950 79892
rect 169668 79704 169720 79756
rect 170266 79908 170318 79960
rect 170818 79908 170870 79960
rect 171002 79908 171054 79960
rect 170358 79840 170410 79892
rect 170542 79840 170594 79892
rect 170404 79704 170456 79756
rect 170312 79636 170364 79688
rect 170772 79772 170824 79824
rect 170910 79772 170962 79824
rect 169208 79568 169260 79620
rect 169484 79568 169536 79620
rect 169852 79568 169904 79620
rect 170036 79568 170088 79620
rect 170496 79568 170548 79620
rect 171278 79908 171330 79960
rect 171646 79908 171698 79960
rect 171738 79908 171790 79960
rect 171830 79908 171882 79960
rect 171922 79908 171974 79960
rect 171462 79840 171514 79892
rect 171416 79704 171468 79756
rect 171508 79636 171560 79688
rect 171140 79568 171192 79620
rect 171692 79772 171744 79824
rect 171784 79704 171836 79756
rect 172106 79908 172158 79960
rect 171784 79568 171836 79620
rect 169024 79500 169076 79552
rect 170772 79500 170824 79552
rect 169300 79432 169352 79484
rect 171968 79704 172020 79756
rect 172060 79704 172112 79756
rect 178132 80112 178184 80164
rect 252560 80112 252612 80164
rect 172382 79908 172434 79960
rect 172842 79908 172894 79960
rect 173026 79908 173078 79960
rect 173118 79908 173170 79960
rect 173302 79908 173354 79960
rect 173578 79908 173630 79960
rect 173670 79908 173722 79960
rect 173762 79908 173814 79960
rect 173946 79908 173998 79960
rect 172474 79840 172526 79892
rect 172566 79840 172618 79892
rect 172336 79704 172388 79756
rect 172428 79636 172480 79688
rect 172152 79568 172204 79620
rect 172934 79772 172986 79824
rect 172888 79636 172940 79688
rect 172796 79568 172848 79620
rect 173716 79772 173768 79824
rect 173164 79636 173216 79688
rect 173256 79568 173308 79620
rect 174038 79840 174090 79892
rect 173992 79704 174044 79756
rect 173900 79636 173952 79688
rect 173348 79500 173400 79552
rect 172888 79432 172940 79484
rect 124128 79160 124180 79212
rect 155868 79228 155920 79280
rect 162124 79228 162176 79280
rect 171600 79364 171652 79416
rect 165160 79296 165212 79348
rect 165528 79296 165580 79348
rect 173900 79296 173952 79348
rect 117964 79092 118016 79144
rect 149060 79092 149112 79144
rect 149704 79092 149756 79144
rect 119068 79024 119120 79076
rect 151084 79092 151136 79144
rect 155776 79092 155828 79144
rect 158812 79092 158864 79144
rect 163504 79092 163556 79144
rect 150992 79024 151044 79076
rect 173440 79228 173492 79280
rect 174498 79908 174550 79960
rect 174314 79840 174366 79892
rect 174406 79840 174458 79892
rect 174176 79568 174228 79620
rect 174498 79772 174550 79824
rect 177856 80044 177908 80096
rect 186504 80044 186556 80096
rect 302240 80044 302292 80096
rect 174682 79908 174734 79960
rect 174958 79840 175010 79892
rect 175510 79908 175562 79960
rect 175694 79840 175746 79892
rect 175878 79840 175930 79892
rect 177948 79976 178000 80028
rect 178040 79976 178092 80028
rect 176246 79908 176298 79960
rect 176338 79908 176390 79960
rect 178684 79908 178736 79960
rect 175464 79772 175516 79824
rect 177074 79840 177126 79892
rect 177764 79840 177816 79892
rect 176292 79772 176344 79824
rect 176522 79772 176574 79824
rect 177258 79772 177310 79824
rect 177856 79772 177908 79824
rect 199476 79772 199528 79824
rect 174544 79636 174596 79688
rect 174452 79568 174504 79620
rect 175924 79704 175976 79756
rect 176476 79636 176528 79688
rect 175280 79568 175332 79620
rect 175648 79568 175700 79620
rect 198004 79704 198056 79756
rect 178132 79568 178184 79620
rect 197636 79568 197688 79620
rect 174728 79432 174780 79484
rect 175004 79432 175056 79484
rect 178316 79500 178368 79552
rect 193956 79500 194008 79552
rect 194508 79500 194560 79552
rect 176936 79432 176988 79484
rect 178224 79432 178276 79484
rect 238760 79432 238812 79484
rect 177396 79364 177448 79416
rect 189908 79364 189960 79416
rect 175188 79296 175240 79348
rect 178040 79296 178092 79348
rect 181904 79296 181956 79348
rect 191288 79296 191340 79348
rect 194508 79296 194560 79348
rect 448520 79296 448572 79348
rect 175832 79228 175884 79280
rect 202328 79228 202380 79280
rect 173532 79160 173584 79212
rect 203708 79160 203760 79212
rect 166172 79092 166224 79144
rect 178408 79092 178460 79144
rect 171140 79024 171192 79076
rect 173256 79024 173308 79076
rect 174544 79024 174596 79076
rect 174820 79024 174872 79076
rect 175832 79024 175884 79076
rect 176752 79024 176804 79076
rect 177212 79024 177264 79076
rect 180156 79092 180208 79144
rect 183744 79092 183796 79144
rect 285680 79092 285732 79144
rect 376760 79024 376812 79076
rect 119252 78956 119304 79008
rect 151544 78956 151596 79008
rect 153108 78956 153160 79008
rect 154672 78956 154724 79008
rect 180156 78956 180208 79008
rect 198096 78956 198148 79008
rect 483020 78956 483072 79008
rect 116492 78888 116544 78940
rect 148140 78888 148192 78940
rect 121092 78820 121144 78872
rect 125600 78820 125652 78872
rect 129556 78820 129608 78872
rect 142160 78820 142212 78872
rect 147956 78820 148008 78872
rect 161664 78820 161716 78872
rect 166172 78820 166224 78872
rect 171600 78888 171652 78940
rect 178040 78888 178092 78940
rect 179328 78888 179380 78940
rect 195244 78888 195296 78940
rect 500960 78888 501012 78940
rect 179972 78820 180024 78872
rect 198004 78820 198056 78872
rect 523132 78820 523184 78872
rect 130660 78752 130712 78804
rect 144920 78752 144972 78804
rect 166264 78752 166316 78804
rect 167000 78752 167052 78804
rect 176200 78752 176252 78804
rect 178684 78752 178736 78804
rect 197636 78752 197688 78804
rect 525800 78752 525852 78804
rect 142068 78684 142120 78736
rect 149520 78684 149572 78736
rect 150164 78684 150216 78736
rect 160192 78684 160244 78736
rect 195428 78684 195480 78736
rect 200764 78684 200816 78736
rect 201408 78684 201460 78736
rect 536840 78684 536892 78736
rect 132316 78616 132368 78668
rect 135260 78616 135312 78668
rect 135904 78616 135956 78668
rect 136732 78616 136784 78668
rect 136916 78616 136968 78668
rect 137100 78616 137152 78668
rect 137744 78616 137796 78668
rect 141240 78616 141292 78668
rect 141516 78616 141568 78668
rect 102140 78548 102192 78600
rect 102876 78548 102928 78600
rect 133880 78548 133932 78600
rect 137284 78548 137336 78600
rect 137836 78548 137888 78600
rect 142436 78616 142488 78668
rect 143908 78616 143960 78668
rect 150072 78616 150124 78668
rect 157984 78616 158036 78668
rect 158444 78616 158496 78668
rect 162032 78616 162084 78668
rect 162400 78616 162452 78668
rect 141976 78548 142028 78600
rect 142712 78548 142764 78600
rect 162952 78548 163004 78600
rect 163228 78548 163280 78600
rect 164424 78548 164476 78600
rect 165528 78548 165580 78600
rect 75920 78480 75972 78532
rect 106832 78480 106884 78532
rect 107200 78480 107252 78532
rect 137376 78480 137428 78532
rect 137744 78480 137796 78532
rect 141516 78480 141568 78532
rect 141700 78480 141752 78532
rect 157616 78480 157668 78532
rect 161664 78480 161716 78532
rect 164240 78480 164292 78532
rect 164884 78480 164936 78532
rect 175188 78616 175240 78668
rect 177028 78616 177080 78668
rect 206284 78616 206336 78668
rect 174084 78548 174136 78600
rect 178960 78548 179012 78600
rect 179328 78548 179380 78600
rect 206468 78548 206520 78600
rect 168472 78480 168524 78532
rect 193588 78480 193640 78532
rect 194508 78480 194560 78532
rect 60740 78276 60792 78328
rect 107108 78412 107160 78464
rect 137192 78412 137244 78464
rect 144184 78412 144236 78464
rect 152372 78412 152424 78464
rect 166264 78412 166316 78464
rect 167644 78412 167696 78464
rect 177396 78412 177448 78464
rect 179972 78412 180024 78464
rect 183468 78412 183520 78464
rect 206192 78412 206244 78464
rect 107016 78344 107068 78396
rect 107200 78344 107252 78396
rect 135996 78344 136048 78396
rect 137560 78344 137612 78396
rect 142620 78344 142672 78396
rect 148140 78344 148192 78396
rect 148876 78344 148928 78396
rect 157432 78344 157484 78396
rect 157708 78344 157760 78396
rect 163964 78344 164016 78396
rect 166172 78344 166224 78396
rect 168288 78344 168340 78396
rect 202236 78344 202288 78396
rect 57980 78208 58032 78260
rect 108488 78208 108540 78260
rect 135720 78276 135772 78328
rect 138112 78276 138164 78328
rect 138756 78276 138808 78328
rect 140136 78276 140188 78328
rect 140504 78276 140556 78328
rect 146576 78276 146628 78328
rect 171876 78276 171928 78328
rect 183008 78276 183060 78328
rect 204812 78276 204864 78328
rect 122472 78208 122524 78260
rect 148324 78208 148376 78260
rect 149336 78208 149388 78260
rect 183560 78208 183612 78260
rect 46940 78140 46992 78192
rect 107200 78140 107252 78192
rect 34520 78072 34572 78124
rect 100760 78072 100812 78124
rect 20720 78004 20772 78056
rect 102140 78004 102192 78056
rect 2780 77936 2832 77988
rect 108580 78072 108632 78124
rect 130936 78140 130988 78192
rect 130844 78072 130896 78124
rect 137652 78140 137704 78192
rect 139860 78140 139912 78192
rect 140228 78140 140280 78192
rect 159824 78140 159876 78192
rect 167276 78140 167328 78192
rect 170036 78140 170088 78192
rect 132684 78072 132736 78124
rect 142436 78072 142488 78124
rect 152004 78072 152056 78124
rect 152556 78072 152608 78124
rect 156144 78072 156196 78124
rect 163044 78072 163096 78124
rect 172428 78140 172480 78192
rect 255964 78140 256016 78192
rect 106924 78004 106976 78056
rect 129924 78004 129976 78056
rect 130384 78004 130436 78056
rect 150164 78004 150216 78056
rect 160100 78004 160152 78056
rect 161112 78004 161164 78056
rect 337384 78072 337436 78124
rect 393320 78004 393372 78056
rect 122840 77936 122892 77988
rect 148416 77936 148468 77988
rect 148600 77936 148652 77988
rect 148876 77936 148928 77988
rect 169668 77936 169720 77988
rect 400864 77936 400916 77988
rect 130936 77868 130988 77920
rect 132684 77868 132736 77920
rect 137836 77868 137888 77920
rect 146760 77868 146812 77920
rect 166724 77868 166776 77920
rect 182824 77868 182876 77920
rect 131212 77800 131264 77852
rect 132132 77800 132184 77852
rect 141976 77800 142028 77852
rect 161940 77800 161992 77852
rect 168656 77800 168708 77852
rect 171876 77800 171928 77852
rect 180708 77800 180760 77852
rect 183008 77800 183060 77852
rect 100760 77732 100812 77784
rect 101496 77732 101548 77784
rect 134984 77732 135036 77784
rect 146944 77732 146996 77784
rect 147404 77732 147456 77784
rect 157064 77732 157116 77784
rect 157432 77732 157484 77784
rect 165804 77732 165856 77784
rect 181628 77732 181680 77784
rect 133972 77664 134024 77716
rect 140044 77664 140096 77716
rect 142712 77664 142764 77716
rect 143264 77664 143316 77716
rect 165436 77664 165488 77716
rect 181904 77664 181956 77716
rect 106832 77596 106884 77648
rect 136732 77596 136784 77648
rect 147772 77596 147824 77648
rect 148508 77596 148560 77648
rect 166448 77596 166500 77648
rect 178776 77596 178828 77648
rect 131672 77528 131724 77580
rect 142252 77528 142304 77580
rect 143080 77528 143132 77580
rect 143264 77528 143316 77580
rect 143448 77528 143500 77580
rect 144184 77528 144236 77580
rect 148324 77528 148376 77580
rect 148600 77528 148652 77580
rect 146760 77460 146812 77512
rect 147312 77460 147364 77512
rect 165528 77460 165580 77512
rect 180340 77460 180392 77512
rect 134340 77392 134392 77444
rect 134800 77392 134852 77444
rect 140780 77392 140832 77444
rect 141240 77392 141292 77444
rect 134800 77256 134852 77308
rect 136916 77256 136968 77308
rect 140504 77256 140556 77308
rect 142988 77256 143040 77308
rect 143632 77256 143684 77308
rect 143724 77256 143776 77308
rect 143908 77256 143960 77308
rect 145012 77256 145064 77308
rect 146116 77256 146168 77308
rect 126980 77188 127032 77240
rect 127624 77188 127676 77240
rect 129648 77188 129700 77240
rect 136640 77188 136692 77240
rect 137192 77188 137244 77240
rect 151268 77188 151320 77240
rect 151820 77256 151872 77308
rect 162308 77256 162360 77308
rect 163596 77256 163648 77308
rect 170864 77256 170916 77308
rect 171140 77256 171192 77308
rect 177028 77256 177080 77308
rect 177672 77256 177724 77308
rect 194508 77256 194560 77308
rect 269764 77256 269816 77308
rect 196716 77188 196768 77240
rect 119712 77120 119764 77172
rect 153476 77120 153528 77172
rect 162308 77120 162360 77172
rect 169760 77120 169812 77172
rect 203156 77120 203208 77172
rect 115664 77052 115716 77104
rect 66260 76644 66312 76696
rect 104072 76984 104124 77036
rect 137468 76984 137520 77036
rect 155408 77052 155460 77104
rect 187424 77052 187476 77104
rect 188804 77052 188856 77104
rect 148232 76984 148284 77036
rect 171600 76984 171652 77036
rect 191472 76984 191524 77036
rect 191748 76984 191800 77036
rect 117228 76916 117280 76968
rect 148784 76916 148836 76968
rect 154856 76916 154908 76968
rect 184480 76916 184532 76968
rect 120540 76848 120592 76900
rect 115756 76780 115808 76832
rect 59360 76576 59412 76628
rect 108304 76712 108356 76764
rect 106372 76644 106424 76696
rect 131672 76644 131724 76696
rect 151084 76848 151136 76900
rect 156972 76780 157024 76832
rect 157156 76780 157208 76832
rect 172520 76848 172572 76900
rect 173532 76848 173584 76900
rect 184204 76848 184256 76900
rect 200856 76848 200908 76900
rect 224224 76780 224276 76832
rect 151268 76712 151320 76764
rect 247040 76712 247092 76764
rect 146024 76644 146076 76696
rect 151084 76644 151136 76696
rect 153108 76644 153160 76696
rect 253940 76644 253992 76696
rect 134800 76576 134852 76628
rect 150716 76576 150768 76628
rect 150900 76576 150952 76628
rect 52460 76508 52512 76560
rect 135996 76508 136048 76560
rect 150072 76508 150124 76560
rect 181352 76576 181404 76628
rect 191748 76576 191800 76628
rect 353300 76576 353352 76628
rect 162584 76508 162636 76560
rect 389180 76508 389232 76560
rect 123024 76440 123076 76492
rect 141608 76440 141660 76492
rect 114376 76372 114428 76424
rect 141056 76372 141108 76424
rect 177212 76372 177264 76424
rect 207112 76372 207164 76424
rect 115480 76304 115532 76356
rect 149796 76304 149848 76356
rect 169760 76304 169812 76356
rect 170588 76304 170640 76356
rect 173348 76304 173400 76356
rect 184204 76304 184256 76356
rect 131672 76236 131724 76288
rect 139584 76236 139636 76288
rect 164424 76236 164476 76288
rect 165436 76236 165488 76288
rect 173440 76236 173492 76288
rect 173716 76236 173768 76288
rect 129648 76168 129700 76220
rect 141792 76168 141844 76220
rect 143356 76168 143408 76220
rect 144736 76168 144788 76220
rect 165252 76100 165304 76152
rect 165436 76100 165488 76152
rect 145380 76032 145432 76084
rect 146024 76032 146076 76084
rect 173072 75964 173124 76016
rect 173808 75964 173860 76016
rect 174360 75964 174412 76016
rect 175188 75964 175240 76016
rect 184480 75964 184532 76016
rect 289820 75964 289872 76016
rect 111800 75896 111852 75948
rect 113640 75896 113692 75948
rect 114376 75896 114428 75948
rect 134524 75896 134576 75948
rect 134708 75896 134760 75948
rect 173900 75896 173952 75948
rect 174544 75896 174596 75948
rect 177212 75896 177264 75948
rect 177672 75896 177724 75948
rect 188804 75896 188856 75948
rect 296720 75896 296772 75948
rect 118240 75828 118292 75880
rect 145104 75828 145156 75880
rect 148324 75828 148376 75880
rect 168840 75828 168892 75880
rect 169576 75828 169628 75880
rect 105544 75760 105596 75812
rect 139492 75760 139544 75812
rect 161388 75760 161440 75812
rect 195520 75760 195572 75812
rect 113732 75692 113784 75744
rect 146668 75692 146720 75744
rect 156328 75692 156380 75744
rect 156696 75692 156748 75744
rect 190644 75692 190696 75744
rect 113088 75624 113140 75676
rect 145656 75624 145708 75676
rect 146484 75624 146536 75676
rect 180800 75624 180852 75676
rect 114100 75488 114152 75540
rect 120724 75556 120776 75608
rect 135444 75556 135496 75608
rect 148048 75556 148100 75608
rect 181536 75556 181588 75608
rect 104256 75420 104308 75472
rect 120724 75420 120776 75472
rect 134064 75420 134116 75472
rect 134524 75420 134576 75472
rect 147680 75488 147732 75540
rect 198740 75488 198792 75540
rect 147128 75420 147180 75472
rect 187700 75420 187752 75472
rect 114468 75352 114520 75404
rect 145472 75352 145524 75404
rect 148876 75352 148928 75404
rect 201500 75352 201552 75404
rect 96620 75284 96672 75336
rect 108764 75284 108816 75336
rect 140228 75284 140280 75336
rect 173256 75284 173308 75336
rect 453304 75284 453356 75336
rect 81440 75216 81492 75268
rect 138756 75216 138808 75268
rect 149428 75216 149480 75268
rect 150072 75216 150124 75268
rect 163044 75216 163096 75268
rect 163688 75216 163740 75268
rect 172888 75216 172940 75268
rect 506480 75216 506532 75268
rect 27620 75148 27672 75200
rect 100116 75148 100168 75200
rect 141424 75148 141476 75200
rect 163136 75148 163188 75200
rect 164056 75148 164108 75200
rect 172336 75148 172388 75200
rect 511264 75148 511316 75200
rect 114560 75080 114612 75132
rect 115112 75080 115164 75132
rect 121276 75080 121328 75132
rect 147220 75080 147272 75132
rect 167828 75080 167880 75132
rect 192668 75080 192720 75132
rect 132408 75012 132460 75064
rect 114008 74944 114060 74996
rect 146484 74944 146536 74996
rect 155868 74944 155920 74996
rect 156788 74944 156840 74996
rect 190736 74944 190788 74996
rect 173992 74876 174044 74928
rect 174912 74876 174964 74928
rect 145656 74808 145708 74860
rect 145932 74808 145984 74860
rect 173992 74740 174044 74792
rect 174268 74740 174320 74792
rect 165068 74604 165120 74656
rect 178868 74604 178920 74656
rect 121368 74468 121420 74520
rect 131120 74468 131172 74520
rect 132316 74468 132368 74520
rect 143908 74468 143960 74520
rect 144460 74468 144512 74520
rect 145564 74468 145616 74520
rect 145840 74468 145892 74520
rect 154028 74468 154080 74520
rect 154212 74468 154264 74520
rect 157892 74468 157944 74520
rect 158168 74468 158220 74520
rect 192300 74468 192352 74520
rect 110144 74400 110196 74452
rect 144644 74400 144696 74452
rect 161204 74400 161256 74452
rect 164884 74400 164936 74452
rect 167000 74400 167052 74452
rect 200580 74400 200632 74452
rect 115572 74332 115624 74384
rect 112720 74264 112772 74316
rect 146116 74264 146168 74316
rect 111156 74196 111208 74248
rect 143172 74196 143224 74248
rect 153384 74332 153436 74384
rect 154212 74332 154264 74384
rect 188528 74332 188580 74384
rect 160744 74264 160796 74316
rect 161296 74264 161348 74316
rect 171324 74264 171376 74316
rect 172152 74264 172204 74316
rect 175372 74264 175424 74316
rect 176200 74264 176252 74316
rect 205916 74264 205968 74316
rect 149980 74196 150032 74248
rect 203708 74196 203760 74248
rect 104348 74128 104400 74180
rect 134248 74128 134300 74180
rect 135168 74128 135220 74180
rect 136916 74128 136968 74180
rect 137928 74128 137980 74180
rect 152740 74128 152792 74180
rect 262220 74128 262272 74180
rect 116676 74060 116728 74112
rect 145840 74060 145892 74112
rect 154488 74060 154540 74112
rect 284300 74060 284352 74112
rect 118056 73992 118108 74044
rect 144000 73992 144052 74044
rect 144276 73992 144328 74044
rect 144644 73992 144696 74044
rect 155960 73992 156012 74044
rect 297364 73992 297416 74044
rect 119620 73924 119672 73976
rect 99380 73856 99432 73908
rect 140320 73856 140372 73908
rect 144092 73924 144144 73976
rect 149704 73924 149756 73976
rect 159180 73924 159232 73976
rect 347780 73924 347832 73976
rect 145196 73856 145248 73908
rect 153476 73856 153528 73908
rect 269120 73856 269172 73908
rect 269764 73856 269816 73908
rect 465172 73856 465224 73908
rect 78680 73788 78732 73840
rect 138296 73788 138348 73840
rect 151728 73788 151780 73840
rect 248420 73788 248472 73840
rect 255964 73788 256016 73840
rect 456800 73788 456852 73840
rect 119528 73720 119580 73772
rect 144460 73720 144512 73772
rect 153200 73720 153252 73772
rect 154304 73720 154356 73772
rect 171324 73720 171376 73772
rect 171692 73720 171744 73772
rect 175556 73720 175608 73772
rect 176476 73720 176528 73772
rect 206008 73720 206060 73772
rect 124864 73652 124916 73704
rect 125600 73652 125652 73704
rect 132684 73652 132736 73704
rect 133696 73652 133748 73704
rect 172152 73652 172204 73704
rect 194968 73652 195020 73704
rect 114744 73584 114796 73636
rect 149152 73584 149204 73636
rect 149980 73584 150032 73636
rect 168472 73584 168524 73636
rect 169208 73584 169260 73636
rect 166356 73516 166408 73568
rect 183744 73516 183796 73568
rect 145196 73448 145248 73500
rect 145656 73448 145708 73500
rect 164332 73176 164384 73228
rect 164976 73176 165028 73228
rect 118608 73108 118660 73160
rect 152280 73108 152332 73160
rect 163320 73108 163372 73160
rect 163688 73108 163740 73160
rect 167184 73108 167236 73160
rect 208492 73108 208544 73160
rect 109868 73040 109920 73092
rect 143908 73040 143960 73092
rect 147036 73040 147088 73092
rect 168104 73040 168156 73092
rect 202144 73040 202196 73092
rect 102140 72972 102192 73024
rect 102784 72972 102836 73024
rect 135536 72972 135588 73024
rect 155224 72972 155276 73024
rect 155408 72972 155460 73024
rect 190000 72972 190052 73024
rect 105728 72904 105780 72956
rect 139308 72904 139360 72956
rect 163688 72904 163740 72956
rect 198188 72904 198240 72956
rect 108672 72836 108724 72888
rect 140596 72836 140648 72888
rect 159640 72836 159692 72888
rect 189816 72836 189868 72888
rect 111248 72768 111300 72820
rect 142804 72768 142856 72820
rect 146668 72768 146720 72820
rect 180340 72768 180392 72820
rect 181996 72768 182048 72820
rect 204260 72768 204312 72820
rect 327724 73108 327776 73160
rect 579988 73108 580040 73160
rect 220084 72768 220136 72820
rect 111432 72700 111484 72752
rect 143080 72700 143132 72752
rect 156604 72700 156656 72752
rect 311164 72700 311216 72752
rect 85580 72632 85632 72684
rect 105728 72632 105780 72684
rect 119804 72632 119856 72684
rect 144368 72632 144420 72684
rect 157248 72632 157300 72684
rect 318800 72632 318852 72684
rect 43444 72564 43496 72616
rect 102140 72564 102192 72616
rect 122104 72564 122156 72616
rect 123024 72564 123076 72616
rect 124220 72564 124272 72616
rect 140780 72564 140832 72616
rect 157800 72564 157852 72616
rect 324964 72564 325016 72616
rect 67640 72496 67692 72548
rect 137744 72496 137796 72548
rect 158260 72496 158312 72548
rect 332600 72496 332652 72548
rect 14464 72428 14516 72480
rect 111616 72428 111668 72480
rect 130016 72428 130068 72480
rect 131028 72428 131080 72480
rect 132500 72428 132552 72480
rect 133512 72428 133564 72480
rect 167092 72428 167144 72480
rect 168380 72428 168432 72480
rect 168656 72428 168708 72480
rect 375380 72428 375432 72480
rect 104532 72360 104584 72412
rect 129096 72360 129148 72412
rect 161664 72360 161716 72412
rect 179696 72360 179748 72412
rect 180616 72360 180668 72412
rect 171508 72292 171560 72344
rect 172244 72292 172296 72344
rect 178408 72292 178460 72344
rect 181996 72292 182048 72344
rect 156420 72224 156472 72276
rect 181260 72224 181312 72276
rect 152280 72088 152332 72140
rect 152740 72088 152792 72140
rect 160192 72020 160244 72072
rect 160560 72020 160612 72072
rect 181260 71816 181312 71868
rect 304264 71816 304316 71868
rect 107660 71748 107712 71800
rect 108672 71748 108724 71800
rect 118332 71680 118384 71732
rect 151912 71680 151964 71732
rect 152648 71680 152700 71732
rect 157708 71680 157760 71732
rect 158076 71680 158128 71732
rect 158352 71680 158404 71732
rect 158628 71680 158680 71732
rect 159088 71680 159140 71732
rect 159916 71680 159968 71732
rect 3516 71612 3568 71664
rect 8944 71612 8996 71664
rect 116308 71612 116360 71664
rect 151176 71612 151228 71664
rect 159548 71612 159600 71664
rect 161756 71612 161808 71664
rect 162584 71612 162636 71664
rect 180616 71748 180668 71800
rect 322940 71748 322992 71800
rect 183560 71680 183612 71732
rect 204720 71680 204772 71732
rect 194324 71612 194376 71664
rect 121184 71544 121236 71596
rect 152464 71544 152516 71596
rect 161112 71544 161164 71596
rect 195152 71544 195204 71596
rect 102140 71476 102192 71528
rect 102968 71476 103020 71528
rect 134708 71476 134760 71528
rect 135444 71476 135496 71528
rect 136548 71476 136600 71528
rect 141424 71476 141476 71528
rect 142804 71476 142856 71528
rect 160376 71476 160428 71528
rect 162124 71476 162176 71528
rect 162584 71476 162636 71528
rect 196808 71476 196860 71528
rect 112168 71408 112220 71460
rect 142436 71408 142488 71460
rect 143264 71408 143316 71460
rect 159916 71408 159968 71460
rect 193864 71408 193916 71460
rect 105636 71340 105688 71392
rect 135444 71340 135496 71392
rect 142804 71340 142856 71392
rect 143172 71340 143224 71392
rect 161572 71340 161624 71392
rect 196900 71340 196952 71392
rect 107476 71272 107528 71324
rect 135720 71272 135772 71324
rect 102784 71204 102836 71256
rect 106740 71204 106792 71256
rect 53840 71136 53892 71188
rect 113548 71204 113600 71256
rect 142160 71272 142212 71324
rect 143448 71272 143500 71324
rect 172428 71272 172480 71324
rect 200396 71272 200448 71324
rect 158996 71204 159048 71256
rect 193496 71204 193548 71256
rect 112536 71136 112588 71188
rect 138020 71136 138072 71188
rect 139124 71136 139176 71188
rect 142988 71136 143040 71188
rect 143448 71136 143500 71188
rect 158628 71136 158680 71188
rect 191196 71136 191248 71188
rect 31024 71068 31076 71120
rect 102140 71068 102192 71120
rect 116216 71068 116268 71120
rect 128360 71068 128412 71120
rect 129556 71068 129608 71120
rect 158444 71068 158496 71120
rect 191104 71068 191156 71120
rect 204720 71136 204772 71188
rect 217324 71136 217376 71188
rect 336004 71068 336056 71120
rect 31760 71000 31812 71052
rect 133420 71000 133472 71052
rect 160836 71000 160888 71052
rect 192576 71000 192628 71052
rect 367100 71000 367152 71052
rect 174912 70932 174964 70984
rect 204352 70932 204404 70984
rect 162584 70864 162636 70916
rect 186412 70864 186464 70916
rect 158076 70796 158128 70848
rect 192760 70796 192812 70848
rect 159640 70456 159692 70508
rect 160008 70456 160060 70508
rect 168380 70388 168432 70440
rect 169116 70388 169168 70440
rect 192116 70388 192168 70440
rect 192300 70388 192352 70440
rect 100300 70320 100352 70372
rect 134156 70320 134208 70372
rect 166724 70320 166776 70372
rect 200672 70320 200724 70372
rect 102140 70252 102192 70304
rect 103060 70252 103112 70304
rect 137008 70252 137060 70304
rect 165252 70252 165304 70304
rect 199384 70252 199436 70304
rect 105912 70184 105964 70236
rect 139584 70184 139636 70236
rect 165712 70184 165764 70236
rect 166356 70184 166408 70236
rect 200488 70184 200540 70236
rect 100392 70116 100444 70168
rect 132500 70116 132552 70168
rect 165528 70116 165580 70168
rect 199752 70116 199804 70168
rect 102232 70048 102284 70100
rect 103244 70048 103296 70100
rect 133604 70048 133656 70100
rect 164056 70048 164108 70100
rect 197728 70048 197780 70100
rect 116768 69980 116820 70032
rect 138204 69980 138256 70032
rect 164608 69980 164660 70032
rect 199016 69980 199068 70032
rect 164516 69912 164568 69964
rect 165252 69912 165304 69964
rect 62120 69844 62172 69896
rect 102140 69844 102192 69896
rect 103520 69844 103572 69896
rect 105912 69844 105964 69896
rect 163136 69844 163188 69896
rect 163964 69844 164016 69896
rect 85672 69776 85724 69828
rect 138112 69776 138164 69828
rect 163228 69776 163280 69828
rect 164056 69776 164108 69828
rect 164700 69844 164752 69896
rect 165528 69844 165580 69896
rect 196532 69912 196584 69964
rect 168932 69844 168984 69896
rect 169392 69844 169444 69896
rect 171048 69844 171100 69896
rect 199108 69844 199160 69896
rect 167276 69776 167328 69828
rect 354680 69776 354732 69828
rect 18604 69708 18656 69760
rect 102232 69708 102284 69760
rect 147128 69708 147180 69760
rect 185584 69708 185636 69760
rect 199016 69708 199068 69760
rect 199292 69708 199344 69760
rect 412640 69708 412692 69760
rect 45560 69640 45612 69692
rect 135260 69640 135312 69692
rect 148232 69640 148284 69692
rect 144000 69572 144052 69624
rect 147128 69572 147180 69624
rect 168748 69572 168800 69624
rect 169484 69572 169536 69624
rect 176936 69572 176988 69624
rect 191932 69640 191984 69692
rect 192116 69640 192168 69692
rect 199108 69640 199160 69692
rect 199660 69640 199712 69692
rect 498200 69640 498252 69692
rect 146392 69504 146444 69556
rect 179420 69504 179472 69556
rect 196624 69572 196676 69624
rect 195152 69504 195204 69556
rect 153752 69368 153804 69420
rect 181168 69368 181220 69420
rect 195152 69028 195204 69080
rect 529940 69028 529992 69080
rect 116124 68960 116176 69012
rect 118516 68892 118568 68944
rect 106004 68824 106056 68876
rect 138664 68824 138716 68876
rect 140780 68824 140832 68876
rect 142160 68824 142212 68876
rect 110236 68756 110288 68808
rect 142252 68756 142304 68808
rect 142712 68756 142764 68808
rect 144460 68960 144512 69012
rect 146300 68960 146352 69012
rect 150624 68960 150676 69012
rect 151176 68960 151228 69012
rect 167368 68960 167420 69012
rect 168012 68960 168064 69012
rect 201960 68960 202012 69012
rect 150624 68824 150676 68876
rect 152556 68892 152608 68944
rect 161756 68892 161808 68944
rect 162492 68892 162544 68944
rect 168840 68892 168892 68944
rect 169576 68892 169628 68944
rect 203616 68892 203668 68944
rect 161572 68824 161624 68876
rect 162400 68824 162452 68876
rect 169484 68824 169536 68876
rect 203432 68824 203484 68876
rect 169392 68756 169444 68808
rect 203524 68756 203576 68808
rect 104440 68688 104492 68740
rect 104624 68688 104676 68740
rect 135720 68688 135772 68740
rect 183836 68688 183888 68740
rect 203064 68688 203116 68740
rect 204168 68688 204220 68740
rect 114284 68620 114336 68672
rect 142344 68620 142396 68672
rect 142896 68620 142948 68672
rect 163044 68620 163096 68672
rect 188252 68620 188304 68672
rect 111156 68552 111208 68604
rect 112260 68552 112312 68604
rect 180708 68552 180760 68604
rect 182180 68552 182232 68604
rect 176752 68484 176804 68536
rect 201408 68552 201460 68604
rect 120080 68416 120132 68468
rect 141608 68416 141660 68468
rect 89720 68348 89772 68400
rect 106004 68348 106056 68400
rect 117320 68348 117372 68400
rect 141148 68348 141200 68400
rect 48320 68280 48372 68332
rect 104624 68280 104676 68332
rect 113180 68280 113232 68332
rect 140964 68280 141016 68332
rect 204168 68280 204220 68332
rect 464344 68280 464396 68332
rect 188252 67668 188304 67720
rect 402980 67668 403032 67720
rect 201408 67600 201460 67652
rect 552664 67600 552716 67652
rect 106004 67532 106056 67584
rect 137100 67532 137152 67584
rect 146024 67532 146076 67584
rect 148416 67532 148468 67584
rect 155132 67532 155184 67584
rect 189172 67532 189224 67584
rect 104532 67464 104584 67516
rect 134800 67464 134852 67516
rect 72424 66920 72476 66972
rect 106004 66920 106056 66972
rect 35164 66852 35216 66904
rect 104532 66852 104584 66904
rect 189172 66852 189224 66904
rect 295340 66852 295392 66904
rect 102140 66172 102192 66224
rect 103152 66172 103204 66224
rect 137192 66172 137244 66224
rect 157340 66172 157392 66224
rect 192300 66172 192352 66224
rect 193128 66172 193180 66224
rect 159364 66104 159416 66156
rect 188068 66104 188120 66156
rect 177120 66036 177172 66088
rect 197544 66036 197596 66088
rect 148784 65560 148836 65612
rect 207020 65560 207072 65612
rect 58624 65492 58676 65544
rect 102140 65492 102192 65544
rect 193128 65492 193180 65544
rect 324320 65492 324372 65544
rect 188620 64948 188672 65000
rect 346400 64948 346452 65000
rect 197544 64880 197596 64932
rect 574744 64880 574796 64932
rect 102140 64812 102192 64864
rect 106096 64812 106148 64864
rect 139860 64812 139912 64864
rect 160468 64812 160520 64864
rect 194876 64812 194928 64864
rect 108948 64744 109000 64796
rect 138480 64744 138532 64796
rect 169024 64744 169076 64796
rect 202972 64744 203024 64796
rect 149796 64268 149848 64320
rect 224960 64268 225012 64320
rect 84844 64200 84896 64252
rect 108948 64200 109000 64252
rect 194876 64200 194928 64252
rect 358820 64200 358872 64252
rect 35900 64132 35952 64184
rect 134340 64132 134392 64184
rect 147312 64132 147364 64184
rect 183560 64132 183612 64184
rect 202972 64132 203024 64184
rect 472624 64132 472676 64184
rect 140044 63520 140096 63572
rect 142988 63520 143040 63572
rect 146116 63520 146168 63572
rect 147220 63520 147272 63572
rect 104716 63452 104768 63504
rect 132776 63452 132828 63504
rect 159456 63452 159508 63504
rect 193404 63452 193456 63504
rect 144368 63044 144420 63096
rect 149796 63044 149848 63096
rect 150256 62840 150308 62892
rect 227720 62840 227772 62892
rect 10324 62772 10376 62824
rect 104716 62772 104768 62824
rect 147404 62772 147456 62824
rect 190460 62772 190512 62824
rect 193404 62772 193456 62824
rect 349160 62772 349212 62824
rect 139400 62296 139452 62348
rect 142804 62296 142856 62348
rect 102232 62024 102284 62076
rect 103428 62024 103480 62076
rect 134432 62024 134484 62076
rect 26240 61412 26292 61464
rect 102232 61412 102284 61464
rect 44824 61344 44876 61396
rect 135628 61344 135680 61396
rect 154764 61208 154816 61260
rect 155224 61208 155276 61260
rect 99472 60664 99524 60716
rect 100576 60664 100628 60716
rect 132684 60664 132736 60716
rect 166172 60664 166224 60716
rect 197452 60664 197504 60716
rect 197820 60664 197872 60716
rect 162952 60596 163004 60648
rect 189356 60596 189408 60648
rect 151912 60120 151964 60172
rect 263600 60120 263652 60172
rect 197452 60052 197504 60104
rect 396080 60052 396132 60104
rect 22744 59984 22796 60036
rect 99472 59984 99524 60036
rect 145932 59984 145984 60036
rect 147312 59984 147364 60036
rect 189356 59984 189408 60036
rect 398840 59984 398892 60036
rect 110420 59848 110472 59900
rect 115020 59848 115072 59900
rect 3516 59304 3568 59356
rect 111064 59304 111116 59356
rect 146392 58760 146444 58812
rect 186320 58760 186372 58812
rect 154028 58692 154080 58744
rect 281540 58692 281592 58744
rect 60832 58624 60884 58676
rect 137376 58624 137428 58676
rect 144276 58624 144328 58676
rect 156604 58624 156656 58676
rect 169300 58624 169352 58676
rect 467840 58624 467892 58676
rect 100760 57876 100812 57928
rect 101680 57876 101732 57928
rect 134524 57876 134576 57928
rect 168472 57876 168524 57928
rect 203340 57876 203392 57928
rect 204168 57876 204220 57928
rect 159272 57808 159324 57860
rect 194140 57808 194192 57860
rect 194508 57808 194560 57860
rect 149980 57400 150032 57452
rect 215300 57400 215352 57452
rect 152004 57332 152056 57384
rect 255320 57332 255372 57384
rect 194508 57264 194560 57316
rect 345020 57264 345072 57316
rect 22100 57196 22152 57248
rect 100760 57196 100812 57248
rect 204168 57196 204220 57248
rect 473452 57196 473504 57248
rect 99472 56516 99524 56568
rect 100668 56516 100720 56568
rect 132960 56516 133012 56568
rect 162860 56516 162912 56568
rect 197636 56516 197688 56568
rect 88340 55904 88392 55956
rect 138756 55904 138808 55956
rect 12440 55836 12492 55888
rect 99472 55836 99524 55888
rect 197636 55836 197688 55888
rect 394700 55836 394752 55888
rect 113824 55156 113876 55208
rect 140136 55156 140188 55208
rect 168380 55156 168432 55208
rect 202880 55156 202932 55208
rect 202880 54476 202932 54528
rect 468484 54476 468536 54528
rect 468576 54476 468628 54528
rect 581092 54476 581144 54528
rect 138664 53796 138716 53848
rect 142436 53796 142488 53848
rect 100484 53728 100536 53780
rect 132868 53728 132920 53780
rect 143632 53388 143684 53440
rect 147680 53388 147732 53440
rect 147864 53184 147916 53236
rect 197452 53184 197504 53236
rect 95240 53116 95292 53168
rect 139768 53116 139820 53168
rect 151544 53116 151596 53168
rect 237380 53116 237432 53168
rect 9680 53048 9732 53100
rect 100484 53048 100536 53100
rect 176016 53048 176068 53100
rect 556160 53048 556212 53100
rect 148140 51756 148192 51808
rect 211160 51756 211212 51808
rect 93952 51688 94004 51740
rect 105544 51688 105596 51740
rect 145840 51688 145892 51740
rect 168472 51688 168524 51740
rect 177488 51688 177540 51740
rect 578240 51688 578292 51740
rect 100760 51008 100812 51060
rect 101864 51008 101916 51060
rect 134616 51008 134668 51060
rect 147588 50396 147640 50448
rect 191840 50396 191892 50448
rect 30380 50328 30432 50380
rect 100760 50328 100812 50380
rect 164976 50328 165028 50380
rect 368480 50328 368532 50380
rect 148692 49240 148744 49292
rect 201592 49240 201644 49292
rect 150072 49036 150124 49088
rect 218152 49036 218204 49088
rect 171416 48968 171468 49020
rect 499580 48968 499632 49020
rect 152740 47676 152792 47728
rect 256700 47676 256752 47728
rect 166264 47608 166316 47660
rect 444380 47608 444432 47660
rect 174728 47540 174780 47592
rect 542360 47540 542412 47592
rect 148600 46248 148652 46300
rect 204260 46248 204312 46300
rect 144920 46180 144972 46232
rect 167000 46180 167052 46232
rect 167920 46180 167972 46232
rect 449900 46180 449952 46232
rect 135260 45568 135312 45620
rect 142344 45568 142396 45620
rect 167828 44956 167880 45008
rect 458180 44956 458232 45008
rect 175280 44888 175332 44940
rect 560300 44888 560352 44940
rect 177580 44820 177632 44872
rect 571984 44820 572036 44872
rect 149152 43596 149204 43648
rect 216680 43596 216732 43648
rect 162124 43528 162176 43580
rect 361580 43528 361632 43580
rect 164424 43460 164476 43512
rect 426440 43460 426492 43512
rect 63500 43392 63552 43444
rect 136640 43392 136692 43444
rect 172244 43392 172296 43444
rect 502340 43392 502392 43444
rect 150532 42304 150584 42356
rect 233240 42304 233292 42356
rect 155408 42236 155460 42288
rect 292672 42236 292724 42288
rect 158168 42168 158220 42220
rect 328460 42168 328512 42220
rect 172152 42100 172204 42152
rect 498292 42100 498344 42152
rect 70400 42032 70452 42084
rect 136916 42032 136968 42084
rect 174820 42032 174872 42084
rect 538864 42032 538916 42084
rect 155500 40944 155552 40996
rect 300860 40944 300912 40996
rect 156696 40876 156748 40928
rect 309140 40876 309192 40928
rect 166356 40808 166408 40860
rect 427820 40808 427872 40860
rect 167092 40740 167144 40792
rect 462320 40740 462372 40792
rect 74540 40672 74592 40724
rect 138204 40672 138256 40724
rect 173532 40672 173584 40724
rect 516140 40672 516192 40724
rect 152648 39584 152700 39636
rect 251180 39584 251232 39636
rect 163504 39516 163556 39568
rect 340972 39516 341024 39568
rect 169392 39448 169444 39500
rect 470600 39448 470652 39500
rect 170588 39380 170640 39432
rect 481640 39380 481692 39432
rect 77392 39312 77444 39364
rect 138296 39312 138348 39364
rect 174084 39312 174136 39364
rect 534080 39312 534132 39364
rect 154212 38156 154264 38208
rect 267832 38156 267884 38208
rect 161204 38088 161256 38140
rect 372620 38088 372672 38140
rect 170680 38020 170732 38072
rect 488540 38020 488592 38072
rect 173624 37952 173676 38004
rect 528560 37952 528612 38004
rect 13820 37884 13872 37936
rect 132500 37884 132552 37936
rect 176200 37884 176252 37936
rect 552020 37884 552072 37936
rect 147772 36864 147824 36916
rect 208400 36864 208452 36916
rect 149060 36796 149112 36848
rect 222200 36796 222252 36848
rect 156788 36728 156840 36780
rect 303620 36728 303672 36780
rect 165620 36660 165672 36712
rect 440332 36660 440384 36712
rect 175832 36592 175884 36644
rect 558920 36592 558972 36644
rect 104164 36524 104216 36576
rect 140412 36524 140464 36576
rect 177672 36524 177724 36576
rect 571340 36524 571392 36576
rect 153292 35436 153344 35488
rect 276020 35436 276072 35488
rect 158076 35368 158128 35420
rect 321560 35368 321612 35420
rect 165160 35300 165212 35352
rect 418160 35300 418212 35352
rect 170772 35232 170824 35284
rect 491300 35232 491352 35284
rect 38660 35164 38712 35216
rect 136364 35164 136416 35216
rect 145656 35164 145708 35216
rect 165620 35164 165672 35216
rect 177764 35164 177816 35216
rect 576860 35164 576912 35216
rect 155592 34008 155644 34060
rect 299572 34008 299624 34060
rect 162308 33940 162360 33992
rect 385040 33940 385092 33992
rect 169668 33872 169720 33924
rect 474740 33872 474792 33924
rect 170864 33804 170916 33856
rect 490012 33804 490064 33856
rect 175924 33736 175976 33788
rect 563704 33736 563756 33788
rect 148508 32648 148560 32700
rect 205640 32648 205692 32700
rect 150900 32580 150952 32632
rect 236000 32580 236052 32632
rect 161112 32512 161164 32564
rect 357440 32512 357492 32564
rect 173716 32444 173768 32496
rect 531412 32444 531464 32496
rect 176660 32376 176712 32428
rect 582380 32376 582432 32428
rect 156880 31220 156932 31272
rect 317420 31220 317472 31272
rect 164332 31152 164384 31204
rect 420920 31152 420972 31204
rect 169484 31084 169536 31136
rect 466460 31084 466512 31136
rect 177304 31016 177356 31068
rect 554780 31016 554832 31068
rect 151268 29860 151320 29912
rect 242992 29860 243044 29912
rect 157984 29792 158036 29844
rect 332692 29792 332744 29844
rect 161296 29724 161348 29776
rect 365812 29724 365864 29776
rect 166448 29656 166500 29708
rect 441620 29656 441672 29708
rect 171324 29588 171376 29640
rect 506572 29588 506624 29640
rect 159732 28432 159784 28484
rect 339500 28432 339552 28484
rect 163872 28364 163924 28416
rect 397460 28364 397512 28416
rect 169576 28296 169628 28348
rect 477500 28296 477552 28348
rect 52552 28228 52604 28280
rect 135444 28228 135496 28280
rect 171232 28228 171284 28280
rect 509240 28228 509292 28280
rect 153200 27140 153252 27192
rect 282920 27140 282972 27192
rect 162400 27072 162452 27124
rect 374092 27072 374144 27124
rect 165344 27004 165396 27056
rect 425060 27004 425112 27056
rect 171876 26936 171928 26988
rect 513380 26936 513432 26988
rect 35992 26868 36044 26920
rect 134248 26868 134300 26920
rect 174912 26868 174964 26920
rect 535460 26868 535512 26920
rect 156972 25780 157024 25832
rect 310520 25780 310572 25832
rect 163780 25712 163832 25764
rect 391940 25712 391992 25764
rect 181628 25644 181680 25696
rect 436100 25644 436152 25696
rect 172612 25576 172664 25628
rect 520280 25576 520332 25628
rect 145748 25508 145800 25560
rect 171784 25508 171836 25560
rect 175004 25508 175056 25560
rect 546500 25508 546552 25560
rect 157064 24352 157116 24404
rect 314660 24352 314712 24404
rect 165252 24284 165304 24336
rect 409880 24284 409932 24336
rect 182824 24216 182876 24268
rect 443000 24216 443052 24268
rect 172520 24148 172572 24200
rect 527180 24148 527232 24200
rect 40040 24080 40092 24132
rect 135352 24080 135404 24132
rect 145564 24080 145616 24132
rect 164884 24080 164936 24132
rect 176292 24080 176344 24132
rect 564532 24080 564584 24132
rect 144184 23468 144236 23520
rect 144920 23468 144972 23520
rect 150164 22992 150216 23044
rect 219440 22992 219492 23044
rect 157156 22924 157208 22976
rect 316132 22924 316184 22976
rect 164240 22856 164292 22908
rect 416780 22856 416832 22908
rect 168196 22788 168248 22840
rect 460940 22788 460992 22840
rect 173992 22720 174044 22772
rect 538220 22720 538272 22772
rect 157432 21632 157484 21684
rect 329840 21632 329892 21684
rect 157524 21564 157576 21616
rect 336740 21564 336792 21616
rect 337384 21564 337436 21616
rect 471980 21564 472032 21616
rect 158720 21496 158772 21548
rect 343640 21496 343692 21548
rect 159824 21428 159876 21480
rect 350540 21428 350592 21480
rect 178868 21360 178920 21412
rect 422300 21360 422352 21412
rect 286324 20612 286376 20664
rect 579988 20612 580040 20664
rect 154396 20204 154448 20256
rect 280160 20204 280212 20256
rect 155224 20136 155276 20188
rect 287060 20136 287112 20188
rect 155684 20068 155736 20120
rect 293960 20068 294012 20120
rect 161940 20000 161992 20052
rect 379520 20000 379572 20052
rect 155776 19932 155828 19984
rect 291200 19932 291252 19984
rect 291844 19932 291896 19984
rect 518900 19932 518952 19984
rect 153016 18844 153068 18896
rect 266360 18844 266412 18896
rect 160284 18776 160336 18828
rect 357532 18776 357584 18828
rect 166816 18708 166868 18760
rect 431960 18708 432012 18760
rect 176384 18640 176436 18692
rect 567200 18640 567252 18692
rect 177948 18572 178000 18624
rect 574100 18572 574152 18624
rect 151176 17484 151228 17536
rect 234712 17484 234764 17536
rect 180432 17416 180484 17468
rect 415492 17416 415544 17468
rect 168104 17348 168156 17400
rect 445760 17348 445812 17400
rect 168012 17280 168064 17332
rect 448612 17280 448664 17332
rect 171968 17212 172020 17264
rect 503720 17212 503772 17264
rect 152832 16056 152884 16108
rect 259552 16056 259604 16108
rect 160100 15988 160152 16040
rect 361120 15988 361172 16040
rect 160192 15920 160244 15972
rect 364616 15920 364668 15972
rect 400864 15920 400916 15972
rect 478880 15920 478932 15972
rect 166632 15852 166684 15904
rect 432052 15852 432104 15904
rect 153936 14696 153988 14748
rect 276112 14696 276164 14748
rect 158536 14628 158588 14680
rect 324412 14628 324464 14680
rect 178776 14560 178828 14612
rect 407212 14560 407264 14612
rect 163964 14492 164016 14544
rect 407120 14492 407172 14544
rect 172060 14424 172112 14476
rect 511264 14424 511316 14476
rect 152464 13268 152516 13320
rect 258264 13268 258316 13320
rect 156512 13200 156564 13252
rect 307944 13200 307996 13252
rect 164056 13132 164108 13184
rect 398932 13132 398984 13184
rect 170956 13064 171008 13116
rect 493048 13064 493100 13116
rect 152556 11908 152608 11960
rect 252376 11908 252428 11960
rect 160008 11840 160060 11892
rect 349252 11840 349304 11892
rect 166724 11772 166776 11824
rect 439136 11772 439188 11824
rect 175096 11704 175148 11756
rect 548616 11704 548668 11756
rect 201500 11636 201552 11688
rect 202696 11636 202748 11688
rect 234620 11636 234672 11688
rect 235816 11636 235868 11688
rect 259460 11636 259512 11688
rect 260656 11636 260708 11688
rect 151636 10548 151688 10600
rect 245200 10548 245252 10600
rect 159916 10480 159968 10532
rect 342904 10480 342956 10532
rect 162676 10412 162728 10464
rect 386696 10412 386748 10464
rect 166908 10344 166960 10396
rect 435088 10344 435140 10396
rect 176568 10276 176620 10328
rect 563060 10276 563112 10328
rect 150808 9188 150860 9240
rect 241704 9188 241756 9240
rect 161388 9120 161440 9172
rect 371700 9120 371752 9172
rect 164148 9052 164200 9104
rect 404820 9052 404872 9104
rect 168288 8984 168340 9036
rect 456892 8984 456944 9036
rect 176476 8916 176528 8968
rect 556160 8916 556212 8968
rect 150348 7828 150400 7880
rect 227536 7828 227588 7880
rect 162492 7760 162544 7812
rect 378876 7760 378928 7812
rect 162032 7692 162084 7744
rect 390652 7692 390704 7744
rect 169760 7624 169812 7676
rect 482836 7624 482888 7676
rect 24216 7556 24268 7608
rect 134156 7556 134208 7608
rect 173900 7556 173952 7608
rect 545488 7556 545540 7608
rect 576124 6808 576176 6860
rect 580172 6808 580224 6860
rect 153844 6400 153896 6452
rect 272432 6400 272484 6452
rect 158628 6332 158680 6384
rect 336280 6332 336332 6384
rect 165436 6264 165488 6316
rect 411904 6264 411956 6316
rect 165528 6196 165580 6248
rect 414296 6196 414348 6248
rect 87972 6128 88024 6180
rect 138020 6128 138072 6180
rect 143540 6128 143592 6180
rect 155408 6128 155460 6180
rect 173808 6128 173860 6180
rect 525432 6128 525484 6180
rect 154120 5040 154172 5092
rect 273628 5040 273680 5092
rect 162584 4972 162636 5024
rect 382372 4972 382424 5024
rect 180156 4904 180208 4956
rect 429660 4904 429712 4956
rect 138848 4836 138900 4888
rect 142252 4836 142304 4888
rect 170312 4836 170364 4888
rect 486424 4836 486476 4888
rect 175188 4768 175240 4820
rect 541992 4768 542044 4820
rect 572 4088 624 4140
rect 7564 4088 7616 4140
rect 73804 4088 73856 4140
rect 75184 4088 75236 4140
rect 103336 4088 103388 4140
rect 104164 4088 104216 4140
rect 146944 4088 146996 4140
rect 147404 4088 147456 4140
rect 149704 4088 149756 4140
rect 151820 4088 151872 4140
rect 196624 4088 196676 4140
rect 203892 4088 203944 4140
rect 304264 4088 304316 4140
rect 309048 4088 309100 4140
rect 450544 4088 450596 4140
rect 451004 4088 451056 4140
rect 6460 4020 6512 4072
rect 7656 4020 7708 4072
rect 180340 4020 180392 4072
rect 186136 4020 186188 4072
rect 189816 4020 189868 4072
rect 193220 4020 193272 4072
rect 193864 4020 193916 4072
rect 196808 4020 196860 4072
rect 203708 4020 203760 4072
rect 223948 4020 224000 4072
rect 224224 4020 224276 4072
rect 240508 4020 240560 4072
rect 164884 3952 164936 4004
rect 168380 3952 168432 4004
rect 181444 3952 181496 4004
rect 226340 3952 226392 4004
rect 276020 3952 276072 4004
rect 276756 3952 276808 4004
rect 299572 3952 299624 4004
rect 300768 3952 300820 4004
rect 147128 3884 147180 3936
rect 150624 3884 150676 3936
rect 155868 3884 155920 3936
rect 306748 3884 306800 3936
rect 311164 3884 311216 3936
rect 312636 3884 312688 3936
rect 44272 3816 44324 3868
rect 46204 3816 46256 3868
rect 69112 3816 69164 3868
rect 65524 3748 65576 3800
rect 19432 3612 19484 3664
rect 21364 3612 21416 3664
rect 43076 3612 43128 3664
rect 44824 3612 44876 3664
rect 51356 3612 51408 3664
rect 54484 3612 54536 3664
rect 70308 3612 70360 3664
rect 72424 3612 72476 3664
rect 122288 3816 122340 3868
rect 127624 3816 127676 3868
rect 147220 3816 147272 3868
rect 163688 3816 163740 3868
rect 178684 3816 178736 3868
rect 401324 3816 401376 3868
rect 111616 3748 111668 3800
rect 131764 3748 131816 3800
rect 148324 3748 148376 3800
rect 164884 3748 164936 3800
rect 170404 3748 170456 3800
rect 174268 3748 174320 3800
rect 183468 3748 183520 3800
rect 200304 3748 200356 3800
rect 200764 3748 200816 3800
rect 210976 3748 211028 3800
rect 220084 3748 220136 3800
rect 447416 3748 447468 3800
rect 453396 3748 453448 3800
rect 497096 3748 497148 3800
rect 129832 3680 129884 3732
rect 131028 3680 131080 3732
rect 143540 3680 143592 3732
rect 148416 3680 148468 3732
rect 170772 3680 170824 3732
rect 179236 3680 179288 3732
rect 137284 3612 137336 3664
rect 147036 3612 147088 3664
rect 149520 3612 149572 3664
rect 7656 3544 7708 3596
rect 129924 3544 129976 3596
rect 130936 3544 130988 3596
rect 4068 3476 4120 3528
rect 4804 3476 4856 3528
rect 5264 3476 5316 3528
rect 8760 3408 8812 3460
rect 10324 3408 10376 3460
rect 17040 3408 17092 3460
rect 18604 3408 18656 3460
rect 20628 3408 20680 3460
rect 27620 3340 27672 3392
rect 28540 3340 28592 3392
rect 33600 3340 33652 3392
rect 35164 3340 35216 3392
rect 41880 3340 41932 3392
rect 43444 3340 43496 3392
rect 52460 3340 52512 3392
rect 53380 3340 53432 3392
rect 60740 3340 60792 3392
rect 61660 3340 61712 3392
rect 85580 3340 85632 3392
rect 86500 3340 86552 3392
rect 91560 3340 91612 3392
rect 93124 3340 93176 3392
rect 93860 3340 93912 3392
rect 94780 3340 94832 3392
rect 101036 3340 101088 3392
rect 102784 3340 102836 3392
rect 109316 3340 109368 3392
rect 111156 3340 111208 3392
rect 119896 3340 119948 3392
rect 120724 3340 120776 3392
rect 15936 3272 15988 3324
rect 17224 3272 17276 3324
rect 83280 3272 83332 3324
rect 84844 3272 84896 3324
rect 123484 3272 123536 3324
rect 124864 3272 124916 3324
rect 126980 3476 127032 3528
rect 128360 3476 128412 3528
rect 129372 3476 129424 3528
rect 130016 3476 130068 3528
rect 137652 3476 137704 3528
rect 138664 3476 138716 3528
rect 128176 3408 128228 3460
rect 130384 3408 130436 3460
rect 131856 3340 131908 3392
rect 147312 3544 147364 3596
rect 171968 3612 172020 3664
rect 180248 3680 180300 3732
rect 454500 3680 454552 3732
rect 143448 3476 143500 3528
rect 144736 3476 144788 3528
rect 162492 3544 162544 3596
rect 171876 3544 171928 3596
rect 177856 3544 177908 3596
rect 182088 3612 182140 3664
rect 480536 3612 480588 3664
rect 486516 3612 486568 3664
rect 518348 3612 518400 3664
rect 487620 3544 487672 3596
rect 489920 3544 489972 3596
rect 490748 3544 490800 3596
rect 504364 3544 504416 3596
rect 505376 3544 505428 3596
rect 506480 3544 506532 3596
rect 507308 3544 507360 3596
rect 520924 3544 520976 3596
rect 524236 3544 524288 3596
rect 525064 3544 525116 3596
rect 533712 3544 533764 3596
rect 151084 3476 151136 3528
rect 171784 3476 171836 3528
rect 173164 3476 173216 3528
rect 179328 3476 179380 3528
rect 531320 3476 531372 3528
rect 538864 3476 538916 3528
rect 539600 3476 539652 3528
rect 545764 3476 545816 3528
rect 551468 3476 551520 3528
rect 552756 3476 552808 3528
rect 572720 3544 572772 3596
rect 574744 3544 574796 3596
rect 576308 3544 576360 3596
rect 567844 3476 567896 3528
rect 569132 3476 569184 3528
rect 131948 3272 132000 3324
rect 132960 3272 133012 3324
rect 141424 3272 141476 3324
rect 147404 3272 147456 3324
rect 156604 3340 156656 3392
rect 157800 3340 157852 3392
rect 175464 3408 175516 3460
rect 176660 3340 176712 3392
rect 180340 3340 180392 3392
rect 581000 3408 581052 3460
rect 185584 3340 185636 3392
rect 189724 3340 189776 3392
rect 217324 3340 217376 3392
rect 218060 3340 218112 3392
rect 229744 3340 229796 3392
rect 231032 3340 231084 3392
rect 324412 3340 324464 3392
rect 325608 3340 325660 3392
rect 332600 3340 332652 3392
rect 333888 3340 333940 3392
rect 349252 3340 349304 3392
rect 350448 3340 350500 3392
rect 357532 3340 357584 3392
rect 358728 3340 358780 3392
rect 364984 3340 365036 3392
rect 367008 3340 367060 3392
rect 374092 3340 374144 3392
rect 375288 3340 375340 3392
rect 382280 3340 382332 3392
rect 383568 3340 383620 3392
rect 390560 3340 390612 3392
rect 391848 3340 391900 3392
rect 398932 3340 398984 3392
rect 400128 3340 400180 3392
rect 400956 3340 401008 3392
rect 402520 3340 402572 3392
rect 407212 3340 407264 3392
rect 408408 3340 408460 3392
rect 414664 3340 414716 3392
rect 416688 3340 416740 3392
rect 418804 3340 418856 3392
rect 420184 3340 420236 3392
rect 423680 3340 423732 3392
rect 424968 3340 425020 3392
rect 432604 3340 432656 3392
rect 434444 3340 434496 3392
rect 440240 3340 440292 3392
rect 441528 3340 441580 3392
rect 448612 3340 448664 3392
rect 449808 3340 449860 3392
rect 456800 3340 456852 3392
rect 458088 3340 458140 3392
rect 464344 3340 464396 3392
rect 466276 3340 466328 3392
rect 468484 3340 468536 3392
rect 469864 3340 469916 3392
rect 472624 3340 472676 3392
rect 473452 3340 473504 3392
rect 315304 3272 315356 3324
rect 317328 3272 317380 3324
rect 431960 3272 432012 3324
rect 433248 3272 433300 3324
rect 1676 3204 1728 3256
rect 8944 3204 8996 3256
rect 136456 3204 136508 3256
rect 140044 3204 140096 3256
rect 18236 3136 18288 3188
rect 22744 3136 22796 3188
rect 30104 3136 30156 3188
rect 31024 3136 31076 3188
rect 38384 3136 38436 3188
rect 39304 3136 39356 3188
rect 125876 3136 125928 3188
rect 131120 3136 131172 3188
rect 181536 3136 181588 3188
rect 184940 3136 184992 3188
rect 324964 3136 325016 3188
rect 326804 3136 326856 3188
rect 336004 3136 336056 3188
rect 342168 3136 342220 3188
rect 382924 3136 382976 3188
rect 384764 3136 384816 3188
rect 451004 3136 451056 3188
rect 452108 3136 452160 3188
rect 511356 3136 511408 3188
rect 514760 3136 514812 3188
rect 56048 3000 56100 3052
rect 58624 3000 58676 3052
rect 118792 3000 118844 3052
rect 122104 3000 122156 3052
rect 297364 3000 297416 3052
rect 298468 3000 298520 3052
rect 514024 3000 514076 3052
rect 515956 3000 516008 3052
rect 563704 3000 563756 3052
rect 565636 3000 565688 3052
rect 571984 3000 572036 3052
rect 573916 3000 573968 3052
rect 12348 2932 12400 2984
rect 14464 2932 14516 2984
rect 149796 2864 149848 2916
rect 154212 2864 154264 2916
rect 454684 2864 454736 2916
rect 455696 2864 455748 2916
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40052 703582 40356 703610
rect 8128 700466 8156 703520
rect 8116 700460 8168 700466
rect 8116 700402 8168 700408
rect 24320 699718 24348 703520
rect 24308 699712 24360 699718
rect 24308 699654 24360 699660
rect 25504 699712 25556 699718
rect 25504 699654 25556 699660
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3330 671256 3386 671265
rect 3330 671191 3386 671200
rect 3344 670818 3372 671191
rect 3332 670812 3384 670818
rect 3332 670754 3384 670760
rect 3330 580000 3386 580009
rect 3330 579935 3386 579944
rect 3344 579698 3372 579935
rect 3332 579692 3384 579698
rect 3332 579634 3384 579640
rect 3238 566944 3294 566953
rect 3238 566879 3294 566888
rect 3252 565894 3280 566879
rect 3240 565888 3292 565894
rect 3240 565830 3292 565836
rect 3330 553888 3386 553897
rect 3330 553823 3386 553832
rect 3344 553450 3372 553823
rect 3332 553444 3384 553450
rect 3332 553386 3384 553392
rect 2778 527912 2834 527921
rect 2778 527847 2834 527856
rect 2792 527202 2820 527847
rect 2780 527196 2832 527202
rect 2780 527138 2832 527144
rect 3054 501800 3110 501809
rect 3054 501735 3110 501744
rect 3068 501022 3096 501735
rect 3056 501016 3108 501022
rect 3056 500958 3108 500964
rect 3054 475688 3110 475697
rect 3054 475623 3110 475632
rect 3068 474774 3096 475623
rect 3056 474768 3108 474774
rect 3056 474710 3108 474716
rect 3146 449576 3202 449585
rect 3146 449511 3202 449520
rect 3160 448594 3188 449511
rect 3148 448588 3200 448594
rect 3148 448530 3200 448536
rect 2870 410544 2926 410553
rect 2870 410479 2926 410488
rect 2884 409902 2912 410479
rect 2872 409896 2924 409902
rect 2872 409838 2924 409844
rect 3146 358456 3202 358465
rect 3146 358391 3202 358400
rect 3160 357474 3188 358391
rect 3148 357468 3200 357474
rect 3148 357410 3200 357416
rect 3330 345400 3386 345409
rect 3330 345335 3386 345344
rect 3344 345098 3372 345335
rect 3332 345092 3384 345098
rect 3332 345034 3384 345040
rect 3330 319288 3386 319297
rect 3330 319223 3386 319232
rect 3344 318850 3372 319223
rect 3332 318844 3384 318850
rect 3332 318786 3384 318792
rect 3054 267200 3110 267209
rect 3054 267135 3110 267144
rect 3068 266422 3096 267135
rect 3056 266416 3108 266422
rect 3056 266358 3108 266364
rect 3436 265674 3464 684247
rect 3514 658200 3570 658209
rect 3514 658135 3516 658144
rect 3568 658135 3570 658144
rect 7564 658164 7616 658170
rect 3516 658106 3568 658112
rect 7564 658106 7616 658112
rect 3516 632120 3568 632126
rect 3514 632088 3516 632097
rect 3568 632088 3570 632097
rect 3514 632023 3570 632032
rect 3514 619168 3570 619177
rect 3514 619103 3570 619112
rect 3528 618322 3556 619103
rect 3516 618316 3568 618322
rect 3516 618258 3568 618264
rect 3514 606112 3570 606121
rect 3514 606047 3570 606056
rect 3528 605878 3556 606047
rect 3516 605872 3568 605878
rect 3516 605814 3568 605820
rect 4804 527196 4856 527202
rect 4804 527138 4856 527144
rect 3514 514856 3570 514865
rect 3514 514791 3516 514800
rect 3568 514791 3570 514800
rect 3516 514762 3568 514768
rect 3514 462632 3570 462641
rect 3514 462567 3570 462576
rect 3528 462398 3556 462567
rect 3516 462392 3568 462398
rect 3516 462334 3568 462340
rect 3514 423600 3570 423609
rect 3514 423535 3570 423544
rect 3528 422346 3556 423535
rect 3516 422340 3568 422346
rect 3516 422282 3568 422288
rect 3516 397520 3568 397526
rect 3514 397488 3516 397497
rect 3568 397488 3570 397497
rect 3514 397423 3570 397432
rect 3514 371376 3570 371385
rect 3514 371311 3516 371320
rect 3568 371311 3570 371320
rect 3516 371282 3568 371288
rect 3514 306232 3570 306241
rect 3514 306167 3570 306176
rect 3528 305046 3556 306167
rect 3516 305040 3568 305046
rect 3516 304982 3568 304988
rect 3514 293176 3570 293185
rect 3514 293111 3570 293120
rect 3528 292602 3556 293111
rect 3516 292596 3568 292602
rect 3516 292538 3568 292544
rect 3424 265668 3476 265674
rect 3424 265610 3476 265616
rect 4816 264246 4844 527138
rect 7576 273970 7604 658106
rect 10324 514820 10376 514826
rect 10324 514762 10376 514768
rect 8944 371340 8996 371346
rect 8944 371282 8996 371288
rect 7564 273964 7616 273970
rect 7564 273906 7616 273912
rect 8956 269890 8984 371282
rect 10336 275330 10364 514762
rect 13084 409896 13136 409902
rect 13084 409838 13136 409844
rect 13096 286346 13124 409838
rect 13084 286340 13136 286346
rect 13084 286282 13136 286288
rect 25516 284986 25544 699654
rect 25504 284980 25556 284986
rect 25504 284922 25556 284928
rect 40052 276690 40080 703582
rect 40328 703474 40356 703582
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218072 703582 218836 703610
rect 40512 703474 40540 703520
rect 40328 703446 40540 703474
rect 72988 700602 73016 703520
rect 89180 700670 89208 703520
rect 89168 700664 89220 700670
rect 89168 700606 89220 700612
rect 72976 700596 73028 700602
rect 72976 700538 73028 700544
rect 105464 699718 105492 703520
rect 137848 699718 137876 703520
rect 154132 702434 154160 703520
rect 170324 702434 170352 703520
rect 153304 702406 154160 702434
rect 169772 702406 170352 702434
rect 153200 700392 153252 700398
rect 153200 700334 153252 700340
rect 149704 700324 149756 700330
rect 149704 700266 149756 700272
rect 105452 699712 105504 699718
rect 105452 699654 105504 699660
rect 106924 699712 106976 699718
rect 106924 699654 106976 699660
rect 137836 699712 137888 699718
rect 137836 699654 137888 699660
rect 140044 699712 140096 699718
rect 140044 699654 140096 699660
rect 40040 276684 40092 276690
rect 40040 276626 40092 276632
rect 10324 275324 10376 275330
rect 10324 275266 10376 275272
rect 8944 269884 8996 269890
rect 8944 269826 8996 269832
rect 106936 268462 106964 699654
rect 138020 430636 138072 430642
rect 138020 430578 138072 430584
rect 135536 324352 135588 324358
rect 135536 324294 135588 324300
rect 134524 271924 134576 271930
rect 134524 271866 134576 271872
rect 106924 268456 106976 268462
rect 106924 268398 106976 268404
rect 114284 264988 114336 264994
rect 114284 264930 114336 264936
rect 4804 264240 4856 264246
rect 4804 264182 4856 264188
rect 114192 263900 114244 263906
rect 114192 263842 114244 263848
rect 112444 263084 112496 263090
rect 112444 263026 112496 263032
rect 3424 262948 3476 262954
rect 3424 262890 3476 262896
rect 2780 215280 2832 215286
rect 2780 215222 2832 215228
rect 2792 214985 2820 215222
rect 2778 214976 2834 214985
rect 2778 214911 2834 214920
rect 3436 201929 3464 262890
rect 111064 262812 111116 262818
rect 111064 262754 111116 262760
rect 3516 262472 3568 262478
rect 3516 262414 3568 262420
rect 3528 254153 3556 262414
rect 4804 261248 4856 261254
rect 4804 261190 4856 261196
rect 3514 254144 3570 254153
rect 3514 254079 3570 254088
rect 3516 241120 3568 241126
rect 3514 241088 3516 241097
rect 3568 241088 3570 241097
rect 3514 241023 3570 241032
rect 4816 215286 4844 261190
rect 7564 260364 7616 260370
rect 7564 260306 7616 260312
rect 7576 241126 7604 260306
rect 7564 241120 7616 241126
rect 7564 241062 7616 241068
rect 4804 215280 4856 215286
rect 4804 215222 4856 215228
rect 3422 201920 3478 201929
rect 3422 201855 3478 201864
rect 109958 200696 110014 200705
rect 109958 200631 110014 200640
rect 107198 200288 107254 200297
rect 107198 200223 107254 200232
rect 105634 200152 105690 200161
rect 105634 200087 105690 200096
rect 103242 199880 103298 199889
rect 103242 199815 103298 199824
rect 100668 194404 100720 194410
rect 100668 194346 100720 194352
rect 100576 190188 100628 190194
rect 100576 190130 100628 190136
rect 3424 189032 3476 189038
rect 3424 188974 3476 188980
rect 3436 188873 3464 188974
rect 3422 188864 3478 188873
rect 3422 188799 3478 188808
rect 3422 162888 3478 162897
rect 3422 162823 3478 162832
rect 3436 151814 3464 162823
rect 3436 151786 3556 151814
rect 3422 149832 3478 149841
rect 3422 149767 3478 149776
rect 3436 149122 3464 149767
rect 3424 149116 3476 149122
rect 3424 149058 3476 149064
rect 3528 146266 3556 151786
rect 100208 148844 100260 148850
rect 100208 148786 100260 148792
rect 100116 148368 100168 148374
rect 100116 148310 100168 148316
rect 3516 146260 3568 146266
rect 3516 146202 3568 146208
rect 3424 142316 3476 142322
rect 3424 142258 3476 142264
rect 3148 111784 3200 111790
rect 3148 111726 3200 111732
rect 3160 110673 3188 111726
rect 3146 110664 3202 110673
rect 3146 110599 3202 110608
rect 2780 77988 2832 77994
rect 2780 77930 2832 77936
rect 2792 16574 2820 77930
rect 2792 16546 2912 16574
rect 572 4140 624 4146
rect 572 4082 624 4088
rect 584 480 612 4082
rect 1676 3256 1728 3262
rect 1676 3198 1728 3204
rect 1688 480 1716 3198
rect 2884 480 2912 16546
rect 3436 6497 3464 142258
rect 8944 141024 8996 141030
rect 8944 140966 8996 140972
rect 3516 137964 3568 137970
rect 3516 137906 3568 137912
rect 3528 136785 3556 137906
rect 3514 136776 3570 136785
rect 3514 136711 3570 136720
rect 4802 76528 4858 76537
rect 4802 76463 4858 76472
rect 3516 71664 3568 71670
rect 3514 71632 3516 71641
rect 3568 71632 3570 71641
rect 3514 71567 3570 71576
rect 3516 59356 3568 59362
rect 3516 59298 3568 59304
rect 3528 58585 3556 59298
rect 3514 58576 3570 58585
rect 3514 58511 3570 58520
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 4816 3534 4844 76463
rect 7562 75168 7618 75177
rect 7562 75103 7618 75112
rect 7576 4146 7604 75103
rect 8956 71670 8984 140966
rect 31022 139496 31078 139505
rect 31022 139431 31078 139440
rect 31036 111790 31064 139431
rect 31024 111784 31076 111790
rect 31024 111726 31076 111732
rect 71780 80708 71832 80714
rect 71780 80650 71832 80656
rect 60740 78328 60792 78334
rect 60740 78270 60792 78276
rect 57980 78260 58032 78266
rect 57980 78202 58032 78208
rect 46940 78192 46992 78198
rect 46940 78134 46992 78140
rect 34520 78124 34572 78130
rect 34520 78066 34572 78072
rect 20720 78056 20772 78062
rect 20720 77998 20772 78004
rect 14464 72480 14516 72486
rect 11058 72448 11114 72457
rect 14464 72422 14516 72428
rect 11058 72383 11114 72392
rect 8944 71664 8996 71670
rect 8944 71606 8996 71612
rect 8942 68232 8998 68241
rect 8942 68167 8998 68176
rect 7654 65512 7710 65521
rect 7654 65447 7710 65456
rect 7564 4140 7616 4146
rect 7564 4082 7616 4088
rect 7668 4078 7696 65447
rect 6460 4072 6512 4078
rect 6460 4014 6512 4020
rect 7656 4072 7708 4078
rect 7656 4014 7708 4020
rect 4068 3528 4120 3534
rect 4068 3470 4120 3476
rect 4804 3528 4856 3534
rect 4804 3470 4856 3476
rect 5264 3528 5316 3534
rect 5264 3470 5316 3476
rect 4080 480 4108 3470
rect 5276 480 5304 3470
rect 6472 480 6500 4014
rect 7656 3596 7708 3602
rect 7656 3538 7708 3544
rect 7668 480 7696 3538
rect 8760 3460 8812 3466
rect 8760 3402 8812 3408
rect 8772 480 8800 3402
rect 8956 3262 8984 68167
rect 10324 62824 10376 62830
rect 10324 62766 10376 62772
rect 9680 53100 9732 53106
rect 9680 53042 9732 53048
rect 8944 3256 8996 3262
rect 8944 3198 8996 3204
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9692 354 9720 53042
rect 10336 3466 10364 62766
rect 11072 16574 11100 72383
rect 12440 55888 12492 55894
rect 12440 55830 12492 55836
rect 12452 16574 12480 55830
rect 13820 37936 13872 37942
rect 13820 37878 13872 37884
rect 13832 16574 13860 37878
rect 11072 16546 11192 16574
rect 12452 16546 13584 16574
rect 13832 16546 14320 16574
rect 10324 3460 10376 3466
rect 10324 3402 10376 3408
rect 11164 480 11192 16546
rect 12348 2984 12400 2990
rect 12348 2926 12400 2932
rect 12360 480 12388 2926
rect 13556 480 13584 16546
rect 9926 354 10038 480
rect 9692 326 10038 354
rect 9926 -960 10038 326
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14292 354 14320 16546
rect 14476 2990 14504 72422
rect 18604 69760 18656 69766
rect 18604 69702 18656 69708
rect 17222 33824 17278 33833
rect 17222 33759 17278 33768
rect 17040 3460 17092 3466
rect 17040 3402 17092 3408
rect 15936 3324 15988 3330
rect 15936 3266 15988 3272
rect 14464 2984 14516 2990
rect 14464 2926 14516 2932
rect 15948 480 15976 3266
rect 17052 480 17080 3402
rect 17236 3330 17264 33759
rect 18616 3466 18644 69702
rect 20732 16574 20760 77998
rect 27620 75200 27672 75206
rect 27620 75142 27672 75148
rect 21362 73808 21418 73817
rect 21362 73743 21418 73752
rect 20732 16546 21312 16574
rect 19432 3664 19484 3670
rect 19432 3606 19484 3612
rect 18604 3460 18656 3466
rect 18604 3402 18656 3408
rect 17224 3324 17276 3330
rect 17224 3266 17276 3272
rect 18236 3188 18288 3194
rect 18236 3130 18288 3136
rect 18248 480 18276 3130
rect 19444 480 19472 3606
rect 21284 3482 21312 16546
rect 21376 3670 21404 73743
rect 24858 66872 24914 66881
rect 24858 66807 24914 66816
rect 22744 60036 22796 60042
rect 22744 59978 22796 59984
rect 22100 57248 22152 57254
rect 22100 57190 22152 57196
rect 22112 16574 22140 57190
rect 22112 16546 22600 16574
rect 21364 3664 21416 3670
rect 21364 3606 21416 3612
rect 20628 3460 20680 3466
rect 21284 3454 21864 3482
rect 20628 3402 20680 3408
rect 20640 480 20668 3402
rect 21836 480 21864 3454
rect 14710 354 14822 480
rect 14292 326 14822 354
rect 14710 -960 14822 326
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22572 354 22600 16546
rect 22756 3194 22784 59978
rect 24872 16574 24900 66807
rect 26240 61464 26292 61470
rect 26240 61406 26292 61412
rect 24872 16546 25360 16574
rect 24216 7608 24268 7614
rect 24216 7550 24268 7556
rect 22744 3188 22796 3194
rect 22744 3130 22796 3136
rect 24228 480 24256 7550
rect 25332 480 25360 16546
rect 22990 354 23102 480
rect 22572 326 23102 354
rect 22990 -960 23102 326
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26252 354 26280 61406
rect 27632 3398 27660 75142
rect 31024 71120 31076 71126
rect 31024 71062 31076 71068
rect 27710 51776 27766 51785
rect 27710 51711 27766 51720
rect 27620 3392 27672 3398
rect 27620 3334 27672 3340
rect 27724 480 27752 51711
rect 30380 50380 30432 50386
rect 30380 50322 30432 50328
rect 30392 16574 30420 50322
rect 30392 16546 30880 16574
rect 28540 3392 28592 3398
rect 28540 3334 28592 3340
rect 26486 354 26598 480
rect 26252 326 26598 354
rect 26486 -960 26598 326
rect 27682 -960 27794 480
rect 28552 354 28580 3334
rect 30104 3188 30156 3194
rect 30104 3130 30156 3136
rect 30116 480 30144 3130
rect 28878 354 28990 480
rect 28552 326 28990 354
rect 28878 -960 28990 326
rect 30074 -960 30186 480
rect 30852 354 30880 16546
rect 31036 3194 31064 71062
rect 31760 71052 31812 71058
rect 31760 70994 31812 71000
rect 31772 16574 31800 70994
rect 31772 16546 31984 16574
rect 31024 3188 31076 3194
rect 31024 3130 31076 3136
rect 31270 354 31382 480
rect 30852 326 31382 354
rect 31956 354 31984 16546
rect 33600 3392 33652 3398
rect 33600 3334 33652 3340
rect 33612 480 33640 3334
rect 32374 354 32486 480
rect 31956 326 32486 354
rect 31270 -960 31382 326
rect 32374 -960 32486 326
rect 33570 -960 33682 480
rect 34532 354 34560 78066
rect 43444 72616 43496 72622
rect 43444 72558 43496 72564
rect 35164 66904 35216 66910
rect 35164 66846 35216 66852
rect 35176 3398 35204 66846
rect 35900 64184 35952 64190
rect 35900 64126 35952 64132
rect 35912 6914 35940 64126
rect 39302 48920 39358 48929
rect 39302 48855 39358 48864
rect 38660 35216 38712 35222
rect 38660 35158 38712 35164
rect 35992 26920 36044 26926
rect 35992 26862 36044 26868
rect 36004 16574 36032 26862
rect 38672 16574 38700 35158
rect 36004 16546 36768 16574
rect 38672 16546 39160 16574
rect 35912 6886 36032 6914
rect 35164 3392 35216 3398
rect 35164 3334 35216 3340
rect 36004 480 36032 6886
rect 34766 354 34878 480
rect 34532 326 34878 354
rect 34766 -960 34878 326
rect 35962 -960 36074 480
rect 36740 354 36768 16546
rect 38384 3188 38436 3194
rect 38384 3130 38436 3136
rect 38396 480 38424 3130
rect 37158 354 37270 480
rect 36740 326 37270 354
rect 37158 -960 37270 326
rect 38354 -960 38466 480
rect 39132 354 39160 16546
rect 39316 3194 39344 48855
rect 40040 24132 40092 24138
rect 40040 24074 40092 24080
rect 40052 16574 40080 24074
rect 40052 16546 40264 16574
rect 39304 3188 39356 3194
rect 39304 3130 39356 3136
rect 39550 354 39662 480
rect 39132 326 39662 354
rect 40236 354 40264 16546
rect 43076 3664 43128 3670
rect 43076 3606 43128 3612
rect 41880 3392 41932 3398
rect 41880 3334 41932 3340
rect 41892 480 41920 3334
rect 43088 480 43116 3606
rect 43456 3398 43484 72558
rect 45560 69692 45612 69698
rect 45560 69634 45612 69640
rect 44824 61396 44876 61402
rect 44824 61338 44876 61344
rect 44178 47560 44234 47569
rect 44178 47495 44234 47504
rect 44192 16574 44220 47495
rect 44192 16546 44772 16574
rect 44272 3868 44324 3874
rect 44272 3810 44324 3816
rect 43444 3392 43496 3398
rect 43444 3334 43496 3340
rect 44284 480 44312 3810
rect 44744 490 44772 16546
rect 44836 3670 44864 61338
rect 45572 16574 45600 69634
rect 46202 64152 46258 64161
rect 46202 64087 46258 64096
rect 45572 16546 46152 16574
rect 44824 3664 44876 3670
rect 44824 3606 44876 3612
rect 46124 3482 46152 16546
rect 46216 3874 46244 64087
rect 46952 16574 46980 78134
rect 52460 76560 52512 76566
rect 52460 76502 52512 76508
rect 48320 68332 48372 68338
rect 48320 68274 48372 68280
rect 48332 16574 48360 68274
rect 49698 46200 49754 46209
rect 49698 46135 49754 46144
rect 49712 16574 49740 46135
rect 46952 16546 47440 16574
rect 48332 16546 48544 16574
rect 49712 16546 50200 16574
rect 46204 3868 46256 3874
rect 46204 3810 46256 3816
rect 46124 3454 46704 3482
rect 40654 354 40766 480
rect 40236 326 40766 354
rect 39550 -960 39662 326
rect 40654 -960 40766 326
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 44744 462 45140 490
rect 46676 480 46704 3454
rect 45112 354 45140 462
rect 45438 354 45550 480
rect 45112 326 45550 354
rect 45438 -960 45550 326
rect 46634 -960 46746 480
rect 47412 354 47440 16546
rect 47830 354 47942 480
rect 47412 326 47942 354
rect 48516 354 48544 16546
rect 50172 480 50200 16546
rect 51356 3664 51408 3670
rect 51356 3606 51408 3612
rect 51368 480 51396 3606
rect 52472 3398 52500 76502
rect 54482 73944 54538 73953
rect 54482 73879 54538 73888
rect 53840 71188 53892 71194
rect 53840 71130 53892 71136
rect 52552 28280 52604 28286
rect 52552 28222 52604 28228
rect 52460 3392 52512 3398
rect 52460 3334 52512 3340
rect 52564 480 52592 28222
rect 53852 16574 53880 71130
rect 53852 16546 54432 16574
rect 54404 3482 54432 16546
rect 54496 3670 54524 73879
rect 56598 54496 56654 54505
rect 56598 54431 56654 54440
rect 56612 16574 56640 54431
rect 57992 16574 58020 78202
rect 59360 76628 59412 76634
rect 59360 76570 59412 76576
rect 58624 65544 58676 65550
rect 58624 65486 58676 65492
rect 56612 16546 56824 16574
rect 57992 16546 58480 16574
rect 54484 3664 54536 3670
rect 54484 3606 54536 3612
rect 54404 3454 54984 3482
rect 53380 3392 53432 3398
rect 53380 3334 53432 3340
rect 48934 354 49046 480
rect 48516 326 49046 354
rect 47830 -960 47942 326
rect 48934 -960 49046 326
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53392 354 53420 3334
rect 54956 480 54984 3454
rect 56048 3052 56100 3058
rect 56048 2994 56100 3000
rect 56060 480 56088 2994
rect 53718 354 53830 480
rect 53392 326 53830 354
rect 53718 -960 53830 326
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 56796 354 56824 16546
rect 58452 480 58480 16546
rect 58636 3058 58664 65486
rect 58624 3052 58676 3058
rect 58624 2994 58676 3000
rect 57214 354 57326 480
rect 56796 326 57326 354
rect 57214 -960 57326 326
rect 58410 -960 58522 480
rect 59372 354 59400 76570
rect 60752 3398 60780 78270
rect 66260 76696 66312 76702
rect 66260 76638 66312 76644
rect 62120 69896 62172 69902
rect 62120 69838 62172 69844
rect 60832 58676 60884 58682
rect 60832 58618 60884 58624
rect 60740 3392 60792 3398
rect 60740 3334 60792 3340
rect 60844 480 60872 58618
rect 62132 16574 62160 69838
rect 63500 43444 63552 43450
rect 63500 43386 63552 43392
rect 63512 16574 63540 43386
rect 66272 16574 66300 76638
rect 67640 72548 67692 72554
rect 67640 72490 67692 72496
rect 62132 16546 63264 16574
rect 63512 16546 64368 16574
rect 66272 16546 66760 16574
rect 61660 3392 61712 3398
rect 61660 3334 61712 3340
rect 59606 354 59718 480
rect 59372 326 59718 354
rect 59606 -960 59718 326
rect 60802 -960 60914 480
rect 61672 354 61700 3334
rect 63236 480 63264 16546
rect 64340 480 64368 16546
rect 65524 3800 65576 3806
rect 65524 3742 65576 3748
rect 65536 480 65564 3742
rect 66732 480 66760 16546
rect 61998 354 62110 480
rect 61672 326 62110 354
rect 61998 -960 62110 326
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67652 354 67680 72490
rect 70400 42084 70452 42090
rect 70400 42026 70452 42032
rect 70412 16574 70440 42026
rect 71792 16574 71820 80650
rect 75920 78532 75972 78538
rect 75920 78474 75972 78480
rect 72424 66972 72476 66978
rect 72424 66914 72476 66920
rect 70412 16546 71544 16574
rect 71792 16546 72372 16574
rect 69112 3868 69164 3874
rect 69112 3810 69164 3816
rect 69124 480 69152 3810
rect 70308 3664 70360 3670
rect 70308 3606 70360 3612
rect 70320 480 70348 3606
rect 71516 480 71544 16546
rect 72344 3482 72372 16546
rect 72436 3670 72464 66914
rect 75182 62792 75238 62801
rect 75182 62727 75238 62736
rect 74540 40724 74592 40730
rect 74540 40666 74592 40672
rect 74552 16574 74580 40666
rect 74552 16546 75040 16574
rect 73804 4140 73856 4146
rect 73804 4082 73856 4088
rect 72424 3664 72476 3670
rect 72424 3606 72476 3612
rect 72344 3454 72648 3482
rect 72620 480 72648 3454
rect 73816 480 73844 4082
rect 75012 480 75040 16546
rect 75196 4146 75224 62727
rect 75184 4140 75236 4146
rect 75184 4082 75236 4088
rect 67886 354 67998 480
rect 67652 326 67998 354
rect 67886 -960 67998 326
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 75932 354 75960 78474
rect 96620 75336 96672 75342
rect 96620 75278 96672 75284
rect 81440 75268 81492 75274
rect 81440 75210 81492 75216
rect 78680 73840 78732 73846
rect 78680 73782 78732 73788
rect 77298 57216 77354 57225
rect 77298 57151 77354 57160
rect 77312 6914 77340 57151
rect 77392 39364 77444 39370
rect 77392 39306 77444 39312
rect 77404 16574 77432 39306
rect 78692 16574 78720 73782
rect 80058 67008 80114 67017
rect 80058 66943 80114 66952
rect 80072 16574 80100 66943
rect 81452 16574 81480 75210
rect 85580 72684 85632 72690
rect 85580 72626 85632 72632
rect 84844 64252 84896 64258
rect 84844 64194 84896 64200
rect 84198 59936 84254 59945
rect 84198 59871 84254 59880
rect 77404 16546 78168 16574
rect 78692 16546 79272 16574
rect 80072 16546 80928 16574
rect 81452 16546 81664 16574
rect 77312 6886 77432 6914
rect 77404 480 77432 6886
rect 76166 354 76278 480
rect 75932 326 76278 354
rect 76166 -960 76278 326
rect 77362 -960 77474 480
rect 78140 354 78168 16546
rect 78558 354 78670 480
rect 78140 326 78670 354
rect 79244 354 79272 16546
rect 80900 480 80928 16546
rect 79662 354 79774 480
rect 79244 326 79774 354
rect 78558 -960 78670 326
rect 79662 -960 79774 326
rect 80858 -960 80970 480
rect 81636 354 81664 16546
rect 83280 3324 83332 3330
rect 83280 3266 83332 3272
rect 83292 480 83320 3266
rect 82054 354 82166 480
rect 81636 326 82166 354
rect 82054 -960 82166 326
rect 83250 -960 83362 480
rect 84212 354 84240 59871
rect 84856 3330 84884 64194
rect 85592 3398 85620 72626
rect 85672 69828 85724 69834
rect 85672 69770 85724 69776
rect 85580 3392 85632 3398
rect 85580 3334 85632 3340
rect 84844 3324 84896 3330
rect 84844 3266 84896 3272
rect 85684 480 85712 69770
rect 89720 68400 89772 68406
rect 89720 68342 89772 68348
rect 88340 55956 88392 55962
rect 88340 55898 88392 55904
rect 88352 16574 88380 55898
rect 89732 16574 89760 68342
rect 93858 65784 93914 65793
rect 93858 65719 93914 65728
rect 93122 65648 93178 65657
rect 93122 65583 93178 65592
rect 92478 62928 92534 62937
rect 92478 62863 92534 62872
rect 88352 16546 89208 16574
rect 89732 16546 89944 16574
rect 87972 6180 88024 6186
rect 87972 6122 88024 6128
rect 86500 3392 86552 3398
rect 86500 3334 86552 3340
rect 84446 354 84558 480
rect 84212 326 84558 354
rect 84446 -960 84558 326
rect 85642 -960 85754 480
rect 86512 354 86540 3334
rect 87984 480 88012 6122
rect 89180 480 89208 16546
rect 86838 354 86950 480
rect 86512 326 86950 354
rect 86838 -960 86950 326
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 89916 354 89944 16546
rect 91560 3392 91612 3398
rect 91560 3334 91612 3340
rect 91572 480 91600 3334
rect 90334 354 90446 480
rect 89916 326 90446 354
rect 90334 -960 90446 326
rect 91530 -960 91642 480
rect 92492 354 92520 62863
rect 93136 3398 93164 65583
rect 93872 3398 93900 65719
rect 95240 53168 95292 53174
rect 95240 53110 95292 53116
rect 93952 51740 94004 51746
rect 93952 51682 94004 51688
rect 93124 3392 93176 3398
rect 93124 3334 93176 3340
rect 93860 3392 93912 3398
rect 93860 3334 93912 3340
rect 93964 480 93992 51682
rect 95252 16574 95280 53110
rect 96632 16574 96660 75278
rect 100128 75206 100156 148310
rect 100116 75200 100168 75206
rect 100116 75142 100168 75148
rect 100220 74361 100248 148786
rect 100392 148776 100444 148782
rect 100392 148718 100444 148724
rect 100300 148504 100352 148510
rect 100300 148446 100352 148452
rect 100206 74352 100262 74361
rect 100206 74287 100262 74296
rect 99380 73908 99432 73914
rect 99380 73850 99432 73856
rect 97998 58576 98054 58585
rect 97998 58511 98054 58520
rect 98012 16574 98040 58511
rect 99392 16574 99420 73850
rect 100220 73817 100248 74287
rect 100206 73808 100262 73817
rect 100206 73743 100262 73752
rect 100312 70378 100340 148446
rect 100300 70372 100352 70378
rect 100300 70314 100352 70320
rect 100404 70174 100432 148718
rect 100482 148336 100538 148345
rect 100482 148271 100538 148280
rect 100392 70168 100444 70174
rect 100392 70110 100444 70116
rect 99472 60716 99524 60722
rect 99472 60658 99524 60664
rect 99484 60042 99512 60658
rect 99472 60036 99524 60042
rect 99472 59978 99524 59984
rect 99472 56568 99524 56574
rect 99472 56510 99524 56516
rect 99484 55894 99512 56510
rect 99472 55888 99524 55894
rect 99472 55830 99524 55836
rect 100496 53786 100524 148271
rect 100588 60722 100616 190130
rect 100576 60716 100628 60722
rect 100576 60658 100628 60664
rect 100680 56574 100708 194346
rect 102048 193996 102100 194002
rect 102048 193938 102100 193944
rect 101956 191276 102008 191282
rect 101956 191218 102008 191224
rect 101864 190120 101916 190126
rect 101864 190062 101916 190068
rect 101588 189984 101640 189990
rect 101588 189926 101640 189932
rect 101600 84194 101628 189926
rect 101772 189916 101824 189922
rect 101772 189858 101824 189864
rect 101680 189848 101732 189854
rect 101680 189790 101732 189796
rect 101508 84166 101628 84194
rect 100760 78124 100812 78130
rect 100760 78066 100812 78072
rect 100772 77790 100800 78066
rect 101508 77790 101536 84166
rect 100760 77784 100812 77790
rect 100760 77726 100812 77732
rect 101496 77784 101548 77790
rect 101496 77726 101548 77732
rect 101692 57934 101720 189790
rect 100760 57928 100812 57934
rect 100760 57870 100812 57876
rect 101680 57928 101732 57934
rect 101680 57870 101732 57876
rect 100772 57254 100800 57870
rect 100760 57248 100812 57254
rect 100760 57190 100812 57196
rect 100668 56568 100720 56574
rect 100668 56510 100720 56516
rect 100484 53780 100536 53786
rect 100484 53722 100536 53728
rect 100496 53106 100524 53722
rect 100484 53100 100536 53106
rect 100484 53042 100536 53048
rect 101784 52465 101812 189858
rect 100758 52456 100814 52465
rect 100758 52391 100814 52400
rect 101770 52456 101826 52465
rect 101770 52391 101826 52400
rect 100772 51785 100800 52391
rect 100758 51776 100814 51785
rect 100758 51711 100814 51720
rect 101876 51066 101904 190062
rect 100760 51060 100812 51066
rect 100760 51002 100812 51008
rect 101864 51060 101916 51066
rect 101864 51002 101916 51008
rect 100772 50386 100800 51002
rect 100760 50380 100812 50386
rect 100760 50322 100812 50328
rect 100758 49600 100814 49609
rect 100758 49535 100814 49544
rect 100772 48929 100800 49535
rect 100758 48920 100814 48929
rect 100758 48855 100814 48864
rect 101968 48249 101996 191218
rect 102060 49609 102088 193938
rect 103060 192568 103112 192574
rect 103060 192510 103112 192516
rect 102784 186992 102836 186998
rect 102784 186934 102836 186940
rect 102692 148640 102744 148646
rect 102692 148582 102744 148588
rect 102140 78600 102192 78606
rect 102140 78542 102192 78548
rect 102152 78062 102180 78542
rect 102140 78056 102192 78062
rect 102140 77998 102192 78004
rect 102140 73024 102192 73030
rect 102140 72966 102192 72972
rect 102152 72622 102180 72966
rect 102140 72616 102192 72622
rect 102140 72558 102192 72564
rect 102140 71528 102192 71534
rect 102140 71470 102192 71476
rect 102152 71126 102180 71470
rect 102140 71120 102192 71126
rect 102140 71062 102192 71068
rect 102140 70304 102192 70310
rect 102140 70246 102192 70252
rect 102152 69902 102180 70246
rect 102232 70100 102284 70106
rect 102232 70042 102284 70048
rect 102140 69896 102192 69902
rect 102140 69838 102192 69844
rect 102244 69766 102272 70042
rect 102232 69760 102284 69766
rect 102232 69702 102284 69708
rect 102140 66224 102192 66230
rect 102140 66166 102192 66172
rect 102152 65550 102180 66166
rect 102140 65544 102192 65550
rect 102140 65486 102192 65492
rect 102140 64864 102192 64870
rect 102140 64806 102192 64812
rect 102230 64832 102286 64841
rect 102046 49600 102102 49609
rect 102046 49535 102102 49544
rect 100758 48240 100814 48249
rect 100758 48175 100814 48184
rect 101954 48240 102010 48249
rect 101954 48175 102010 48184
rect 100772 47569 100800 48175
rect 100758 47560 100814 47569
rect 100758 47495 100814 47504
rect 102152 16574 102180 64806
rect 102230 64767 102286 64776
rect 102244 64161 102272 64767
rect 102230 64152 102286 64161
rect 102230 64087 102286 64096
rect 102232 62076 102284 62082
rect 102232 62018 102284 62024
rect 102244 61470 102272 62018
rect 102232 61464 102284 61470
rect 102232 61406 102284 61412
rect 102704 46889 102732 148582
rect 102796 73030 102824 186934
rect 102876 184204 102928 184210
rect 102876 184146 102928 184152
rect 102888 78606 102916 184146
rect 102968 176996 103020 177002
rect 102968 176938 103020 176944
rect 102876 78600 102928 78606
rect 102876 78542 102928 78548
rect 102784 73024 102836 73030
rect 102784 72966 102836 72972
rect 102980 71534 103008 176938
rect 102968 71528 103020 71534
rect 102968 71470 103020 71476
rect 102784 71256 102836 71262
rect 102784 71198 102836 71204
rect 102230 46880 102286 46889
rect 102230 46815 102286 46824
rect 102690 46880 102746 46889
rect 102690 46815 102746 46824
rect 102244 46209 102272 46815
rect 102230 46200 102286 46209
rect 102230 46135 102286 46144
rect 95252 16546 95832 16574
rect 96632 16546 97488 16574
rect 98012 16546 98224 16574
rect 99392 16546 99880 16574
rect 102152 16546 102272 16574
rect 94780 3392 94832 3398
rect 94780 3334 94832 3340
rect 92726 354 92838 480
rect 92492 326 92838 354
rect 92726 -960 92838 326
rect 93922 -960 94034 480
rect 94792 354 94820 3334
rect 95118 354 95230 480
rect 94792 326 95230 354
rect 95804 354 95832 16546
rect 97460 480 97488 16546
rect 96222 354 96334 480
rect 95804 326 96334 354
rect 95118 -960 95230 326
rect 96222 -960 96334 326
rect 97418 -960 97530 480
rect 98196 354 98224 16546
rect 99852 480 99880 16546
rect 101036 3392 101088 3398
rect 101036 3334 101088 3340
rect 101048 480 101076 3334
rect 102244 480 102272 16546
rect 102796 3398 102824 71198
rect 103072 70310 103100 192510
rect 103152 192500 103204 192506
rect 103152 192442 103204 192448
rect 103060 70304 103112 70310
rect 103060 70246 103112 70252
rect 103164 66230 103192 192442
rect 103256 70106 103284 199815
rect 104440 199504 104492 199510
rect 104440 199446 104492 199452
rect 104452 194410 104480 199446
rect 105544 195288 105596 195294
rect 105544 195230 105596 195236
rect 104806 195120 104862 195129
rect 104806 195055 104862 195064
rect 104440 194404 104492 194410
rect 104440 194346 104492 194352
rect 104254 192808 104310 192817
rect 104254 192743 104310 192752
rect 103336 192704 103388 192710
rect 103336 192646 103388 192652
rect 103244 70100 103296 70106
rect 103244 70042 103296 70048
rect 103152 66224 103204 66230
rect 103152 66166 103204 66172
rect 103348 64841 103376 192646
rect 104072 192636 104124 192642
rect 104072 192578 104124 192584
rect 103428 185768 103480 185774
rect 103428 185710 103480 185716
rect 103334 64832 103390 64841
rect 103334 64767 103390 64776
rect 103440 62082 103468 185710
rect 103980 148572 104032 148578
rect 103980 148514 104032 148520
rect 103520 69896 103572 69902
rect 103520 69838 103572 69844
rect 103428 62076 103480 62082
rect 103428 62018 103480 62024
rect 103532 16574 103560 69838
rect 103886 60616 103942 60625
rect 103886 60551 103942 60560
rect 103900 59945 103928 60551
rect 103886 59936 103942 59945
rect 103886 59871 103942 59880
rect 103992 55185 104020 148514
rect 104084 77042 104112 192578
rect 104164 181620 104216 181626
rect 104164 181562 104216 181568
rect 104072 77036 104124 77042
rect 104072 76978 104124 76984
rect 104176 76265 104204 181562
rect 104162 76256 104218 76265
rect 104162 76191 104218 76200
rect 104268 75478 104296 192743
rect 104820 189990 104848 195055
rect 104808 189984 104860 189990
rect 104808 189926 104860 189932
rect 104808 189780 104860 189786
rect 104808 189722 104860 189728
rect 104438 186552 104494 186561
rect 104438 186487 104494 186496
rect 104348 185564 104400 185570
rect 104348 185506 104400 185512
rect 104256 75472 104308 75478
rect 104256 75414 104308 75420
rect 104360 74186 104388 185506
rect 104348 74180 104400 74186
rect 104348 74122 104400 74128
rect 104452 68746 104480 186487
rect 104624 185632 104676 185638
rect 104624 185574 104676 185580
rect 104532 182572 104584 182578
rect 104532 182514 104584 182520
rect 104544 72418 104572 182514
rect 104532 72412 104584 72418
rect 104532 72354 104584 72360
rect 104636 70666 104664 185574
rect 104716 176452 104768 176458
rect 104716 176394 104768 176400
rect 104544 70638 104664 70666
rect 104440 68740 104492 68746
rect 104440 68682 104492 68688
rect 104544 67522 104572 70638
rect 104624 68740 104676 68746
rect 104624 68682 104676 68688
rect 104636 68338 104664 68682
rect 104624 68332 104676 68338
rect 104624 68274 104676 68280
rect 104532 67516 104584 67522
rect 104532 67458 104584 67464
rect 104544 66910 104572 67458
rect 104532 66904 104584 66910
rect 104532 66846 104584 66852
rect 104728 63510 104756 176394
rect 104716 63504 104768 63510
rect 104716 63446 104768 63452
rect 104728 62830 104756 63446
rect 104716 62824 104768 62830
rect 104716 62766 104768 62772
rect 104820 60625 104848 189722
rect 105556 75818 105584 195230
rect 105544 75812 105596 75818
rect 105544 75754 105596 75760
rect 104806 60616 104862 60625
rect 104806 60551 104862 60560
rect 103978 55176 104034 55185
rect 103978 55111 104034 55120
rect 103992 54505 104020 55111
rect 103978 54496 104034 54505
rect 103978 54431 104034 54440
rect 104898 54496 104954 54505
rect 104898 54431 104954 54440
rect 104164 36576 104216 36582
rect 104164 36518 104216 36524
rect 103532 16546 104112 16574
rect 103336 4140 103388 4146
rect 103336 4082 103388 4088
rect 102784 3392 102836 3398
rect 102784 3334 102836 3340
rect 103348 480 103376 4082
rect 98614 354 98726 480
rect 98196 326 98726 354
rect 98614 -960 98726 326
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104084 354 104112 16546
rect 104176 4146 104204 36518
rect 104912 16574 104940 54431
rect 105556 51746 105584 75754
rect 105648 71398 105676 200087
rect 106924 199912 106976 199918
rect 106924 199854 106976 199860
rect 105912 196784 105964 196790
rect 105912 196726 105964 196732
rect 105728 195492 105780 195498
rect 105728 195434 105780 195440
rect 105740 72962 105768 195434
rect 105820 185700 105872 185706
rect 105820 185642 105872 185648
rect 105728 72956 105780 72962
rect 105728 72898 105780 72904
rect 105740 72690 105768 72898
rect 105728 72684 105780 72690
rect 105728 72626 105780 72632
rect 105636 71392 105688 71398
rect 105636 71334 105688 71340
rect 105832 68218 105860 185642
rect 105924 70242 105952 196726
rect 106004 195560 106056 195566
rect 106004 195502 106056 195508
rect 105912 70236 105964 70242
rect 105912 70178 105964 70184
rect 105924 69902 105952 70178
rect 105912 69896 105964 69902
rect 105912 69838 105964 69844
rect 106016 68882 106044 195502
rect 106832 195356 106884 195362
rect 106832 195298 106884 195304
rect 106096 193860 106148 193866
rect 106096 193802 106148 193808
rect 106004 68876 106056 68882
rect 106004 68818 106056 68824
rect 106016 68406 106044 68818
rect 106004 68400 106056 68406
rect 106004 68342 106056 68348
rect 105832 68190 106044 68218
rect 106016 67590 106044 68190
rect 106004 67584 106056 67590
rect 106004 67526 106056 67532
rect 106016 66978 106044 67526
rect 106004 66972 106056 66978
rect 106004 66914 106056 66920
rect 106108 64870 106136 193802
rect 106738 192536 106794 192545
rect 106738 192471 106794 192480
rect 106188 190256 106240 190262
rect 106188 190198 106240 190204
rect 106096 64864 106148 64870
rect 106096 64806 106148 64812
rect 106200 57905 106228 190198
rect 106752 79558 106780 192471
rect 106844 79898 106872 195298
rect 106832 79892 106884 79898
rect 106832 79834 106884 79840
rect 106740 79552 106792 79558
rect 106740 79494 106792 79500
rect 106844 79370 106872 79834
rect 106752 79342 106872 79370
rect 106372 76696 106424 76702
rect 106372 76638 106424 76644
rect 106384 64874 106412 76638
rect 106752 71262 106780 79342
rect 106832 78532 106884 78538
rect 106832 78474 106884 78480
rect 106844 77654 106872 78474
rect 106936 78062 106964 199854
rect 107016 184408 107068 184414
rect 107016 184350 107068 184356
rect 107028 78402 107056 184350
rect 107108 174276 107160 174282
rect 107108 174218 107160 174224
rect 107120 78470 107148 174218
rect 107212 78538 107240 200223
rect 108762 198112 108818 198121
rect 108762 198047 108818 198056
rect 108672 192908 108724 192914
rect 108672 192850 108724 192856
rect 107568 190324 107620 190330
rect 107568 190266 107620 190272
rect 107384 189712 107436 189718
rect 107384 189654 107436 189660
rect 107292 186244 107344 186250
rect 107292 186186 107344 186192
rect 107200 78532 107252 78538
rect 107200 78474 107252 78480
rect 107108 78464 107160 78470
rect 107108 78406 107160 78412
rect 107016 78396 107068 78402
rect 107016 78338 107068 78344
rect 107200 78396 107252 78402
rect 107200 78338 107252 78344
rect 107212 78198 107240 78338
rect 107200 78192 107252 78198
rect 107200 78134 107252 78140
rect 106924 78056 106976 78062
rect 106924 77998 106976 78004
rect 106832 77648 106884 77654
rect 106832 77590 106884 77596
rect 107304 74225 107332 186186
rect 107290 74216 107346 74225
rect 107290 74151 107346 74160
rect 106740 71256 106792 71262
rect 106740 71198 106792 71204
rect 107396 67561 107424 189654
rect 107474 185872 107530 185881
rect 107474 185807 107530 185816
rect 107488 71330 107516 185807
rect 107476 71324 107528 71330
rect 107476 71266 107528 71272
rect 107382 67552 107438 67561
rect 107382 67487 107438 67496
rect 106292 64846 106412 64874
rect 105818 57896 105874 57905
rect 105818 57831 105874 57840
rect 106186 57896 106242 57905
rect 106186 57831 106242 57840
rect 105832 57225 105860 57831
rect 105818 57216 105874 57225
rect 105818 57151 105874 57160
rect 105544 51740 105596 51746
rect 105544 51682 105596 51688
rect 106292 16574 106320 64846
rect 107580 59265 107608 190266
rect 108302 186824 108358 186833
rect 108302 186759 108358 186768
rect 108212 178492 108264 178498
rect 108212 178434 108264 178440
rect 108120 148912 108172 148918
rect 108120 148854 108172 148860
rect 107660 71800 107712 71806
rect 107660 71742 107712 71748
rect 107566 59256 107622 59265
rect 107566 59191 107622 59200
rect 107580 58585 107608 59191
rect 107566 58576 107622 58585
rect 107566 58511 107622 58520
rect 107672 16574 107700 71742
rect 108132 63481 108160 148854
rect 108224 80850 108252 178434
rect 108212 80844 108264 80850
rect 108212 80786 108264 80792
rect 108224 80714 108252 80786
rect 108212 80708 108264 80714
rect 108212 80650 108264 80656
rect 108316 76770 108344 186759
rect 108580 185224 108632 185230
rect 108580 185166 108632 185172
rect 108396 185020 108448 185026
rect 108396 184962 108448 184968
rect 108408 80986 108436 184962
rect 108488 182164 108540 182170
rect 108488 182106 108540 182112
rect 108396 80980 108448 80986
rect 108396 80922 108448 80928
rect 108500 78266 108528 182106
rect 108488 78260 108540 78266
rect 108488 78202 108540 78208
rect 108592 78130 108620 185166
rect 108580 78124 108632 78130
rect 108580 78066 108632 78072
rect 108304 76764 108356 76770
rect 108304 76706 108356 76712
rect 108684 72894 108712 192850
rect 108776 75342 108804 198047
rect 109776 195424 109828 195430
rect 109776 195366 109828 195372
rect 108948 193724 109000 193730
rect 108948 193666 109000 193672
rect 108856 189644 108908 189650
rect 108856 189586 108908 189592
rect 108764 75336 108816 75342
rect 108764 75278 108816 75284
rect 108672 72888 108724 72894
rect 108672 72830 108724 72836
rect 108684 71806 108712 72830
rect 108672 71800 108724 71806
rect 108672 71742 108724 71748
rect 108868 66201 108896 189586
rect 108854 66192 108910 66201
rect 108854 66127 108910 66136
rect 108960 64802 108988 193666
rect 109684 191140 109736 191146
rect 109684 191082 109736 191088
rect 109696 79762 109724 191082
rect 109684 79756 109736 79762
rect 109684 79698 109736 79704
rect 109788 79354 109816 195366
rect 109868 191208 109920 191214
rect 109868 191150 109920 191156
rect 109776 79348 109828 79354
rect 109776 79290 109828 79296
rect 109880 73098 109908 191150
rect 109972 79422 110000 200631
rect 110144 196852 110196 196858
rect 110144 196794 110196 196800
rect 110052 190460 110104 190466
rect 110052 190402 110104 190408
rect 109960 79416 110012 79422
rect 109960 79358 110012 79364
rect 109868 73092 109920 73098
rect 109868 73034 109920 73040
rect 110064 68377 110092 190402
rect 110156 74458 110184 196794
rect 110236 195628 110288 195634
rect 110236 195570 110288 195576
rect 110144 74452 110196 74458
rect 110144 74394 110196 74400
rect 110248 68814 110276 195570
rect 110972 192976 111024 192982
rect 110972 192918 111024 192924
rect 110328 192364 110380 192370
rect 110328 192306 110380 192312
rect 110236 68808 110288 68814
rect 110236 68750 110288 68756
rect 110050 68368 110106 68377
rect 110050 68303 110106 68312
rect 108948 64796 109000 64802
rect 108948 64738 109000 64744
rect 108960 64258 108988 64738
rect 108948 64252 109000 64258
rect 108948 64194 109000 64200
rect 108118 63472 108174 63481
rect 108118 63407 108174 63416
rect 108132 62937 108160 63407
rect 110340 63345 110368 192306
rect 110880 190392 110932 190398
rect 110880 190334 110932 190340
rect 110892 79626 110920 190334
rect 110880 79620 110932 79626
rect 110880 79562 110932 79568
rect 110984 79490 111012 192918
rect 111076 147014 111104 262754
rect 112352 261112 112404 261118
rect 112352 261054 112404 261060
rect 111616 199028 111668 199034
rect 111616 198970 111668 198976
rect 111432 196920 111484 196926
rect 111432 196862 111484 196868
rect 111248 195764 111300 195770
rect 111248 195706 111300 195712
rect 111156 195696 111208 195702
rect 111156 195638 111208 195644
rect 111064 147008 111116 147014
rect 111064 146950 111116 146956
rect 111064 141092 111116 141098
rect 111064 141034 111116 141040
rect 110972 79484 111024 79490
rect 110972 79426 111024 79432
rect 110326 63336 110382 63345
rect 110326 63271 110382 63280
rect 108118 62928 108174 62937
rect 108118 62863 108174 62872
rect 110340 62801 110368 63271
rect 110326 62792 110382 62801
rect 110326 62727 110382 62736
rect 110420 59900 110472 59906
rect 110420 59842 110472 59848
rect 110432 16574 110460 59842
rect 111076 59362 111104 141034
rect 111168 74254 111196 195638
rect 111156 74248 111208 74254
rect 111156 74190 111208 74196
rect 111260 72826 111288 195706
rect 111340 191344 111392 191350
rect 111340 191286 111392 191292
rect 111248 72820 111300 72826
rect 111248 72762 111300 72768
rect 111352 68785 111380 191286
rect 111444 72758 111472 196862
rect 111524 190052 111576 190058
rect 111524 189994 111576 190000
rect 111432 72752 111484 72758
rect 111432 72694 111484 72700
rect 111338 68776 111394 68785
rect 111338 68711 111394 68720
rect 111156 68604 111208 68610
rect 111156 68546 111208 68552
rect 111064 59356 111116 59362
rect 111064 59298 111116 59304
rect 104912 16546 105768 16574
rect 106292 16546 106504 16574
rect 107672 16546 108160 16574
rect 110432 16546 110552 16574
rect 104164 4140 104216 4146
rect 104164 4082 104216 4088
rect 105740 480 105768 16546
rect 104502 354 104614 480
rect 104084 326 104614 354
rect 104502 -960 104614 326
rect 105698 -960 105810 480
rect 106476 354 106504 16546
rect 108132 480 108160 16546
rect 109316 3392 109368 3398
rect 109316 3334 109368 3340
rect 109328 480 109356 3334
rect 110524 480 110552 16546
rect 111168 3398 111196 68546
rect 111536 65657 111564 189994
rect 111628 72486 111656 198970
rect 111706 198656 111762 198665
rect 111706 198591 111762 198600
rect 111616 72480 111668 72486
rect 111616 72422 111668 72428
rect 111720 71369 111748 198591
rect 112168 148980 112220 148986
rect 112168 148922 112220 148928
rect 111800 75948 111852 75954
rect 111800 75890 111852 75896
rect 111706 71360 111762 71369
rect 111706 71295 111762 71304
rect 111522 65648 111578 65657
rect 111522 65583 111578 65592
rect 111812 16574 111840 75890
rect 112180 71466 112208 148922
rect 112364 146062 112392 261054
rect 112352 146056 112404 146062
rect 112352 145998 112404 146004
rect 112352 145580 112404 145586
rect 112352 145522 112404 145528
rect 112260 141568 112312 141574
rect 112260 141510 112312 141516
rect 112272 76809 112300 141510
rect 112258 76800 112314 76809
rect 112258 76735 112314 76744
rect 112168 71460 112220 71466
rect 112168 71402 112220 71408
rect 112272 68610 112300 76735
rect 112260 68604 112312 68610
rect 112260 68546 112312 68552
rect 112364 67017 112392 145522
rect 112456 144226 112484 263026
rect 113824 260908 113876 260914
rect 113824 260850 113876 260856
rect 112996 199368 113048 199374
rect 112996 199310 113048 199316
rect 112628 196648 112680 196654
rect 112628 196590 112680 196596
rect 112536 189576 112588 189582
rect 112536 189518 112588 189524
rect 112444 144220 112496 144226
rect 112444 144162 112496 144168
rect 112548 71194 112576 189518
rect 112640 77217 112668 196590
rect 112812 194268 112864 194274
rect 112812 194210 112864 194216
rect 112720 194132 112772 194138
rect 112720 194074 112772 194080
rect 112626 77208 112682 77217
rect 112626 77143 112682 77152
rect 112732 74322 112760 194074
rect 112720 74316 112772 74322
rect 112720 74258 112772 74264
rect 112824 71233 112852 194210
rect 112902 191040 112958 191049
rect 112902 190975 112958 190984
rect 112810 71224 112866 71233
rect 112536 71188 112588 71194
rect 112810 71159 112866 71168
rect 112536 71130 112588 71136
rect 112916 68513 112944 190975
rect 113008 75721 113036 199310
rect 113088 198960 113140 198966
rect 113088 198902 113140 198908
rect 112994 75712 113050 75721
rect 113100 75682 113128 198902
rect 113548 148232 113600 148238
rect 113548 148174 113600 148180
rect 113456 146940 113508 146946
rect 113456 146882 113508 146888
rect 112994 75647 113050 75656
rect 113088 75676 113140 75682
rect 113088 75618 113140 75624
rect 113468 75313 113496 146882
rect 113454 75304 113510 75313
rect 113454 75239 113510 75248
rect 113560 71262 113588 148174
rect 113836 146198 113864 260850
rect 113916 259956 113968 259962
rect 113916 259898 113968 259904
rect 113824 146192 113876 146198
rect 113824 146134 113876 146140
rect 113640 144764 113692 144770
rect 113640 144706 113692 144712
rect 113652 75954 113680 144706
rect 113732 144288 113784 144294
rect 113732 144230 113784 144236
rect 113640 75948 113692 75954
rect 113640 75890 113692 75896
rect 113744 75750 113772 144230
rect 113928 141710 113956 259898
rect 114100 194200 114152 194206
rect 114100 194142 114152 194148
rect 114008 194064 114060 194070
rect 114008 194006 114060 194012
rect 113916 141704 113968 141710
rect 113916 141646 113968 141652
rect 113916 139460 113968 139466
rect 113916 139402 113968 139408
rect 113732 75744 113784 75750
rect 113732 75686 113784 75692
rect 113548 71256 113600 71262
rect 113548 71198 113600 71204
rect 113928 70281 113956 139402
rect 114020 75002 114048 194006
rect 114112 75546 114140 194142
rect 114204 144702 114232 263842
rect 114296 146130 114324 264930
rect 119160 264444 119212 264450
rect 119160 264386 119212 264392
rect 118148 264308 118200 264314
rect 118148 264250 118200 264256
rect 117136 264172 117188 264178
rect 117136 264114 117188 264120
rect 117044 264036 117096 264042
rect 117044 263978 117096 263984
rect 115204 263016 115256 263022
rect 115204 262958 115256 262964
rect 115112 259480 115164 259486
rect 115112 259422 115164 259428
rect 114374 199472 114430 199481
rect 114374 199407 114430 199416
rect 114284 146124 114336 146130
rect 114284 146066 114336 146072
rect 114284 144832 114336 144838
rect 114284 144774 114336 144780
rect 114192 144696 114244 144702
rect 114192 144638 114244 144644
rect 114100 75540 114152 75546
rect 114100 75482 114152 75488
rect 114008 74996 114060 75002
rect 114008 74938 114060 74944
rect 113914 70272 113970 70281
rect 113914 70207 113970 70216
rect 114296 68678 114324 144774
rect 114388 77081 114416 199407
rect 114468 199096 114520 199102
rect 114468 199038 114520 199044
rect 114374 77072 114430 77081
rect 114374 77007 114430 77016
rect 114376 76424 114428 76430
rect 114376 76366 114428 76372
rect 114388 75954 114416 76366
rect 114376 75948 114428 75954
rect 114376 75890 114428 75896
rect 114480 75410 114508 199038
rect 114836 145784 114888 145790
rect 114836 145726 114888 145732
rect 114744 145648 114796 145654
rect 114744 145590 114796 145596
rect 114468 75404 114520 75410
rect 114468 75346 114520 75352
rect 114560 75132 114612 75138
rect 114560 75074 114612 75080
rect 114284 68672 114336 68678
rect 114284 68614 114336 68620
rect 112902 68504 112958 68513
rect 112902 68439 112958 68448
rect 113180 68332 113232 68338
rect 113180 68274 113232 68280
rect 112350 67008 112406 67017
rect 112350 66943 112406 66952
rect 113192 16574 113220 68274
rect 113824 55208 113876 55214
rect 113824 55150 113876 55156
rect 113836 55049 113864 55150
rect 113822 55040 113878 55049
rect 113822 54975 113878 54984
rect 113836 54505 113864 54975
rect 113822 54496 113878 54505
rect 113822 54431 113878 54440
rect 114572 16574 114600 75074
rect 114756 73642 114784 145590
rect 114848 79830 114876 145726
rect 114928 145716 114980 145722
rect 114928 145658 114980 145664
rect 114836 79824 114888 79830
rect 114836 79766 114888 79772
rect 114744 73636 114796 73642
rect 114744 73578 114796 73584
rect 114940 71777 114968 145658
rect 115124 145450 115152 259422
rect 115216 145518 115244 262958
rect 116952 262744 117004 262750
rect 116952 262686 117004 262692
rect 116768 261180 116820 261186
rect 116768 261122 116820 261128
rect 116584 260024 116636 260030
rect 116584 259966 116636 259972
rect 115388 259888 115440 259894
rect 115388 259830 115440 259836
rect 115296 259548 115348 259554
rect 115296 259490 115348 259496
rect 115204 145512 115256 145518
rect 115204 145454 115256 145460
rect 115112 145444 115164 145450
rect 115112 145386 115164 145392
rect 115308 141846 115336 259490
rect 115296 141840 115348 141846
rect 115296 141782 115348 141788
rect 115400 141506 115428 259830
rect 115756 199300 115808 199306
rect 115756 199242 115808 199248
rect 115664 197668 115716 197674
rect 115664 197610 115716 197616
rect 115480 196716 115532 196722
rect 115480 196658 115532 196664
rect 115388 141500 115440 141506
rect 115388 141442 115440 141448
rect 115018 139224 115074 139233
rect 115018 139159 115074 139168
rect 115032 80238 115060 139159
rect 115110 138952 115166 138961
rect 115110 138887 115166 138896
rect 115020 80232 115072 80238
rect 115020 80174 115072 80180
rect 114926 71768 114982 71777
rect 114926 71703 114982 71712
rect 115032 59906 115060 80174
rect 115124 75138 115152 138887
rect 115492 76362 115520 196658
rect 115570 193896 115626 193905
rect 115570 193831 115626 193840
rect 115480 76356 115532 76362
rect 115480 76298 115532 76304
rect 115112 75132 115164 75138
rect 115112 75074 115164 75080
rect 115584 74390 115612 193831
rect 115676 77110 115704 197610
rect 115664 77104 115716 77110
rect 115664 77046 115716 77052
rect 115768 76838 115796 199242
rect 115848 194336 115900 194342
rect 115848 194278 115900 194284
rect 115756 76832 115808 76838
rect 115756 76774 115808 76780
rect 115572 74384 115624 74390
rect 115572 74326 115624 74332
rect 115860 68649 115888 194278
rect 116308 148436 116360 148442
rect 116308 148378 116360 148384
rect 116214 146976 116270 146985
rect 116214 146911 116270 146920
rect 116124 144900 116176 144906
rect 116124 144842 116176 144848
rect 116136 69018 116164 144842
rect 116228 71126 116256 146911
rect 116320 71670 116348 148378
rect 116596 144634 116624 259966
rect 116676 259820 116728 259826
rect 116676 259762 116728 259768
rect 116584 144628 116636 144634
rect 116584 144570 116636 144576
rect 116688 142186 116716 259762
rect 116780 143342 116808 261122
rect 116860 192432 116912 192438
rect 116860 192374 116912 192380
rect 116768 143336 116820 143342
rect 116768 143278 116820 143284
rect 116676 142180 116728 142186
rect 116676 142122 116728 142128
rect 116676 140480 116728 140486
rect 116676 140422 116728 140428
rect 116584 140412 116636 140418
rect 116584 140354 116636 140360
rect 116400 140140 116452 140146
rect 116400 140082 116452 140088
rect 116412 80782 116440 140082
rect 116492 140072 116544 140078
rect 116492 140014 116544 140020
rect 116400 80776 116452 80782
rect 116400 80718 116452 80724
rect 116504 78946 116532 140014
rect 116492 78940 116544 78946
rect 116492 78882 116544 78888
rect 116596 76945 116624 140354
rect 116582 76936 116638 76945
rect 116582 76871 116638 76880
rect 116688 74118 116716 140422
rect 116766 138816 116822 138825
rect 116766 138751 116822 138760
rect 116676 74112 116728 74118
rect 116676 74054 116728 74060
rect 116308 71664 116360 71670
rect 116308 71606 116360 71612
rect 116216 71120 116268 71126
rect 116216 71062 116268 71068
rect 116780 70038 116808 138751
rect 116872 74089 116900 192374
rect 116964 141778 116992 262686
rect 117056 143138 117084 263978
rect 117044 143132 117096 143138
rect 117044 143074 117096 143080
rect 116952 141772 117004 141778
rect 116952 141714 117004 141720
rect 117148 141642 117176 264114
rect 118056 262880 118108 262886
rect 118056 262822 118108 262828
rect 117964 262676 118016 262682
rect 117964 262618 118016 262624
rect 117872 262404 117924 262410
rect 117872 262346 117924 262352
rect 117228 199164 117280 199170
rect 117228 199106 117280 199112
rect 117136 141636 117188 141642
rect 117136 141578 117188 141584
rect 117240 76974 117268 199106
rect 117884 166326 117912 262346
rect 117872 166320 117924 166326
rect 117872 166262 117924 166268
rect 117688 148708 117740 148714
rect 117688 148650 117740 148656
rect 117700 80714 117728 148650
rect 117884 143410 117912 166262
rect 117976 145994 118004 262618
rect 117964 145988 118016 145994
rect 117964 145930 118016 145936
rect 117964 145852 118016 145858
rect 117964 145794 118016 145800
rect 117872 143404 117924 143410
rect 117872 143346 117924 143352
rect 117870 140312 117926 140321
rect 117870 140247 117926 140256
rect 117780 140208 117832 140214
rect 117780 140150 117832 140156
rect 117688 80708 117740 80714
rect 117688 80650 117740 80656
rect 117792 80209 117820 140150
rect 117778 80200 117834 80209
rect 117778 80135 117834 80144
rect 117884 79694 117912 140247
rect 117872 79688 117924 79694
rect 117872 79630 117924 79636
rect 117976 79150 118004 145794
rect 118068 143274 118096 262822
rect 118056 143268 118108 143274
rect 118056 143210 118108 143216
rect 118160 143002 118188 264250
rect 118332 263764 118384 263770
rect 118332 263706 118384 263712
rect 118240 259752 118292 259758
rect 118240 259694 118292 259700
rect 118252 259593 118280 259694
rect 118238 259584 118294 259593
rect 118238 259519 118294 259528
rect 118240 197056 118292 197062
rect 118240 196998 118292 197004
rect 118148 142996 118200 143002
rect 118148 142938 118200 142944
rect 118056 136332 118108 136338
rect 118056 136274 118108 136280
rect 117964 79144 118016 79150
rect 117964 79086 118016 79092
rect 117228 76968 117280 76974
rect 117228 76910 117280 76916
rect 116858 74080 116914 74089
rect 118068 74050 118096 136274
rect 118252 75886 118280 196998
rect 118344 142118 118372 263706
rect 118424 199232 118476 199238
rect 118424 199174 118476 199180
rect 118332 142112 118384 142118
rect 118332 142054 118384 142060
rect 118332 139664 118384 139670
rect 118332 139606 118384 139612
rect 118240 75880 118292 75886
rect 118240 75822 118292 75828
rect 116858 74015 116914 74024
rect 118056 74044 118108 74050
rect 118056 73986 118108 73992
rect 118344 71738 118372 139606
rect 118436 75585 118464 199174
rect 118606 198928 118662 198937
rect 118606 198863 118662 198872
rect 118516 193928 118568 193934
rect 118516 193870 118568 193876
rect 118422 75576 118478 75585
rect 118422 75511 118478 75520
rect 118332 71732 118384 71738
rect 118332 71674 118384 71680
rect 116768 70032 116820 70038
rect 116768 69974 116820 69980
rect 116124 69012 116176 69018
rect 116124 68954 116176 68960
rect 118528 68950 118556 193870
rect 118620 73166 118648 198863
rect 119068 145920 119120 145926
rect 119068 145862 119120 145868
rect 118700 141160 118752 141166
rect 118700 141102 118752 141108
rect 118712 137970 118740 141102
rect 118700 137964 118752 137970
rect 118700 137906 118752 137912
rect 119080 79082 119108 145862
rect 119172 143041 119200 264386
rect 134536 264178 134564 271866
rect 133972 264172 134024 264178
rect 133972 264114 134024 264120
rect 134524 264172 134576 264178
rect 134524 264114 134576 264120
rect 119804 264104 119856 264110
rect 119804 264046 119856 264052
rect 119620 263968 119672 263974
rect 119620 263910 119672 263916
rect 119436 262540 119488 262546
rect 119436 262482 119488 262488
rect 119344 259684 119396 259690
rect 119344 259626 119396 259632
rect 119252 259616 119304 259622
rect 119252 259558 119304 259564
rect 119264 144430 119292 259558
rect 119252 144424 119304 144430
rect 119252 144366 119304 144372
rect 119158 143032 119214 143041
rect 119158 142967 119214 142976
rect 119356 142769 119384 259626
rect 119448 144498 119476 262482
rect 119528 262336 119580 262342
rect 119528 262278 119580 262284
rect 119436 144492 119488 144498
rect 119436 144434 119488 144440
rect 119342 142760 119398 142769
rect 119342 142695 119398 142704
rect 119540 141914 119568 262278
rect 119632 142934 119660 263910
rect 119816 143206 119844 264046
rect 121000 263832 121052 263838
rect 121000 263774 121052 263780
rect 120908 263628 120960 263634
rect 120908 263570 120960 263576
rect 120632 262608 120684 262614
rect 120632 262550 120684 262556
rect 120540 261044 120592 261050
rect 120540 260986 120592 260992
rect 120354 198248 120410 198257
rect 120354 198183 120410 198192
rect 119986 196752 120042 196761
rect 119986 196687 120042 196696
rect 119896 195900 119948 195906
rect 119896 195842 119948 195848
rect 119804 143200 119856 143206
rect 119804 143142 119856 143148
rect 119620 142928 119672 142934
rect 119620 142870 119672 142876
rect 119712 142724 119764 142730
rect 119712 142666 119764 142672
rect 119528 141908 119580 141914
rect 119528 141850 119580 141856
rect 119528 140684 119580 140690
rect 119528 140626 119580 140632
rect 119344 140276 119396 140282
rect 119344 140218 119396 140224
rect 119250 138544 119306 138553
rect 119250 138479 119306 138488
rect 119068 79076 119120 79082
rect 119068 79018 119120 79024
rect 119264 79014 119292 138479
rect 119356 79286 119384 140218
rect 119344 79280 119396 79286
rect 119344 79222 119396 79228
rect 119252 79008 119304 79014
rect 119252 78950 119304 78956
rect 119540 73778 119568 140626
rect 119620 140004 119672 140010
rect 119620 139946 119672 139952
rect 119632 73982 119660 139946
rect 119724 77178 119752 142666
rect 119804 140752 119856 140758
rect 119804 140694 119856 140700
rect 119712 77172 119764 77178
rect 119712 77114 119764 77120
rect 119620 73976 119672 73982
rect 119620 73918 119672 73924
rect 119528 73772 119580 73778
rect 119528 73714 119580 73720
rect 118608 73160 118660 73166
rect 118608 73102 118660 73108
rect 119816 72690 119844 140694
rect 119908 72865 119936 195842
rect 120000 73001 120028 196687
rect 120368 195770 120396 198183
rect 120356 195764 120408 195770
rect 120356 195706 120408 195712
rect 120170 194848 120226 194857
rect 120170 194783 120226 194792
rect 120184 189582 120212 194783
rect 120172 189576 120224 189582
rect 120172 189518 120224 189524
rect 120552 189038 120580 260986
rect 120540 189032 120592 189038
rect 120540 188974 120592 188980
rect 120540 144560 120592 144566
rect 120540 144502 120592 144508
rect 120552 76906 120580 144502
rect 120644 144362 120672 262550
rect 120816 259412 120868 259418
rect 120816 259354 120868 259360
rect 120722 199064 120778 199073
rect 120722 198999 120778 199008
rect 120632 144356 120684 144362
rect 120632 144298 120684 144304
rect 120736 79529 120764 198999
rect 120828 141982 120856 259354
rect 120920 142905 120948 263570
rect 120906 142896 120962 142905
rect 121012 142866 121040 263774
rect 121092 263696 121144 263702
rect 121092 263638 121144 263644
rect 121104 143070 121132 263638
rect 131212 263084 131264 263090
rect 131212 263026 131264 263032
rect 133696 263084 133748 263090
rect 133696 263026 133748 263032
rect 129740 262812 129792 262818
rect 129740 262754 129792 262760
rect 128452 262744 128504 262750
rect 127898 262712 127954 262721
rect 128452 262686 128504 262692
rect 127898 262647 127954 262656
rect 125140 262336 125192 262342
rect 125140 262278 125192 262284
rect 126242 262304 126298 262313
rect 121184 262268 121236 262274
rect 121184 262210 121236 262216
rect 121092 143064 121144 143070
rect 121092 143006 121144 143012
rect 120906 142831 120962 142840
rect 121000 142860 121052 142866
rect 121000 142802 121052 142808
rect 121196 142050 121224 262210
rect 123484 260092 123536 260098
rect 123484 260034 123536 260040
rect 123496 259894 123524 260034
rect 125152 259978 125180 262278
rect 126242 262239 126298 262248
rect 126980 262268 127032 262274
rect 126256 259978 126284 262239
rect 126980 262210 127032 262216
rect 126992 259978 127020 262210
rect 127912 259978 127940 262647
rect 128464 259978 128492 262686
rect 129752 259978 129780 262754
rect 130108 262404 130160 262410
rect 130108 262346 130160 262352
rect 130120 259978 130148 262346
rect 131120 261180 131172 261186
rect 131120 261122 131172 261128
rect 130660 260908 130712 260914
rect 130660 260850 130712 260856
rect 125152 259950 125488 259978
rect 126256 259950 126592 259978
rect 126992 259950 127144 259978
rect 127360 259962 127696 259978
rect 127348 259956 127696 259962
rect 127400 259950 127696 259956
rect 127912 259950 128248 259978
rect 128464 259950 128800 259978
rect 129752 259950 129904 259978
rect 130120 259950 130456 259978
rect 127348 259898 127400 259904
rect 123484 259888 123536 259894
rect 130672 259842 130700 260850
rect 131132 260302 131160 261122
rect 131120 260296 131172 260302
rect 131120 260238 131172 260244
rect 131224 259978 131252 263026
rect 132592 263016 132644 263022
rect 132592 262958 132644 262964
rect 132040 260296 132092 260302
rect 132040 260238 132092 260244
rect 132052 259978 132080 260238
rect 131224 259950 131560 259978
rect 132052 259950 132112 259978
rect 132604 259842 132632 262958
rect 133144 262880 133196 262886
rect 133144 262822 133196 262828
rect 133156 261322 133184 262822
rect 133708 262585 133736 263026
rect 133788 263016 133840 263022
rect 133788 262958 133840 262964
rect 133800 262818 133828 262958
rect 133788 262812 133840 262818
rect 133788 262754 133840 262760
rect 133326 262576 133382 262585
rect 133326 262511 133382 262520
rect 133694 262576 133750 262585
rect 133694 262511 133750 262520
rect 133144 261316 133196 261322
rect 133144 261258 133196 261264
rect 133340 259842 133368 262511
rect 133696 261316 133748 261322
rect 133696 261258 133748 261264
rect 133708 259978 133736 261258
rect 133984 259978 134012 264114
rect 135352 264036 135404 264042
rect 135352 263978 135404 263984
rect 135168 261112 135220 261118
rect 135168 261054 135220 261060
rect 135180 259978 135208 261054
rect 133708 259950 133768 259978
rect 133984 259950 134320 259978
rect 134872 259950 135208 259978
rect 135364 259978 135392 263978
rect 135548 259978 135576 324294
rect 135904 311908 135956 311914
rect 135904 311850 135956 311856
rect 135916 264994 135944 311850
rect 135996 298172 136048 298178
rect 135996 298114 136048 298120
rect 135904 264988 135956 264994
rect 135904 264930 135956 264936
rect 135916 263922 135944 264930
rect 136008 264042 136036 298114
rect 137284 282192 137336 282198
rect 137284 282134 137336 282140
rect 137192 264308 137244 264314
rect 137192 264250 137244 264256
rect 135996 264036 136048 264042
rect 135996 263978 136048 263984
rect 137100 264036 137152 264042
rect 137100 263978 137152 263984
rect 135916 263894 136128 263922
rect 136100 259978 136128 263894
rect 137112 263770 137140 263978
rect 137204 263770 137232 264250
rect 137296 263906 137324 282134
rect 137284 263900 137336 263906
rect 137284 263842 137336 263848
rect 137100 263764 137152 263770
rect 137100 263706 137152 263712
rect 137192 263764 137244 263770
rect 137192 263706 137244 263712
rect 135364 259950 135424 259978
rect 135548 259950 135976 259978
rect 136100 259950 136528 259978
rect 135548 259894 135576 259950
rect 123484 259830 123536 259836
rect 124232 259826 124384 259842
rect 124220 259820 124384 259826
rect 124272 259814 124384 259820
rect 130672 259814 131008 259842
rect 132604 259814 132664 259842
rect 133216 259814 133368 259842
rect 135536 259888 135588 259894
rect 137204 259842 137232 263706
rect 137296 259978 137324 263842
rect 138032 260817 138060 430578
rect 138664 404388 138716 404394
rect 138664 404330 138716 404336
rect 138676 264110 138704 404330
rect 140056 271182 140084 699654
rect 146576 696992 146628 696998
rect 146576 696934 146628 696940
rect 144920 643136 144972 643142
rect 144920 643078 144972 643084
rect 143724 590708 143776 590714
rect 143724 590650 143776 590656
rect 142160 536852 142212 536858
rect 142160 536794 142212 536800
rect 140136 418192 140188 418198
rect 140136 418134 140188 418140
rect 140044 271176 140096 271182
rect 140044 271118 140096 271124
rect 140148 265033 140176 418134
rect 140228 351960 140280 351966
rect 140228 351902 140280 351908
rect 140134 265024 140190 265033
rect 140134 264959 140190 264968
rect 139768 264376 139820 264382
rect 139768 264318 139820 264324
rect 138664 264104 138716 264110
rect 138664 264046 138716 264052
rect 138296 263560 138348 263566
rect 138296 263502 138348 263508
rect 138308 260953 138336 263502
rect 138294 260944 138350 260953
rect 138294 260879 138350 260888
rect 138018 260808 138074 260817
rect 138018 260743 138074 260752
rect 138032 260409 138060 260743
rect 138018 260400 138074 260409
rect 138018 260335 138074 260344
rect 137296 259950 137632 259978
rect 138308 259842 138336 260879
rect 138676 259978 138704 264046
rect 139780 263702 139808 264318
rect 139768 263696 139820 263702
rect 139768 263638 139820 263644
rect 138938 260808 138994 260817
rect 138938 260743 138994 260752
rect 138952 259978 138980 260743
rect 140148 259978 140176 264959
rect 140240 263770 140268 351902
rect 141424 283620 141476 283626
rect 141424 283562 141476 283568
rect 141056 267028 141108 267034
rect 141056 266970 141108 266976
rect 141068 264042 141096 266970
rect 141056 264036 141108 264042
rect 141056 263978 141108 263984
rect 140228 263764 140280 263770
rect 140228 263706 140280 263712
rect 140320 263696 140372 263702
rect 140320 263638 140372 263644
rect 138676 259950 138736 259978
rect 138952 259950 139288 259978
rect 139840 259950 140176 259978
rect 140332 259978 140360 263638
rect 140332 259950 140392 259978
rect 141068 259842 141096 263978
rect 141436 262449 141464 283562
rect 141608 265736 141660 265742
rect 141608 265678 141660 265684
rect 141620 263974 141648 265678
rect 141608 263968 141660 263974
rect 141608 263910 141660 263916
rect 141422 262440 141478 262449
rect 141422 262375 141478 262384
rect 141436 259978 141464 262375
rect 141620 259978 141648 263910
rect 142172 259978 142200 536794
rect 142252 524476 142304 524482
rect 142252 524418 142304 524424
rect 142264 260137 142292 524418
rect 143632 263832 143684 263838
rect 143632 263774 143684 263780
rect 142250 260128 142306 260137
rect 142250 260063 142306 260072
rect 143124 260128 143180 260137
rect 143124 260063 143180 260072
rect 141436 259950 141496 259978
rect 141620 259950 142048 259978
rect 142172 259950 142600 259978
rect 143138 259964 143166 260063
rect 143644 259978 143672 263774
rect 143736 260273 143764 590650
rect 143816 576904 143868 576910
rect 143816 576846 143868 576852
rect 143828 260817 143856 576846
rect 144184 563100 144236 563106
rect 144184 563042 144236 563048
rect 144196 263838 144224 563042
rect 144184 263832 144236 263838
rect 144184 263774 144236 263780
rect 143814 260808 143870 260817
rect 143814 260743 143870 260752
rect 144458 260808 144514 260817
rect 144458 260743 144514 260752
rect 143722 260264 143778 260273
rect 143722 260199 143778 260208
rect 143736 260114 143764 260199
rect 143736 260086 143856 260114
rect 143828 259978 143856 260086
rect 144472 259978 144500 260743
rect 144932 260273 144960 643078
rect 145564 616888 145616 616894
rect 145564 616830 145616 616836
rect 145576 264450 145604 616830
rect 145564 264444 145616 264450
rect 145564 264386 145616 264392
rect 144918 260264 144974 260273
rect 144918 260199 144974 260208
rect 144550 259992 144606 260001
rect 143644 259950 143704 259978
rect 143828 259950 144256 259978
rect 144472 259950 144550 259978
rect 135536 259830 135588 259836
rect 137080 259814 137232 259842
rect 138184 259814 138336 259842
rect 140944 259814 141096 259842
rect 142172 259826 142200 259950
rect 145576 259978 145604 264386
rect 146392 263220 146444 263226
rect 146392 263162 146444 263168
rect 146404 262682 146432 263162
rect 146392 262676 146444 262682
rect 146392 262618 146444 262624
rect 145884 260264 145940 260273
rect 145884 260199 145940 260208
rect 144606 259950 144808 259978
rect 145360 259950 145604 259978
rect 145898 259964 145926 260199
rect 144550 259927 144606 259936
rect 144564 259867 144592 259927
rect 146404 259842 146432 262618
rect 146588 260234 146616 696934
rect 148324 683188 148376 683194
rect 148324 683130 148376 683136
rect 146944 670744 146996 670750
rect 146944 670686 146996 670692
rect 146956 263809 146984 670686
rect 147036 630692 147088 630698
rect 147036 630634 147088 630640
rect 146942 263800 146998 263809
rect 146942 263735 146998 263744
rect 146576 260228 146628 260234
rect 146576 260170 146628 260176
rect 142160 259820 142212 259826
rect 124220 259762 124272 259768
rect 125690 259720 125746 259729
rect 125746 259678 126040 259706
rect 125690 259655 125746 259664
rect 130856 259593 130884 259814
rect 146404 259814 146464 259842
rect 142160 259762 142212 259768
rect 146588 259758 146616 260170
rect 146956 259978 146984 263735
rect 147048 263226 147076 630634
rect 147680 268388 147732 268394
rect 147680 268330 147732 268336
rect 147036 263220 147088 263226
rect 147036 263162 147088 263168
rect 147692 260234 147720 268330
rect 148336 262857 148364 683130
rect 149244 278044 149296 278050
rect 149244 277986 149296 277992
rect 149152 269816 149204 269822
rect 149152 269758 149204 269764
rect 149164 263634 149192 269758
rect 149152 263628 149204 263634
rect 149152 263570 149204 263576
rect 148322 262848 148378 262857
rect 148322 262783 148378 262792
rect 147542 260228 147594 260234
rect 147542 260170 147594 260176
rect 147680 260228 147732 260234
rect 147680 260170 147732 260176
rect 146956 259950 147016 259978
rect 147554 259964 147582 260170
rect 146576 259752 146628 259758
rect 146576 259694 146628 259700
rect 147692 259690 147720 260170
rect 148336 259978 148364 262783
rect 149256 260545 149284 277986
rect 149716 262546 149744 700266
rect 152464 501016 152516 501022
rect 152464 500958 152516 500964
rect 151820 280220 151872 280226
rect 151820 280162 151872 280168
rect 151084 279472 151136 279478
rect 151084 279414 151136 279420
rect 151096 263673 151124 279414
rect 151082 263664 151138 263673
rect 149980 263628 150032 263634
rect 151082 263599 151138 263608
rect 149980 263570 150032 263576
rect 149704 262540 149756 262546
rect 149704 262482 149756 262488
rect 149242 260536 149298 260545
rect 149242 260471 149298 260480
rect 149256 260250 149284 260471
rect 148646 260228 148698 260234
rect 148646 260170 148698 260176
rect 149210 260222 149284 260250
rect 148120 259950 148364 259978
rect 148658 259964 148686 260170
rect 149210 259964 149238 260222
rect 149716 259978 149744 262482
rect 149992 259978 150020 263570
rect 150438 262848 150494 262857
rect 150438 262783 150494 262792
rect 150452 262614 150480 262783
rect 150440 262608 150492 262614
rect 150440 262550 150492 262556
rect 151096 259978 151124 263599
rect 151832 263498 151860 280162
rect 152476 272542 152504 500958
rect 152464 272536 152516 272542
rect 152464 272478 152516 272484
rect 151910 270600 151966 270609
rect 151910 270535 151966 270544
rect 151820 263492 151872 263498
rect 151820 263434 151872 263440
rect 151358 262848 151414 262857
rect 151358 262783 151414 262792
rect 149716 259950 149776 259978
rect 149992 259950 150328 259978
rect 150880 259950 151124 259978
rect 151372 259978 151400 262783
rect 151924 259978 151952 270535
rect 152188 263492 152240 263498
rect 152188 263434 152240 263440
rect 152200 259978 152228 263434
rect 153014 262984 153070 262993
rect 153014 262919 153070 262928
rect 153028 259978 153056 262919
rect 153212 260234 153240 700334
rect 153304 265130 153332 702406
rect 157340 700732 157392 700738
rect 157340 700674 157392 700680
rect 157248 700528 157300 700534
rect 157248 700470 157300 700476
rect 154578 276040 154634 276049
rect 154578 275975 154634 275984
rect 153384 274712 153436 274718
rect 153384 274654 153436 274660
rect 153292 265124 153344 265130
rect 153292 265066 153344 265072
rect 153200 260228 153252 260234
rect 153200 260170 153252 260176
rect 151372 259950 151432 259978
rect 151924 259950 151984 259978
rect 152200 259950 152536 259978
rect 153028 259950 153088 259978
rect 147680 259684 147732 259690
rect 147680 259626 147732 259632
rect 153212 259622 153240 260170
rect 153396 259978 153424 274654
rect 154592 267734 154620 275975
rect 155960 273284 156012 273290
rect 155960 273226 156012 273232
rect 155972 267734 156000 273226
rect 154592 267706 155448 267734
rect 155972 267706 156552 267734
rect 155224 263628 155276 263634
rect 155224 263570 155276 263576
rect 155040 262540 155092 262546
rect 155040 262482 155092 262488
rect 154166 260228 154218 260234
rect 154166 260170 154218 260176
rect 153396 259950 153640 259978
rect 154178 259964 154206 260170
rect 155052 259978 155080 262482
rect 154744 259950 155080 259978
rect 155236 259978 155264 263570
rect 155420 259978 155448 267706
rect 156328 264988 156380 264994
rect 156328 264930 156380 264936
rect 156340 259978 156368 264930
rect 156524 259978 156552 267706
rect 157260 264994 157288 700470
rect 157248 264988 157300 264994
rect 157248 264930 157300 264936
rect 157352 260438 157380 700674
rect 160744 700664 160796 700670
rect 160744 700606 160796 700612
rect 160100 700596 160152 700602
rect 160100 700538 160152 700544
rect 157616 605124 157668 605130
rect 157616 605066 157668 605072
rect 157340 260432 157392 260438
rect 157340 260374 157392 260380
rect 157352 259978 157380 260374
rect 157628 260234 157656 605066
rect 158720 271176 158772 271182
rect 158720 271118 158772 271124
rect 158352 262608 158404 262614
rect 158352 262550 158404 262556
rect 157616 260228 157668 260234
rect 157616 260170 157668 260176
rect 158364 259978 158392 262550
rect 158582 260228 158634 260234
rect 158582 260170 158634 260176
rect 155236 259950 155296 259978
rect 155420 259950 155848 259978
rect 156340 259950 156400 259978
rect 156524 259950 156952 259978
rect 157352 259950 157504 259978
rect 158056 259950 158392 259978
rect 158594 259706 158622 260170
rect 158732 259978 158760 271118
rect 158812 265124 158864 265130
rect 158812 265066 158864 265072
rect 158824 264994 158852 265066
rect 158812 264988 158864 264994
rect 158812 264930 158864 264936
rect 159640 264988 159692 264994
rect 159640 264930 159692 264936
rect 159652 259978 159680 264930
rect 160112 260273 160140 700538
rect 160192 268456 160244 268462
rect 160192 268398 160244 268404
rect 160098 260264 160154 260273
rect 160098 260199 160154 260208
rect 160204 259978 160232 268398
rect 160756 265130 160784 700606
rect 162124 700460 162176 700466
rect 162124 700402 162176 700408
rect 161480 276684 161532 276690
rect 161480 276626 161532 276632
rect 160744 265124 160796 265130
rect 160744 265066 160796 265072
rect 161296 265124 161348 265130
rect 161296 265066 161348 265072
rect 160788 260264 160844 260273
rect 160788 260199 160844 260208
rect 158732 259950 159496 259978
rect 159652 259950 159712 259978
rect 160204 259950 160600 259978
rect 158720 259752 158772 259758
rect 158594 259700 158720 259706
rect 158594 259694 158772 259700
rect 158594 259692 158760 259694
rect 158608 259678 158760 259692
rect 159468 259690 159496 259950
rect 160572 259826 160600 259950
rect 160560 259820 160612 259826
rect 160560 259762 160612 259768
rect 160802 259706 160830 260199
rect 161308 259978 161336 265066
rect 161308 259950 161368 259978
rect 161492 259842 161520 276626
rect 162136 262449 162164 700402
rect 164884 670812 164936 670818
rect 164884 670754 164936 670760
rect 164240 632120 164292 632126
rect 164240 632062 164292 632068
rect 163504 284980 163556 284986
rect 163504 284922 163556 284928
rect 163516 267734 163544 284922
rect 163596 273964 163648 273970
rect 163596 273906 163648 273912
rect 163424 267706 163544 267734
rect 163608 267734 163636 273906
rect 163608 267706 163728 267734
rect 163424 265033 163452 267706
rect 163504 265668 163556 265674
rect 163504 265610 163556 265616
rect 163410 265024 163466 265033
rect 163410 264959 163466 264968
rect 162122 262440 162178 262449
rect 162122 262375 162178 262384
rect 162136 259978 162164 262375
rect 163424 259978 163452 264959
rect 163516 260273 163544 265610
rect 163700 262585 163728 267706
rect 163686 262576 163742 262585
rect 163686 262511 163742 262520
rect 163502 260264 163558 260273
rect 163502 260199 163558 260208
rect 162136 259950 162472 259978
rect 163024 259950 163452 259978
rect 163516 259978 163544 260199
rect 163700 259978 163728 262511
rect 164252 260001 164280 632062
rect 164896 265198 164924 670754
rect 166264 618316 166316 618322
rect 166264 618258 166316 618264
rect 165620 579692 165672 579698
rect 165620 579634 165672 579640
rect 164884 265192 164936 265198
rect 164884 265134 164936 265140
rect 164238 259992 164294 260001
rect 163516 259950 163576 259978
rect 163700 259950 164128 259978
rect 164896 259978 164924 265134
rect 165632 260234 165660 579634
rect 166276 265169 166304 618258
rect 166356 605872 166408 605878
rect 166356 605814 166408 605820
rect 166262 265160 166318 265169
rect 166262 265095 166318 265104
rect 166078 263256 166134 263265
rect 166078 263191 166134 263200
rect 166092 262721 166120 263191
rect 166078 262712 166134 262721
rect 166078 262647 166134 262656
rect 165620 260228 165672 260234
rect 165620 260170 165672 260176
rect 164680 259950 164924 259978
rect 165066 259992 165122 260001
rect 164238 259927 164294 259936
rect 166092 259978 166120 262647
rect 165122 259950 165232 259978
rect 165784 259950 166120 259978
rect 166276 259978 166304 265095
rect 166368 263265 166396 605814
rect 169772 605130 169800 702406
rect 202800 700738 202828 703520
rect 202788 700732 202840 700738
rect 202788 700674 202840 700680
rect 169760 605124 169812 605130
rect 169760 605066 169812 605072
rect 167644 565888 167696 565894
rect 167644 565830 167696 565836
rect 167656 265305 167684 565830
rect 167736 553444 167788 553450
rect 167736 553386 167788 553392
rect 167642 265296 167698 265305
rect 167642 265231 167698 265240
rect 166354 263256 166410 263265
rect 166354 263191 166410 263200
rect 167550 263120 167606 263129
rect 167550 263055 167606 263064
rect 166862 260228 166914 260234
rect 166862 260170 166914 260176
rect 166874 259978 166902 260170
rect 167564 259978 167592 263055
rect 166276 259950 166336 259978
rect 166874 259964 167040 259978
rect 166888 259950 167040 259964
rect 167440 259950 167592 259978
rect 167656 259978 167684 265231
rect 167748 263129 167776 553386
rect 180064 510672 180116 510678
rect 180064 510614 180116 510620
rect 169760 474768 169812 474774
rect 169760 474710 169812 474716
rect 169116 275324 169168 275330
rect 169116 275266 169168 275272
rect 169024 272536 169076 272542
rect 169024 272478 169076 272484
rect 168380 264240 168432 264246
rect 168380 264182 168432 264188
rect 168392 263702 168420 264182
rect 168380 263696 168432 263702
rect 168380 263638 168432 263644
rect 167734 263120 167790 263129
rect 167734 263055 167790 263064
rect 168392 259978 168420 263638
rect 169036 262682 169064 272478
rect 169128 265334 169156 275266
rect 169116 265328 169168 265334
rect 169116 265270 169168 265276
rect 169576 265328 169628 265334
rect 169576 265270 169628 265276
rect 169024 262676 169076 262682
rect 169024 262618 169076 262624
rect 169036 259978 169064 262618
rect 169588 259978 169616 265270
rect 169772 259978 169800 474710
rect 171784 462392 171836 462398
rect 171784 462334 171836 462340
rect 170404 448588 170456 448594
rect 170404 448530 170456 448536
rect 170416 262750 170444 448530
rect 171140 422340 171192 422346
rect 171140 422282 171192 422288
rect 170404 262744 170456 262750
rect 170404 262686 170456 262692
rect 170174 260228 170226 260234
rect 170174 260170 170226 260176
rect 170186 259978 170214 260170
rect 167656 259950 167992 259978
rect 168392 259950 168544 259978
rect 169036 259950 169096 259978
rect 169588 259950 169648 259978
rect 169772 259964 170214 259978
rect 170416 259978 170444 262686
rect 171046 260264 171102 260273
rect 171046 260199 171102 260208
rect 171060 260001 171088 260199
rect 171152 260166 171180 422282
rect 171796 267734 171824 462334
rect 178684 456816 178736 456822
rect 178684 456758 178736 456764
rect 171876 397520 171928 397526
rect 171876 397462 171928 397468
rect 171704 267706 171824 267734
rect 171888 267734 171916 397462
rect 174544 357468 174596 357474
rect 174544 357410 174596 357416
rect 173900 345092 173952 345098
rect 173900 345034 173952 345040
rect 173164 286340 173216 286346
rect 173164 286282 173216 286288
rect 172520 269884 172572 269890
rect 172520 269826 172572 269832
rect 171888 267706 172008 267734
rect 171704 265810 171732 267706
rect 171692 265804 171744 265810
rect 171692 265746 171744 265752
rect 171140 260160 171192 260166
rect 171140 260102 171192 260108
rect 171046 259992 171102 260001
rect 169772 259950 170200 259964
rect 170416 259950 170752 259978
rect 165066 259927 165122 259936
rect 167012 259894 167040 259950
rect 171704 259978 171732 265746
rect 171980 265538 172008 267706
rect 171968 265532 172020 265538
rect 171968 265474 172020 265480
rect 171830 260160 171882 260166
rect 171830 260102 171882 260108
rect 171304 259950 171732 259978
rect 171842 259964 171870 260102
rect 171980 259978 172008 265474
rect 172532 260166 172560 269826
rect 173176 265470 173204 286282
rect 173164 265464 173216 265470
rect 173164 265406 173216 265412
rect 172520 260160 172572 260166
rect 172520 260102 172572 260108
rect 173176 259978 173204 265406
rect 173486 260160 173538 260166
rect 173486 260102 173538 260108
rect 171980 259950 172408 259978
rect 172960 259950 173204 259978
rect 173498 259964 173526 260102
rect 173912 259978 173940 345034
rect 173992 318844 174044 318850
rect 173992 318786 174044 318792
rect 174004 260166 174032 318786
rect 174556 265402 174584 357410
rect 175924 305040 175976 305046
rect 175924 304982 175976 304988
rect 175936 265606 175964 304982
rect 176016 292596 176068 292602
rect 176016 292538 176068 292544
rect 176028 265674 176056 292538
rect 176660 266416 176712 266422
rect 176660 266358 176712 266364
rect 176108 265804 176160 265810
rect 176108 265746 176160 265752
rect 176016 265668 176068 265674
rect 176016 265610 176068 265616
rect 175924 265600 175976 265606
rect 175924 265542 175976 265548
rect 174544 265396 174596 265402
rect 174544 265338 174596 265344
rect 173992 260160 174044 260166
rect 173992 260102 174044 260108
rect 174556 259978 174584 265338
rect 175832 265260 175884 265266
rect 175832 265202 175884 265208
rect 175188 260500 175240 260506
rect 175188 260442 175240 260448
rect 175200 260250 175228 260442
rect 175154 260222 175228 260250
rect 175154 260166 175182 260222
rect 175142 260160 175194 260166
rect 175142 260102 175194 260108
rect 173912 259950 174400 259978
rect 174556 259950 174616 259978
rect 175154 259964 175182 260102
rect 175844 259978 175872 265202
rect 175720 259950 175872 259978
rect 175936 259978 175964 265542
rect 176028 265266 176056 265610
rect 176120 265266 176148 265746
rect 176016 265260 176068 265266
rect 176016 265202 176068 265208
rect 176108 265260 176160 265266
rect 176108 265202 176160 265208
rect 176672 263770 176700 266358
rect 178696 264314 178724 456758
rect 180076 265742 180104 510614
rect 181444 484424 181496 484430
rect 181444 484366 181496 484372
rect 181456 267034 181484 484366
rect 192484 470620 192536 470626
rect 192484 470562 192536 470568
rect 185584 378208 185636 378214
rect 185584 378150 185636 378156
rect 185596 282198 185624 378150
rect 192496 283626 192524 470562
rect 192484 283620 192536 283626
rect 192484 283562 192536 283568
rect 185584 282192 185636 282198
rect 185584 282134 185636 282140
rect 186412 280832 186464 280838
rect 186412 280774 186464 280780
rect 186424 280226 186452 280774
rect 186412 280220 186464 280226
rect 186412 280162 186464 280168
rect 181444 267028 181496 267034
rect 181444 266970 181496 266976
rect 180064 265736 180116 265742
rect 180064 265678 180116 265684
rect 178684 264308 178736 264314
rect 178684 264250 178736 264256
rect 176660 263764 176712 263770
rect 176660 263706 176712 263712
rect 176672 259978 176700 263706
rect 178776 262948 178828 262954
rect 178776 262890 178828 262896
rect 180432 262948 180484 262954
rect 180432 262890 180484 262896
rect 178132 262880 178184 262886
rect 178132 262822 178184 262828
rect 177764 262472 177816 262478
rect 177764 262414 177816 262420
rect 177776 260982 177804 262414
rect 178144 261254 178172 262822
rect 178132 261248 178184 261254
rect 178132 261190 178184 261196
rect 177764 260976 177816 260982
rect 177764 260918 177816 260924
rect 177028 260364 177080 260370
rect 177028 260306 177080 260312
rect 177040 259978 177068 260306
rect 177776 259978 177804 260918
rect 178144 259978 178172 261190
rect 178684 261180 178736 261186
rect 178684 261122 178736 261128
rect 178696 261050 178724 261122
rect 178788 261050 178816 262890
rect 178684 261044 178736 261050
rect 178684 260986 178736 260992
rect 178776 261044 178828 261050
rect 178776 260986 178828 260992
rect 179512 261044 179564 261050
rect 179512 260986 179564 260992
rect 178696 259978 178724 260986
rect 179524 259978 179552 260986
rect 180444 259978 180472 262890
rect 180616 262472 180668 262478
rect 180616 262414 180668 262420
rect 175936 259950 176272 259978
rect 176672 259950 176824 259978
rect 177040 259950 177712 259978
rect 177776 259950 177928 259978
rect 178144 259950 178480 259978
rect 178696 259950 179032 259978
rect 179524 259950 179584 259978
rect 180136 259950 180472 259978
rect 180628 259978 180656 262414
rect 183192 262404 183244 262410
rect 183192 262346 183244 262352
rect 182088 262268 182140 262274
rect 182088 262210 182140 262216
rect 181536 261384 181588 261390
rect 181536 261326 181588 261332
rect 180890 260264 180946 260273
rect 180890 260199 180946 260208
rect 180628 259950 180688 259978
rect 171046 259927 171102 259936
rect 167000 259888 167052 259894
rect 162122 259856 162178 259865
rect 161492 259814 162122 259842
rect 167000 259830 167052 259836
rect 162122 259791 162178 259800
rect 160926 259720 160982 259729
rect 160802 259692 160926 259706
rect 159456 259684 159508 259690
rect 160816 259678 160926 259692
rect 160926 259655 160982 259664
rect 159456 259626 159508 259632
rect 174372 259622 174400 259950
rect 153200 259616 153252 259622
rect 130842 259584 130898 259593
rect 123496 259542 123832 259570
rect 124600 259554 124936 259570
rect 124588 259548 124936 259554
rect 123496 259418 123524 259542
rect 124640 259542 124936 259548
rect 129016 259542 129352 259570
rect 124588 259490 124640 259496
rect 129016 259486 129044 259542
rect 153200 259558 153252 259564
rect 174360 259616 174412 259622
rect 174360 259558 174412 259564
rect 177684 259554 177712 259950
rect 180904 259729 180932 260199
rect 181548 259978 181576 261326
rect 182100 259978 182128 262210
rect 182640 260364 182692 260370
rect 182640 260306 182692 260312
rect 182652 259978 182680 260306
rect 183204 259978 183232 262346
rect 184848 260908 184900 260914
rect 184848 260850 184900 260856
rect 184860 259978 184888 260850
rect 181240 259950 181576 259978
rect 181792 259950 182128 259978
rect 182344 259950 182680 259978
rect 182896 259950 183232 259978
rect 184552 259950 184888 259978
rect 184940 260024 184992 260030
rect 184940 259966 184992 259972
rect 180890 259720 180946 259729
rect 180890 259655 180946 259664
rect 184952 259622 184980 259966
rect 184940 259616 184992 259622
rect 130842 259519 130898 259528
rect 177672 259548 177724 259554
rect 184000 259542 184336 259570
rect 185398 259584 185454 259593
rect 184940 259558 184992 259564
rect 185104 259554 185348 259570
rect 185104 259548 185360 259554
rect 185104 259542 185308 259548
rect 177672 259490 177724 259496
rect 184308 259486 184336 259542
rect 186042 259584 186098 259593
rect 185454 259542 185656 259570
rect 185398 259519 185454 259528
rect 186098 259542 186208 259570
rect 186042 259519 186098 259528
rect 185308 259490 185360 259496
rect 129004 259480 129056 259486
rect 129004 259422 129056 259428
rect 184296 259480 184348 259486
rect 184296 259422 184348 259428
rect 123484 259412 123536 259418
rect 123484 259354 123536 259360
rect 183652 259344 183704 259350
rect 183448 259292 183652 259298
rect 183448 259286 183704 259292
rect 183448 259270 183692 259286
rect 131304 199912 131356 199918
rect 132040 199912 132092 199918
rect 131304 199854 131356 199860
rect 131670 199880 131726 199889
rect 123482 199744 123538 199753
rect 123482 199679 123538 199688
rect 122748 198280 122800 198286
rect 122748 198222 122800 198228
rect 122104 191412 122156 191418
rect 122104 191354 122156 191360
rect 121368 185360 121420 185366
rect 121368 185302 121420 185308
rect 121276 183796 121328 183802
rect 121276 183738 121328 183744
rect 121184 142044 121236 142050
rect 121184 141986 121236 141992
rect 120816 141976 120868 141982
rect 120816 141918 120868 141924
rect 121184 141432 121236 141438
rect 121184 141374 121236 141380
rect 120816 140616 120868 140622
rect 120816 140558 120868 140564
rect 120828 136338 120856 140558
rect 120908 140344 120960 140350
rect 120908 140286 120960 140292
rect 120816 136332 120868 136338
rect 120816 136274 120868 136280
rect 120920 80918 120948 140286
rect 121000 139732 121052 139738
rect 121000 139674 121052 139680
rect 120908 80912 120960 80918
rect 120908 80854 120960 80860
rect 120722 79520 120778 79529
rect 120722 79455 120778 79464
rect 120540 76900 120592 76906
rect 120540 76842 120592 76848
rect 120724 75608 120776 75614
rect 120724 75550 120776 75556
rect 120736 75478 120764 75550
rect 120724 75472 120776 75478
rect 121012 75449 121040 139674
rect 121092 79620 121144 79626
rect 121092 79562 121144 79568
rect 121104 78878 121132 79562
rect 121092 78872 121144 78878
rect 121092 78814 121144 78820
rect 120724 75414 120776 75420
rect 120998 75440 121054 75449
rect 120998 75375 121054 75384
rect 119986 72992 120042 73001
rect 119986 72927 120042 72936
rect 119894 72856 119950 72865
rect 119894 72791 119950 72800
rect 119804 72684 119856 72690
rect 119804 72626 119856 72632
rect 118516 68944 118568 68950
rect 118516 68886 118568 68892
rect 115846 68640 115902 68649
rect 115846 68575 115902 68584
rect 120080 68468 120132 68474
rect 120080 68410 120132 68416
rect 117320 68400 117372 68406
rect 115938 68368 115994 68377
rect 117320 68342 117372 68348
rect 115938 68303 115994 68312
rect 115020 59900 115072 59906
rect 115020 59842 115072 59848
rect 115952 16574 115980 68303
rect 111812 16546 112392 16574
rect 113192 16546 114048 16574
rect 114572 16546 114784 16574
rect 115952 16546 116440 16574
rect 111616 3800 111668 3806
rect 111616 3742 111668 3748
rect 111156 3392 111208 3398
rect 111156 3334 111208 3340
rect 111628 480 111656 3742
rect 106894 354 107006 480
rect 106476 326 107006 354
rect 106894 -960 107006 326
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112364 354 112392 16546
rect 114020 480 114048 16546
rect 112782 354 112894 480
rect 112364 326 112894 354
rect 112782 -960 112894 326
rect 113978 -960 114090 480
rect 114756 354 114784 16546
rect 116412 480 116440 16546
rect 115174 354 115286 480
rect 114756 326 115286 354
rect 115174 -960 115286 326
rect 116370 -960 116482 480
rect 117332 354 117360 68342
rect 120092 16574 120120 68410
rect 121012 64874 121040 75375
rect 121196 71602 121224 141374
rect 121288 75138 121316 183738
rect 121276 75132 121328 75138
rect 121276 75074 121328 75080
rect 121380 74526 121408 185302
rect 122116 139466 122144 191354
rect 122380 149048 122432 149054
rect 122380 148990 122432 148996
rect 122196 148164 122248 148170
rect 122196 148106 122248 148112
rect 122104 139460 122156 139466
rect 122104 139402 122156 139408
rect 121920 139392 121972 139398
rect 121918 139360 121920 139369
rect 121972 139360 121974 139369
rect 121918 139295 121974 139304
rect 122208 139233 122236 148106
rect 122194 139224 122250 139233
rect 122194 139159 122250 139168
rect 122392 138553 122420 148990
rect 122760 139369 122788 198222
rect 123496 140729 123524 199679
rect 131316 199617 131344 199854
rect 132374 199900 132402 200124
rect 132040 199854 132092 199860
rect 132144 199872 132402 199900
rect 131670 199815 131726 199824
rect 131948 199844 132000 199850
rect 131684 199714 131712 199815
rect 131948 199786 132000 199792
rect 131672 199708 131724 199714
rect 131672 199650 131724 199656
rect 131302 199608 131358 199617
rect 131302 199543 131358 199552
rect 126244 198824 126296 198830
rect 126244 198766 126296 198772
rect 125048 192296 125100 192302
rect 125048 192238 125100 192244
rect 123576 190936 123628 190942
rect 123576 190878 123628 190884
rect 123482 140720 123538 140729
rect 123482 140655 123538 140664
rect 123588 140010 123616 190878
rect 124128 186924 124180 186930
rect 124128 186866 124180 186872
rect 123666 148472 123722 148481
rect 123666 148407 123722 148416
rect 123576 140004 123628 140010
rect 123576 139946 123628 139952
rect 123680 139398 123708 148407
rect 123944 148300 123996 148306
rect 123944 148242 123996 148248
rect 123760 141976 123812 141982
rect 123760 141918 123812 141924
rect 123772 139890 123800 141918
rect 123772 139876 123832 139890
rect 123772 139862 123846 139876
rect 123818 139482 123846 139862
rect 123956 139670 123984 148242
rect 123944 139664 123996 139670
rect 123944 139606 123996 139612
rect 123818 139468 124076 139482
rect 123832 139466 124076 139468
rect 123832 139460 124088 139466
rect 123832 139454 124036 139460
rect 124036 139402 124088 139408
rect 123668 139392 123720 139398
rect 122746 139360 122802 139369
rect 122746 139295 122802 139304
rect 122930 139360 122986 139369
rect 124140 139369 124168 186866
rect 124220 142180 124272 142186
rect 124220 142122 124272 142128
rect 124232 141137 124260 142122
rect 124588 141840 124640 141846
rect 124588 141782 124640 141788
rect 124218 141128 124274 141137
rect 124218 141063 124274 141072
rect 124232 139890 124260 141063
rect 124232 139862 124384 139890
rect 124600 139754 124628 141782
rect 124600 139726 124936 139754
rect 125060 139738 125088 192238
rect 125598 143440 125654 143449
rect 125598 143375 125654 143384
rect 125612 142254 125640 143375
rect 125690 142624 125746 142633
rect 125690 142559 125746 142568
rect 125600 142248 125652 142254
rect 125600 142190 125652 142196
rect 125140 141908 125192 141914
rect 125140 141850 125192 141856
rect 125152 141001 125180 141850
rect 125138 140992 125194 141001
rect 125138 140927 125194 140936
rect 125152 139890 125180 140927
rect 125704 139890 125732 142559
rect 126256 140554 126284 198766
rect 131026 198520 131082 198529
rect 131026 198455 131082 198464
rect 129648 197940 129700 197946
rect 129648 197882 129700 197888
rect 128268 194744 128320 194750
rect 128268 194686 128320 194692
rect 127900 194540 127952 194546
rect 127900 194482 127952 194488
rect 127716 190732 127768 190738
rect 127716 190674 127768 190680
rect 126336 188896 126388 188902
rect 126336 188838 126388 188844
rect 126244 140548 126296 140554
rect 126244 140490 126296 140496
rect 126348 140418 126376 188838
rect 127624 188012 127676 188018
rect 127624 187954 127676 187960
rect 126888 184340 126940 184346
rect 126888 184282 126940 184288
rect 126520 142248 126572 142254
rect 126520 142190 126572 142196
rect 126336 140412 126388 140418
rect 126336 140354 126388 140360
rect 126532 139890 126560 142190
rect 125152 139862 125488 139890
rect 125704 139862 126192 139890
rect 126532 139862 126592 139890
rect 125048 139732 125100 139738
rect 124876 139482 124904 139726
rect 125048 139674 125100 139680
rect 126164 139602 126192 139862
rect 126152 139596 126204 139602
rect 126152 139538 126204 139544
rect 125048 139528 125100 139534
rect 124876 139476 125048 139482
rect 124876 139470 125100 139476
rect 124876 139454 125088 139470
rect 126900 139369 126928 184282
rect 127636 147674 127664 187954
rect 127544 147646 127664 147674
rect 126978 145888 127034 145897
rect 126978 145823 127034 145832
rect 126992 142225 127020 145823
rect 126978 142216 127034 142225
rect 126978 142151 127034 142160
rect 127072 142044 127124 142050
rect 127072 141986 127124 141992
rect 126980 141704 127032 141710
rect 126980 141646 127032 141652
rect 126992 140826 127020 141646
rect 127084 140962 127112 141986
rect 127072 140956 127124 140962
rect 127072 140898 127124 140904
rect 126980 140820 127032 140826
rect 126980 140762 127032 140768
rect 127084 139890 127112 140898
rect 127544 140690 127572 147646
rect 127624 140820 127676 140826
rect 127624 140762 127676 140768
rect 127532 140684 127584 140690
rect 127532 140626 127584 140632
rect 127636 139890 127664 140762
rect 127728 140622 127756 190674
rect 127808 185156 127860 185162
rect 127808 185098 127860 185104
rect 127820 140758 127848 185098
rect 127912 142730 127940 194482
rect 128280 193730 128308 194686
rect 128268 193724 128320 193730
rect 128268 193666 128320 193672
rect 129004 180396 129056 180402
rect 129004 180338 129056 180344
rect 129016 144770 129044 180338
rect 129556 145444 129608 145450
rect 129556 145386 129608 145392
rect 129004 144764 129056 144770
rect 129004 144706 129056 144712
rect 129568 143546 129596 145386
rect 129556 143540 129608 143546
rect 129556 143482 129608 143488
rect 127900 142724 127952 142730
rect 127900 142666 127952 142672
rect 128174 142216 128230 142225
rect 128174 142151 128230 142160
rect 127808 140752 127860 140758
rect 127808 140694 127860 140700
rect 127716 140616 127768 140622
rect 127716 140558 127768 140564
rect 128188 139890 128216 142151
rect 129004 141772 129056 141778
rect 129004 141714 129056 141720
rect 129016 140894 129044 141714
rect 129004 140888 129056 140894
rect 129004 140830 129056 140836
rect 129016 139890 129044 140830
rect 129568 139890 129596 143482
rect 127084 139862 127144 139890
rect 127636 139862 127696 139890
rect 128188 139862 128248 139890
rect 128800 139862 129044 139890
rect 129352 139862 129596 139890
rect 129660 139369 129688 197882
rect 131040 196790 131068 198455
rect 131960 198014 131988 199786
rect 132052 198082 132080 199854
rect 132040 198076 132092 198082
rect 132040 198018 132092 198024
rect 131948 198008 132000 198014
rect 131948 197950 132000 197956
rect 131028 196784 131080 196790
rect 131028 196726 131080 196732
rect 131948 193724 132000 193730
rect 131948 193666 132000 193672
rect 130476 193656 130528 193662
rect 130476 193598 130528 193604
rect 130384 187468 130436 187474
rect 130384 187410 130436 187416
rect 130200 147008 130252 147014
rect 130200 146950 130252 146956
rect 130212 146334 130240 146950
rect 130200 146328 130252 146334
rect 130200 146270 130252 146276
rect 130212 144242 130240 146270
rect 130396 144838 130424 187410
rect 130488 144906 130516 193598
rect 131764 191004 131816 191010
rect 131764 190946 131816 190952
rect 130752 146192 130804 146198
rect 130752 146134 130804 146140
rect 130568 145512 130620 145518
rect 130568 145454 130620 145460
rect 130476 144900 130528 144906
rect 130476 144842 130528 144848
rect 130384 144832 130436 144838
rect 130384 144774 130436 144780
rect 130028 144214 130240 144242
rect 130028 139890 130056 144214
rect 130108 143404 130160 143410
rect 130108 143346 130160 143352
rect 129904 139862 130056 139890
rect 130120 139890 130148 143346
rect 130580 142526 130608 145454
rect 130568 142520 130620 142526
rect 130568 142462 130620 142468
rect 130658 141944 130714 141953
rect 130658 141879 130714 141888
rect 130672 141681 130700 141879
rect 130658 141672 130714 141681
rect 130658 141607 130714 141616
rect 130764 139890 130792 146134
rect 131776 146062 131804 190946
rect 131856 188964 131908 188970
rect 131856 188906 131908 188912
rect 131028 146056 131080 146062
rect 131028 145998 131080 146004
rect 131764 146056 131816 146062
rect 131764 145998 131816 146004
rect 131040 142730 131068 145998
rect 131868 145874 131896 188906
rect 131684 145846 131896 145874
rect 131488 144220 131540 144226
rect 131488 144162 131540 144168
rect 131028 142724 131080 142730
rect 131028 142666 131080 142672
rect 130120 139862 130456 139890
rect 130764 139862 131008 139890
rect 131500 139754 131528 144162
rect 131684 141574 131712 145846
rect 131854 145752 131910 145761
rect 131854 145687 131910 145696
rect 131868 143342 131896 145687
rect 131856 143336 131908 143342
rect 131856 143278 131908 143284
rect 131672 141568 131724 141574
rect 131672 141510 131724 141516
rect 131960 140026 131988 193666
rect 132144 185745 132172 199872
rect 132466 199832 132494 200124
rect 132558 199918 132586 200124
rect 132546 199912 132598 199918
rect 132546 199854 132598 199860
rect 132374 199804 132494 199832
rect 132374 199730 132402 199804
rect 132374 199702 132448 199730
rect 132316 198552 132368 198558
rect 132316 198494 132368 198500
rect 132328 197849 132356 198494
rect 132314 197840 132370 197849
rect 132314 197775 132370 197784
rect 132130 185736 132186 185745
rect 132130 185671 132186 185680
rect 132420 185609 132448 199702
rect 132650 199628 132678 200124
rect 132742 199923 132770 200124
rect 132728 199914 132784 199923
rect 132728 199849 132784 199858
rect 132834 199850 132862 200124
rect 132926 199923 132954 200124
rect 132912 199914 132968 199923
rect 132822 199844 132874 199850
rect 132912 199849 132968 199858
rect 132822 199786 132874 199792
rect 133018 199696 133046 200124
rect 132604 199600 132678 199628
rect 132972 199668 133046 199696
rect 132500 198076 132552 198082
rect 132500 198018 132552 198024
rect 132406 185600 132462 185609
rect 132406 185535 132462 185544
rect 132512 185230 132540 198018
rect 132500 185224 132552 185230
rect 132500 185166 132552 185172
rect 132604 181626 132632 199600
rect 132868 198008 132920 198014
rect 132774 197976 132830 197985
rect 132868 197950 132920 197956
rect 132774 197911 132830 197920
rect 132788 185745 132816 197911
rect 132880 186153 132908 197950
rect 132866 186144 132922 186153
rect 132866 186079 132922 186088
rect 132774 185736 132830 185745
rect 132774 185671 132830 185680
rect 132866 185328 132922 185337
rect 132866 185263 132922 185272
rect 132592 181620 132644 181626
rect 132592 181562 132644 181568
rect 132592 181484 132644 181490
rect 132592 181426 132644 181432
rect 132604 148345 132632 181426
rect 132684 174140 132736 174146
rect 132684 174082 132736 174088
rect 132696 148782 132724 174082
rect 132880 148850 132908 185263
rect 132972 176458 133000 199668
rect 133110 199628 133138 200124
rect 133064 199600 133138 199628
rect 133064 181490 133092 199600
rect 133202 199594 133230 200124
rect 133294 199696 133322 200124
rect 133386 199764 133414 200124
rect 133478 199923 133506 200124
rect 133464 199914 133520 199923
rect 133464 199849 133520 199858
rect 133386 199736 133460 199764
rect 133294 199668 133368 199696
rect 133202 199566 133276 199594
rect 133248 185201 133276 199566
rect 133234 185192 133290 185201
rect 133234 185127 133290 185136
rect 133340 182578 133368 199668
rect 133432 199646 133460 199736
rect 133420 199640 133472 199646
rect 133570 199628 133598 200124
rect 133662 199782 133690 200124
rect 133754 199782 133782 200124
rect 133846 199850 133874 200124
rect 133938 199923 133966 200124
rect 133924 199914 133980 199923
rect 133834 199844 133886 199850
rect 133924 199849 133980 199858
rect 134030 199850 134058 200124
rect 134122 199918 134150 200124
rect 134110 199912 134162 199918
rect 134110 199854 134162 199860
rect 133834 199786 133886 199792
rect 134018 199844 134070 199850
rect 134018 199786 134070 199792
rect 133650 199776 133702 199782
rect 133650 199718 133702 199724
rect 133742 199776 133794 199782
rect 134214 199764 134242 200124
rect 134306 199918 134334 200124
rect 134294 199912 134346 199918
rect 134398 199889 134426 200124
rect 134294 199854 134346 199860
rect 134384 199880 134440 199889
rect 134384 199815 134440 199824
rect 134490 199764 134518 200124
rect 134214 199736 134288 199764
rect 133742 199718 133794 199724
rect 134064 199708 134116 199714
rect 134064 199650 134116 199656
rect 133788 199640 133840 199646
rect 133570 199600 133736 199628
rect 133420 199582 133472 199588
rect 133604 199504 133656 199510
rect 133604 199446 133656 199452
rect 133510 197976 133566 197985
rect 133510 197911 133566 197920
rect 133328 182572 133380 182578
rect 133328 182514 133380 182520
rect 133052 181484 133104 181490
rect 133052 181426 133104 181432
rect 132960 176452 133012 176458
rect 132960 176394 133012 176400
rect 133524 174146 133552 197911
rect 133616 189854 133644 199446
rect 133604 189848 133656 189854
rect 133604 189790 133656 189796
rect 133708 185609 133736 199600
rect 133788 199582 133840 199588
rect 133800 190194 133828 199582
rect 133880 199572 133932 199578
rect 133880 199514 133932 199520
rect 133892 198393 133920 199514
rect 133970 199336 134026 199345
rect 133970 199271 134026 199280
rect 133878 198384 133934 198393
rect 133878 198319 133934 198328
rect 133984 198098 134012 199271
rect 133892 198070 134012 198098
rect 133788 190188 133840 190194
rect 133788 190130 133840 190136
rect 133892 185745 133920 198070
rect 133972 197804 134024 197810
rect 133972 197746 134024 197752
rect 133984 189922 134012 197746
rect 133972 189916 134024 189922
rect 133972 189858 134024 189864
rect 133878 185736 133934 185745
rect 133878 185671 133934 185680
rect 133694 185600 133750 185609
rect 133694 185535 133750 185544
rect 134076 184210 134104 199650
rect 134154 197704 134210 197713
rect 134154 197639 134210 197648
rect 134168 194594 134196 197639
rect 134260 197577 134288 199736
rect 134444 199736 134518 199764
rect 134340 199504 134392 199510
rect 134340 199446 134392 199452
rect 134352 198393 134380 199446
rect 134338 198384 134394 198393
rect 134338 198319 134394 198328
rect 134338 197976 134394 197985
rect 134338 197911 134394 197920
rect 134246 197568 134302 197577
rect 134246 197503 134302 197512
rect 134168 194566 134288 194594
rect 134260 185774 134288 194566
rect 134352 191282 134380 197911
rect 134444 197810 134472 199736
rect 134582 199696 134610 200124
rect 134674 199764 134702 200124
rect 134766 199923 134794 200124
rect 134752 199914 134808 199923
rect 134752 199849 134808 199858
rect 134858 199782 134886 200124
rect 134846 199776 134898 199782
rect 134674 199736 134748 199764
rect 134536 199668 134610 199696
rect 134536 197849 134564 199668
rect 134522 197840 134578 197849
rect 134432 197804 134484 197810
rect 134522 197775 134578 197784
rect 134432 197746 134484 197752
rect 134524 197532 134576 197538
rect 134524 197474 134576 197480
rect 134340 191276 134392 191282
rect 134340 191218 134392 191224
rect 134338 186144 134394 186153
rect 134338 186079 134394 186088
rect 134248 185768 134300 185774
rect 134248 185710 134300 185716
rect 134246 185600 134302 185609
rect 134246 185535 134302 185544
rect 134064 184204 134116 184210
rect 134064 184146 134116 184152
rect 133512 174140 133564 174146
rect 133512 174082 133564 174088
rect 132868 148844 132920 148850
rect 132868 148786 132920 148792
rect 132684 148776 132736 148782
rect 132684 148718 132736 148724
rect 134260 148510 134288 185535
rect 134248 148504 134300 148510
rect 134248 148446 134300 148452
rect 134352 148374 134380 186079
rect 134536 185638 134564 197474
rect 134720 195974 134748 199736
rect 134846 199718 134898 199724
rect 134950 199628 134978 200124
rect 135042 199918 135070 200124
rect 135134 199923 135162 200124
rect 135030 199912 135082 199918
rect 135030 199854 135082 199860
rect 135120 199914 135176 199923
rect 135226 199918 135254 200124
rect 135318 199923 135346 200124
rect 135120 199849 135176 199858
rect 135214 199912 135266 199918
rect 135214 199854 135266 199860
rect 135304 199914 135360 199923
rect 135304 199849 135360 199858
rect 135410 199850 135438 200124
rect 135502 199918 135530 200124
rect 135594 199918 135622 200124
rect 135686 199918 135714 200124
rect 135490 199912 135542 199918
rect 135490 199854 135542 199860
rect 135582 199912 135634 199918
rect 135582 199854 135634 199860
rect 135674 199912 135726 199918
rect 135674 199854 135726 199860
rect 135778 199850 135806 200124
rect 135870 199923 135898 200124
rect 135856 199914 135912 199923
rect 135962 199918 135990 200124
rect 135398 199844 135450 199850
rect 135398 199786 135450 199792
rect 135766 199844 135818 199850
rect 135856 199849 135912 199858
rect 135950 199912 136002 199918
rect 135950 199854 136002 199860
rect 135766 199786 135818 199792
rect 135260 199776 135312 199782
rect 135180 199736 135260 199764
rect 134904 199600 134978 199628
rect 135076 199640 135128 199646
rect 134798 197840 134854 197849
rect 134798 197775 134854 197784
rect 134628 195946 134748 195974
rect 134524 185632 134576 185638
rect 134524 185574 134576 185580
rect 134628 177002 134656 195946
rect 134812 190126 134840 197775
rect 134904 197538 134932 199600
rect 135076 199582 135128 199588
rect 134982 198384 135038 198393
rect 134982 198319 135038 198328
rect 134892 197532 134944 197538
rect 134892 197474 134944 197480
rect 134800 190120 134852 190126
rect 134800 190062 134852 190068
rect 134996 185609 135024 198319
rect 134982 185600 135038 185609
rect 134982 185535 135038 185544
rect 135088 185473 135116 199582
rect 135180 185570 135208 199736
rect 135260 199718 135312 199724
rect 136054 199730 136082 200124
rect 136146 199850 136174 200124
rect 136238 199850 136266 200124
rect 136330 199850 136358 200124
rect 136422 199918 136450 200124
rect 136514 199918 136542 200124
rect 136606 199923 136634 200124
rect 136410 199912 136462 199918
rect 136410 199854 136462 199860
rect 136502 199912 136554 199918
rect 136502 199854 136554 199860
rect 136592 199914 136648 199923
rect 136134 199844 136186 199850
rect 136134 199786 136186 199792
rect 136226 199844 136278 199850
rect 136226 199786 136278 199792
rect 136318 199844 136370 199850
rect 136592 199849 136648 199858
rect 136318 199786 136370 199792
rect 136548 199776 136600 199782
rect 135444 199708 135496 199714
rect 135444 199650 135496 199656
rect 135536 199708 135588 199714
rect 135536 199650 135588 199656
rect 135812 199708 135864 199714
rect 136054 199702 136220 199730
rect 136698 199730 136726 200124
rect 136790 199850 136818 200124
rect 136882 199918 136910 200124
rect 136974 199918 137002 200124
rect 137066 199918 137094 200124
rect 137158 199923 137186 200124
rect 136870 199912 136922 199918
rect 136870 199854 136922 199860
rect 136962 199912 137014 199918
rect 136962 199854 137014 199860
rect 137054 199912 137106 199918
rect 137054 199854 137106 199860
rect 137144 199914 137200 199923
rect 137250 199918 137278 200124
rect 137342 199923 137370 200124
rect 136778 199844 136830 199850
rect 137144 199849 137200 199858
rect 137238 199912 137290 199918
rect 137238 199854 137290 199860
rect 137328 199914 137384 199923
rect 137328 199849 137384 199858
rect 136778 199786 136830 199792
rect 136548 199718 136600 199724
rect 136192 199696 136220 199702
rect 136456 199708 136508 199714
rect 136192 199668 136312 199696
rect 135812 199650 135864 199656
rect 135260 199640 135312 199646
rect 135312 199600 135392 199628
rect 135260 199582 135312 199588
rect 135258 199336 135314 199345
rect 135258 199271 135314 199280
rect 135272 194002 135300 199271
rect 135364 197849 135392 199600
rect 135350 197840 135406 197849
rect 135350 197775 135406 197784
rect 135260 193996 135312 194002
rect 135260 193938 135312 193944
rect 135456 192817 135484 199650
rect 135442 192808 135498 192817
rect 135442 192743 135498 192752
rect 135548 186998 135576 199650
rect 135720 199640 135772 199646
rect 135720 199582 135772 199588
rect 135536 186992 135588 186998
rect 135536 186934 135588 186940
rect 135732 186289 135760 199582
rect 135824 192710 135852 199650
rect 135996 199640 136048 199646
rect 135996 199582 136048 199588
rect 136088 199640 136140 199646
rect 136088 199582 136140 199588
rect 135904 199572 135956 199578
rect 135904 199514 135956 199520
rect 135812 192704 135864 192710
rect 135812 192646 135864 192652
rect 135718 186280 135774 186289
rect 135718 186215 135774 186224
rect 135168 185564 135220 185570
rect 135168 185506 135220 185512
rect 135074 185464 135130 185473
rect 135074 185399 135130 185408
rect 135916 183161 135944 199514
rect 136008 197849 136036 199582
rect 136100 198393 136128 199582
rect 136180 199572 136232 199578
rect 136180 199514 136232 199520
rect 136086 198384 136142 198393
rect 136086 198319 136142 198328
rect 136088 198076 136140 198082
rect 136088 198018 136140 198024
rect 135994 197840 136050 197849
rect 135994 197775 136050 197784
rect 136100 184414 136128 198018
rect 136088 184408 136140 184414
rect 136088 184350 136140 184356
rect 135902 183152 135958 183161
rect 135902 183087 135958 183096
rect 136192 179042 136220 199514
rect 136284 198082 136312 199668
rect 136456 199650 136508 199656
rect 136468 199617 136496 199650
rect 136454 199608 136510 199617
rect 136454 199543 136510 199552
rect 136456 199504 136508 199510
rect 136456 199446 136508 199452
rect 136364 199436 136416 199442
rect 136364 199378 136416 199384
rect 136376 198898 136404 199378
rect 136364 198892 136416 198898
rect 136364 198834 136416 198840
rect 136272 198076 136324 198082
rect 136272 198018 136324 198024
rect 136270 197976 136326 197985
rect 136270 197911 136326 197920
rect 135628 179036 135680 179042
rect 135628 178978 135680 178984
rect 136180 179036 136232 179042
rect 136180 178978 136232 178984
rect 134616 176996 134668 177002
rect 134616 176938 134668 176944
rect 135640 148646 135668 178978
rect 136284 174282 136312 197911
rect 136468 186250 136496 199446
rect 136560 199209 136588 199718
rect 136652 199702 136726 199730
rect 136916 199776 136968 199782
rect 137330 199776 137382 199782
rect 136916 199718 136968 199724
rect 137204 199724 137330 199730
rect 137204 199718 137382 199724
rect 136652 199510 136680 199702
rect 136732 199640 136784 199646
rect 136732 199582 136784 199588
rect 136640 199504 136692 199510
rect 136640 199446 136692 199452
rect 136546 199200 136602 199209
rect 136546 199135 136602 199144
rect 136744 199016 136772 199582
rect 136560 198988 136772 199016
rect 136560 186318 136588 198988
rect 136640 198892 136692 198898
rect 136640 198834 136692 198840
rect 136652 186697 136680 198834
rect 136928 195974 136956 199718
rect 137100 199708 137152 199714
rect 137100 199650 137152 199656
rect 137204 199702 137370 199718
rect 137008 199640 137060 199646
rect 137008 199582 137060 199588
rect 136836 195946 136956 195974
rect 136638 186688 136694 186697
rect 136638 186623 136694 186632
rect 136548 186312 136600 186318
rect 136548 186254 136600 186260
rect 136456 186244 136508 186250
rect 136456 186186 136508 186192
rect 136836 182170 136864 195946
rect 137020 186833 137048 199582
rect 137006 186824 137062 186833
rect 137006 186759 137062 186768
rect 137112 185609 137140 199650
rect 137204 186561 137232 199702
rect 137284 199640 137336 199646
rect 137434 199628 137462 200124
rect 137284 199582 137336 199588
rect 137388 199600 137462 199628
rect 137190 186552 137246 186561
rect 137190 186487 137246 186496
rect 137192 186312 137244 186318
rect 137192 186254 137244 186260
rect 137098 185600 137154 185609
rect 137098 185535 137154 185544
rect 136824 182164 136876 182170
rect 136824 182106 136876 182112
rect 136272 174276 136324 174282
rect 136272 174218 136324 174224
rect 137008 173596 137060 173602
rect 137008 173538 137060 173544
rect 135628 148640 135680 148646
rect 135628 148582 135680 148588
rect 134340 148368 134392 148374
rect 132590 148336 132646 148345
rect 134340 148310 134392 148316
rect 132590 148271 132646 148280
rect 137020 147665 137048 173538
rect 137204 148578 137232 186254
rect 137296 185706 137324 199582
rect 137284 185700 137336 185706
rect 137284 185642 137336 185648
rect 137388 173602 137416 199600
rect 137526 199594 137554 200124
rect 137618 199918 137646 200124
rect 137606 199912 137658 199918
rect 137606 199854 137658 199860
rect 137710 199764 137738 200124
rect 137802 199918 137830 200124
rect 137894 199923 137922 200124
rect 137790 199912 137842 199918
rect 137790 199854 137842 199860
rect 137880 199914 137936 199923
rect 137986 199918 138014 200124
rect 138078 199923 138106 200124
rect 137880 199849 137936 199858
rect 137974 199912 138026 199918
rect 137974 199854 138026 199860
rect 138064 199914 138120 199923
rect 138064 199849 138120 199858
rect 138170 199764 138198 200124
rect 138262 199918 138290 200124
rect 138354 199918 138382 200124
rect 138446 199923 138474 200124
rect 138250 199912 138302 199918
rect 138250 199854 138302 199860
rect 138342 199912 138394 199918
rect 138342 199854 138394 199860
rect 138432 199914 138488 199923
rect 138432 199849 138488 199858
rect 137710 199736 137784 199764
rect 138170 199736 138244 199764
rect 137526 199566 137600 199594
rect 137468 199504 137520 199510
rect 137468 199446 137520 199452
rect 137572 199458 137600 199566
rect 137480 192506 137508 199446
rect 137572 199430 137692 199458
rect 137664 192642 137692 199430
rect 137652 192636 137704 192642
rect 137652 192578 137704 192584
rect 137468 192500 137520 192506
rect 137468 192442 137520 192448
rect 137756 185026 137784 199736
rect 137928 199708 137980 199714
rect 137928 199650 137980 199656
rect 138020 199708 138072 199714
rect 138020 199650 138072 199656
rect 137836 198892 137888 198898
rect 137836 198834 137888 198840
rect 137848 195362 137876 198834
rect 137836 195356 137888 195362
rect 137836 195298 137888 195304
rect 137744 185020 137796 185026
rect 137744 184962 137796 184968
rect 137940 178498 137968 199650
rect 138032 199617 138060 199650
rect 138018 199608 138074 199617
rect 138018 199543 138074 199552
rect 138020 199504 138072 199510
rect 138020 199446 138072 199452
rect 138032 192574 138060 199446
rect 138020 192568 138072 192574
rect 138020 192510 138072 192516
rect 138018 192400 138074 192409
rect 138018 192335 138020 192344
rect 138072 192335 138074 192344
rect 138020 192306 138072 192312
rect 137928 178492 137980 178498
rect 137928 178434 137980 178440
rect 137376 173596 137428 173602
rect 137376 173538 137428 173544
rect 138216 172514 138244 199736
rect 138538 199730 138566 200124
rect 138492 199702 138566 199730
rect 138296 199640 138348 199646
rect 138296 199582 138348 199588
rect 138308 190262 138336 199582
rect 138388 199572 138440 199578
rect 138388 199514 138440 199520
rect 138296 190256 138348 190262
rect 138296 190198 138348 190204
rect 138400 177177 138428 199514
rect 138492 190097 138520 199702
rect 138630 199628 138658 200124
rect 138722 199918 138750 200124
rect 138710 199912 138762 199918
rect 138710 199854 138762 199860
rect 138814 199764 138842 200124
rect 138584 199600 138658 199628
rect 138768 199736 138842 199764
rect 138478 190088 138534 190097
rect 138478 190023 138534 190032
rect 138584 189718 138612 199600
rect 138662 196888 138718 196897
rect 138662 196823 138718 196832
rect 138676 195566 138704 196823
rect 138664 195560 138716 195566
rect 138664 195502 138716 195508
rect 138662 195392 138718 195401
rect 138662 195327 138718 195336
rect 138676 192914 138704 195327
rect 138768 194750 138796 199736
rect 138906 199696 138934 200124
rect 138860 199668 138934 199696
rect 138998 199696 139026 200124
rect 139090 199764 139118 200124
rect 139182 199923 139210 200124
rect 139168 199914 139224 199923
rect 139274 199918 139302 200124
rect 139366 199923 139394 200124
rect 139168 199849 139224 199858
rect 139262 199912 139314 199918
rect 139262 199854 139314 199860
rect 139352 199914 139408 199923
rect 139352 199849 139408 199858
rect 139090 199736 139164 199764
rect 138998 199668 139072 199696
rect 138756 194744 138808 194750
rect 138756 194686 138808 194692
rect 138664 192908 138716 192914
rect 138664 192850 138716 192856
rect 138860 189786 138888 199668
rect 138938 199200 138994 199209
rect 138938 199135 138994 199144
rect 138952 198898 138980 199135
rect 138940 198892 138992 198898
rect 138940 198834 138992 198840
rect 138938 198384 138994 198393
rect 138938 198319 138994 198328
rect 138952 191010 138980 198319
rect 138940 191004 138992 191010
rect 138940 190946 138992 190952
rect 138938 189816 138994 189825
rect 138848 189780 138900 189786
rect 138938 189751 138994 189760
rect 138848 189722 138900 189728
rect 138572 189712 138624 189718
rect 138572 189654 138624 189660
rect 138952 189650 138980 189751
rect 138940 189644 138992 189650
rect 138940 189586 138992 189592
rect 138386 177168 138442 177177
rect 138386 177103 138442 177112
rect 139044 175001 139072 199668
rect 139136 195498 139164 199736
rect 139458 199730 139486 200124
rect 139550 199923 139578 200124
rect 139536 199914 139592 199923
rect 139642 199918 139670 200124
rect 139734 199923 139762 200124
rect 139536 199849 139592 199858
rect 139630 199912 139682 199918
rect 139630 199854 139682 199860
rect 139720 199914 139776 199923
rect 139720 199849 139776 199858
rect 139412 199702 139486 199730
rect 139584 199776 139636 199782
rect 139826 199764 139854 200124
rect 139918 199918 139946 200124
rect 139906 199912 139958 199918
rect 139906 199854 139958 199860
rect 139584 199718 139636 199724
rect 139780 199736 139854 199764
rect 139216 199640 139268 199646
rect 139216 199582 139268 199588
rect 139124 195492 139176 195498
rect 139124 195434 139176 195440
rect 139228 186289 139256 199582
rect 139412 190058 139440 199702
rect 139596 195294 139624 199718
rect 139584 195288 139636 195294
rect 139584 195230 139636 195236
rect 139400 190052 139452 190058
rect 139400 189994 139452 190000
rect 139214 186280 139270 186289
rect 139214 186215 139270 186224
rect 139122 185736 139178 185745
rect 139122 185671 139178 185680
rect 139136 183802 139164 185671
rect 139124 183796 139176 183802
rect 139124 183738 139176 183744
rect 139780 179353 139808 199736
rect 139860 199640 139912 199646
rect 140010 199628 140038 200124
rect 140102 199764 140130 200124
rect 140194 199923 140222 200124
rect 140180 199914 140236 199923
rect 140180 199849 140236 199858
rect 140286 199764 140314 200124
rect 140102 199736 140176 199764
rect 139860 199582 139912 199588
rect 139964 199600 140038 199628
rect 139872 198121 139900 199582
rect 139858 198112 139914 198121
rect 139858 198047 139914 198056
rect 139858 195800 139914 195809
rect 139858 195735 139914 195744
rect 139872 191418 139900 195735
rect 139860 191412 139912 191418
rect 139860 191354 139912 191360
rect 139964 190330 139992 199600
rect 140044 199504 140096 199510
rect 140044 199446 140096 199452
rect 140056 199306 140084 199446
rect 140044 199300 140096 199306
rect 140044 199242 140096 199248
rect 139952 190324 140004 190330
rect 139952 190266 140004 190272
rect 140148 186289 140176 199736
rect 140240 199736 140314 199764
rect 140240 193866 140268 199736
rect 140378 199696 140406 200124
rect 140470 199923 140498 200124
rect 140456 199914 140512 199923
rect 140456 199849 140512 199858
rect 140562 199764 140590 200124
rect 140332 199668 140406 199696
rect 140516 199736 140590 199764
rect 140332 198121 140360 199668
rect 140412 199436 140464 199442
rect 140412 199378 140464 199384
rect 140424 199345 140452 199378
rect 140410 199336 140466 199345
rect 140410 199271 140466 199280
rect 140318 198112 140374 198121
rect 140318 198047 140374 198056
rect 140228 193860 140280 193866
rect 140228 193802 140280 193808
rect 140516 189689 140544 199736
rect 140654 199696 140682 200124
rect 140746 199923 140774 200124
rect 140732 199914 140788 199923
rect 140838 199918 140866 200124
rect 140732 199849 140788 199858
rect 140826 199912 140878 199918
rect 140826 199854 140878 199860
rect 140780 199776 140832 199782
rect 140780 199718 140832 199724
rect 140608 199668 140682 199696
rect 140502 189680 140558 189689
rect 140502 189615 140558 189624
rect 139858 186280 139914 186289
rect 139858 186215 139914 186224
rect 140134 186280 140190 186289
rect 140134 186215 140190 186224
rect 139766 179344 139822 179353
rect 139766 179279 139822 179288
rect 139030 174992 139086 175001
rect 139030 174927 139086 174936
rect 138216 172486 138520 172514
rect 138492 151814 138520 172486
rect 138308 151786 138520 151814
rect 137192 148572 137244 148578
rect 137192 148514 137244 148520
rect 137006 147656 137062 147665
rect 137006 147591 137062 147600
rect 132408 146124 132460 146130
rect 132408 146066 132460 146072
rect 132224 146056 132276 146062
rect 132224 145998 132276 146004
rect 132040 143404 132092 143410
rect 132040 143346 132092 143352
rect 131684 139998 131988 140026
rect 131500 139726 131560 139754
rect 131684 139369 131712 139998
rect 132052 139890 132080 143346
rect 132052 139862 132112 139890
rect 132236 139369 132264 145998
rect 132420 142798 132448 146066
rect 137284 144696 137336 144702
rect 137284 144638 137336 144644
rect 132866 143304 132922 143313
rect 132866 143239 132922 143248
rect 133420 143268 133472 143274
rect 132408 142792 132460 142798
rect 132408 142734 132460 142740
rect 132500 142520 132552 142526
rect 132500 142462 132552 142468
rect 132512 139890 132540 142462
rect 132880 139890 132908 143239
rect 133420 143210 133472 143216
rect 133432 139890 133460 143210
rect 135260 143132 135312 143138
rect 135260 143074 135312 143080
rect 134524 142724 134576 142730
rect 134524 142666 134576 142672
rect 133972 141636 134024 141642
rect 133972 141578 134024 141584
rect 133984 139890 134012 141578
rect 134536 139890 134564 142666
rect 135272 139890 135300 143074
rect 136732 142996 136784 143002
rect 136732 142938 136784 142944
rect 136180 142792 136232 142798
rect 136180 142734 136232 142740
rect 135628 141500 135680 141506
rect 135628 141442 135680 141448
rect 135640 139890 135668 141442
rect 136192 139890 136220 142734
rect 136744 139890 136772 142938
rect 137296 139890 137324 144638
rect 138020 143336 138072 143342
rect 138020 143278 138072 143284
rect 138032 139890 138060 143278
rect 132512 139862 132664 139890
rect 132880 139862 133216 139890
rect 133432 139862 133768 139890
rect 133984 139862 134320 139890
rect 134536 139862 134872 139890
rect 135272 139862 135424 139890
rect 135640 139862 135976 139890
rect 136192 139862 136528 139890
rect 136744 139862 137080 139890
rect 137296 139862 137632 139890
rect 138032 139862 138184 139890
rect 138308 139369 138336 151786
rect 139872 148918 139900 186215
rect 140608 185609 140636 199668
rect 140688 199572 140740 199578
rect 140688 199514 140740 199520
rect 140700 192982 140728 199514
rect 140688 192976 140740 192982
rect 140688 192918 140740 192924
rect 140792 188970 140820 199718
rect 140930 199696 140958 200124
rect 141022 199764 141050 200124
rect 141114 199918 141142 200124
rect 141102 199912 141154 199918
rect 141102 199854 141154 199860
rect 141206 199764 141234 200124
rect 141298 199923 141326 200124
rect 141284 199914 141340 199923
rect 141284 199849 141340 199858
rect 141022 199736 141096 199764
rect 140930 199668 141004 199696
rect 140872 199504 140924 199510
rect 140872 199446 140924 199452
rect 140780 188964 140832 188970
rect 140780 188906 140832 188912
rect 140594 185600 140650 185609
rect 140594 185535 140650 185544
rect 140884 180402 140912 199446
rect 140976 185337 141004 199668
rect 141068 185473 141096 199736
rect 141160 199736 141234 199764
rect 141160 185638 141188 199736
rect 141390 199696 141418 200124
rect 141482 199764 141510 200124
rect 141574 199918 141602 200124
rect 141666 199918 141694 200124
rect 141758 199923 141786 200124
rect 141562 199912 141614 199918
rect 141562 199854 141614 199860
rect 141654 199912 141706 199918
rect 141654 199854 141706 199860
rect 141744 199914 141800 199923
rect 141850 199918 141878 200124
rect 141744 199849 141800 199858
rect 141838 199912 141890 199918
rect 141838 199854 141890 199860
rect 141942 199764 141970 200124
rect 141482 199736 141556 199764
rect 141390 199668 141464 199696
rect 141332 199164 141384 199170
rect 141332 199106 141384 199112
rect 141344 191282 141372 199106
rect 141332 191276 141384 191282
rect 141332 191218 141384 191224
rect 141436 190466 141464 199668
rect 141424 190460 141476 190466
rect 141424 190402 141476 190408
rect 141528 186266 141556 199736
rect 141896 199736 141970 199764
rect 141608 199708 141660 199714
rect 141608 199650 141660 199656
rect 141620 192545 141648 199650
rect 141700 199640 141752 199646
rect 141700 199582 141752 199588
rect 141606 192536 141662 192545
rect 141606 192471 141662 192480
rect 141712 192302 141740 199582
rect 141792 199504 141844 199510
rect 141792 199446 141844 199452
rect 141804 198121 141832 199446
rect 141790 198112 141846 198121
rect 141790 198047 141846 198056
rect 141700 192296 141752 192302
rect 141700 192238 141752 192244
rect 141896 190398 141924 199736
rect 142034 199696 142062 200124
rect 142126 199764 142154 200124
rect 142218 199918 142246 200124
rect 142310 199923 142338 200124
rect 142206 199912 142258 199918
rect 142206 199854 142258 199860
rect 142296 199914 142352 199923
rect 142402 199918 142430 200124
rect 142494 199923 142522 200124
rect 142296 199849 142352 199858
rect 142390 199912 142442 199918
rect 142390 199854 142442 199860
rect 142480 199914 142536 199923
rect 142480 199849 142536 199858
rect 142586 199764 142614 200124
rect 142678 199923 142706 200124
rect 142664 199914 142720 199923
rect 142770 199918 142798 200124
rect 142664 199849 142720 199858
rect 142758 199912 142810 199918
rect 142758 199854 142810 199860
rect 142126 199736 142200 199764
rect 141988 199668 142062 199696
rect 141884 190392 141936 190398
rect 141884 190334 141936 190340
rect 141436 186238 141556 186266
rect 141148 185632 141200 185638
rect 141148 185574 141200 185580
rect 141054 185464 141110 185473
rect 141054 185399 141110 185408
rect 140962 185328 141018 185337
rect 140962 185263 141018 185272
rect 140872 180396 140924 180402
rect 140872 180338 140924 180344
rect 139860 148912 139912 148918
rect 139860 148854 139912 148860
rect 141146 144528 141202 144537
rect 141146 144463 141202 144472
rect 138938 143984 138994 143993
rect 138938 143919 138994 143928
rect 138388 143200 138440 143206
rect 138388 143142 138440 143148
rect 138400 139890 138428 143142
rect 138952 139890 138980 143919
rect 140044 143064 140096 143070
rect 140044 143006 140096 143012
rect 139490 140040 139546 140049
rect 139490 139975 139546 139984
rect 139504 139890 139532 139975
rect 140056 139890 140084 143006
rect 140780 142180 140832 142186
rect 140780 142122 140832 142128
rect 140792 139890 140820 142122
rect 141160 139890 141188 144463
rect 141436 141681 141464 186238
rect 141516 185632 141568 185638
rect 141988 185609 142016 199668
rect 141516 185574 141568 185580
rect 141974 185600 142030 185609
rect 141422 141672 141478 141681
rect 141422 141607 141478 141616
rect 141528 141273 141556 185574
rect 141974 185535 142030 185544
rect 142172 185366 142200 199736
rect 142540 199736 142614 199764
rect 142712 199776 142764 199782
rect 142436 199708 142488 199714
rect 142436 199650 142488 199656
rect 142252 199640 142304 199646
rect 142252 199582 142304 199588
rect 142264 195634 142292 199582
rect 142448 198966 142476 199650
rect 142436 198960 142488 198966
rect 142436 198902 142488 198908
rect 142342 198520 142398 198529
rect 142342 198455 142398 198464
rect 142356 197674 142384 198455
rect 142434 198112 142490 198121
rect 142434 198047 142490 198056
rect 142344 197668 142396 197674
rect 142344 197610 142396 197616
rect 142252 195628 142304 195634
rect 142252 195570 142304 195576
rect 142448 185570 142476 198047
rect 142540 195430 142568 199736
rect 142862 199764 142890 200124
rect 142712 199718 142764 199724
rect 142816 199736 142890 199764
rect 142618 199200 142674 199209
rect 142618 199135 142674 199144
rect 142632 198898 142660 199135
rect 142620 198892 142672 198898
rect 142620 198834 142672 198840
rect 142528 195424 142580 195430
rect 142528 195366 142580 195372
rect 142724 185688 142752 199718
rect 142816 187474 142844 199736
rect 142954 199696 142982 200124
rect 143046 199923 143074 200124
rect 143032 199914 143088 199923
rect 143138 199918 143166 200124
rect 143230 199918 143258 200124
rect 143032 199849 143088 199858
rect 143126 199912 143178 199918
rect 143126 199854 143178 199860
rect 143218 199912 143270 199918
rect 143218 199854 143270 199860
rect 143172 199776 143224 199782
rect 142908 199668 142982 199696
rect 143078 199744 143134 199753
rect 143322 199764 143350 200124
rect 143414 199918 143442 200124
rect 143506 199918 143534 200124
rect 143402 199912 143454 199918
rect 143402 199854 143454 199860
rect 143494 199912 143546 199918
rect 143494 199854 143546 199860
rect 143598 199764 143626 200124
rect 143690 199918 143718 200124
rect 143678 199912 143730 199918
rect 143678 199854 143730 199860
rect 143782 199764 143810 200124
rect 143172 199718 143224 199724
rect 143276 199736 143350 199764
rect 143552 199736 143626 199764
rect 143736 199736 143810 199764
rect 143078 199679 143134 199688
rect 142908 196926 142936 199668
rect 142896 196920 142948 196926
rect 142896 196862 142948 196868
rect 143092 191350 143120 199679
rect 143184 195702 143212 199718
rect 143172 195696 143224 195702
rect 143172 195638 143224 195644
rect 143080 191344 143132 191350
rect 143080 191286 143132 191292
rect 142804 187468 142856 187474
rect 142804 187410 142856 187416
rect 142540 185660 142752 185688
rect 142436 185564 142488 185570
rect 142436 185506 142488 185512
rect 142160 185360 142212 185366
rect 142160 185302 142212 185308
rect 142436 178492 142488 178498
rect 142436 178434 142488 178440
rect 142066 171048 142122 171057
rect 142066 170983 142122 170992
rect 142080 161537 142108 170983
rect 142066 161528 142122 161537
rect 142066 161463 142122 161472
rect 142066 161392 142122 161401
rect 142066 161327 142122 161336
rect 142080 151881 142108 161327
rect 142066 151872 142122 151881
rect 142066 151807 142122 151816
rect 142066 151736 142122 151745
rect 142066 151671 142122 151680
rect 141700 142928 141752 142934
rect 141700 142870 141752 142876
rect 141514 141264 141570 141273
rect 141514 141199 141570 141208
rect 141712 139890 141740 142870
rect 142080 142361 142108 151671
rect 142448 148238 142476 178434
rect 142436 148232 142488 148238
rect 142436 148174 142488 148180
rect 142540 145586 142568 185660
rect 142986 185600 143042 185609
rect 142712 185564 142764 185570
rect 142986 185535 143042 185544
rect 142712 185506 142764 185512
rect 142724 146946 142752 185506
rect 143000 148986 143028 185535
rect 143276 178498 143304 199736
rect 143356 199640 143408 199646
rect 143356 199582 143408 199588
rect 143368 192273 143396 199582
rect 143448 199572 143500 199578
rect 143448 199514 143500 199520
rect 143354 192264 143410 192273
rect 143354 192199 143410 192208
rect 143460 192137 143488 199514
rect 143446 192128 143502 192137
rect 143446 192063 143502 192072
rect 143552 191865 143580 199736
rect 143632 199640 143684 199646
rect 143632 199582 143684 199588
rect 143538 191856 143594 191865
rect 143538 191791 143594 191800
rect 143644 191185 143672 199582
rect 143630 191176 143686 191185
rect 143630 191111 143686 191120
rect 143736 188018 143764 199736
rect 143874 199696 143902 200124
rect 143828 199668 143902 199696
rect 143828 190641 143856 199668
rect 143966 199628 143994 200124
rect 144058 199918 144086 200124
rect 144046 199912 144098 199918
rect 144046 199854 144098 199860
rect 144150 199764 144178 200124
rect 144242 199918 144270 200124
rect 144334 199918 144362 200124
rect 144230 199912 144282 199918
rect 144230 199854 144282 199860
rect 144322 199912 144374 199918
rect 144322 199854 144374 199860
rect 143920 199600 143994 199628
rect 144104 199736 144178 199764
rect 144426 199764 144454 200124
rect 144518 199923 144546 200124
rect 144504 199914 144560 199923
rect 144504 199849 144560 199858
rect 144610 199764 144638 200124
rect 144702 199923 144730 200124
rect 144688 199914 144744 199923
rect 144688 199849 144744 199858
rect 144794 199764 144822 200124
rect 144886 199918 144914 200124
rect 144874 199912 144926 199918
rect 144874 199854 144926 199860
rect 144978 199764 145006 200124
rect 144426 199736 144500 199764
rect 144610 199736 144684 199764
rect 143920 199170 143948 199600
rect 144000 199504 144052 199510
rect 144000 199446 144052 199452
rect 143908 199164 143960 199170
rect 143908 199106 143960 199112
rect 144012 190738 144040 199446
rect 144000 190732 144052 190738
rect 144000 190674 144052 190680
rect 143814 190632 143870 190641
rect 143814 190567 143870 190576
rect 144104 190505 144132 199736
rect 144276 199708 144328 199714
rect 144276 199650 144328 199656
rect 144184 199640 144236 199646
rect 144184 199582 144236 199588
rect 144196 191146 144224 199582
rect 144184 191140 144236 191146
rect 144184 191082 144236 191088
rect 144090 190496 144146 190505
rect 144090 190431 144146 190440
rect 143724 188012 143776 188018
rect 143724 187954 143776 187960
rect 144288 185162 144316 199650
rect 144472 190777 144500 199736
rect 144552 199572 144604 199578
rect 144552 199514 144604 199520
rect 144564 192438 144592 199514
rect 144656 196858 144684 199736
rect 144748 199736 144822 199764
rect 144932 199736 145006 199764
rect 144644 196852 144696 196858
rect 144644 196794 144696 196800
rect 144552 192432 144604 192438
rect 144552 192374 144604 192380
rect 144748 191049 144776 199736
rect 144828 199640 144880 199646
rect 144828 199582 144880 199588
rect 144840 199034 144868 199582
rect 144828 199028 144880 199034
rect 144828 198970 144880 198976
rect 144734 191040 144790 191049
rect 144734 190975 144790 190984
rect 144458 190768 144514 190777
rect 144458 190703 144514 190712
rect 144276 185156 144328 185162
rect 144276 185098 144328 185104
rect 144932 184346 144960 199736
rect 145070 199696 145098 200124
rect 145162 199730 145190 200124
rect 145254 199850 145282 200124
rect 145346 199850 145374 200124
rect 145438 199918 145466 200124
rect 145530 199918 145558 200124
rect 145426 199912 145478 199918
rect 145426 199854 145478 199860
rect 145518 199912 145570 199918
rect 145518 199854 145570 199860
rect 145242 199844 145294 199850
rect 145242 199786 145294 199792
rect 145334 199844 145386 199850
rect 145334 199786 145386 199792
rect 145622 199764 145650 200124
rect 145714 199923 145742 200124
rect 145700 199914 145756 199923
rect 145806 199918 145834 200124
rect 145700 199849 145756 199858
rect 145794 199912 145846 199918
rect 145794 199854 145846 199860
rect 145748 199776 145800 199782
rect 145622 199736 145696 199764
rect 145162 199702 145236 199730
rect 145024 199668 145098 199696
rect 145024 194138 145052 199668
rect 145208 197062 145236 199702
rect 145288 199708 145340 199714
rect 145288 199650 145340 199656
rect 145380 199708 145432 199714
rect 145380 199650 145432 199656
rect 145196 197056 145248 197062
rect 145196 196998 145248 197004
rect 145012 194132 145064 194138
rect 145012 194074 145064 194080
rect 145300 190942 145328 199650
rect 145288 190936 145340 190942
rect 145288 190878 145340 190884
rect 145392 186017 145420 199650
rect 145564 199640 145616 199646
rect 145564 199582 145616 199588
rect 145576 198830 145604 199582
rect 145564 198824 145616 198830
rect 145564 198766 145616 198772
rect 145668 192953 145696 199736
rect 145898 199764 145926 200124
rect 145990 199918 146018 200124
rect 145978 199912 146030 199918
rect 145978 199854 146030 199860
rect 146082 199764 146110 200124
rect 145748 199718 145800 199724
rect 145852 199736 145926 199764
rect 146036 199736 146110 199764
rect 145654 192944 145710 192953
rect 145654 192879 145710 192888
rect 145760 190369 145788 199718
rect 145852 194274 145880 199736
rect 145840 194268 145892 194274
rect 145840 194210 145892 194216
rect 145746 190360 145802 190369
rect 145746 190295 145802 190304
rect 146036 188902 146064 199736
rect 146174 199696 146202 200124
rect 146266 199764 146294 200124
rect 146358 199923 146386 200124
rect 146344 199914 146400 199923
rect 146344 199849 146400 199858
rect 146450 199764 146478 200124
rect 146266 199736 146340 199764
rect 146128 199668 146202 199696
rect 146128 198801 146156 199668
rect 146114 198792 146170 198801
rect 146114 198727 146170 198736
rect 146024 188896 146076 188902
rect 146024 188838 146076 188844
rect 145378 186008 145434 186017
rect 145378 185943 145434 185952
rect 144920 184340 144972 184346
rect 144920 184282 144972 184288
rect 145564 179036 145616 179042
rect 145564 178978 145616 178984
rect 143264 178492 143316 178498
rect 143264 178434 143316 178440
rect 145196 175908 145248 175914
rect 145196 175850 145248 175856
rect 142988 148980 143040 148986
rect 142988 148922 143040 148928
rect 142712 146940 142764 146946
rect 142712 146882 142764 146888
rect 145208 145586 145236 175850
rect 145576 145654 145604 178978
rect 146312 175914 146340 199736
rect 146404 199736 146478 199764
rect 146404 194070 146432 199736
rect 146542 199696 146570 200124
rect 146634 199764 146662 200124
rect 146726 199923 146754 200124
rect 146712 199914 146768 199923
rect 146712 199849 146768 199858
rect 146818 199764 146846 200124
rect 146910 199923 146938 200124
rect 146896 199914 146952 199923
rect 146896 199849 146952 199858
rect 147002 199764 147030 200124
rect 147094 199923 147122 200124
rect 147080 199914 147136 199923
rect 147080 199849 147136 199858
rect 147186 199764 147214 200124
rect 146634 199736 146708 199764
rect 146496 199668 146570 199696
rect 146392 194064 146444 194070
rect 146392 194006 146444 194012
rect 146300 175908 146352 175914
rect 146300 175850 146352 175856
rect 146496 152590 146524 199668
rect 146680 191457 146708 199736
rect 146772 199736 146846 199764
rect 146956 199736 147030 199764
rect 147140 199736 147214 199764
rect 147278 199764 147306 200124
rect 147370 199918 147398 200124
rect 147358 199912 147410 199918
rect 147358 199854 147410 199860
rect 147462 199764 147490 200124
rect 147554 199918 147582 200124
rect 147542 199912 147594 199918
rect 147542 199854 147594 199860
rect 147646 199764 147674 200124
rect 147278 199736 147352 199764
rect 146666 191448 146722 191457
rect 146666 191383 146722 191392
rect 146772 184210 146800 199736
rect 146956 194206 146984 199736
rect 146944 194200 146996 194206
rect 146944 194142 146996 194148
rect 147140 189961 147168 199736
rect 147126 189952 147182 189961
rect 147126 189887 147182 189896
rect 146760 184204 146812 184210
rect 146760 184146 146812 184152
rect 147324 181937 147352 199736
rect 147416 199736 147490 199764
rect 147600 199736 147674 199764
rect 147738 199764 147766 200124
rect 147830 199923 147858 200124
rect 147816 199914 147872 199923
rect 147816 199849 147872 199858
rect 147738 199736 147812 199764
rect 147310 181928 147366 181937
rect 147310 181863 147366 181872
rect 147416 180538 147444 199736
rect 147496 199504 147548 199510
rect 147496 199446 147548 199452
rect 147508 186289 147536 199446
rect 147600 196654 147628 199736
rect 147680 199640 147732 199646
rect 147680 199582 147732 199588
rect 147588 196648 147640 196654
rect 147588 196590 147640 196596
rect 147692 191321 147720 199582
rect 147678 191312 147734 191321
rect 147678 191247 147734 191256
rect 147494 186280 147550 186289
rect 147494 186215 147550 186224
rect 147588 182708 147640 182714
rect 147588 182650 147640 182656
rect 146852 180532 146904 180538
rect 146852 180474 146904 180480
rect 147404 180532 147456 180538
rect 147404 180474 147456 180480
rect 146758 179344 146814 179353
rect 146758 179279 146814 179288
rect 146484 152584 146536 152590
rect 146484 152526 146536 152532
rect 146300 145988 146352 145994
rect 146300 145930 146352 145936
rect 145564 145648 145616 145654
rect 145564 145590 145616 145596
rect 142528 145580 142580 145586
rect 142528 145522 142580 145528
rect 145196 145580 145248 145586
rect 145196 145522 145248 145528
rect 142802 144800 142858 144809
rect 142802 144735 142858 144744
rect 142252 144628 142304 144634
rect 142252 144570 142304 144576
rect 142066 142352 142122 142361
rect 142066 142287 142122 142296
rect 142264 139890 142292 144570
rect 142816 139890 142844 144735
rect 144458 144664 144514 144673
rect 144458 144599 144514 144608
rect 143540 142860 143592 142866
rect 143540 142802 143592 142808
rect 143552 139890 143580 142802
rect 143906 141808 143962 141817
rect 143906 141743 143962 141752
rect 143920 139890 143948 141743
rect 144472 139890 144500 144599
rect 145562 144392 145618 144401
rect 145562 144327 145618 144336
rect 145102 143032 145158 143041
rect 145102 142967 145158 142976
rect 145116 139890 145144 142967
rect 145576 139890 145604 144327
rect 146312 139890 146340 145930
rect 146666 143168 146722 143177
rect 146666 143103 146722 143112
rect 146680 139890 146708 143103
rect 146772 140146 146800 179279
rect 146864 140214 146892 180474
rect 146944 177200 146996 177206
rect 146944 177142 146996 177148
rect 146956 140282 146984 177142
rect 147600 145654 147628 182650
rect 147784 177206 147812 199736
rect 147922 199628 147950 200124
rect 148014 199764 148042 200124
rect 148106 199918 148134 200124
rect 148198 199923 148226 200124
rect 148094 199912 148146 199918
rect 148094 199854 148146 199860
rect 148184 199914 148240 199923
rect 148290 199918 148318 200124
rect 148184 199849 148240 199858
rect 148278 199912 148330 199918
rect 148278 199854 148330 199860
rect 148140 199776 148192 199782
rect 148014 199736 148088 199764
rect 147922 199600 147996 199628
rect 147772 177200 147824 177206
rect 147772 177142 147824 177148
rect 147968 172514 147996 199600
rect 148060 190913 148088 199736
rect 148382 199764 148410 200124
rect 148140 199718 148192 199724
rect 148336 199736 148410 199764
rect 148046 190904 148102 190913
rect 148046 190839 148102 190848
rect 148152 187241 148180 199718
rect 148232 199572 148284 199578
rect 148232 199514 148284 199520
rect 148244 194342 148272 199514
rect 148232 194336 148284 194342
rect 148232 194278 148284 194284
rect 148138 187232 148194 187241
rect 148138 187167 148194 187176
rect 148336 186930 148364 199736
rect 148474 199696 148502 200124
rect 148428 199668 148502 199696
rect 148428 199102 148456 199668
rect 148566 199628 148594 200124
rect 148658 199918 148686 200124
rect 148750 199918 148778 200124
rect 148842 199918 148870 200124
rect 148934 199918 148962 200124
rect 149026 199923 149054 200124
rect 148646 199912 148698 199918
rect 148646 199854 148698 199860
rect 148738 199912 148790 199918
rect 148738 199854 148790 199860
rect 148830 199912 148882 199918
rect 148830 199854 148882 199860
rect 148922 199912 148974 199918
rect 148922 199854 148974 199860
rect 149012 199914 149068 199923
rect 149118 199918 149146 200124
rect 149210 199918 149238 200124
rect 149302 199923 149330 200124
rect 149012 199849 149068 199858
rect 149106 199912 149158 199918
rect 149106 199854 149158 199860
rect 149198 199912 149250 199918
rect 149198 199854 149250 199860
rect 149288 199914 149344 199923
rect 149394 199918 149422 200124
rect 149288 199849 149344 199858
rect 149382 199912 149434 199918
rect 149382 199854 149434 199860
rect 148692 199776 148744 199782
rect 148692 199718 148744 199724
rect 148784 199776 148836 199782
rect 149060 199776 149112 199782
rect 148784 199718 148836 199724
rect 148966 199744 149022 199753
rect 148520 199600 148594 199628
rect 148416 199096 148468 199102
rect 148416 199038 148468 199044
rect 148324 186924 148376 186930
rect 148324 186866 148376 186872
rect 148520 186266 148548 199600
rect 148704 199238 148732 199718
rect 148692 199232 148744 199238
rect 148692 199174 148744 199180
rect 148152 186238 148548 186266
rect 148048 184204 148100 184210
rect 148048 184146 148100 184152
rect 147876 172486 147996 172514
rect 147876 152522 147904 172486
rect 147864 152516 147916 152522
rect 147864 152458 147916 152464
rect 147588 145648 147640 145654
rect 147588 145590 147640 145596
rect 148060 144294 148088 184146
rect 148048 144288 148100 144294
rect 147218 144256 147274 144265
rect 148048 144230 148100 144236
rect 147218 144191 147274 144200
rect 146944 140276 146996 140282
rect 146944 140218 146996 140224
rect 146852 140208 146904 140214
rect 146852 140150 146904 140156
rect 146760 140140 146812 140146
rect 146760 140082 146812 140088
rect 147232 139890 147260 144191
rect 147770 144120 147826 144129
rect 147770 144055 147826 144064
rect 147784 139890 147812 144055
rect 148152 140350 148180 186238
rect 148796 186182 148824 199718
rect 148876 199708 148928 199714
rect 149060 199718 149112 199724
rect 149152 199776 149204 199782
rect 149152 199718 149204 199724
rect 149244 199776 149296 199782
rect 149486 199764 149514 200124
rect 149244 199718 149296 199724
rect 149440 199736 149514 199764
rect 149578 199764 149606 200124
rect 149670 199918 149698 200124
rect 149658 199912 149710 199918
rect 149658 199854 149710 199860
rect 149762 199764 149790 200124
rect 149578 199736 149652 199764
rect 148966 199679 149022 199688
rect 148876 199650 148928 199656
rect 148888 186289 148916 199650
rect 148980 199481 149008 199679
rect 148966 199472 149022 199481
rect 148966 199407 149022 199416
rect 148874 186280 148930 186289
rect 148874 186215 148930 186224
rect 148968 186244 149020 186250
rect 148968 186186 149020 186192
rect 148324 186176 148376 186182
rect 148324 186118 148376 186124
rect 148784 186176 148836 186182
rect 148784 186118 148836 186124
rect 148336 151814 148364 186118
rect 148244 151786 148364 151814
rect 148140 140344 148192 140350
rect 148140 140286 148192 140292
rect 148244 140078 148272 151786
rect 148980 149734 149008 186186
rect 149072 179042 149100 199718
rect 149164 198286 149192 199718
rect 149152 198280 149204 198286
rect 149152 198222 149204 198228
rect 149256 193769 149284 199718
rect 149336 199708 149388 199714
rect 149336 199650 149388 199656
rect 149242 193760 149298 193769
rect 149242 193695 149298 193704
rect 149348 191264 149376 199650
rect 149440 194313 149468 199736
rect 149520 199640 149572 199646
rect 149520 199582 149572 199588
rect 149532 196722 149560 199582
rect 149624 197985 149652 199736
rect 149716 199736 149790 199764
rect 149610 197976 149666 197985
rect 149610 197911 149666 197920
rect 149520 196716 149572 196722
rect 149520 196658 149572 196664
rect 149426 194304 149482 194313
rect 149426 194239 149482 194248
rect 149716 193905 149744 199736
rect 149854 199714 149882 200124
rect 149946 199764 149974 200124
rect 150038 199918 150066 200124
rect 150130 199918 150158 200124
rect 150026 199912 150078 199918
rect 150026 199854 150078 199860
rect 150118 199912 150170 199918
rect 150118 199854 150170 199860
rect 150222 199764 150250 200124
rect 150314 199923 150342 200124
rect 150300 199914 150356 199923
rect 150300 199849 150356 199858
rect 150406 199782 150434 200124
rect 149946 199736 150020 199764
rect 149842 199708 149894 199714
rect 149842 199650 149894 199656
rect 149888 199504 149940 199510
rect 149888 199446 149940 199452
rect 149702 193896 149758 193905
rect 149702 193831 149758 193840
rect 149256 191236 149376 191264
rect 149060 179036 149112 179042
rect 149060 178978 149112 178984
rect 148968 149728 149020 149734
rect 148968 149670 149020 149676
rect 149256 145858 149284 191236
rect 149334 191176 149390 191185
rect 149334 191111 149390 191120
rect 149348 152658 149376 191111
rect 149612 185632 149664 185638
rect 149900 185609 149928 199446
rect 149612 185574 149664 185580
rect 149886 185600 149942 185609
rect 149520 182028 149572 182034
rect 149520 181970 149572 181976
rect 149336 152652 149388 152658
rect 149336 152594 149388 152600
rect 149244 145852 149296 145858
rect 149244 145794 149296 145800
rect 149532 145790 149560 181970
rect 149520 145784 149572 145790
rect 149520 145726 149572 145732
rect 149624 145722 149652 185574
rect 149886 185535 149942 185544
rect 149992 182034 150020 199736
rect 150176 199736 150250 199764
rect 150394 199776 150446 199782
rect 150072 199708 150124 199714
rect 150072 199650 150124 199656
rect 150084 197946 150112 199650
rect 150072 197940 150124 197946
rect 150072 197882 150124 197888
rect 150176 185638 150204 199736
rect 150394 199718 150446 199724
rect 150348 199640 150400 199646
rect 150498 199628 150526 200124
rect 150590 199696 150618 200124
rect 150682 199764 150710 200124
rect 150774 199918 150802 200124
rect 150762 199912 150814 199918
rect 150762 199854 150814 199860
rect 150866 199764 150894 200124
rect 150958 199923 150986 200124
rect 150944 199914 151000 199923
rect 150944 199849 151000 199858
rect 151050 199764 151078 200124
rect 151142 199923 151170 200124
rect 151128 199914 151184 199923
rect 151234 199918 151262 200124
rect 151128 199849 151184 199858
rect 151222 199912 151274 199918
rect 151222 199854 151274 199860
rect 150682 199736 150756 199764
rect 150866 199736 150940 199764
rect 150590 199668 150664 199696
rect 150498 199600 150572 199628
rect 150348 199582 150400 199588
rect 150360 195906 150388 199582
rect 150348 195900 150400 195906
rect 150348 195842 150400 195848
rect 150544 186266 150572 199600
rect 150636 193662 150664 199668
rect 150728 198966 150756 199736
rect 150808 199640 150860 199646
rect 150808 199582 150860 199588
rect 150716 198960 150768 198966
rect 150716 198902 150768 198908
rect 150820 198558 150848 199582
rect 150808 198552 150860 198558
rect 150808 198494 150860 198500
rect 150624 193656 150676 193662
rect 150624 193598 150676 193604
rect 150912 186425 150940 199736
rect 151004 199736 151078 199764
rect 151176 199776 151228 199782
rect 150898 186416 150954 186425
rect 150898 186351 150954 186360
rect 150544 186238 150756 186266
rect 150164 185632 150216 185638
rect 150164 185574 150216 185580
rect 150624 184612 150676 184618
rect 150624 184554 150676 184560
rect 150348 183048 150400 183054
rect 150348 182990 150400 182996
rect 149980 182028 150032 182034
rect 149980 181970 150032 181976
rect 149704 178764 149756 178770
rect 149704 178706 149756 178712
rect 149716 148170 149744 178706
rect 149704 148164 149756 148170
rect 149704 148106 149756 148112
rect 149612 145716 149664 145722
rect 149612 145658 149664 145664
rect 149428 144492 149480 144498
rect 149428 144434 149480 144440
rect 148322 142760 148378 142769
rect 148322 142695 148378 142704
rect 148232 140072 148284 140078
rect 148232 140014 148284 140020
rect 148336 139890 148364 142695
rect 149058 141536 149114 141545
rect 149058 141471 149114 141480
rect 149072 139890 149100 141471
rect 149440 139890 149468 144434
rect 149978 142896 150034 142905
rect 149978 142831 150034 142840
rect 149992 139890 150020 142831
rect 150360 140185 150388 182990
rect 150532 181212 150584 181218
rect 150532 181154 150584 181160
rect 150544 144566 150572 181154
rect 150636 145926 150664 184554
rect 150728 148714 150756 186238
rect 151004 184618 151032 199736
rect 151326 199764 151354 200124
rect 151418 199918 151446 200124
rect 151406 199912 151458 199918
rect 151406 199854 151458 199860
rect 151176 199718 151228 199724
rect 151280 199736 151354 199764
rect 151510 199764 151538 200124
rect 151602 199918 151630 200124
rect 151694 199918 151722 200124
rect 151590 199912 151642 199918
rect 151590 199854 151642 199860
rect 151682 199912 151734 199918
rect 151682 199854 151734 199860
rect 151786 199764 151814 200124
rect 151510 199736 151584 199764
rect 151084 199640 151136 199646
rect 151084 199582 151136 199588
rect 150992 184612 151044 184618
rect 150992 184554 151044 184560
rect 150808 184340 150860 184346
rect 150808 184282 150860 184288
rect 150716 148708 150768 148714
rect 150716 148650 150768 148656
rect 150820 148442 150848 184282
rect 151096 171134 151124 199582
rect 151188 199481 151216 199718
rect 151174 199472 151230 199481
rect 151174 199407 151230 199416
rect 151280 184346 151308 199736
rect 151556 199696 151584 199736
rect 151740 199736 151814 199764
rect 151878 199764 151906 200124
rect 151970 199918 151998 200124
rect 152062 199918 152090 200124
rect 151958 199912 152010 199918
rect 151958 199854 152010 199860
rect 152050 199912 152102 199918
rect 152050 199854 152102 199860
rect 152154 199764 152182 200124
rect 151878 199736 152044 199764
rect 151372 199668 151584 199696
rect 151636 199708 151688 199714
rect 151372 199306 151400 199668
rect 151636 199650 151688 199656
rect 151452 199572 151504 199578
rect 151452 199514 151504 199520
rect 151544 199572 151596 199578
rect 151544 199514 151596 199520
rect 151360 199300 151412 199306
rect 151360 199242 151412 199248
rect 151464 185609 151492 199514
rect 151556 193934 151584 199514
rect 151544 193928 151596 193934
rect 151544 193870 151596 193876
rect 151450 185600 151506 185609
rect 151450 185535 151506 185544
rect 151268 184340 151320 184346
rect 151268 184282 151320 184288
rect 151648 181218 151676 199650
rect 151740 199345 151768 199736
rect 151726 199336 151782 199345
rect 151726 199271 151782 199280
rect 151912 185632 151964 185638
rect 151912 185574 151964 185580
rect 152016 185586 152044 199736
rect 152108 199736 152182 199764
rect 152108 185824 152136 199736
rect 152246 199628 152274 200124
rect 152338 199764 152366 200124
rect 152430 199918 152458 200124
rect 152418 199912 152470 199918
rect 152418 199854 152470 199860
rect 152522 199764 152550 200124
rect 152614 199918 152642 200124
rect 152602 199912 152654 199918
rect 152602 199854 152654 199860
rect 152706 199764 152734 200124
rect 152338 199736 152412 199764
rect 152522 199736 152596 199764
rect 152246 199600 152320 199628
rect 152188 199504 152240 199510
rect 152188 199446 152240 199452
rect 152200 195673 152228 199446
rect 152186 195664 152242 195673
rect 152186 195599 152242 195608
rect 152108 185796 152228 185824
rect 151636 181212 151688 181218
rect 151636 181154 151688 181160
rect 151096 171106 151216 171134
rect 150808 148436 150860 148442
rect 150808 148378 150860 148384
rect 150624 145920 150676 145926
rect 150624 145862 150676 145868
rect 150532 144560 150584 144566
rect 150532 144502 150584 144508
rect 151188 142154 151216 171106
rect 151268 144356 151320 144362
rect 151268 144298 151320 144304
rect 151096 142126 151216 142154
rect 150530 141400 150586 141409
rect 150530 141335 150586 141344
rect 150346 140176 150402 140185
rect 150346 140111 150402 140120
rect 150544 139890 150572 141335
rect 138400 139862 138736 139890
rect 138952 139862 139288 139890
rect 139504 139862 139840 139890
rect 140056 139862 140392 139890
rect 140792 139862 140944 139890
rect 141160 139862 141496 139890
rect 141712 139862 142048 139890
rect 142264 139862 142600 139890
rect 142816 139862 143152 139890
rect 143552 139862 143704 139890
rect 143920 139862 144256 139890
rect 144472 139862 144808 139890
rect 145116 139862 145360 139890
rect 145576 139862 145912 139890
rect 146312 139862 146464 139890
rect 146680 139862 147016 139890
rect 147232 139862 147568 139890
rect 147784 139862 148120 139890
rect 148336 139862 148672 139890
rect 149072 139862 149224 139890
rect 149440 139862 149776 139890
rect 149992 139862 150328 139890
rect 150544 139862 150880 139890
rect 151096 139369 151124 142126
rect 151280 139890 151308 144298
rect 151924 141438 151952 185574
rect 152016 185558 152136 185586
rect 152004 179988 152056 179994
rect 152004 179930 152056 179936
rect 152016 146985 152044 179930
rect 152108 148306 152136 185558
rect 152200 149054 152228 185796
rect 152292 185609 152320 199600
rect 152384 198937 152412 199736
rect 152464 199640 152516 199646
rect 152464 199582 152516 199588
rect 152370 198928 152426 198937
rect 152370 198863 152426 198872
rect 152476 185638 152504 199582
rect 152464 185632 152516 185638
rect 152278 185600 152334 185609
rect 152568 185609 152596 199736
rect 152660 199736 152734 199764
rect 152464 185574 152516 185580
rect 152554 185600 152610 185609
rect 152278 185535 152334 185544
rect 152554 185535 152610 185544
rect 152660 179994 152688 199736
rect 152798 199696 152826 200124
rect 152890 199764 152918 200124
rect 152982 199918 153010 200124
rect 153074 199923 153102 200124
rect 152970 199912 153022 199918
rect 152970 199854 153022 199860
rect 153060 199914 153116 199923
rect 153060 199849 153116 199858
rect 153166 199764 153194 200124
rect 153258 199918 153286 200124
rect 153246 199912 153298 199918
rect 153246 199854 153298 199860
rect 153350 199850 153378 200124
rect 153338 199844 153390 199850
rect 153338 199786 153390 199792
rect 152890 199736 152964 199764
rect 152752 199668 152826 199696
rect 152752 186425 152780 199668
rect 152832 199572 152884 199578
rect 152832 199514 152884 199520
rect 152738 186416 152794 186425
rect 152738 186351 152794 186360
rect 152648 179988 152700 179994
rect 152648 179930 152700 179936
rect 152844 172514 152872 199514
rect 152936 199073 152964 199736
rect 153120 199736 153194 199764
rect 153442 199764 153470 200124
rect 153534 199918 153562 200124
rect 153626 199918 153654 200124
rect 153522 199912 153574 199918
rect 153522 199854 153574 199860
rect 153614 199912 153666 199918
rect 153614 199854 153666 199860
rect 153568 199776 153620 199782
rect 153442 199736 153516 199764
rect 152922 199064 152978 199073
rect 152922 198999 152978 199008
rect 153120 196761 153148 199736
rect 153200 199504 153252 199510
rect 153200 199446 153252 199452
rect 153292 199504 153344 199510
rect 153292 199446 153344 199452
rect 153212 198830 153240 199446
rect 153200 198824 153252 198830
rect 153200 198766 153252 198772
rect 153106 196752 153162 196761
rect 153106 196687 153162 196696
rect 153304 194546 153332 199446
rect 153384 199436 153436 199442
rect 153384 199378 153436 199384
rect 153292 194540 153344 194546
rect 153292 194482 153344 194488
rect 153396 192506 153424 199378
rect 153488 194954 153516 199736
rect 153718 199764 153746 200124
rect 153810 199923 153838 200124
rect 153796 199914 153852 199923
rect 153796 199849 153852 199858
rect 153902 199764 153930 200124
rect 153994 199918 154022 200124
rect 154086 199918 154114 200124
rect 154178 199918 154206 200124
rect 154270 199918 154298 200124
rect 153982 199912 154034 199918
rect 153982 199854 154034 199860
rect 154074 199912 154126 199918
rect 154074 199854 154126 199860
rect 154166 199912 154218 199918
rect 154166 199854 154218 199860
rect 154258 199912 154310 199918
rect 154258 199854 154310 199860
rect 153718 199736 153792 199764
rect 153568 199718 153620 199724
rect 153476 194948 153528 194954
rect 153476 194890 153528 194896
rect 153384 192500 153436 192506
rect 153384 192442 153436 192448
rect 153290 186280 153346 186289
rect 153290 186215 153346 186224
rect 152660 172486 152872 172514
rect 152188 149048 152240 149054
rect 152188 148990 152240 148996
rect 152096 148300 152148 148306
rect 152096 148242 152148 148248
rect 152002 146976 152058 146985
rect 152002 146911 152058 146920
rect 152278 142760 152334 142769
rect 152278 142695 152334 142704
rect 151912 141432 151964 141438
rect 151912 141374 151964 141380
rect 152292 139890 152320 142695
rect 152660 142154 152688 172486
rect 153304 145625 153332 186215
rect 153384 185632 153436 185638
rect 153384 185574 153436 185580
rect 153396 149841 153424 185574
rect 153580 178770 153608 199718
rect 153660 199640 153712 199646
rect 153660 199582 153712 199588
rect 153672 186289 153700 199582
rect 153764 196625 153792 199736
rect 153856 199736 153930 199764
rect 154120 199776 154172 199782
rect 153750 196616 153806 196625
rect 153750 196551 153806 196560
rect 153856 186425 153884 199736
rect 154120 199718 154172 199724
rect 154212 199776 154264 199782
rect 154362 199764 154390 200124
rect 154454 199923 154482 200124
rect 154440 199914 154496 199923
rect 154546 199918 154574 200124
rect 154638 199918 154666 200124
rect 154440 199849 154496 199858
rect 154534 199912 154586 199918
rect 154534 199854 154586 199860
rect 154626 199912 154678 199918
rect 154626 199854 154678 199860
rect 154488 199776 154540 199782
rect 154362 199736 154436 199764
rect 154212 199718 154264 199724
rect 154028 199708 154080 199714
rect 154028 199650 154080 199656
rect 154040 196761 154068 199650
rect 154026 196752 154082 196761
rect 154026 196687 154082 196696
rect 153842 186416 153898 186425
rect 153842 186351 153898 186360
rect 153658 186280 153714 186289
rect 153658 186215 153714 186224
rect 153936 185700 153988 185706
rect 153936 185642 153988 185648
rect 153568 178764 153620 178770
rect 153568 178706 153620 178712
rect 153382 149832 153438 149841
rect 153382 149767 153438 149776
rect 153290 145616 153346 145625
rect 153290 145551 153346 145560
rect 153108 144356 153160 144362
rect 153108 144298 153160 144304
rect 151280 139862 151432 139890
rect 151984 139862 152320 139890
rect 152384 142126 152688 142154
rect 152384 139369 152412 142126
rect 152830 141400 152886 141409
rect 152830 141335 152886 141344
rect 152844 139890 152872 141335
rect 153120 140162 153148 144298
rect 153842 142896 153898 142905
rect 153842 142831 153898 142840
rect 152536 139862 152872 139890
rect 153074 140134 153148 140162
rect 153074 139876 153102 140134
rect 153856 139890 153884 142831
rect 153948 140185 153976 185642
rect 154132 185638 154160 199718
rect 154120 185632 154172 185638
rect 154224 185609 154252 199718
rect 154304 199640 154356 199646
rect 154304 199582 154356 199588
rect 154316 197305 154344 199582
rect 154302 197296 154358 197305
rect 154302 197231 154358 197240
rect 154408 185706 154436 199736
rect 154488 199718 154540 199724
rect 154580 199776 154632 199782
rect 154730 199764 154758 200124
rect 154580 199718 154632 199724
rect 154684 199736 154758 199764
rect 154500 197266 154528 199718
rect 154488 197260 154540 197266
rect 154488 197202 154540 197208
rect 154592 196897 154620 199718
rect 154578 196888 154634 196897
rect 154578 196823 154634 196832
rect 154684 193730 154712 199736
rect 154822 199696 154850 200124
rect 154914 199918 154942 200124
rect 155006 199923 155034 200124
rect 154902 199912 154954 199918
rect 154902 199854 154954 199860
rect 154992 199914 155048 199923
rect 155098 199918 155126 200124
rect 155190 199918 155218 200124
rect 155282 199918 155310 200124
rect 154992 199849 155048 199858
rect 155086 199912 155138 199918
rect 155086 199854 155138 199860
rect 155178 199912 155230 199918
rect 155178 199854 155230 199860
rect 155270 199912 155322 199918
rect 155270 199854 155322 199860
rect 155132 199776 155184 199782
rect 155132 199718 155184 199724
rect 155224 199776 155276 199782
rect 155224 199718 155276 199724
rect 154776 199668 154850 199696
rect 154776 196518 154804 199668
rect 155040 199640 155092 199646
rect 155040 199582 155092 199588
rect 154764 196512 154816 196518
rect 154764 196454 154816 196460
rect 155052 194041 155080 199582
rect 155144 198626 155172 199718
rect 155132 198620 155184 198626
rect 155132 198562 155184 198568
rect 155038 194032 155094 194041
rect 155038 193967 155094 193976
rect 154672 193724 154724 193730
rect 154672 193666 154724 193672
rect 154856 186448 154908 186454
rect 154856 186390 154908 186396
rect 154488 185836 154540 185842
rect 154488 185778 154540 185784
rect 154396 185700 154448 185706
rect 154396 185642 154448 185648
rect 154120 185574 154172 185580
rect 154210 185600 154266 185609
rect 154210 185535 154266 185544
rect 154500 145722 154528 185778
rect 154764 185632 154816 185638
rect 154764 185574 154816 185580
rect 154488 145716 154540 145722
rect 154488 145658 154540 145664
rect 154028 144424 154080 144430
rect 154028 144366 154080 144372
rect 153934 140176 153990 140185
rect 153934 140111 153990 140120
rect 153640 139862 153884 139890
rect 154040 139890 154068 144366
rect 154776 140321 154804 185574
rect 154868 149705 154896 186390
rect 155236 182714 155264 199718
rect 155374 199696 155402 200124
rect 155466 199764 155494 200124
rect 155558 199918 155586 200124
rect 155650 199923 155678 200124
rect 155546 199912 155598 199918
rect 155546 199854 155598 199860
rect 155636 199914 155692 199923
rect 155636 199849 155692 199858
rect 155742 199764 155770 200124
rect 155466 199736 155540 199764
rect 155328 199668 155402 199696
rect 155328 197606 155356 199668
rect 155408 199572 155460 199578
rect 155408 199514 155460 199520
rect 155316 197600 155368 197606
rect 155316 197542 155368 197548
rect 155420 185609 155448 199514
rect 155512 186454 155540 199736
rect 155696 199736 155770 199764
rect 155592 199572 155644 199578
rect 155592 199514 155644 199520
rect 155500 186448 155552 186454
rect 155500 186390 155552 186396
rect 155500 185700 155552 185706
rect 155500 185642 155552 185648
rect 155406 185600 155462 185609
rect 155406 185535 155462 185544
rect 155224 182708 155276 182714
rect 155224 182650 155276 182656
rect 154854 149696 154910 149705
rect 154854 149631 154910 149640
rect 155406 143032 155462 143041
rect 155406 142967 155462 142976
rect 155040 142860 155092 142866
rect 155040 142802 155092 142808
rect 154762 140312 154818 140321
rect 154762 140247 154818 140256
rect 155052 139890 155080 142802
rect 155420 139890 155448 142967
rect 154040 139862 154192 139890
rect 154744 139862 155080 139890
rect 155296 139862 155448 139890
rect 155512 139398 155540 185642
rect 155604 171134 155632 199514
rect 155696 185638 155724 199736
rect 155834 199696 155862 200124
rect 155926 199764 155954 200124
rect 156018 199923 156046 200124
rect 156004 199914 156060 199923
rect 156004 199849 156060 199858
rect 156110 199764 156138 200124
rect 156202 199918 156230 200124
rect 156294 199918 156322 200124
rect 156386 199918 156414 200124
rect 156478 199923 156506 200124
rect 156190 199912 156242 199918
rect 156190 199854 156242 199860
rect 156282 199912 156334 199918
rect 156282 199854 156334 199860
rect 156374 199912 156426 199918
rect 156374 199854 156426 199860
rect 156464 199914 156520 199923
rect 156464 199849 156520 199858
rect 156236 199776 156288 199782
rect 155926 199753 156000 199764
rect 155926 199744 156014 199753
rect 155926 199736 155958 199744
rect 155788 199668 155862 199696
rect 156110 199736 156184 199764
rect 155958 199679 156014 199688
rect 155788 185706 155816 199668
rect 156156 193186 156184 199736
rect 156236 199718 156288 199724
rect 156328 199776 156380 199782
rect 156570 199764 156598 200124
rect 156328 199718 156380 199724
rect 156524 199736 156598 199764
rect 156662 199764 156690 200124
rect 156754 199918 156782 200124
rect 156742 199912 156794 199918
rect 156742 199854 156794 199860
rect 156846 199764 156874 200124
rect 156662 199753 156736 199764
rect 156662 199744 156750 199753
rect 156662 199736 156694 199744
rect 156248 195906 156276 199718
rect 156236 195900 156288 195906
rect 156236 195842 156288 195848
rect 156144 193180 156196 193186
rect 156144 193122 156196 193128
rect 156050 186280 156106 186289
rect 156050 186215 156106 186224
rect 155776 185700 155828 185706
rect 155776 185642 155828 185648
rect 155684 185632 155736 185638
rect 155684 185574 155736 185580
rect 155604 171106 155724 171134
rect 155132 139392 155184 139398
rect 123668 139334 123720 139340
rect 124126 139360 124182 139369
rect 122930 139295 122986 139304
rect 124126 139295 124182 139304
rect 126886 139360 126942 139369
rect 126886 139295 126942 139304
rect 129646 139360 129702 139369
rect 129646 139295 129702 139304
rect 131670 139360 131726 139369
rect 131670 139295 131726 139304
rect 132222 139360 132278 139369
rect 132222 139295 132278 139304
rect 138294 139360 138350 139369
rect 138294 139295 138350 139304
rect 151082 139360 151138 139369
rect 151082 139295 151138 139304
rect 152370 139360 152426 139369
rect 152370 139295 152426 139304
rect 155130 139360 155132 139369
rect 155500 139392 155552 139398
rect 155184 139360 155186 139369
rect 155696 139369 155724 171106
rect 156064 150385 156092 186215
rect 156144 185632 156196 185638
rect 156144 185574 156196 185580
rect 156156 152561 156184 185574
rect 156340 183054 156368 199718
rect 156420 199708 156472 199714
rect 156420 199650 156472 199656
rect 156432 192953 156460 199650
rect 156418 192944 156474 192953
rect 156418 192879 156474 192888
rect 156328 183048 156380 183054
rect 156328 182990 156380 182996
rect 156524 171134 156552 199736
rect 156694 199679 156750 199688
rect 156800 199736 156874 199764
rect 156938 199764 156966 200124
rect 157030 199918 157058 200124
rect 157122 199918 157150 200124
rect 157214 199923 157242 200124
rect 157018 199912 157070 199918
rect 157018 199854 157070 199860
rect 157110 199912 157162 199918
rect 157110 199854 157162 199860
rect 157200 199914 157256 199923
rect 157200 199849 157256 199858
rect 157064 199776 157116 199782
rect 156938 199736 157012 199764
rect 156696 199640 156748 199646
rect 156696 199582 156748 199588
rect 156708 197198 156736 199582
rect 156696 197192 156748 197198
rect 156696 197134 156748 197140
rect 156800 185570 156828 199736
rect 156984 185609 157012 199736
rect 157306 199764 157334 200124
rect 157398 199918 157426 200124
rect 157386 199912 157438 199918
rect 157386 199854 157438 199860
rect 157490 199764 157518 200124
rect 157582 199918 157610 200124
rect 157674 199918 157702 200124
rect 157766 199918 157794 200124
rect 157570 199912 157622 199918
rect 157570 199854 157622 199860
rect 157662 199912 157714 199918
rect 157662 199854 157714 199860
rect 157754 199912 157806 199918
rect 157754 199854 157806 199860
rect 157064 199718 157116 199724
rect 157154 199744 157210 199753
rect 157076 185638 157104 199718
rect 157306 199736 157380 199764
rect 157490 199736 157564 199764
rect 157154 199679 157156 199688
rect 157208 199679 157210 199688
rect 157156 199650 157208 199656
rect 157352 195634 157380 199736
rect 157340 195628 157392 195634
rect 157340 195570 157392 195576
rect 157536 193089 157564 199736
rect 157858 199730 157886 200124
rect 157950 199918 157978 200124
rect 158042 199923 158070 200124
rect 157938 199912 157990 199918
rect 157938 199854 157990 199860
rect 158028 199914 158084 199923
rect 158028 199849 158084 199858
rect 158134 199764 158162 200124
rect 158088 199736 158162 199764
rect 157708 199708 157760 199714
rect 157858 199702 158024 199730
rect 157708 199650 157760 199656
rect 157720 199594 157748 199650
rect 157892 199640 157944 199646
rect 157720 199566 157840 199594
rect 157892 199582 157944 199588
rect 157708 199504 157760 199510
rect 157708 199446 157760 199452
rect 157720 196654 157748 199446
rect 157708 196648 157760 196654
rect 157708 196590 157760 196596
rect 157522 193080 157578 193089
rect 157522 193015 157578 193024
rect 157812 186250 157840 199566
rect 157800 186244 157852 186250
rect 157800 186186 157852 186192
rect 157064 185632 157116 185638
rect 156970 185600 157026 185609
rect 156788 185564 156840 185570
rect 157064 185574 157116 185580
rect 157524 185632 157576 185638
rect 157524 185574 157576 185580
rect 156970 185535 157026 185544
rect 157248 185564 157300 185570
rect 156788 185506 156840 185512
rect 157248 185506 157300 185512
rect 156248 171106 156552 171134
rect 156142 152552 156198 152561
rect 156142 152487 156198 152496
rect 156050 150376 156106 150385
rect 156050 150311 156106 150320
rect 156248 150249 156276 171106
rect 156234 150240 156290 150249
rect 156234 150175 156290 150184
rect 157260 147121 157288 185506
rect 157432 179852 157484 179858
rect 157432 179794 157484 179800
rect 157246 147112 157302 147121
rect 157246 147047 157302 147056
rect 157444 145790 157472 179794
rect 157536 152697 157564 185574
rect 157904 179858 157932 199582
rect 157996 196994 158024 199702
rect 157984 196988 158036 196994
rect 157984 196930 158036 196936
rect 158088 195294 158116 199736
rect 158226 199696 158254 200124
rect 158318 199923 158346 200124
rect 158304 199914 158360 199923
rect 158410 199918 158438 200124
rect 158304 199849 158360 199858
rect 158398 199912 158450 199918
rect 158398 199854 158450 199860
rect 158352 199776 158404 199782
rect 158502 199764 158530 200124
rect 158594 199923 158622 200124
rect 158580 199914 158636 199923
rect 158580 199849 158636 199858
rect 158686 199764 158714 200124
rect 158778 199918 158806 200124
rect 158766 199912 158818 199918
rect 158766 199854 158818 199860
rect 158870 199764 158898 200124
rect 158962 199918 158990 200124
rect 158950 199912 159002 199918
rect 158950 199854 159002 199860
rect 159054 199764 159082 200124
rect 158352 199718 158404 199724
rect 158456 199736 158530 199764
rect 158640 199736 158714 199764
rect 158824 199736 158898 199764
rect 159008 199736 159082 199764
rect 158180 199668 158254 199696
rect 158076 195288 158128 195294
rect 158076 195230 158128 195236
rect 158180 185881 158208 199668
rect 158260 199572 158312 199578
rect 158260 199514 158312 199520
rect 158272 186289 158300 199514
rect 158364 195362 158392 199718
rect 158352 195356 158404 195362
rect 158352 195298 158404 195304
rect 158258 186280 158314 186289
rect 158258 186215 158314 186224
rect 158166 185872 158222 185881
rect 158166 185807 158222 185816
rect 158456 185638 158484 199736
rect 158536 199368 158588 199374
rect 158536 199310 158588 199316
rect 158444 185632 158496 185638
rect 158444 185574 158496 185580
rect 157892 179852 157944 179858
rect 157892 179794 157944 179800
rect 157522 152688 157578 152697
rect 157522 152623 157578 152632
rect 158548 145858 158576 199310
rect 158640 199170 158668 199736
rect 158824 199696 158852 199736
rect 158732 199668 158852 199696
rect 158628 199164 158680 199170
rect 158628 199106 158680 199112
rect 158732 185609 158760 199668
rect 158904 199640 158956 199646
rect 158904 199582 158956 199588
rect 158812 199572 158864 199578
rect 158812 199514 158864 199520
rect 158824 185842 158852 199514
rect 158916 196586 158944 199582
rect 158904 196580 158956 196586
rect 158904 196522 158956 196528
rect 159008 192488 159036 199736
rect 159146 199696 159174 200124
rect 159100 199668 159174 199696
rect 159238 199696 159266 200124
rect 159330 199764 159358 200124
rect 159422 199918 159450 200124
rect 159514 199918 159542 200124
rect 159410 199912 159462 199918
rect 159410 199854 159462 199860
rect 159502 199912 159554 199918
rect 159502 199854 159554 199860
rect 159456 199776 159508 199782
rect 159330 199736 159404 199764
rect 159238 199668 159312 199696
rect 159100 192681 159128 199668
rect 159180 199572 159232 199578
rect 159180 199514 159232 199520
rect 159086 192672 159142 192681
rect 159086 192607 159142 192616
rect 159008 192460 159128 192488
rect 158904 186312 158956 186318
rect 158904 186254 158956 186260
rect 158812 185836 158864 185842
rect 158812 185778 158864 185784
rect 158812 185700 158864 185706
rect 158812 185642 158864 185648
rect 158718 185600 158774 185609
rect 158718 185535 158774 185544
rect 158536 145852 158588 145858
rect 158536 145794 158588 145800
rect 157432 145784 157484 145790
rect 158824 145761 158852 185642
rect 158916 152930 158944 186254
rect 158996 175228 159048 175234
rect 158996 175170 159048 175176
rect 159008 152998 159036 175170
rect 159100 153134 159128 192460
rect 159192 179489 159220 199514
rect 159284 195770 159312 199668
rect 159272 195764 159324 195770
rect 159272 195706 159324 195712
rect 159178 179480 159234 179489
rect 159178 179415 159234 179424
rect 159376 175234 159404 199736
rect 159606 199764 159634 200124
rect 159698 199923 159726 200124
rect 159684 199914 159740 199923
rect 159684 199849 159740 199858
rect 159790 199764 159818 200124
rect 159456 199718 159508 199724
rect 159560 199736 159634 199764
rect 159744 199736 159818 199764
rect 159468 196790 159496 199718
rect 159456 196784 159508 196790
rect 159456 196726 159508 196732
rect 159560 186318 159588 199736
rect 159744 197554 159772 199736
rect 159882 199696 159910 200124
rect 159652 197526 159772 197554
rect 159836 199668 159910 199696
rect 159652 195838 159680 197526
rect 159640 195832 159692 195838
rect 159640 195774 159692 195780
rect 159548 186312 159600 186318
rect 159548 186254 159600 186260
rect 159836 185706 159864 199668
rect 159974 199628 160002 200124
rect 160066 199764 160094 200124
rect 160158 199923 160186 200124
rect 160144 199914 160200 199923
rect 160144 199849 160200 199858
rect 160250 199850 160278 200124
rect 160342 199918 160370 200124
rect 160434 199918 160462 200124
rect 160330 199912 160382 199918
rect 160330 199854 160382 199860
rect 160422 199912 160474 199918
rect 160422 199854 160474 199860
rect 160238 199844 160290 199850
rect 160238 199786 160290 199792
rect 160526 199764 160554 200124
rect 160618 199918 160646 200124
rect 160606 199912 160658 199918
rect 160606 199854 160658 199860
rect 160710 199764 160738 200124
rect 160066 199736 160140 199764
rect 160526 199736 160600 199764
rect 159928 199600 160002 199628
rect 159824 185700 159876 185706
rect 159824 185642 159876 185648
rect 159364 175228 159416 175234
rect 159364 175170 159416 175176
rect 159928 172514 159956 199600
rect 160112 195498 160140 199736
rect 160192 199708 160244 199714
rect 160192 199650 160244 199656
rect 160100 195492 160152 195498
rect 160100 195434 160152 195440
rect 160008 186652 160060 186658
rect 160008 186594 160060 186600
rect 159836 172486 159956 172514
rect 159088 153128 159140 153134
rect 159088 153070 159140 153076
rect 158996 152992 159048 152998
rect 158996 152934 159048 152940
rect 158904 152924 158956 152930
rect 158904 152866 158956 152872
rect 157432 145726 157484 145732
rect 158810 145752 158866 145761
rect 158810 145687 158866 145696
rect 158352 144560 158404 144566
rect 158352 144502 158404 144508
rect 157800 144492 157852 144498
rect 157800 144434 157852 144440
rect 156696 144424 156748 144430
rect 156696 144366 156748 144372
rect 155868 142180 155920 142186
rect 155868 142122 155920 142128
rect 155880 140162 155908 142122
rect 155834 140134 155908 140162
rect 155834 139876 155862 140134
rect 156708 139890 156736 144366
rect 157706 144120 157762 144129
rect 157706 144055 157762 144064
rect 157246 143168 157302 143177
rect 157246 143103 157302 143112
rect 157260 139890 157288 143103
rect 157720 142866 157748 144055
rect 157708 142860 157760 142866
rect 157708 142802 157760 142808
rect 157340 142180 157392 142186
rect 157340 142122 157392 142128
rect 157352 142089 157380 142122
rect 157338 142080 157394 142089
rect 157338 142015 157394 142024
rect 157812 139890 157840 144434
rect 158364 139890 158392 144502
rect 158628 142860 158680 142866
rect 158628 142802 158680 142808
rect 158640 140162 158668 142802
rect 159456 142180 159508 142186
rect 159836 142154 159864 172486
rect 159916 144288 159968 144294
rect 159916 144230 159968 144236
rect 159456 142122 159508 142128
rect 159560 142126 159864 142154
rect 156400 139862 156736 139890
rect 156952 139862 157288 139890
rect 157504 139862 157840 139890
rect 158056 139862 158392 139890
rect 158594 140134 158668 140162
rect 158594 139876 158622 140134
rect 159468 139890 159496 142122
rect 159160 139862 159496 139890
rect 159560 139369 159588 142126
rect 159928 139890 159956 144230
rect 159712 139862 159956 139890
rect 160020 139369 160048 186594
rect 160204 186153 160232 199650
rect 160284 199640 160336 199646
rect 160468 199640 160520 199646
rect 160284 199582 160336 199588
rect 160374 199608 160430 199617
rect 160296 196858 160324 199582
rect 160468 199582 160520 199588
rect 160374 199543 160430 199552
rect 160284 196852 160336 196858
rect 160284 196794 160336 196800
rect 160388 195430 160416 199543
rect 160376 195424 160428 195430
rect 160376 195366 160428 195372
rect 160480 186402 160508 199582
rect 160388 186374 160508 186402
rect 160190 186144 160246 186153
rect 160190 186079 160246 186088
rect 160100 185632 160152 185638
rect 160100 185574 160152 185580
rect 160112 140078 160140 185574
rect 160284 185020 160336 185026
rect 160284 184962 160336 184968
rect 160192 181484 160244 181490
rect 160192 181426 160244 181432
rect 160204 145926 160232 181426
rect 160296 153066 160324 184962
rect 160388 153202 160416 186374
rect 160466 186280 160522 186289
rect 160466 186215 160522 186224
rect 160376 153196 160428 153202
rect 160376 153138 160428 153144
rect 160284 153060 160336 153066
rect 160284 153002 160336 153008
rect 160480 152454 160508 186215
rect 160572 178537 160600 199736
rect 160664 199736 160738 199764
rect 160664 185026 160692 199736
rect 160802 199696 160830 200124
rect 160894 199923 160922 200124
rect 160880 199914 160936 199923
rect 160880 199849 160936 199858
rect 160986 199850 161014 200124
rect 160974 199844 161026 199850
rect 160974 199786 161026 199792
rect 161078 199730 161106 200124
rect 161170 199782 161198 200124
rect 161262 199782 161290 200124
rect 161354 199923 161382 200124
rect 161340 199914 161396 199923
rect 161340 199849 161396 199858
rect 160756 199668 160830 199696
rect 160928 199708 160980 199714
rect 160652 185020 160704 185026
rect 160652 184962 160704 184968
rect 160558 178528 160614 178537
rect 160558 178463 160614 178472
rect 160756 177993 160784 199668
rect 160928 199650 160980 199656
rect 161032 199702 161106 199730
rect 161158 199776 161210 199782
rect 161158 199718 161210 199724
rect 161250 199776 161302 199782
rect 161250 199718 161302 199724
rect 160836 199572 160888 199578
rect 160836 199514 160888 199520
rect 160848 181801 160876 199514
rect 160940 185638 160968 199650
rect 160928 185632 160980 185638
rect 161032 185609 161060 199702
rect 161446 199696 161474 200124
rect 161538 199850 161566 200124
rect 161630 199923 161658 200124
rect 161616 199914 161672 199923
rect 161526 199844 161578 199850
rect 161616 199849 161672 199858
rect 161526 199786 161578 199792
rect 161400 199668 161474 199696
rect 161570 199744 161626 199753
rect 161570 199679 161626 199688
rect 161296 199572 161348 199578
rect 161296 199514 161348 199520
rect 160928 185574 160980 185580
rect 161018 185600 161074 185609
rect 161018 185535 161074 185544
rect 160834 181792 160890 181801
rect 160834 181727 160890 181736
rect 161308 181490 161336 199514
rect 161400 191690 161428 199668
rect 161480 199572 161532 199578
rect 161480 199514 161532 199520
rect 161388 191684 161440 191690
rect 161388 191626 161440 191632
rect 161388 185632 161440 185638
rect 161388 185574 161440 185580
rect 161296 181484 161348 181490
rect 161296 181426 161348 181432
rect 161296 179172 161348 179178
rect 161296 179114 161348 179120
rect 160742 177984 160798 177993
rect 160742 177919 160798 177928
rect 161308 171193 161336 179114
rect 161294 171184 161350 171193
rect 161294 171119 161350 171128
rect 161294 171048 161350 171057
rect 161294 170983 161350 170992
rect 161308 161537 161336 170983
rect 161294 161528 161350 161537
rect 161294 161463 161350 161472
rect 161294 161392 161350 161401
rect 161294 161327 161350 161336
rect 160468 152448 160520 152454
rect 160468 152390 160520 152396
rect 161308 151881 161336 161327
rect 161294 151872 161350 151881
rect 161294 151807 161350 151816
rect 161294 151736 161350 151745
rect 161294 151671 161350 151680
rect 160192 145920 160244 145926
rect 160192 145862 160244 145868
rect 160926 145616 160982 145625
rect 160926 145551 160982 145560
rect 160560 142928 160612 142934
rect 160560 142870 160612 142876
rect 160100 140072 160152 140078
rect 160100 140014 160152 140020
rect 160572 139890 160600 142870
rect 160744 141432 160796 141438
rect 160744 141374 160796 141380
rect 160264 139862 160600 139890
rect 160756 139890 160784 141374
rect 160940 139890 160968 145551
rect 161308 142361 161336 151671
rect 161400 151094 161428 185574
rect 161388 151088 161440 151094
rect 161388 151030 161440 151036
rect 161492 148782 161520 199514
rect 161584 195566 161612 199679
rect 161722 199628 161750 200124
rect 161814 199764 161842 200124
rect 161906 199918 161934 200124
rect 161998 199918 162026 200124
rect 162090 199923 162118 200124
rect 161894 199912 161946 199918
rect 161894 199854 161946 199860
rect 161986 199912 162038 199918
rect 161986 199854 162038 199860
rect 162076 199914 162132 199923
rect 162182 199918 162210 200124
rect 162274 199918 162302 200124
rect 162366 199918 162394 200124
rect 162458 199918 162486 200124
rect 162550 199918 162578 200124
rect 162642 199923 162670 200124
rect 162076 199849 162132 199858
rect 162170 199912 162222 199918
rect 162170 199854 162222 199860
rect 162262 199912 162314 199918
rect 162262 199854 162314 199860
rect 162354 199912 162406 199918
rect 162354 199854 162406 199860
rect 162446 199912 162498 199918
rect 162446 199854 162498 199860
rect 162538 199912 162590 199918
rect 162538 199854 162590 199860
rect 162628 199914 162684 199923
rect 162628 199849 162684 199858
rect 161940 199776 161992 199782
rect 161814 199736 161888 199764
rect 161676 199600 161750 199628
rect 161572 195560 161624 195566
rect 161572 195502 161624 195508
rect 161676 193361 161704 199600
rect 161662 193352 161718 193361
rect 161662 193287 161718 193296
rect 161572 186312 161624 186318
rect 161572 186254 161624 186260
rect 161584 148986 161612 186254
rect 161664 179988 161716 179994
rect 161664 179930 161716 179936
rect 161676 152318 161704 179930
rect 161860 172514 161888 199736
rect 162584 199776 162636 199782
rect 162122 199744 162178 199753
rect 161940 199718 161992 199724
rect 161952 196722 161980 199718
rect 162044 199702 162122 199730
rect 161940 196716 161992 196722
rect 161940 196658 161992 196664
rect 162044 186318 162072 199702
rect 162734 199764 162762 200124
rect 162826 199918 162854 200124
rect 162814 199912 162866 199918
rect 162814 199854 162866 199860
rect 162918 199782 162946 200124
rect 163010 199889 163038 200124
rect 162996 199880 163052 199889
rect 163102 199850 163130 200124
rect 163194 199850 163222 200124
rect 163286 199923 163314 200124
rect 163272 199914 163328 199923
rect 163378 199918 163406 200124
rect 162996 199815 163052 199824
rect 163090 199844 163142 199850
rect 163090 199786 163142 199792
rect 163182 199844 163234 199850
rect 163272 199849 163328 199858
rect 163366 199912 163418 199918
rect 163470 199889 163498 200124
rect 163562 199918 163590 200124
rect 163654 199918 163682 200124
rect 163746 199923 163774 200124
rect 163550 199912 163602 199918
rect 163366 199854 163418 199860
rect 163456 199880 163512 199889
rect 163550 199854 163602 199860
rect 163642 199912 163694 199918
rect 163642 199854 163694 199860
rect 163732 199914 163788 199923
rect 163732 199849 163788 199858
rect 163838 199850 163866 200124
rect 163456 199815 163512 199824
rect 163826 199844 163878 199850
rect 163182 199786 163234 199792
rect 163826 199786 163878 199792
rect 162584 199718 162636 199724
rect 162688 199736 162762 199764
rect 162906 199776 162958 199782
rect 162122 199679 162178 199688
rect 162216 199708 162268 199714
rect 162216 199650 162268 199656
rect 162308 199708 162360 199714
rect 162308 199650 162360 199656
rect 162492 199708 162544 199714
rect 162492 199650 162544 199656
rect 162124 199640 162176 199646
rect 162124 199582 162176 199588
rect 162032 186312 162084 186318
rect 162032 186254 162084 186260
rect 162136 179178 162164 199582
rect 162228 197130 162256 199650
rect 162216 197124 162268 197130
rect 162216 197066 162268 197072
rect 162216 192500 162268 192506
rect 162216 192442 162268 192448
rect 162124 179172 162176 179178
rect 162124 179114 162176 179120
rect 161768 172486 161888 172514
rect 161768 152386 161796 172486
rect 161756 152380 161808 152386
rect 161756 152322 161808 152328
rect 161664 152312 161716 152318
rect 161664 152254 161716 152260
rect 161572 148980 161624 148986
rect 161572 148922 161624 148928
rect 161480 148776 161532 148782
rect 161480 148718 161532 148724
rect 162228 145994 162256 192442
rect 162320 179994 162348 199650
rect 162398 199608 162454 199617
rect 162398 199543 162454 199552
rect 162412 199306 162440 199543
rect 162400 199300 162452 199306
rect 162400 199242 162452 199248
rect 162504 186289 162532 199650
rect 162596 193322 162624 199718
rect 162584 193316 162636 193322
rect 162584 193258 162636 193264
rect 162688 186425 162716 199736
rect 162906 199718 162958 199724
rect 163688 199776 163740 199782
rect 163688 199718 163740 199724
rect 163778 199744 163834 199753
rect 163136 199708 163188 199714
rect 163136 199650 163188 199656
rect 163412 199708 163464 199714
rect 163412 199650 163464 199656
rect 163044 199640 163096 199646
rect 163044 199582 163096 199588
rect 162952 199572 163004 199578
rect 162952 199514 163004 199520
rect 162766 198384 162822 198393
rect 162766 198319 162822 198328
rect 162674 186416 162730 186425
rect 162674 186351 162730 186360
rect 162490 186280 162546 186289
rect 162490 186215 162546 186224
rect 162308 179988 162360 179994
rect 162308 179930 162360 179936
rect 162780 179081 162808 198319
rect 162964 198257 162992 199514
rect 162950 198248 163006 198257
rect 162860 198212 162912 198218
rect 162950 198183 163006 198192
rect 162860 198154 162912 198160
rect 162872 192545 162900 198154
rect 162950 198112 163006 198121
rect 162950 198047 163006 198056
rect 162858 192536 162914 192545
rect 162858 192471 162914 192480
rect 162766 179072 162822 179081
rect 162766 179007 162822 179016
rect 162964 149054 162992 198047
rect 163056 197334 163084 199582
rect 163044 197328 163096 197334
rect 163044 197270 163096 197276
rect 163148 186538 163176 199650
rect 163320 199572 163372 199578
rect 163320 199514 163372 199520
rect 163332 198218 163360 199514
rect 163320 198212 163372 198218
rect 163320 198154 163372 198160
rect 163318 198112 163374 198121
rect 163318 198047 163374 198056
rect 163228 197804 163280 197810
rect 163228 197746 163280 197752
rect 163240 186969 163268 197746
rect 163226 186960 163282 186969
rect 163226 186895 163282 186904
rect 163226 186824 163282 186833
rect 163226 186759 163282 186768
rect 163056 186510 163176 186538
rect 162952 149048 163004 149054
rect 162952 148990 163004 148996
rect 163056 148850 163084 186510
rect 163136 179172 163188 179178
rect 163136 179114 163188 179120
rect 163044 148844 163096 148850
rect 163044 148786 163096 148792
rect 163148 148345 163176 179114
rect 163240 152862 163268 186759
rect 163332 186425 163360 198047
rect 163424 186998 163452 199650
rect 163504 199640 163556 199646
rect 163504 199582 163556 199588
rect 163412 186992 163464 186998
rect 163412 186934 163464 186940
rect 163318 186416 163374 186425
rect 163318 186351 163374 186360
rect 163516 186153 163544 199582
rect 163596 199572 163648 199578
rect 163596 199514 163648 199520
rect 163608 197810 163636 199514
rect 163596 197804 163648 197810
rect 163596 197746 163648 197752
rect 163700 196926 163728 199718
rect 163930 199730 163958 200124
rect 164022 199918 164050 200124
rect 164114 199918 164142 200124
rect 164206 199918 164234 200124
rect 164298 199918 164326 200124
rect 164390 199918 164418 200124
rect 164482 199918 164510 200124
rect 164010 199912 164062 199918
rect 164010 199854 164062 199860
rect 164102 199912 164154 199918
rect 164102 199854 164154 199860
rect 164194 199912 164246 199918
rect 164194 199854 164246 199860
rect 164286 199912 164338 199918
rect 164286 199854 164338 199860
rect 164378 199912 164430 199918
rect 164378 199854 164430 199860
rect 164470 199912 164522 199918
rect 164470 199854 164522 199860
rect 164574 199850 164602 200124
rect 164562 199844 164614 199850
rect 164562 199786 164614 199792
rect 164666 199764 164694 200124
rect 164758 199923 164786 200124
rect 164744 199914 164800 199923
rect 164850 199918 164878 200124
rect 164942 199918 164970 200124
rect 165034 199918 165062 200124
rect 165126 199918 165154 200124
rect 165218 199923 165246 200124
rect 164744 199849 164800 199858
rect 164838 199912 164890 199918
rect 164838 199854 164890 199860
rect 164930 199912 164982 199918
rect 164930 199854 164982 199860
rect 165022 199912 165074 199918
rect 165022 199854 165074 199860
rect 165114 199912 165166 199918
rect 165114 199854 165166 199860
rect 165204 199914 165260 199923
rect 165204 199849 165260 199858
rect 164792 199776 164844 199782
rect 164666 199753 164740 199764
rect 164666 199744 164754 199753
rect 164666 199736 164698 199744
rect 163930 199702 164004 199730
rect 163778 199679 163834 199688
rect 163688 196920 163740 196926
rect 163688 196862 163740 196868
rect 163502 186144 163558 186153
rect 163502 186079 163558 186088
rect 163792 179178 163820 199679
rect 163872 199504 163924 199510
rect 163872 199446 163924 199452
rect 163780 179172 163832 179178
rect 163780 179114 163832 179120
rect 163884 172514 163912 199446
rect 163976 187338 164004 199702
rect 164056 199708 164108 199714
rect 164056 199650 164108 199656
rect 164148 199708 164200 199714
rect 164148 199650 164200 199656
rect 164424 199708 164476 199714
rect 164424 199650 164476 199656
rect 164516 199708 164568 199714
rect 165310 199764 165338 200124
rect 164792 199718 164844 199724
rect 165264 199736 165338 199764
rect 164698 199679 164754 199688
rect 164516 199650 164568 199656
rect 163964 187332 164016 187338
rect 163964 187274 164016 187280
rect 164068 186289 164096 199650
rect 164160 192574 164188 199650
rect 164240 199640 164292 199646
rect 164240 199582 164292 199588
rect 164148 192568 164200 192574
rect 164148 192510 164200 192516
rect 164054 186280 164110 186289
rect 164054 186215 164110 186224
rect 164148 185700 164200 185706
rect 164148 185642 164200 185648
rect 163792 172486 163912 172514
rect 163228 152856 163280 152862
rect 163228 152798 163280 152804
rect 163792 151814 163820 172486
rect 163792 151786 164004 151814
rect 163134 148336 163190 148345
rect 163134 148271 163190 148280
rect 162216 145988 162268 145994
rect 162216 145930 162268 145936
rect 162950 145888 163006 145897
rect 162950 145823 163006 145832
rect 162492 144628 162544 144634
rect 162492 144570 162544 144576
rect 162214 143304 162270 143313
rect 162214 143239 162270 143248
rect 161294 142352 161350 142361
rect 161294 142287 161350 142296
rect 162228 139890 162256 143239
rect 162504 142186 162532 144570
rect 162766 144256 162822 144265
rect 162766 144191 162822 144200
rect 162492 142180 162544 142186
rect 162492 142122 162544 142128
rect 162780 139890 162808 144191
rect 160756 139862 160816 139890
rect 160940 139862 161368 139890
rect 161920 139862 162256 139890
rect 162472 139862 162808 139890
rect 162964 139890 162992 145823
rect 163870 143440 163926 143449
rect 163870 143375 163926 143384
rect 163884 139890 163912 143375
rect 162964 139862 163024 139890
rect 163576 139862 163912 139890
rect 163976 139369 164004 151786
rect 164160 147082 164188 185642
rect 164252 182918 164280 199582
rect 164436 183433 164464 199650
rect 164422 183424 164478 183433
rect 164422 183359 164478 183368
rect 164424 183320 164476 183326
rect 164424 183262 164476 183268
rect 164240 182912 164292 182918
rect 164240 182854 164292 182860
rect 164240 182776 164292 182782
rect 164240 182718 164292 182724
rect 164252 148374 164280 182718
rect 164332 175772 164384 175778
rect 164332 175714 164384 175720
rect 164344 148578 164372 175714
rect 164436 148918 164464 183262
rect 164528 152794 164556 199650
rect 164700 199572 164752 199578
rect 164700 199514 164752 199520
rect 164606 198112 164662 198121
rect 164606 198047 164662 198056
rect 164620 186425 164648 198047
rect 164712 193254 164740 199514
rect 164700 193248 164752 193254
rect 164700 193190 164752 193196
rect 164606 186416 164662 186425
rect 164606 186351 164662 186360
rect 164608 182912 164660 182918
rect 164608 182854 164660 182860
rect 164516 152788 164568 152794
rect 164516 152730 164568 152736
rect 164620 152726 164648 182854
rect 164804 175778 164832 199718
rect 164884 199708 164936 199714
rect 164884 199650 164936 199656
rect 164976 199708 165028 199714
rect 164976 199650 165028 199656
rect 165068 199708 165120 199714
rect 165264 199696 165292 199736
rect 165068 199650 165120 199656
rect 165218 199668 165292 199696
rect 164896 186289 164924 199650
rect 164988 193050 165016 199650
rect 164976 193044 165028 193050
rect 164976 192986 165028 192992
rect 164882 186280 164938 186289
rect 164882 186215 164938 186224
rect 165080 182782 165108 199650
rect 165218 199594 165246 199668
rect 165218 199566 165292 199594
rect 165264 192817 165292 199566
rect 165402 199560 165430 200124
rect 165494 199918 165522 200124
rect 165482 199912 165534 199918
rect 165482 199854 165534 199860
rect 165586 199696 165614 200124
rect 165678 199850 165706 200124
rect 165666 199844 165718 199850
rect 165666 199786 165718 199792
rect 165770 199730 165798 200124
rect 165862 199918 165890 200124
rect 165850 199912 165902 199918
rect 165850 199854 165902 199860
rect 165954 199730 165982 200124
rect 166046 199918 166074 200124
rect 166138 199918 166166 200124
rect 166230 199918 166258 200124
rect 166322 199918 166350 200124
rect 166034 199912 166086 199918
rect 166034 199854 166086 199860
rect 166126 199912 166178 199918
rect 166126 199854 166178 199860
rect 166218 199912 166270 199918
rect 166218 199854 166270 199860
rect 166310 199912 166362 199918
rect 166310 199854 166362 199860
rect 165770 199702 165844 199730
rect 165586 199668 165660 199696
rect 165482 199640 165534 199646
rect 165534 199588 165568 199594
rect 165482 199582 165568 199588
rect 165494 199566 165568 199582
rect 165356 199532 165430 199560
rect 165250 192808 165306 192817
rect 165250 192743 165306 192752
rect 165356 183326 165384 199532
rect 165436 199436 165488 199442
rect 165436 199378 165488 199384
rect 165448 199073 165476 199378
rect 165434 199064 165490 199073
rect 165434 198999 165490 199008
rect 165344 183320 165396 183326
rect 165344 183262 165396 183268
rect 165068 182776 165120 182782
rect 165068 182718 165120 182724
rect 165540 178537 165568 199566
rect 165632 189106 165660 199668
rect 165712 199640 165764 199646
rect 165712 199582 165764 199588
rect 165620 189100 165672 189106
rect 165620 189042 165672 189048
rect 165724 185473 165752 199582
rect 165816 190505 165844 199702
rect 165908 199702 165982 199730
rect 166262 199744 166318 199753
rect 166080 199708 166132 199714
rect 165802 190496 165858 190505
rect 165802 190431 165858 190440
rect 165908 185586 165936 199702
rect 166080 199650 166132 199656
rect 166172 199708 166224 199714
rect 166414 199730 166442 200124
rect 166506 199918 166534 200124
rect 166494 199912 166546 199918
rect 166494 199854 166546 199860
rect 166414 199702 166488 199730
rect 166262 199679 166318 199688
rect 166172 199650 166224 199656
rect 165988 199640 166040 199646
rect 165988 199582 166040 199588
rect 166000 185745 166028 199582
rect 166092 192302 166120 199650
rect 166080 192296 166132 192302
rect 166080 192238 166132 192244
rect 165986 185736 166042 185745
rect 165986 185671 166042 185680
rect 165816 185558 165936 185586
rect 165710 185464 165766 185473
rect 165710 185399 165766 185408
rect 165710 185328 165766 185337
rect 165710 185263 165766 185272
rect 165526 178528 165582 178537
rect 165526 178463 165582 178472
rect 164792 175772 164844 175778
rect 164792 175714 164844 175720
rect 164608 152720 164660 152726
rect 164608 152662 164660 152668
rect 164424 148912 164476 148918
rect 164424 148854 164476 148860
rect 164332 148572 164384 148578
rect 164332 148514 164384 148520
rect 165724 148481 165752 185263
rect 165816 155718 165844 185558
rect 166184 172514 166212 199650
rect 166276 199578 166304 199679
rect 166356 199640 166408 199646
rect 166356 199582 166408 199588
rect 166264 199572 166316 199578
rect 166264 199514 166316 199520
rect 166264 199368 166316 199374
rect 166264 199310 166316 199316
rect 166276 197062 166304 199310
rect 166264 197056 166316 197062
rect 166264 196998 166316 197004
rect 166368 180305 166396 199582
rect 166460 192098 166488 199702
rect 166598 199696 166626 200124
rect 166690 199850 166718 200124
rect 166782 199850 166810 200124
rect 166874 199918 166902 200124
rect 166862 199912 166914 199918
rect 166966 199889 166994 200124
rect 166862 199854 166914 199860
rect 166952 199880 167008 199889
rect 166678 199844 166730 199850
rect 166678 199786 166730 199792
rect 166770 199844 166822 199850
rect 166952 199815 167008 199824
rect 166770 199786 166822 199792
rect 166908 199776 166960 199782
rect 166814 199744 166870 199753
rect 166908 199718 166960 199724
rect 166598 199668 166672 199696
rect 166814 199679 166816 199688
rect 166540 199572 166592 199578
rect 166540 199514 166592 199520
rect 166448 192092 166500 192098
rect 166448 192034 166500 192040
rect 166354 180296 166410 180305
rect 166354 180231 166410 180240
rect 165908 172486 166212 172514
rect 165804 155712 165856 155718
rect 165804 155654 165856 155660
rect 165908 155514 165936 172486
rect 166552 171134 166580 199514
rect 166644 185609 166672 199668
rect 166868 199679 166870 199688
rect 166816 199650 166868 199656
rect 166724 199640 166776 199646
rect 166724 199582 166776 199588
rect 166736 193866 166764 199582
rect 166724 193860 166776 193866
rect 166724 193802 166776 193808
rect 166920 185745 166948 199718
rect 167058 199696 167086 200124
rect 167150 199850 167178 200124
rect 167242 199918 167270 200124
rect 167230 199912 167282 199918
rect 167230 199854 167282 199860
rect 167138 199844 167190 199850
rect 167138 199786 167190 199792
rect 167334 199764 167362 200124
rect 167426 199918 167454 200124
rect 167518 199918 167546 200124
rect 167610 199918 167638 200124
rect 167414 199912 167466 199918
rect 167414 199854 167466 199860
rect 167506 199912 167558 199918
rect 167506 199854 167558 199860
rect 167598 199912 167650 199918
rect 167598 199854 167650 199860
rect 167334 199736 167408 199764
rect 167058 199668 167132 199696
rect 166998 198112 167054 198121
rect 166998 198047 167054 198056
rect 167012 195974 167040 198047
rect 167000 195968 167052 195974
rect 167000 195910 167052 195916
rect 166906 185736 166962 185745
rect 166906 185671 166962 185680
rect 166630 185600 166686 185609
rect 167104 185586 167132 199668
rect 167276 199640 167328 199646
rect 167276 199582 167328 199588
rect 167184 199572 167236 199578
rect 167184 199514 167236 199520
rect 167196 198898 167224 199514
rect 167184 198892 167236 198898
rect 167184 198834 167236 198840
rect 167288 185706 167316 199582
rect 167276 185700 167328 185706
rect 167276 185642 167328 185648
rect 167104 185558 167224 185586
rect 166630 185535 166686 185544
rect 167092 176996 167144 177002
rect 167092 176938 167144 176944
rect 166552 171106 166856 171134
rect 165896 155508 165948 155514
rect 165896 155450 165948 155456
rect 166828 148646 166856 171106
rect 167104 148714 167132 176938
rect 167196 155242 167224 185558
rect 167276 185564 167328 185570
rect 167276 185506 167328 185512
rect 167288 155650 167316 185506
rect 167276 155644 167328 155650
rect 167276 155586 167328 155592
rect 167380 155582 167408 199736
rect 167550 199744 167606 199753
rect 167702 199730 167730 200124
rect 167606 199702 167730 199730
rect 167550 199679 167606 199688
rect 167460 199572 167512 199578
rect 167794 199560 167822 200124
rect 167886 199889 167914 200124
rect 167978 199918 168006 200124
rect 168070 199923 168098 200124
rect 167966 199912 168018 199918
rect 167872 199880 167928 199889
rect 167966 199854 168018 199860
rect 168056 199914 168112 199923
rect 168056 199849 168112 199858
rect 168162 199850 168190 200124
rect 168254 199923 168282 200124
rect 168240 199914 168296 199923
rect 168346 199918 168374 200124
rect 167872 199815 167928 199824
rect 168150 199844 168202 199850
rect 168240 199849 168296 199858
rect 168334 199912 168386 199918
rect 168334 199854 168386 199860
rect 168150 199786 168202 199792
rect 168438 199764 168466 200124
rect 168530 199918 168558 200124
rect 168622 199923 168650 200124
rect 168518 199912 168570 199918
rect 168518 199854 168570 199860
rect 168608 199914 168664 199923
rect 168714 199918 168742 200124
rect 168608 199849 168664 199858
rect 168702 199912 168754 199918
rect 168702 199854 168754 199860
rect 168806 199764 168834 200124
rect 168898 199923 168926 200124
rect 168884 199914 168940 199923
rect 168990 199918 169018 200124
rect 169082 199918 169110 200124
rect 169174 199918 169202 200124
rect 168884 199849 168940 199858
rect 168978 199912 169030 199918
rect 168978 199854 169030 199860
rect 169070 199912 169122 199918
rect 169070 199854 169122 199860
rect 169162 199912 169214 199918
rect 169162 199854 169214 199860
rect 169266 199764 169294 200124
rect 169358 199918 169386 200124
rect 169450 199918 169478 200124
rect 169542 199923 169570 200124
rect 169346 199912 169398 199918
rect 169346 199854 169398 199860
rect 169438 199912 169490 199918
rect 169438 199854 169490 199860
rect 169528 199914 169584 199923
rect 169528 199849 169584 199858
rect 168102 199744 168158 199753
rect 168392 199736 168466 199764
rect 168760 199753 168834 199764
rect 168746 199744 168834 199753
rect 168102 199679 168158 199688
rect 168288 199708 168340 199714
rect 167794 199532 167868 199560
rect 167460 199514 167512 199520
rect 167472 192778 167500 199514
rect 167644 199368 167696 199374
rect 167644 199310 167696 199316
rect 167552 199300 167604 199306
rect 167552 199242 167604 199248
rect 167460 192772 167512 192778
rect 167460 192714 167512 192720
rect 167564 185609 167592 199242
rect 167656 198257 167684 199310
rect 167642 198248 167698 198257
rect 167642 198183 167698 198192
rect 167644 198144 167696 198150
rect 167644 198086 167696 198092
rect 167550 185600 167606 185609
rect 167656 185570 167684 198086
rect 167734 197840 167790 197849
rect 167734 197775 167790 197784
rect 167748 185745 167776 197775
rect 167840 193934 167868 199532
rect 167920 199436 167972 199442
rect 167920 199378 167972 199384
rect 167932 198218 167960 199378
rect 167920 198212 167972 198218
rect 168116 198200 168144 199679
rect 168288 199650 168340 199656
rect 168196 199640 168248 199646
rect 168196 199582 168248 199588
rect 167920 198154 167972 198160
rect 168024 198172 168144 198200
rect 167918 198112 167974 198121
rect 167918 198047 167974 198056
rect 167828 193928 167880 193934
rect 167828 193870 167880 193876
rect 167734 185736 167790 185745
rect 167734 185671 167790 185680
rect 167550 185535 167606 185544
rect 167644 185564 167696 185570
rect 167644 185506 167696 185512
rect 167368 155576 167420 155582
rect 167368 155518 167420 155524
rect 167184 155236 167236 155242
rect 167184 155178 167236 155184
rect 167092 148708 167144 148714
rect 167092 148650 167144 148656
rect 166816 148640 166868 148646
rect 166816 148582 166868 148588
rect 167932 148510 167960 198047
rect 168024 185609 168052 198172
rect 168102 198112 168158 198121
rect 168102 198047 168158 198056
rect 168116 190738 168144 198047
rect 168104 190732 168156 190738
rect 168104 190674 168156 190680
rect 168010 185600 168066 185609
rect 168010 185535 168066 185544
rect 168208 177002 168236 199582
rect 168300 192234 168328 199650
rect 168288 192228 168340 192234
rect 168288 192170 168340 192176
rect 168392 185638 168420 199736
rect 168802 199736 168834 199744
rect 169036 199736 169294 199764
rect 168746 199679 168802 199688
rect 168932 199708 168984 199714
rect 168932 199650 168984 199656
rect 168748 199640 168800 199646
rect 168748 199582 168800 199588
rect 168472 199572 168524 199578
rect 168472 199514 168524 199520
rect 168380 185632 168432 185638
rect 168380 185574 168432 185580
rect 168196 176996 168248 177002
rect 168196 176938 168248 176944
rect 168484 155310 168512 199514
rect 168760 192846 168788 199582
rect 168748 192840 168800 192846
rect 168748 192782 168800 192788
rect 168944 185688 168972 199650
rect 168576 185660 168972 185688
rect 168576 155378 168604 185660
rect 169036 172514 169064 199736
rect 169634 199730 169662 200124
rect 169726 199923 169754 200124
rect 169712 199914 169768 199923
rect 169712 199849 169768 199858
rect 169818 199850 169846 200124
rect 169806 199844 169858 199850
rect 169806 199786 169858 199792
rect 169588 199702 169662 199730
rect 169758 199744 169814 199753
rect 169208 199640 169260 199646
rect 169208 199582 169260 199588
rect 169300 199640 169352 199646
rect 169300 199582 169352 199588
rect 169116 199572 169168 199578
rect 169116 199514 169168 199520
rect 169128 180033 169156 199514
rect 169220 192710 169248 199582
rect 169208 192704 169260 192710
rect 169208 192646 169260 192652
rect 169206 185872 169262 185881
rect 169206 185807 169262 185816
rect 169114 180024 169170 180033
rect 169114 179959 169170 179968
rect 168668 172486 169064 172514
rect 168668 155446 168696 172486
rect 168656 155440 168708 155446
rect 168656 155382 168708 155388
rect 168564 155372 168616 155378
rect 168564 155314 168616 155320
rect 168472 155304 168524 155310
rect 168472 155246 168524 155252
rect 167920 148504 167972 148510
rect 165710 148472 165766 148481
rect 167920 148446 167972 148452
rect 169220 148442 169248 185807
rect 169312 185745 169340 199582
rect 169392 199572 169444 199578
rect 169392 199514 169444 199520
rect 169404 193905 169432 199514
rect 169390 193896 169446 193905
rect 169390 193831 169446 193840
rect 169298 185736 169354 185745
rect 169298 185671 169354 185680
rect 169588 185609 169616 199702
rect 169910 199696 169938 200124
rect 170002 199918 170030 200124
rect 170094 199918 170122 200124
rect 170186 199918 170214 200124
rect 170278 199918 170306 200124
rect 169990 199912 170042 199918
rect 169990 199854 170042 199860
rect 170082 199912 170134 199918
rect 170082 199854 170134 199860
rect 170174 199912 170226 199918
rect 170174 199854 170226 199860
rect 170266 199912 170318 199918
rect 170266 199854 170318 199860
rect 170370 199764 170398 200124
rect 170462 199918 170490 200124
rect 170554 199923 170582 200124
rect 170450 199912 170502 199918
rect 170450 199854 170502 199860
rect 170540 199914 170596 199923
rect 170540 199849 170596 199858
rect 169758 199679 169814 199688
rect 169668 199640 169720 199646
rect 169668 199582 169720 199588
rect 169680 198218 169708 199582
rect 169772 199442 169800 199679
rect 169864 199668 169938 199696
rect 170034 199744 170090 199753
rect 170034 199679 170036 199688
rect 169760 199436 169812 199442
rect 169760 199378 169812 199384
rect 169668 198212 169720 198218
rect 169668 198154 169720 198160
rect 169864 186561 169892 199668
rect 170088 199679 170090 199688
rect 170324 199736 170398 199764
rect 170646 199764 170674 200124
rect 170738 199918 170766 200124
rect 170830 199918 170858 200124
rect 170922 199918 170950 200124
rect 171014 199923 171042 200124
rect 170726 199912 170778 199918
rect 170726 199854 170778 199860
rect 170818 199912 170870 199918
rect 170818 199854 170870 199860
rect 170910 199912 170962 199918
rect 170910 199854 170962 199860
rect 171000 199914 171056 199923
rect 171106 199918 171134 200124
rect 171198 199923 171226 200124
rect 171000 199849 171056 199858
rect 171094 199912 171146 199918
rect 171094 199854 171146 199860
rect 171184 199914 171240 199923
rect 171290 199918 171318 200124
rect 171382 199918 171410 200124
rect 171474 199918 171502 200124
rect 171184 199849 171240 199858
rect 171278 199912 171330 199918
rect 171278 199854 171330 199860
rect 171370 199912 171422 199918
rect 171370 199854 171422 199860
rect 171462 199912 171514 199918
rect 171566 199889 171594 200124
rect 171658 199918 171686 200124
rect 171750 199918 171778 200124
rect 171842 199918 171870 200124
rect 171934 199918 171962 200124
rect 172026 199918 172054 200124
rect 171646 199912 171698 199918
rect 171462 199854 171514 199860
rect 171552 199880 171608 199889
rect 171646 199854 171698 199860
rect 171738 199912 171790 199918
rect 171738 199854 171790 199860
rect 171830 199912 171882 199918
rect 171830 199854 171882 199860
rect 171922 199912 171974 199918
rect 171922 199854 171974 199860
rect 172014 199912 172066 199918
rect 172014 199854 172066 199860
rect 171552 199815 171608 199824
rect 170772 199776 170824 199782
rect 170646 199753 170720 199764
rect 170494 199744 170550 199753
rect 170036 199650 170088 199656
rect 170128 199640 170180 199646
rect 170128 199582 170180 199588
rect 170220 199640 170272 199646
rect 170220 199582 170272 199588
rect 169944 199572 169996 199578
rect 169944 199514 169996 199520
rect 169956 199034 169984 199514
rect 170036 199504 170088 199510
rect 170036 199446 170088 199452
rect 169944 199028 169996 199034
rect 169944 198970 169996 198976
rect 169942 196480 169998 196489
rect 169942 196415 169998 196424
rect 169956 196110 169984 196415
rect 169944 196104 169996 196110
rect 169944 196046 169996 196052
rect 169942 195936 169998 195945
rect 169942 195871 169998 195880
rect 169956 194002 169984 195871
rect 169944 193996 169996 194002
rect 169944 193938 169996 193944
rect 169850 186552 169906 186561
rect 169850 186487 169906 186496
rect 169852 186312 169904 186318
rect 169852 186254 169904 186260
rect 169760 185632 169812 185638
rect 169574 185600 169630 185609
rect 169760 185574 169812 185580
rect 169574 185535 169630 185544
rect 165710 148407 165766 148416
rect 169208 148436 169260 148442
rect 169208 148378 169260 148384
rect 164240 148368 164292 148374
rect 164240 148310 164292 148316
rect 164148 147076 164200 147082
rect 164148 147018 164200 147024
rect 164238 146024 164294 146033
rect 164238 145959 164294 145968
rect 164146 144528 164202 144537
rect 164146 144463 164202 144472
rect 164160 140162 164188 144463
rect 164114 140134 164188 140162
rect 164114 139876 164142 140134
rect 164252 139890 164280 145959
rect 167734 144664 167790 144673
rect 167734 144599 167790 144608
rect 166630 144392 166686 144401
rect 166630 144327 166686 144336
rect 165528 142996 165580 143002
rect 165528 142938 165580 142944
rect 165540 139890 165568 142938
rect 166078 141536 166134 141545
rect 166078 141471 166134 141480
rect 166092 139890 166120 141471
rect 166644 139890 166672 144327
rect 166908 143064 166960 143070
rect 166908 143006 166960 143012
rect 166920 140162 166948 143006
rect 164252 139862 164680 139890
rect 165232 139862 165568 139890
rect 165784 139862 166120 139890
rect 166336 139862 166672 139890
rect 166874 140134 166948 140162
rect 166874 139876 166902 140134
rect 167748 139890 167776 144599
rect 168840 143132 168892 143138
rect 168840 143074 168892 143080
rect 168852 139890 168880 143074
rect 169392 141500 169444 141506
rect 169392 141442 169444 141448
rect 169404 139890 169432 141442
rect 169772 140758 169800 185574
rect 169864 147529 169892 186254
rect 170048 185586 170076 199446
rect 169956 185558 170076 185586
rect 169850 147520 169906 147529
rect 169850 147455 169906 147464
rect 169956 147354 169984 185558
rect 170140 171134 170168 199582
rect 170232 198257 170260 199582
rect 170218 198248 170274 198257
rect 170218 198183 170274 198192
rect 170324 185638 170352 199736
rect 170646 199744 170734 199753
rect 170646 199736 170678 199744
rect 170494 199679 170550 199688
rect 171048 199776 171100 199782
rect 170772 199718 170824 199724
rect 170862 199744 170918 199753
rect 170678 199679 170734 199688
rect 170508 198801 170536 199679
rect 170588 199640 170640 199646
rect 170588 199582 170640 199588
rect 170494 198792 170550 198801
rect 170494 198727 170550 198736
rect 170600 186289 170628 199582
rect 170680 199572 170732 199578
rect 170680 199514 170732 199520
rect 170586 186280 170642 186289
rect 170586 186215 170642 186224
rect 170312 185632 170364 185638
rect 170312 185574 170364 185580
rect 170692 184929 170720 199514
rect 170784 198121 170812 199718
rect 171600 199776 171652 199782
rect 171048 199718 171100 199724
rect 171138 199744 171194 199753
rect 170862 199679 170918 199688
rect 170770 198112 170826 198121
rect 170770 198047 170826 198056
rect 170876 186318 170904 199679
rect 171060 198150 171088 199718
rect 171506 199744 171562 199753
rect 171138 199679 171194 199688
rect 171324 199708 171376 199714
rect 171048 198144 171100 198150
rect 171048 198086 171100 198092
rect 171152 186640 171180 199679
rect 171324 199650 171376 199656
rect 171416 199708 171468 199714
rect 172118 199730 172146 200124
rect 172210 199918 172238 200124
rect 172198 199912 172250 199918
rect 172198 199854 172250 199860
rect 172302 199764 172330 200124
rect 172394 199918 172422 200124
rect 172382 199912 172434 199918
rect 172382 199854 172434 199860
rect 172486 199764 172514 200124
rect 172578 199918 172606 200124
rect 172670 199918 172698 200124
rect 172762 199918 172790 200124
rect 172566 199912 172618 199918
rect 172566 199854 172618 199860
rect 172658 199912 172710 199918
rect 172658 199854 172710 199860
rect 172750 199912 172802 199918
rect 172750 199854 172802 199860
rect 172302 199736 172376 199764
rect 171600 199718 171652 199724
rect 171506 199679 171562 199688
rect 171416 199650 171468 199656
rect 171232 199640 171284 199646
rect 171232 199582 171284 199588
rect 171244 186658 171272 199582
rect 171336 186726 171364 199650
rect 171324 186720 171376 186726
rect 171324 186662 171376 186668
rect 171060 186612 171180 186640
rect 171232 186652 171284 186658
rect 171060 186318 171088 186612
rect 171232 186594 171284 186600
rect 171428 186504 171456 199650
rect 171520 199442 171548 199679
rect 171508 199436 171560 199442
rect 171508 199378 171560 199384
rect 171612 186658 171640 199718
rect 171876 199708 171928 199714
rect 171876 199650 171928 199656
rect 171968 199708 172020 199714
rect 171968 199650 172020 199656
rect 172072 199702 172146 199730
rect 171692 199640 171744 199646
rect 171692 199582 171744 199588
rect 171600 186652 171652 186658
rect 171600 186594 171652 186600
rect 171152 186476 171456 186504
rect 170864 186312 170916 186318
rect 170864 186254 170916 186260
rect 171048 186312 171100 186318
rect 171048 186254 171100 186260
rect 170678 184920 170734 184929
rect 170678 184855 170734 184864
rect 170048 171106 170168 171134
rect 169944 147348 169996 147354
rect 169944 147290 169996 147296
rect 170048 146946 170076 171106
rect 171152 147393 171180 186476
rect 171704 186402 171732 199582
rect 171784 199572 171836 199578
rect 171784 199514 171836 199520
rect 171428 186374 171732 186402
rect 171232 178288 171284 178294
rect 171232 178230 171284 178236
rect 171244 147490 171272 178230
rect 171324 175228 171376 175234
rect 171324 175170 171376 175176
rect 171232 147484 171284 147490
rect 171232 147426 171284 147432
rect 171336 147422 171364 175170
rect 171324 147416 171376 147422
rect 171138 147384 171194 147393
rect 171324 147358 171376 147364
rect 171138 147319 171194 147328
rect 171428 147286 171456 186374
rect 171508 186312 171560 186318
rect 171508 186254 171560 186260
rect 171520 147558 171548 186254
rect 171796 175234 171824 199514
rect 171888 185609 171916 199650
rect 171980 193118 172008 199650
rect 171968 193112 172020 193118
rect 171968 193054 172020 193060
rect 172072 185609 172100 199702
rect 172152 199640 172204 199646
rect 172152 199582 172204 199588
rect 172244 199640 172296 199646
rect 172244 199582 172296 199588
rect 171874 185600 171930 185609
rect 171874 185535 171930 185544
rect 172058 185600 172114 185609
rect 172058 185535 172114 185544
rect 172164 185201 172192 199582
rect 172256 185745 172284 199582
rect 172242 185736 172298 185745
rect 172242 185671 172298 185680
rect 172150 185192 172206 185201
rect 172150 185127 172206 185136
rect 172348 178294 172376 199736
rect 172440 199736 172514 199764
rect 172854 199764 172882 200124
rect 172946 199918 172974 200124
rect 173038 199918 173066 200124
rect 173130 199918 173158 200124
rect 172934 199912 172986 199918
rect 172934 199854 172986 199860
rect 173026 199912 173078 199918
rect 173026 199854 173078 199860
rect 173118 199912 173170 199918
rect 173222 199889 173250 200124
rect 173314 199918 173342 200124
rect 173302 199912 173354 199918
rect 173118 199854 173170 199860
rect 173208 199880 173264 199889
rect 173406 199889 173434 200124
rect 173302 199854 173354 199860
rect 173392 199880 173448 199889
rect 173208 199815 173264 199824
rect 173392 199815 173448 199824
rect 173072 199776 173124 199782
rect 172854 199736 172928 199764
rect 172440 184074 172468 199736
rect 172612 199708 172664 199714
rect 172612 199650 172664 199656
rect 172704 199708 172756 199714
rect 172756 199668 172836 199696
rect 172704 199650 172756 199656
rect 172624 199594 172652 199650
rect 172624 199566 172744 199594
rect 172612 185632 172664 185638
rect 172612 185574 172664 185580
rect 172428 184068 172480 184074
rect 172428 184010 172480 184016
rect 172520 182028 172572 182034
rect 172520 181970 172572 181976
rect 172336 178288 172388 178294
rect 172336 178230 172388 178236
rect 171784 175228 171836 175234
rect 171784 175170 171836 175176
rect 171508 147552 171560 147558
rect 171508 147494 171560 147500
rect 171416 147280 171468 147286
rect 171416 147222 171468 147228
rect 170036 146940 170088 146946
rect 170036 146882 170088 146888
rect 171048 144764 171100 144770
rect 171048 144706 171100 144712
rect 170496 141636 170548 141642
rect 170496 141578 170548 141584
rect 169760 140752 169812 140758
rect 169760 140694 169812 140700
rect 170508 139890 170536 141578
rect 171060 139890 171088 144706
rect 172428 144696 172480 144702
rect 172428 144638 172480 144644
rect 172152 141704 172204 141710
rect 172152 141646 172204 141652
rect 172164 139890 172192 141646
rect 172440 140162 172468 144638
rect 172532 140622 172560 181970
rect 172624 147014 172652 185574
rect 172716 147150 172744 199566
rect 172808 186386 172836 199668
rect 172900 199646 172928 199736
rect 173072 199718 173124 199724
rect 173164 199776 173216 199782
rect 173498 199764 173526 200124
rect 173590 199918 173618 200124
rect 173682 199918 173710 200124
rect 173578 199912 173630 199918
rect 173578 199854 173630 199860
rect 173670 199912 173722 199918
rect 173670 199854 173722 199860
rect 173268 199753 173526 199764
rect 173164 199718 173216 199724
rect 173254 199744 173526 199753
rect 172888 199640 172940 199646
rect 172888 199582 172940 199588
rect 172980 199572 173032 199578
rect 172980 199514 173032 199520
rect 172888 199504 172940 199510
rect 172888 199446 172940 199452
rect 172900 186522 172928 199446
rect 172888 186516 172940 186522
rect 172888 186458 172940 186464
rect 172796 186380 172848 186386
rect 172796 186322 172848 186328
rect 172992 186266 173020 199514
rect 172808 186238 173020 186266
rect 172808 147218 172836 186238
rect 172886 186144 172942 186153
rect 172886 186079 172942 186088
rect 172900 149870 172928 186079
rect 173084 185337 173112 199718
rect 173176 199594 173204 199718
rect 173310 199736 173526 199744
rect 173624 199776 173676 199782
rect 173774 199730 173802 200124
rect 173866 199918 173894 200124
rect 173958 199918 173986 200124
rect 173854 199912 173906 199918
rect 173854 199854 173906 199860
rect 173946 199912 173998 199918
rect 173946 199854 173998 199860
rect 174050 199764 174078 200124
rect 173624 199718 173676 199724
rect 173254 199679 173310 199688
rect 173348 199640 173400 199646
rect 173176 199566 173296 199594
rect 173348 199582 173400 199588
rect 173164 199436 173216 199442
rect 173164 199378 173216 199384
rect 173176 185609 173204 199378
rect 173268 185638 173296 199566
rect 173256 185632 173308 185638
rect 173162 185600 173218 185609
rect 173360 185609 173388 199582
rect 173438 198792 173494 198801
rect 173438 198727 173494 198736
rect 173452 198082 173480 198727
rect 173440 198076 173492 198082
rect 173440 198018 173492 198024
rect 173440 197600 173492 197606
rect 173440 197542 173492 197548
rect 173452 195022 173480 197542
rect 173440 195016 173492 195022
rect 173440 194958 173492 194964
rect 173256 185574 173308 185580
rect 173346 185600 173402 185609
rect 173162 185535 173218 185544
rect 173346 185535 173402 185544
rect 173070 185328 173126 185337
rect 173070 185263 173126 185272
rect 173636 182034 173664 199718
rect 173728 199702 173802 199730
rect 174004 199736 174078 199764
rect 173900 199708 173952 199714
rect 173728 186017 173756 199702
rect 173900 199650 173952 199656
rect 173808 199232 173860 199238
rect 173808 199174 173860 199180
rect 173820 198966 173848 199174
rect 173808 198960 173860 198966
rect 173808 198902 173860 198908
rect 173714 186008 173770 186017
rect 173714 185943 173770 185952
rect 173624 182028 173676 182034
rect 173624 181970 173676 181976
rect 172888 149864 172940 149870
rect 172888 149806 172940 149812
rect 173072 149660 173124 149666
rect 173072 149602 173124 149608
rect 172796 147212 172848 147218
rect 172796 147154 172848 147160
rect 172704 147144 172756 147150
rect 172704 147086 172756 147092
rect 172612 147008 172664 147014
rect 172612 146950 172664 146956
rect 172520 140616 172572 140622
rect 172520 140558 172572 140564
rect 167440 139862 167776 139890
rect 167992 139874 168328 139890
rect 167992 139868 168340 139874
rect 167992 139862 168288 139868
rect 168544 139862 168880 139890
rect 169096 139862 169432 139890
rect 170200 139862 170536 139890
rect 170752 139862 171088 139890
rect 171856 139862 172192 139890
rect 172394 140134 172468 140162
rect 172394 139876 172422 140134
rect 173084 139890 173112 149602
rect 173912 146169 173940 199650
rect 174004 192982 174032 199736
rect 174142 199696 174170 200124
rect 174234 199764 174262 200124
rect 174326 199923 174354 200124
rect 174312 199914 174368 199923
rect 174418 199918 174446 200124
rect 174312 199849 174368 199858
rect 174406 199912 174458 199918
rect 174406 199854 174458 199860
rect 174510 199764 174538 200124
rect 174602 199918 174630 200124
rect 174590 199912 174642 199918
rect 174590 199854 174642 199860
rect 174694 199764 174722 200124
rect 174786 199918 174814 200124
rect 174774 199912 174826 199918
rect 174878 199889 174906 200124
rect 174774 199854 174826 199860
rect 174864 199880 174920 199889
rect 174864 199815 174920 199824
rect 174970 199764 174998 200124
rect 174234 199736 174400 199764
rect 174510 199736 174584 199764
rect 174694 199736 174768 199764
rect 174142 199668 174216 199696
rect 174084 199368 174136 199374
rect 174084 199310 174136 199316
rect 174096 199034 174124 199310
rect 174084 199028 174136 199034
rect 174084 198970 174136 198976
rect 174188 194206 174216 199668
rect 174268 199640 174320 199646
rect 174268 199582 174320 199588
rect 174176 194200 174228 194206
rect 174176 194142 174228 194148
rect 173992 192976 174044 192982
rect 173992 192918 174044 192924
rect 174084 192500 174136 192506
rect 174084 192442 174136 192448
rect 173992 192432 174044 192438
rect 173992 192374 174044 192380
rect 174004 147257 174032 192374
rect 174096 150278 174124 192442
rect 174280 186454 174308 199582
rect 174372 194070 174400 199736
rect 174556 199560 174584 199736
rect 174464 199532 174584 199560
rect 174360 194064 174412 194070
rect 174360 194006 174412 194012
rect 174268 186448 174320 186454
rect 174268 186390 174320 186396
rect 174464 186266 174492 199532
rect 174636 199504 174688 199510
rect 174636 199446 174688 199452
rect 174544 199436 174596 199442
rect 174544 199378 174596 199384
rect 174556 186289 174584 199378
rect 174188 186238 174492 186266
rect 174542 186280 174598 186289
rect 174084 150272 174136 150278
rect 174084 150214 174136 150220
rect 174188 150113 174216 186238
rect 174542 186215 174598 186224
rect 174648 185706 174676 199446
rect 174740 199034 174768 199736
rect 174832 199736 174998 199764
rect 174728 199028 174780 199034
rect 174728 198970 174780 198976
rect 174832 198801 174860 199736
rect 174912 199640 174964 199646
rect 175062 199594 175090 200124
rect 175154 199918 175182 200124
rect 175246 199918 175274 200124
rect 175142 199912 175194 199918
rect 175142 199854 175194 199860
rect 175234 199912 175286 199918
rect 175234 199854 175286 199860
rect 175188 199776 175240 199782
rect 175186 199744 175188 199753
rect 175338 199764 175366 200124
rect 175430 199923 175458 200124
rect 175416 199914 175472 199923
rect 175416 199849 175472 199858
rect 175522 199764 175550 200124
rect 175240 199744 175242 199753
rect 175186 199679 175242 199688
rect 175292 199736 175366 199764
rect 175476 199753 175550 199764
rect 175462 199744 175550 199753
rect 175292 199646 175320 199736
rect 175518 199736 175550 199744
rect 175614 199696 175642 200124
rect 175706 199850 175734 200124
rect 175798 199918 175826 200124
rect 175786 199912 175838 199918
rect 175786 199854 175838 199860
rect 175694 199844 175746 199850
rect 175694 199786 175746 199792
rect 175890 199730 175918 200124
rect 175982 199889 176010 200124
rect 176074 199918 176102 200124
rect 176166 199918 176194 200124
rect 176258 199918 176286 200124
rect 176062 199912 176114 199918
rect 175968 199880 176024 199889
rect 176062 199854 176114 199860
rect 176154 199912 176206 199918
rect 176154 199854 176206 199860
rect 176246 199912 176298 199918
rect 176350 199889 176378 200124
rect 176442 199918 176470 200124
rect 176534 199923 176562 200124
rect 176430 199912 176482 199918
rect 176246 199854 176298 199860
rect 176336 199880 176392 199889
rect 175968 199815 176024 199824
rect 176430 199854 176482 199860
rect 176520 199914 176576 199923
rect 176520 199849 176576 199858
rect 176336 199815 176392 199824
rect 175462 199679 175518 199688
rect 175568 199668 175642 199696
rect 175740 199708 175792 199714
rect 174912 199582 174964 199588
rect 174818 198792 174874 198801
rect 174818 198727 174874 198736
rect 174820 198620 174872 198626
rect 174820 198562 174872 198568
rect 174832 194886 174860 198562
rect 174820 194880 174872 194886
rect 174820 194822 174872 194828
rect 174728 194064 174780 194070
rect 174728 194006 174780 194012
rect 174636 185700 174688 185706
rect 174636 185642 174688 185648
rect 174740 172514 174768 194006
rect 174924 192506 174952 199582
rect 175016 199566 175090 199594
rect 175280 199640 175332 199646
rect 175280 199582 175332 199588
rect 174912 192500 174964 192506
rect 174912 192442 174964 192448
rect 175016 192438 175044 199566
rect 175568 199560 175596 199668
rect 175740 199650 175792 199656
rect 175844 199702 175918 199730
rect 176292 199776 176344 199782
rect 176626 199764 176654 200124
rect 176718 199918 176746 200124
rect 176810 199918 176838 200124
rect 176902 199923 176930 200124
rect 176706 199912 176758 199918
rect 176706 199854 176758 199860
rect 176798 199912 176850 199918
rect 176798 199854 176850 199860
rect 176888 199914 176944 199923
rect 176994 199918 177022 200124
rect 176888 199849 176944 199858
rect 176982 199912 177034 199918
rect 176982 199854 177034 199860
rect 176844 199776 176896 199782
rect 176626 199736 176700 199764
rect 176292 199718 176344 199724
rect 176016 199708 176068 199714
rect 175384 199532 175596 199560
rect 175648 199572 175700 199578
rect 175004 192432 175056 192438
rect 175004 192374 175056 192380
rect 175280 185632 175332 185638
rect 175280 185574 175332 185580
rect 174372 172486 174768 172514
rect 174174 150104 174230 150113
rect 174174 150039 174230 150048
rect 174372 149977 174400 172486
rect 174358 149968 174414 149977
rect 174358 149903 174414 149912
rect 175292 149802 175320 185574
rect 175384 149938 175412 199532
rect 175648 199514 175700 199520
rect 175556 199436 175608 199442
rect 175556 199378 175608 199384
rect 175464 183116 175516 183122
rect 175464 183058 175516 183064
rect 175476 150006 175504 183058
rect 175568 150074 175596 199378
rect 175660 185881 175688 199514
rect 175646 185872 175702 185881
rect 175646 185807 175702 185816
rect 175752 185745 175780 199650
rect 175738 185736 175794 185745
rect 175738 185671 175794 185680
rect 175844 185638 175872 199702
rect 176016 199650 176068 199656
rect 176200 199708 176252 199714
rect 176200 199650 176252 199656
rect 175832 185632 175884 185638
rect 175832 185574 175884 185580
rect 176028 185473 176056 199650
rect 176014 185464 176070 185473
rect 176014 185399 176070 185408
rect 176212 183122 176240 199650
rect 176304 186289 176332 199718
rect 176384 199708 176436 199714
rect 176384 199650 176436 199656
rect 176290 186280 176346 186289
rect 176290 186215 176346 186224
rect 176200 183116 176252 183122
rect 176200 183058 176252 183064
rect 176396 178090 176424 199650
rect 176672 186561 176700 199736
rect 177086 199764 177114 200124
rect 177178 199918 177206 200124
rect 177166 199912 177218 199918
rect 177166 199854 177218 199860
rect 177270 199764 177298 200124
rect 177362 199918 177390 200124
rect 177350 199912 177402 199918
rect 177350 199854 177402 199860
rect 177454 199764 177482 200124
rect 177086 199736 177160 199764
rect 176844 199718 176896 199724
rect 176750 197976 176806 197985
rect 176750 197911 176806 197920
rect 176764 197577 176792 197911
rect 176750 197568 176806 197577
rect 176750 197503 176806 197512
rect 176856 192914 176884 199718
rect 176936 199708 176988 199714
rect 176936 199650 176988 199656
rect 176844 192908 176896 192914
rect 176844 192850 176896 192856
rect 176658 186552 176714 186561
rect 176658 186487 176714 186496
rect 176844 186312 176896 186318
rect 176844 186254 176896 186260
rect 176752 186244 176804 186250
rect 176752 186186 176804 186192
rect 176660 186176 176712 186182
rect 176660 186118 176712 186124
rect 175648 178084 175700 178090
rect 175648 178026 175700 178032
rect 176384 178084 176436 178090
rect 176384 178026 176436 178032
rect 175660 150210 175688 178026
rect 175648 150204 175700 150210
rect 175648 150146 175700 150152
rect 175556 150068 175608 150074
rect 175556 150010 175608 150016
rect 175464 150000 175516 150006
rect 175464 149942 175516 149948
rect 175372 149932 175424 149938
rect 175372 149874 175424 149880
rect 175280 149796 175332 149802
rect 175280 149738 175332 149744
rect 173990 147248 174046 147257
rect 173990 147183 174046 147192
rect 173898 146160 173954 146169
rect 173898 146095 173954 146104
rect 174360 144832 174412 144838
rect 174360 144774 174412 144780
rect 174372 139890 174400 144774
rect 176568 143404 176620 143410
rect 176568 143346 176620 143352
rect 176016 143336 176068 143342
rect 176016 143278 176068 143284
rect 175188 143200 175240 143206
rect 175188 143142 175240 143148
rect 174728 141568 174780 141574
rect 174728 141510 174780 141516
rect 174740 139890 174768 141510
rect 174818 140312 174874 140321
rect 174818 140247 174874 140256
rect 173084 139862 173512 139890
rect 174064 139862 174400 139890
rect 174616 139862 174768 139890
rect 168288 139810 168340 139816
rect 173256 139800 173308 139806
rect 169648 139738 169800 139754
rect 172960 139748 173256 139754
rect 172960 139742 173308 139748
rect 169648 139732 169812 139738
rect 169648 139726 169760 139732
rect 172960 139726 173296 139742
rect 169760 139674 169812 139680
rect 171600 139664 171652 139670
rect 171304 139612 171600 139618
rect 171304 139606 171652 139612
rect 171304 139590 171640 139606
rect 174832 139505 174860 140247
rect 175200 140162 175228 143142
rect 175154 140134 175228 140162
rect 175154 139876 175182 140134
rect 176028 139890 176056 143278
rect 176580 139890 176608 143346
rect 176672 141273 176700 186118
rect 176764 141681 176792 186186
rect 176856 150346 176884 186254
rect 176844 150340 176896 150346
rect 176844 150282 176896 150288
rect 176948 150142 176976 199650
rect 177132 194070 177160 199736
rect 177224 199736 177298 199764
rect 177408 199736 177482 199764
rect 177120 194064 177172 194070
rect 177120 194006 177172 194012
rect 177224 186318 177252 199736
rect 177408 199730 177436 199736
rect 177362 199702 177436 199730
rect 177362 199696 177390 199702
rect 177546 199696 177574 200124
rect 177638 199918 177666 200124
rect 177626 199912 177678 199918
rect 177626 199854 177678 199860
rect 177764 199912 177816 199918
rect 177764 199854 177816 199860
rect 177316 199668 177390 199696
rect 177500 199668 177574 199696
rect 177212 186312 177264 186318
rect 177212 186254 177264 186260
rect 177316 176633 177344 199668
rect 177500 186250 177528 199668
rect 177488 186244 177540 186250
rect 177488 186186 177540 186192
rect 177776 186182 177804 199854
rect 177856 199844 177908 199850
rect 177856 199786 177908 199792
rect 177868 186289 177896 199786
rect 179052 199640 179104 199646
rect 179052 199582 179104 199588
rect 178960 199436 179012 199442
rect 178960 199378 179012 199384
rect 178868 190732 178920 190738
rect 178868 190674 178920 190680
rect 178776 189100 178828 189106
rect 178776 189042 178828 189048
rect 178684 186992 178736 186998
rect 178684 186934 178736 186940
rect 177854 186280 177910 186289
rect 177854 186215 177910 186224
rect 177764 186176 177816 186182
rect 177764 186118 177816 186124
rect 177302 176624 177358 176633
rect 177302 176559 177358 176568
rect 176936 150136 176988 150142
rect 176936 150078 176988 150084
rect 178592 146872 178644 146878
rect 178592 146814 178644 146820
rect 178040 146124 178092 146130
rect 178040 146066 178092 146072
rect 177672 143472 177724 143478
rect 177672 143414 177724 143420
rect 177120 142792 177172 142798
rect 177120 142734 177172 142740
rect 176750 141672 176806 141681
rect 176750 141607 176806 141616
rect 176658 141264 176714 141273
rect 176658 141199 176714 141208
rect 177132 139890 177160 142734
rect 177684 139890 177712 143414
rect 177948 142656 178000 142662
rect 177948 142598 178000 142604
rect 177960 140162 177988 142598
rect 178052 140690 178080 146066
rect 178132 145512 178184 145518
rect 178132 145454 178184 145460
rect 178040 140684 178092 140690
rect 178040 140626 178092 140632
rect 175720 139862 176056 139890
rect 176272 139862 176608 139890
rect 176824 139862 177160 139890
rect 177376 139862 177712 139890
rect 177914 140134 177988 140162
rect 177914 139876 177942 140134
rect 178144 139890 178172 145454
rect 178604 143410 178632 146814
rect 178592 143404 178644 143410
rect 178592 143346 178644 143352
rect 178696 142154 178724 186934
rect 178788 146962 178816 189042
rect 178880 147098 178908 190674
rect 178972 147234 179000 199378
rect 179064 150414 179092 199582
rect 183192 199368 183244 199374
rect 183192 199310 183244 199316
rect 180248 199164 180300 199170
rect 180248 199106 180300 199112
rect 180800 199164 180852 199170
rect 180800 199106 180852 199112
rect 180156 195832 180208 195838
rect 180156 195774 180208 195780
rect 180064 195696 180116 195702
rect 180064 195638 180116 195644
rect 179052 150408 179104 150414
rect 179052 150350 179104 150356
rect 179328 147620 179380 147626
rect 179328 147562 179380 147568
rect 178972 147206 179092 147234
rect 178880 147070 179000 147098
rect 178788 146934 178908 146962
rect 178696 142126 178816 142154
rect 178590 140720 178646 140729
rect 178590 140655 178646 140664
rect 178684 140684 178736 140690
rect 178144 139862 178480 139890
rect 178604 139874 178632 140655
rect 178684 140626 178736 140632
rect 178696 139890 178724 140626
rect 178788 140418 178816 142126
rect 178776 140412 178828 140418
rect 178776 140354 178828 140360
rect 178880 140282 178908 146934
rect 178972 142154 179000 147070
rect 179064 146266 179092 147206
rect 179052 146260 179104 146266
rect 179052 146202 179104 146208
rect 179064 142730 179092 146202
rect 179052 142724 179104 142730
rect 179052 142666 179104 142672
rect 179340 142662 179368 147562
rect 179788 146260 179840 146266
rect 179788 146202 179840 146208
rect 179604 146056 179656 146062
rect 179604 145998 179656 146004
rect 179512 145444 179564 145450
rect 179512 145386 179564 145392
rect 179420 145376 179472 145382
rect 179420 145318 179472 145324
rect 179432 143478 179460 145318
rect 179420 143472 179472 143478
rect 179420 143414 179472 143420
rect 179524 142798 179552 145386
rect 179512 142792 179564 142798
rect 179512 142734 179564 142740
rect 179328 142656 179380 142662
rect 179328 142598 179380 142604
rect 178972 142126 179276 142154
rect 178868 140276 178920 140282
rect 178868 140218 178920 140224
rect 179248 140146 179276 142126
rect 179616 140162 179644 145998
rect 179800 143342 179828 146202
rect 180076 144906 180104 195638
rect 180168 148238 180196 195774
rect 180156 148232 180208 148238
rect 180156 148174 180208 148180
rect 180064 144900 180116 144906
rect 180064 144842 180116 144848
rect 180260 144786 180288 199106
rect 180430 198928 180486 198937
rect 180430 198863 180486 198872
rect 180340 192840 180392 192846
rect 180340 192782 180392 192788
rect 180352 147665 180380 192782
rect 180444 151814 180472 198863
rect 180444 151786 180564 151814
rect 180338 147656 180394 147665
rect 180338 147591 180394 147600
rect 179892 144758 180288 144786
rect 179788 143336 179840 143342
rect 179788 143278 179840 143284
rect 179892 143154 179920 144758
rect 179236 140140 179288 140146
rect 179236 140082 179288 140088
rect 179570 140134 179644 140162
rect 179708 143126 179920 143154
rect 178592 139868 178644 139874
rect 178696 139862 179032 139890
rect 179570 139876 179598 140134
rect 178592 139810 178644 139816
rect 174818 139496 174874 139505
rect 174818 139431 174874 139440
rect 179708 139369 179736 143126
rect 179788 142724 179840 142730
rect 179788 142666 179840 142672
rect 179800 139890 179828 142666
rect 180156 141840 180208 141846
rect 180156 141782 180208 141788
rect 180168 141166 180196 141782
rect 180156 141160 180208 141166
rect 180156 141102 180208 141108
rect 179800 139862 180136 139890
rect 180430 139768 180486 139777
rect 180430 139703 180486 139712
rect 179878 139632 179934 139641
rect 179878 139567 179880 139576
rect 179932 139567 179934 139576
rect 179880 139538 179932 139544
rect 180444 139534 180472 139703
rect 180432 139528 180484 139534
rect 180432 139470 180484 139476
rect 180536 139369 180564 151786
rect 180616 141160 180668 141166
rect 180616 141102 180668 141108
rect 180628 139890 180656 141102
rect 180812 140321 180840 199106
rect 182824 198756 182876 198762
rect 182824 198698 182876 198704
rect 181536 193180 181588 193186
rect 181536 193122 181588 193128
rect 181444 187332 181496 187338
rect 181444 187274 181496 187280
rect 180892 149116 180944 149122
rect 180892 149058 180944 149064
rect 180798 140312 180854 140321
rect 180798 140247 180854 140256
rect 180904 139890 180932 149058
rect 181456 140554 181484 187274
rect 181548 143478 181576 193122
rect 182088 149592 182140 149598
rect 182088 149534 182140 149540
rect 182100 149122 182128 149534
rect 182088 149116 182140 149122
rect 182088 149058 182140 149064
rect 182454 144936 182510 144945
rect 182454 144871 182510 144880
rect 181536 143472 181588 143478
rect 181536 143414 181588 143420
rect 182272 142044 182324 142050
rect 182272 141986 182324 141992
rect 181444 140548 181496 140554
rect 181444 140490 181496 140496
rect 181442 140312 181498 140321
rect 181442 140247 181498 140256
rect 181456 139890 181484 140247
rect 182086 140176 182142 140185
rect 182086 140111 182142 140120
rect 180628 139862 180688 139890
rect 180904 139862 181240 139890
rect 181456 139862 181792 139890
rect 182100 139466 182128 140111
rect 182178 139904 182234 139913
rect 182284 139890 182312 141986
rect 182468 139890 182496 144871
rect 182836 141030 182864 198698
rect 183204 198014 183232 199310
rect 183192 198008 183244 198014
rect 183192 197950 183244 197956
rect 183100 196104 183152 196110
rect 183100 196046 183152 196052
rect 182916 195968 182968 195974
rect 182916 195910 182968 195916
rect 182824 141024 182876 141030
rect 182824 140966 182876 140972
rect 182928 140978 182956 195910
rect 183112 192846 183140 196046
rect 183468 193316 183520 193322
rect 183468 193258 183520 193264
rect 183100 192840 183152 192846
rect 183100 192782 183152 192788
rect 183480 192506 183508 193258
rect 184112 193248 184164 193254
rect 184112 193190 184164 193196
rect 183468 192500 183520 192506
rect 183468 192442 183520 192448
rect 184124 192438 184152 193190
rect 184112 192432 184164 192438
rect 184112 192374 184164 192380
rect 185584 192296 185636 192302
rect 185584 192238 185636 192244
rect 183008 192092 183060 192098
rect 183008 192034 183060 192040
rect 183020 141114 183048 192034
rect 183100 191684 183152 191690
rect 183100 191626 183152 191632
rect 183112 141982 183140 191626
rect 184388 153128 184440 153134
rect 184388 153070 184440 153076
rect 184204 152312 184256 152318
rect 184204 152254 184256 152260
rect 183468 146192 183520 146198
rect 183468 146134 183520 146140
rect 183480 144945 183508 146134
rect 183466 144936 183522 144945
rect 183466 144871 183522 144880
rect 183100 141976 183152 141982
rect 183100 141918 183152 141924
rect 183020 141086 183232 141114
rect 182836 140842 182864 140966
rect 182928 140950 183140 140978
rect 182836 140814 183048 140842
rect 183020 139890 183048 140814
rect 183112 140214 183140 140950
rect 183100 140208 183152 140214
rect 183100 140150 183152 140156
rect 183204 140049 183232 141086
rect 183190 140040 183246 140049
rect 184216 140010 184244 152254
rect 184296 143336 184348 143342
rect 184296 143278 184348 143284
rect 184308 140865 184336 143278
rect 184400 142118 184428 153070
rect 184480 152992 184532 152998
rect 184480 152934 184532 152940
rect 184388 142112 184440 142118
rect 184388 142054 184440 142060
rect 184492 141137 184520 152934
rect 184572 152448 184624 152454
rect 184572 152390 184624 152396
rect 184584 141914 184612 152390
rect 184664 152380 184716 152386
rect 184664 152322 184716 152328
rect 184676 143274 184704 152322
rect 184756 149728 184808 149734
rect 184756 149670 184808 149676
rect 184664 143268 184716 143274
rect 184664 143210 184716 143216
rect 184572 141908 184624 141914
rect 184572 141850 184624 141856
rect 184478 141128 184534 141137
rect 184478 141063 184534 141072
rect 184294 140856 184350 140865
rect 184294 140791 184350 140800
rect 183190 139975 183246 139984
rect 184204 140004 184256 140010
rect 184204 139946 184256 139952
rect 184308 139890 184336 140791
rect 184768 140049 184796 149670
rect 185308 149048 185360 149054
rect 185308 148990 185360 148996
rect 185032 148300 185084 148306
rect 185032 148242 185084 148248
rect 184848 141772 184900 141778
rect 184848 141714 184900 141720
rect 184860 141098 184888 141714
rect 184848 141092 184900 141098
rect 184848 141034 184900 141040
rect 184754 140040 184810 140049
rect 184754 139975 184810 139984
rect 184860 139890 184888 141034
rect 184938 140584 184994 140593
rect 184938 140519 184994 140528
rect 184952 140298 184980 140519
rect 185044 140457 185072 148242
rect 185030 140448 185086 140457
rect 185030 140383 185086 140392
rect 185030 140312 185086 140321
rect 184952 140270 185030 140298
rect 185030 140247 185086 140256
rect 182234 139862 182344 139890
rect 182468 139862 182896 139890
rect 183020 139862 183448 139890
rect 184000 139862 184336 139890
rect 184552 139862 184888 139890
rect 185044 139890 185072 140247
rect 185320 139913 185348 148990
rect 185596 143585 185624 192238
rect 185676 153196 185728 153202
rect 185676 153138 185728 153144
rect 185582 143576 185638 143585
rect 185582 143511 185638 143520
rect 185584 143404 185636 143410
rect 185584 143346 185636 143352
rect 185596 142322 185624 143346
rect 185584 142316 185636 142322
rect 185584 142258 185636 142264
rect 185306 139904 185362 139913
rect 185044 139862 185104 139890
rect 182178 139839 182234 139848
rect 185596 139890 185624 142258
rect 185688 140622 185716 153138
rect 185768 153060 185820 153066
rect 185768 153002 185820 153008
rect 185676 140616 185728 140622
rect 185676 140558 185728 140564
rect 185596 139862 185656 139890
rect 185306 139839 185362 139848
rect 182088 139460 182140 139466
rect 182088 139402 182140 139408
rect 185780 139398 185808 153002
rect 185860 152924 185912 152930
rect 185860 152866 185912 152872
rect 185872 140350 185900 152866
rect 186320 148980 186372 148986
rect 186320 148922 186372 148928
rect 186332 140865 186360 148922
rect 186424 141409 186452 280162
rect 186688 275324 186740 275330
rect 186688 275266 186740 275272
rect 186700 274718 186728 275266
rect 186504 274712 186556 274718
rect 186504 274654 186556 274660
rect 186688 274712 186740 274718
rect 186688 274654 186740 274660
rect 186516 142905 186544 274654
rect 187700 273964 187752 273970
rect 187700 273906 187752 273912
rect 187712 273290 187740 273906
rect 187700 273284 187752 273290
rect 187700 273226 187752 273232
rect 186594 262984 186650 262993
rect 186594 262919 186650 262928
rect 187148 262948 187200 262954
rect 186608 144362 186636 262919
rect 187148 262890 187200 262896
rect 187056 262268 187108 262274
rect 187056 262210 187108 262216
rect 186964 260160 187016 260166
rect 186964 260102 187016 260108
rect 186870 259992 186926 260001
rect 186870 259927 186926 259936
rect 186688 259888 186740 259894
rect 186688 259830 186740 259836
rect 186596 144356 186648 144362
rect 186596 144298 186648 144304
rect 186700 143070 186728 259830
rect 186780 259820 186832 259826
rect 186780 259762 186832 259768
rect 186688 143064 186740 143070
rect 186688 143006 186740 143012
rect 186792 142934 186820 259762
rect 186884 143449 186912 259927
rect 186976 149666 187004 260102
rect 187068 199170 187096 262210
rect 187160 199442 187188 262890
rect 187240 259548 187292 259554
rect 187240 259490 187292 259496
rect 187252 202881 187280 259490
rect 187238 202872 187294 202881
rect 187238 202807 187294 202816
rect 187240 199776 187292 199782
rect 187240 199718 187292 199724
rect 187148 199436 187200 199442
rect 187148 199378 187200 199384
rect 187056 199164 187108 199170
rect 187056 199106 187108 199112
rect 187056 197260 187108 197266
rect 187056 197202 187108 197208
rect 186964 149660 187016 149666
rect 186964 149602 187016 149608
rect 186962 149152 187018 149161
rect 186962 149087 187018 149096
rect 186870 143440 186926 143449
rect 186870 143375 186926 143384
rect 186780 142928 186832 142934
rect 186502 142896 186558 142905
rect 186780 142870 186832 142876
rect 186502 142831 186558 142840
rect 186976 142769 187004 149087
rect 186962 142760 187018 142769
rect 186962 142695 187018 142704
rect 186410 141400 186466 141409
rect 186410 141335 186466 141344
rect 186318 140856 186374 140865
rect 186318 140791 186374 140800
rect 185950 140448 186006 140457
rect 185950 140383 186006 140392
rect 185860 140344 185912 140350
rect 185860 140286 185912 140292
rect 185964 139890 185992 140383
rect 185964 139862 186208 139890
rect 185768 139392 185820 139398
rect 155500 139334 155552 139340
rect 155682 139360 155738 139369
rect 155130 139295 155186 139304
rect 155682 139295 155738 139304
rect 159546 139360 159602 139369
rect 159546 139295 159602 139304
rect 160006 139360 160062 139369
rect 160006 139295 160062 139304
rect 163962 139360 164018 139369
rect 163962 139295 164018 139304
rect 179694 139360 179750 139369
rect 179694 139295 179750 139304
rect 180522 139360 180578 139369
rect 185768 139334 185820 139340
rect 186412 139392 186464 139398
rect 186412 139334 186464 139340
rect 180522 139295 180578 139304
rect 122378 138544 122434 138553
rect 122378 138479 122434 138488
rect 122944 138014 122972 139295
rect 186424 139233 186452 139334
rect 186410 139224 186466 139233
rect 186410 139159 186466 139168
rect 187068 138145 187096 197202
rect 187252 174593 187280 199718
rect 187238 174584 187294 174593
rect 187238 174519 187294 174528
rect 187712 143177 187740 273226
rect 192300 265668 192352 265674
rect 192300 265610 192352 265616
rect 190460 265056 190512 265062
rect 190460 264998 190512 265004
rect 188252 264240 188304 264246
rect 188252 264182 188304 264188
rect 188264 263634 188292 264182
rect 189264 263696 189316 263702
rect 189264 263638 189316 263644
rect 188252 263628 188304 263634
rect 188252 263570 188304 263576
rect 187976 263492 188028 263498
rect 187976 263434 188028 263440
rect 187988 262546 188016 263434
rect 187976 262540 188028 262546
rect 187976 262482 188028 262488
rect 187988 262313 188016 262482
rect 187974 262304 188030 262313
rect 187974 262239 188030 262248
rect 187792 261112 187844 261118
rect 187792 261054 187844 261060
rect 187804 259418 187832 261054
rect 187974 260128 188030 260137
rect 187974 260063 188030 260072
rect 187884 259956 187936 259962
rect 187884 259898 187936 259904
rect 187792 259412 187844 259418
rect 187792 259354 187844 259360
rect 187792 259276 187844 259282
rect 187792 259218 187844 259224
rect 187698 143168 187754 143177
rect 187698 143103 187754 143112
rect 187804 143041 187832 259218
rect 187790 143032 187846 143041
rect 187790 142967 187846 142976
rect 187896 141710 187924 259898
rect 187988 143002 188016 260063
rect 188158 259856 188214 259865
rect 188158 259791 188214 259800
rect 188068 259752 188120 259758
rect 188068 259694 188120 259700
rect 187976 142996 188028 143002
rect 187976 142938 188028 142944
rect 188080 142866 188108 259694
rect 188172 143313 188200 259791
rect 188264 259434 188292 263570
rect 188434 259720 188490 259729
rect 188434 259655 188490 259664
rect 188264 259406 188384 259434
rect 188252 259344 188304 259350
rect 188252 259286 188304 259292
rect 188264 198762 188292 259286
rect 188356 259282 188384 259406
rect 188344 259276 188396 259282
rect 188344 259218 188396 259224
rect 188342 201784 188398 201793
rect 188342 201719 188398 201728
rect 188252 198756 188304 198762
rect 188252 198698 188304 198704
rect 188252 194948 188304 194954
rect 188252 194890 188304 194896
rect 188158 143304 188214 143313
rect 188158 143239 188214 143248
rect 188068 142860 188120 142866
rect 188068 142802 188120 142808
rect 188160 142248 188212 142254
rect 188160 142190 188212 142196
rect 187884 141704 187936 141710
rect 187884 141646 187936 141652
rect 188172 138718 188200 142190
rect 188160 138712 188212 138718
rect 188160 138654 188212 138660
rect 187054 138136 187110 138145
rect 187054 138071 187110 138080
rect 122760 138009 122972 138014
rect 122746 138000 122972 138009
rect 122802 137986 122972 138000
rect 122746 137935 122802 137944
rect 122746 128480 122802 128489
rect 122746 128415 122802 128424
rect 122760 122913 122788 128415
rect 122746 122904 122802 122913
rect 122746 122839 122802 122848
rect 122746 122768 122802 122777
rect 122746 122703 122802 122712
rect 122760 113257 122788 122703
rect 122746 113248 122802 113257
rect 122746 113183 122802 113192
rect 122746 113112 122802 113121
rect 122746 113047 122802 113056
rect 122760 103601 122788 113047
rect 122746 103592 122802 103601
rect 122746 103527 122802 103536
rect 122746 103456 122802 103465
rect 122746 103391 122802 103400
rect 122760 93945 122788 103391
rect 122746 93936 122802 93945
rect 122746 93871 122802 93880
rect 122746 93800 122802 93809
rect 122746 93735 122802 93744
rect 122760 89729 122788 93735
rect 122746 89720 122802 89729
rect 122746 89655 122802 89664
rect 122470 81424 122526 81433
rect 122470 81359 122526 81368
rect 122484 78266 122512 81359
rect 188160 81252 188212 81258
rect 188160 81194 188212 81200
rect 186502 81016 186558 81025
rect 123484 80980 123536 80986
rect 186502 80951 186558 80960
rect 187146 81016 187202 81025
rect 187146 80951 187202 80960
rect 187422 81016 187478 81025
rect 187422 80951 187478 80960
rect 123484 80922 123536 80928
rect 123496 80714 123524 80922
rect 186412 80912 186464 80918
rect 186412 80854 186464 80860
rect 124036 80844 124088 80850
rect 124036 80786 124088 80792
rect 123484 80708 123536 80714
rect 123484 80650 123536 80656
rect 122838 80336 122894 80345
rect 122838 80271 122894 80280
rect 122472 78260 122524 78266
rect 122472 78202 122524 78208
rect 122852 77994 122880 80271
rect 124048 79898 124076 80786
rect 177762 80744 177818 80753
rect 129832 80708 129884 80714
rect 177652 80702 177762 80730
rect 178406 80744 178462 80753
rect 177762 80679 177818 80688
rect 177856 80708 177908 80714
rect 129832 80650 129884 80656
rect 183664 80714 183876 80730
rect 178406 80679 178462 80688
rect 183652 80708 183888 80714
rect 177856 80650 177908 80656
rect 129844 80102 129872 80650
rect 177764 80640 177816 80646
rect 132038 80608 132094 80617
rect 177868 80617 177896 80650
rect 177764 80582 177816 80588
rect 177854 80608 177910 80617
rect 132038 80543 132094 80552
rect 131946 80472 132002 80481
rect 131946 80407 132002 80416
rect 131762 80336 131818 80345
rect 131762 80271 131818 80280
rect 129832 80096 129884 80102
rect 129832 80038 129884 80044
rect 130844 80096 130896 80102
rect 130844 80038 130896 80044
rect 124036 79892 124088 79898
rect 124036 79834 124088 79840
rect 123484 79756 123536 79762
rect 123484 79698 123536 79704
rect 123024 79620 123076 79626
rect 123024 79562 123076 79568
rect 122840 77988 122892 77994
rect 122840 77930 122892 77936
rect 123036 76498 123064 79562
rect 123496 79422 123524 79698
rect 124126 79656 124182 79665
rect 124126 79591 124182 79600
rect 129096 79620 129148 79626
rect 123484 79416 123536 79422
rect 123484 79358 123536 79364
rect 124140 79218 124168 79591
rect 129096 79562 129148 79568
rect 126980 79552 127032 79558
rect 126980 79494 127032 79500
rect 124128 79212 124180 79218
rect 124128 79154 124180 79160
rect 125600 78872 125652 78878
rect 125600 78814 125652 78820
rect 125612 76673 125640 78814
rect 126992 77246 127020 79494
rect 126980 77240 127032 77246
rect 126980 77182 127032 77188
rect 127624 77240 127676 77246
rect 127624 77182 127676 77188
rect 125598 76664 125654 76673
rect 125598 76599 125654 76608
rect 123024 76492 123076 76498
rect 123024 76434 123076 76440
rect 121368 74520 121420 74526
rect 121368 74462 121420 74468
rect 123036 72622 123064 76434
rect 125612 73710 125640 76599
rect 124864 73704 124916 73710
rect 124864 73646 124916 73652
rect 125600 73704 125652 73710
rect 125600 73646 125652 73652
rect 122104 72616 122156 72622
rect 122104 72558 122156 72564
rect 123024 72616 123076 72622
rect 123024 72558 123076 72564
rect 124220 72616 124272 72622
rect 124220 72558 124272 72564
rect 121184 71596 121236 71602
rect 121184 71538 121236 71544
rect 120736 64846 121040 64874
rect 120092 16546 120672 16574
rect 119896 3392 119948 3398
rect 119896 3334 119948 3340
rect 118792 3052 118844 3058
rect 118792 2994 118844 3000
rect 118804 480 118832 2994
rect 119908 480 119936 3334
rect 117566 354 117678 480
rect 117332 326 117678 354
rect 117566 -960 117678 326
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 120644 354 120672 16546
rect 120736 3398 120764 64846
rect 120724 3392 120776 3398
rect 120724 3334 120776 3340
rect 122116 3058 122144 72558
rect 124232 16574 124260 72558
rect 124232 16546 124720 16574
rect 122288 3868 122340 3874
rect 122288 3810 122340 3816
rect 122104 3052 122156 3058
rect 122104 2994 122156 3000
rect 122300 480 122328 3810
rect 123484 3324 123536 3330
rect 123484 3266 123536 3272
rect 123496 480 123524 3266
rect 124692 480 124720 16546
rect 124876 3330 124904 73646
rect 127636 3874 127664 77182
rect 129108 72418 129136 79562
rect 129556 78872 129608 78878
rect 129556 78814 129608 78820
rect 129096 72412 129148 72418
rect 129096 72354 129148 72360
rect 129568 71126 129596 78814
rect 129648 77240 129700 77246
rect 129648 77182 129700 77188
rect 129660 76226 129688 77182
rect 129648 76220 129700 76226
rect 129648 76162 129700 76168
rect 129738 75304 129794 75313
rect 129738 75239 129794 75248
rect 128360 71120 128412 71126
rect 128360 71062 128412 71068
rect 129556 71120 129608 71126
rect 129556 71062 129608 71068
rect 127624 3868 127676 3874
rect 127624 3810 127676 3816
rect 128372 3534 128400 71062
rect 126980 3528 127032 3534
rect 126980 3470 127032 3476
rect 128360 3528 128412 3534
rect 128360 3470 128412 3476
rect 129372 3528 129424 3534
rect 129372 3470 129424 3476
rect 124864 3324 124916 3330
rect 124864 3266 124916 3272
rect 125876 3188 125928 3194
rect 125876 3130 125928 3136
rect 125888 480 125916 3130
rect 126992 480 127020 3470
rect 128176 3460 128228 3466
rect 128176 3402 128228 3408
rect 128188 480 128216 3402
rect 129384 480 129412 3470
rect 129752 3346 129780 75239
rect 129844 3738 129872 80038
rect 129924 79892 129976 79898
rect 129924 79834 129976 79840
rect 129936 78062 129964 79834
rect 130658 79792 130714 79801
rect 130658 79727 130714 79736
rect 130672 78810 130700 79727
rect 130752 79688 130804 79694
rect 130752 79630 130804 79636
rect 130660 78804 130712 78810
rect 130660 78746 130712 78752
rect 130382 78568 130438 78577
rect 130382 78503 130438 78512
rect 130396 78062 130424 78503
rect 129924 78056 129976 78062
rect 129924 77998 129976 78004
rect 130384 78056 130436 78062
rect 130384 77998 130436 78004
rect 129832 3732 129884 3738
rect 129832 3674 129884 3680
rect 129936 3602 129964 77998
rect 130382 75984 130438 75993
rect 130382 75919 130438 75928
rect 130016 72480 130068 72486
rect 130016 72422 130068 72428
rect 129924 3596 129976 3602
rect 129924 3538 129976 3544
rect 130028 3534 130056 72422
rect 130016 3528 130068 3534
rect 130016 3470 130068 3476
rect 130396 3466 130424 75919
rect 130672 70394 130700 78746
rect 130764 72298 130792 79630
rect 130856 78130 130884 80038
rect 130934 79792 130990 79801
rect 130934 79727 130990 79736
rect 130948 78198 130976 79727
rect 131672 79552 131724 79558
rect 131672 79494 131724 79500
rect 130936 78192 130988 78198
rect 130936 78134 130988 78140
rect 130844 78124 130896 78130
rect 130844 78066 130896 78072
rect 130936 77920 130988 77926
rect 130936 77862 130988 77868
rect 130948 75313 130976 77862
rect 131212 77852 131264 77858
rect 131212 77794 131264 77800
rect 130934 75304 130990 75313
rect 130934 75239 130990 75248
rect 131120 74520 131172 74526
rect 131120 74462 131172 74468
rect 131026 72584 131082 72593
rect 131026 72519 131082 72528
rect 131040 72486 131068 72519
rect 131028 72480 131080 72486
rect 131028 72422 131080 72428
rect 130764 72270 131068 72298
rect 130672 70366 130976 70394
rect 130948 3602 130976 70366
rect 131040 3738 131068 72270
rect 131028 3732 131080 3738
rect 131028 3674 131080 3680
rect 130936 3596 130988 3602
rect 130936 3538 130988 3544
rect 130384 3460 130436 3466
rect 130384 3402 130436 3408
rect 129752 3318 130608 3346
rect 130580 480 130608 3318
rect 131132 3194 131160 74462
rect 131224 16574 131252 77794
rect 131684 77586 131712 79494
rect 131672 77580 131724 77586
rect 131672 77522 131724 77528
rect 131684 76786 131712 77522
rect 131592 76758 131712 76786
rect 131592 75993 131620 76758
rect 131672 76696 131724 76702
rect 131672 76638 131724 76644
rect 131684 76294 131712 76638
rect 131672 76288 131724 76294
rect 131672 76230 131724 76236
rect 131578 75984 131634 75993
rect 131578 75919 131634 75928
rect 131224 16546 131344 16574
rect 131120 3188 131172 3194
rect 131120 3130 131172 3136
rect 121062 354 121174 480
rect 120644 326 121174 354
rect 121062 -960 121174 326
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131316 354 131344 16546
rect 131776 3806 131804 80271
rect 131960 79966 131988 80407
rect 132052 80170 132080 80543
rect 177776 80306 177804 80582
rect 177854 80543 177910 80552
rect 177764 80300 177816 80306
rect 177764 80242 177816 80248
rect 178316 80232 178368 80238
rect 178316 80174 178368 80180
rect 132040 80164 132092 80170
rect 132040 80106 132092 80112
rect 178132 80164 178184 80170
rect 178132 80106 178184 80112
rect 177856 80096 177908 80102
rect 132052 80022 132388 80050
rect 177856 80038 177908 80044
rect 131948 79960 132000 79966
rect 131868 79920 131948 79948
rect 131764 3800 131816 3806
rect 131764 3742 131816 3748
rect 131868 3398 131896 79920
rect 131948 79902 132000 79908
rect 131946 78568 132002 78577
rect 131946 78503 132002 78512
rect 131856 3392 131908 3398
rect 131856 3334 131908 3340
rect 131960 3330 131988 78503
rect 132052 77897 132080 80022
rect 132466 79948 132494 80036
rect 132558 79971 132586 80036
rect 132328 79937 132494 79948
rect 132314 79928 132494 79937
rect 132370 79920 132494 79928
rect 132544 79962 132600 79971
rect 132544 79897 132600 79906
rect 132314 79863 132370 79872
rect 132650 79778 132678 80036
rect 132742 79966 132770 80036
rect 132834 79966 132862 80036
rect 132730 79960 132782 79966
rect 132730 79902 132782 79908
rect 132822 79960 132874 79966
rect 132822 79902 132874 79908
rect 132926 79898 132954 80036
rect 133018 79966 133046 80036
rect 133110 79971 133138 80036
rect 133006 79960 133058 79966
rect 133006 79902 133058 79908
rect 133096 79962 133152 79971
rect 133202 79966 133230 80036
rect 133294 79966 133322 80036
rect 133386 79966 133414 80036
rect 133478 79966 133506 80036
rect 132914 79892 132966 79898
rect 133096 79897 133152 79906
rect 133190 79960 133242 79966
rect 133190 79902 133242 79908
rect 133282 79960 133334 79966
rect 133282 79902 133334 79908
rect 133374 79960 133426 79966
rect 133374 79902 133426 79908
rect 133466 79960 133518 79966
rect 133466 79902 133518 79908
rect 132914 79834 132966 79840
rect 132316 79756 132368 79762
rect 132316 79698 132368 79704
rect 132604 79750 132678 79778
rect 133096 79826 133152 79835
rect 133570 79801 133598 80036
rect 133662 79966 133690 80036
rect 133754 79966 133782 80036
rect 133650 79960 133702 79966
rect 133650 79902 133702 79908
rect 133742 79960 133794 79966
rect 133742 79902 133794 79908
rect 133846 79898 133874 80036
rect 133938 79937 133966 80036
rect 133924 79928 133980 79937
rect 133834 79892 133886 79898
rect 133924 79863 133980 79872
rect 133834 79834 133886 79840
rect 133696 79824 133748 79830
rect 132776 79756 132828 79762
rect 133096 79761 133152 79770
rect 133556 79792 133612 79801
rect 132224 79688 132276 79694
rect 132224 79630 132276 79636
rect 132236 79354 132264 79630
rect 132328 79422 132356 79698
rect 132408 79552 132460 79558
rect 132408 79494 132460 79500
rect 132316 79416 132368 79422
rect 132316 79358 132368 79364
rect 132132 79348 132184 79354
rect 132132 79290 132184 79296
rect 132224 79348 132276 79354
rect 132224 79290 132276 79296
rect 132038 77888 132094 77897
rect 132144 77858 132172 79290
rect 132316 78668 132368 78674
rect 132316 78610 132368 78616
rect 132038 77823 132094 77832
rect 132132 77852 132184 77858
rect 132132 77794 132184 77800
rect 132328 74526 132356 78610
rect 132420 75070 132448 79494
rect 132604 76265 132632 79750
rect 132776 79698 132828 79704
rect 132684 78124 132736 78130
rect 132684 78066 132736 78072
rect 132696 77926 132724 78066
rect 132684 77920 132736 77926
rect 132684 77862 132736 77868
rect 132590 76256 132646 76265
rect 132590 76191 132646 76200
rect 132408 75064 132460 75070
rect 132408 75006 132460 75012
rect 132316 74520 132368 74526
rect 132316 74462 132368 74468
rect 132684 73704 132736 73710
rect 132684 73646 132736 73652
rect 132500 72480 132552 72486
rect 132500 72422 132552 72428
rect 132512 70174 132540 72422
rect 132500 70168 132552 70174
rect 132500 70110 132552 70116
rect 132512 37942 132540 70110
rect 132696 60722 132724 73646
rect 132788 63510 132816 79698
rect 133110 79676 133138 79761
rect 133328 79756 133380 79762
rect 134030 79778 134058 80036
rect 134122 79830 134150 80036
rect 133696 79766 133748 79772
rect 133556 79727 133612 79736
rect 133328 79698 133380 79704
rect 132880 79648 133138 79676
rect 133236 79688 133288 79694
rect 132776 63504 132828 63510
rect 132776 63446 132828 63452
rect 132684 60716 132736 60722
rect 132684 60658 132736 60664
rect 132880 53786 132908 79648
rect 133236 79630 133288 79636
rect 133248 77897 133276 79630
rect 133234 77888 133290 77897
rect 133234 77823 133290 77832
rect 133248 72457 133276 77823
rect 133234 72448 133290 72457
rect 133234 72383 133290 72392
rect 133340 67634 133368 79698
rect 133512 79688 133564 79694
rect 133512 79630 133564 79636
rect 133604 79688 133656 79694
rect 133604 79630 133656 79636
rect 133418 77888 133474 77897
rect 133418 77823 133474 77832
rect 133432 71058 133460 77823
rect 133524 72486 133552 79630
rect 133512 72480 133564 72486
rect 133512 72422 133564 72428
rect 133420 71052 133472 71058
rect 133420 70994 133472 71000
rect 133616 70106 133644 79630
rect 133708 73710 133736 79766
rect 133788 79756 133840 79762
rect 133788 79698 133840 79704
rect 133984 79750 134058 79778
rect 134110 79824 134162 79830
rect 134110 79766 134162 79772
rect 133800 74361 133828 79698
rect 133984 79676 134012 79750
rect 134214 79676 134242 80036
rect 134306 79898 134334 80036
rect 134398 79966 134426 80036
rect 134386 79960 134438 79966
rect 134490 79937 134518 80036
rect 134386 79902 134438 79908
rect 134476 79928 134532 79937
rect 134294 79892 134346 79898
rect 134582 79898 134610 80036
rect 134476 79863 134532 79872
rect 134570 79892 134622 79898
rect 134294 79834 134346 79840
rect 134570 79834 134622 79840
rect 134432 79824 134484 79830
rect 134338 79792 134394 79801
rect 134432 79766 134484 79772
rect 134338 79727 134340 79736
rect 134392 79727 134394 79736
rect 134340 79698 134392 79704
rect 133892 79648 134012 79676
rect 134168 79648 134242 79676
rect 133892 78606 133920 79648
rect 134064 79620 134116 79626
rect 134064 79562 134116 79568
rect 133880 78600 133932 78606
rect 133880 78542 133932 78548
rect 133972 77716 134024 77722
rect 133972 77658 134024 77664
rect 133984 77625 134012 77658
rect 133970 77616 134026 77625
rect 133970 77551 134026 77560
rect 134076 75478 134104 79562
rect 134064 75472 134116 75478
rect 134064 75414 134116 75420
rect 133786 74352 133842 74361
rect 133786 74287 133842 74296
rect 133696 73704 133748 73710
rect 133696 73646 133748 73652
rect 134168 70378 134196 79648
rect 134340 77444 134392 77450
rect 134340 77386 134392 77392
rect 134248 74180 134300 74186
rect 134248 74122 134300 74128
rect 134156 70372 134208 70378
rect 134156 70314 134208 70320
rect 133604 70100 133656 70106
rect 133604 70042 133656 70048
rect 132972 67606 133368 67634
rect 132972 56574 133000 67606
rect 133878 67008 133934 67017
rect 133878 66943 133934 66952
rect 132960 56568 133012 56574
rect 132960 56510 133012 56516
rect 132868 53780 132920 53786
rect 132868 53722 132920 53728
rect 132500 37936 132552 37942
rect 132500 37878 132552 37884
rect 131948 3324 132000 3330
rect 131948 3266 132000 3272
rect 132960 3324 133012 3330
rect 132960 3266 133012 3272
rect 132972 480 133000 3266
rect 131734 354 131846 480
rect 131316 326 131846 354
rect 131734 -960 131846 326
rect 132930 -960 133042 480
rect 133892 354 133920 66943
rect 134168 7614 134196 70314
rect 134260 26926 134288 74122
rect 134352 64190 134380 77386
rect 134340 64184 134392 64190
rect 134340 64126 134392 64132
rect 134444 62082 134472 79766
rect 134674 79744 134702 80036
rect 134536 79716 134702 79744
rect 134766 79744 134794 80036
rect 134858 79903 134886 80036
rect 134844 79894 134900 79903
rect 134844 79829 134900 79838
rect 134766 79716 134840 79744
rect 134536 75954 134564 79716
rect 134812 79665 134840 79716
rect 134950 79676 134978 80036
rect 135042 79830 135070 80036
rect 135134 79898 135162 80036
rect 135226 79898 135254 80036
rect 135318 79898 135346 80036
rect 135410 79966 135438 80036
rect 135398 79960 135450 79966
rect 135398 79902 135450 79908
rect 135122 79892 135174 79898
rect 135122 79834 135174 79840
rect 135214 79892 135266 79898
rect 135214 79834 135266 79840
rect 135306 79892 135358 79898
rect 135306 79834 135358 79840
rect 135030 79824 135082 79830
rect 135502 79812 135530 80036
rect 135030 79766 135082 79772
rect 135456 79784 135530 79812
rect 135168 79756 135220 79762
rect 135168 79698 135220 79704
rect 134614 79656 134670 79665
rect 134614 79591 134670 79600
rect 134798 79656 134854 79665
rect 134798 79591 134854 79600
rect 134904 79648 134978 79676
rect 134524 75948 134576 75954
rect 134524 75890 134576 75896
rect 134524 75472 134576 75478
rect 134524 75414 134576 75420
rect 134432 62076 134484 62082
rect 134432 62018 134484 62024
rect 134536 57934 134564 75414
rect 134524 57928 134576 57934
rect 134524 57870 134576 57876
rect 134628 51066 134656 79591
rect 134800 79552 134852 79558
rect 134800 79494 134852 79500
rect 134812 78577 134840 79494
rect 134798 78568 134854 78577
rect 134798 78503 134854 78512
rect 134812 77450 134840 78503
rect 134800 77444 134852 77450
rect 134800 77386 134852 77392
rect 134800 77308 134852 77314
rect 134800 77250 134852 77256
rect 134812 76634 134840 77250
rect 134800 76628 134852 76634
rect 134800 76570 134852 76576
rect 134708 75948 134760 75954
rect 134708 75890 134760 75896
rect 134720 71534 134748 75890
rect 134708 71528 134760 71534
rect 134708 71470 134760 71476
rect 134904 67634 134932 79648
rect 135180 79642 135208 79698
rect 135076 79620 135128 79626
rect 135180 79614 135300 79642
rect 135076 79562 135128 79568
rect 134984 79552 135036 79558
rect 134984 79494 135036 79500
rect 134996 77790 135024 79494
rect 134984 77784 135036 77790
rect 134984 77726 135036 77732
rect 135088 73953 135116 79562
rect 135272 78792 135300 79614
rect 135180 78764 135300 78792
rect 135180 74186 135208 78764
rect 135260 78668 135312 78674
rect 135260 78610 135312 78616
rect 135168 74180 135220 74186
rect 135168 74122 135220 74128
rect 135074 73944 135130 73953
rect 135074 73879 135130 73888
rect 135272 69698 135300 78610
rect 135456 75614 135484 79784
rect 135594 79744 135622 80036
rect 135686 79898 135714 80036
rect 135778 79937 135806 80036
rect 135870 79966 135898 80036
rect 135858 79960 135910 79966
rect 135764 79928 135820 79937
rect 135674 79892 135726 79898
rect 135858 79902 135910 79908
rect 135962 79898 135990 80036
rect 135764 79863 135820 79872
rect 135950 79892 136002 79898
rect 135674 79834 135726 79840
rect 135950 79834 136002 79840
rect 135812 79824 135864 79830
rect 135812 79766 135864 79772
rect 135902 79792 135958 79801
rect 135548 79716 135622 79744
rect 135444 75608 135496 75614
rect 135444 75550 135496 75556
rect 135456 71774 135484 75550
rect 135548 73030 135576 79716
rect 135626 79656 135682 79665
rect 135626 79591 135628 79600
rect 135680 79591 135682 79600
rect 135720 79620 135772 79626
rect 135628 79562 135680 79568
rect 135720 79562 135772 79568
rect 135536 73024 135588 73030
rect 135536 72966 135588 72972
rect 135364 71746 135484 71774
rect 135260 69692 135312 69698
rect 135260 69634 135312 69640
rect 134812 67606 134932 67634
rect 134812 67522 134840 67606
rect 134800 67516 134852 67522
rect 134800 67458 134852 67464
rect 134616 51060 134668 51066
rect 134616 51002 134668 51008
rect 135260 45620 135312 45626
rect 135260 45562 135312 45568
rect 134248 26920 134300 26926
rect 134248 26862 134300 26868
rect 134156 7608 134208 7614
rect 134156 7550 134208 7556
rect 135272 480 135300 45562
rect 135364 24138 135392 71746
rect 135444 71528 135496 71534
rect 135444 71470 135496 71476
rect 135456 71398 135484 71470
rect 135444 71392 135496 71398
rect 135444 71334 135496 71340
rect 135456 28286 135484 71334
rect 135640 61402 135668 79562
rect 135732 78334 135760 79562
rect 135720 78328 135772 78334
rect 135720 78270 135772 78276
rect 135718 77888 135774 77897
rect 135718 77823 135774 77832
rect 135732 71330 135760 77823
rect 135824 76537 135852 79766
rect 136054 79744 136082 80036
rect 135902 79727 135904 79736
rect 135956 79727 135958 79736
rect 135904 79698 135956 79704
rect 136008 79716 136082 79744
rect 135916 78674 135944 79698
rect 135904 78668 135956 78674
rect 135904 78610 135956 78616
rect 136008 78402 136036 79716
rect 136146 79676 136174 80036
rect 136238 79744 136266 80036
rect 136330 79898 136358 80036
rect 136318 79892 136370 79898
rect 136318 79834 136370 79840
rect 136422 79812 136450 80036
rect 136514 79971 136542 80036
rect 136500 79962 136556 79971
rect 136500 79897 136556 79906
rect 136422 79784 136496 79812
rect 136238 79716 136404 79744
rect 136100 79648 136174 79676
rect 135996 78396 136048 78402
rect 135996 78338 136048 78344
rect 135994 77616 136050 77625
rect 135994 77551 136050 77560
rect 136008 76566 136036 77551
rect 135996 76560 136048 76566
rect 135810 76528 135866 76537
rect 135996 76502 136048 76508
rect 135810 76463 135866 76472
rect 135720 71324 135772 71330
rect 135720 71266 135772 71272
rect 136100 70394 136128 79648
rect 136272 79620 136324 79626
rect 136272 79562 136324 79568
rect 136180 79552 136232 79558
rect 136180 79494 136232 79500
rect 136192 78577 136220 79494
rect 136178 78568 136234 78577
rect 136178 78503 136234 78512
rect 135732 70366 136128 70394
rect 135732 68746 135760 70366
rect 135720 68740 135772 68746
rect 135720 68682 135772 68688
rect 136192 67634 136220 78503
rect 136284 74225 136312 79562
rect 136376 78724 136404 79716
rect 136468 78792 136496 79784
rect 136606 79744 136634 80036
rect 136698 79812 136726 80036
rect 136790 79966 136818 80036
rect 136882 79966 136910 80036
rect 136778 79960 136830 79966
rect 136778 79902 136830 79908
rect 136870 79960 136922 79966
rect 136974 79937 137002 80036
rect 136870 79902 136922 79908
rect 136960 79928 137016 79937
rect 137066 79898 137094 80036
rect 136960 79863 137016 79872
rect 137054 79892 137106 79898
rect 137054 79834 137106 79840
rect 137158 79830 137186 80036
rect 137250 79966 137278 80036
rect 137238 79960 137290 79966
rect 137238 79902 137290 79908
rect 137342 79835 137370 80036
rect 137434 79966 137462 80036
rect 137422 79960 137474 79966
rect 137422 79902 137474 79908
rect 137146 79824 137198 79830
rect 136698 79784 136772 79812
rect 136606 79716 136680 79744
rect 136652 79665 136680 79716
rect 136638 79656 136694 79665
rect 136638 79591 136694 79600
rect 136744 78792 136772 79784
rect 137146 79766 137198 79772
rect 137328 79826 137384 79835
rect 137008 79756 137060 79762
rect 137328 79761 137384 79770
rect 137526 79778 137554 80036
rect 137618 79966 137646 80036
rect 137606 79960 137658 79966
rect 137606 79902 137658 79908
rect 137710 79812 137738 80036
rect 137664 79784 137738 79812
rect 137526 79750 137600 79778
rect 137008 79698 137060 79704
rect 136916 79688 136968 79694
rect 136822 79656 136878 79665
rect 136916 79630 136968 79636
rect 136822 79591 136878 79600
rect 136468 78764 136588 78792
rect 136376 78696 136496 78724
rect 136270 74216 136326 74225
rect 136270 74151 136326 74160
rect 136468 73817 136496 78696
rect 136454 73808 136510 73817
rect 136454 73743 136510 73752
rect 136560 71534 136588 78764
rect 136652 78764 136772 78792
rect 136652 77246 136680 78764
rect 136732 78668 136784 78674
rect 136732 78610 136784 78616
rect 136744 78577 136772 78610
rect 136730 78568 136786 78577
rect 136730 78503 136786 78512
rect 136730 77888 136786 77897
rect 136730 77823 136786 77832
rect 136744 77654 136772 77823
rect 136732 77648 136784 77654
rect 136732 77590 136784 77596
rect 136640 77240 136692 77246
rect 136640 77182 136692 77188
rect 136548 71528 136600 71534
rect 136548 71470 136600 71476
rect 136836 70394 136864 79591
rect 136928 78674 136956 79630
rect 136916 78668 136968 78674
rect 136916 78610 136968 78616
rect 136914 78568 136970 78577
rect 136914 78503 136970 78512
rect 136928 77314 136956 78503
rect 136916 77308 136968 77314
rect 136916 77250 136968 77256
rect 136916 74180 136968 74186
rect 136916 74122 136968 74128
rect 136744 70366 136864 70394
rect 136192 67606 136404 67634
rect 135628 61396 135680 61402
rect 135628 61338 135680 61344
rect 136376 35222 136404 67606
rect 136744 64874 136772 70366
rect 136652 64846 136772 64874
rect 136652 43450 136680 64846
rect 136640 43444 136692 43450
rect 136640 43386 136692 43392
rect 136928 42090 136956 74122
rect 137020 70310 137048 79698
rect 137376 79688 137428 79694
rect 137098 79656 137154 79665
rect 137098 79591 137154 79600
rect 137282 79656 137338 79665
rect 137572 79676 137600 79750
rect 137376 79630 137428 79636
rect 137480 79648 137600 79676
rect 137282 79591 137284 79600
rect 137112 79506 137140 79591
rect 137336 79591 137338 79600
rect 137284 79562 137336 79568
rect 137388 79506 137416 79630
rect 137112 79478 137416 79506
rect 137100 78668 137152 78674
rect 137100 78610 137152 78616
rect 137008 70304 137060 70310
rect 137008 70246 137060 70252
rect 137112 67590 137140 78610
rect 137284 78600 137336 78606
rect 137190 78568 137246 78577
rect 137284 78542 137336 78548
rect 137190 78503 137246 78512
rect 137204 78470 137232 78503
rect 137192 78464 137244 78470
rect 137192 78406 137244 78412
rect 137192 77240 137244 77246
rect 137192 77182 137244 77188
rect 137100 67584 137152 67590
rect 137100 67526 137152 67532
rect 137204 66230 137232 77182
rect 137192 66224 137244 66230
rect 137192 66166 137244 66172
rect 136916 42084 136968 42090
rect 136916 42026 136968 42032
rect 136364 35216 136416 35222
rect 136364 35158 136416 35164
rect 135444 28280 135496 28286
rect 135444 28222 135496 28228
rect 135352 24132 135404 24138
rect 135352 24074 135404 24080
rect 137296 3670 137324 78542
rect 137388 78538 137416 79478
rect 137376 78532 137428 78538
rect 137376 78474 137428 78480
rect 137480 77042 137508 79648
rect 137560 79552 137612 79558
rect 137560 79494 137612 79500
rect 137572 78577 137600 79494
rect 137558 78568 137614 78577
rect 137558 78503 137614 78512
rect 137560 78396 137612 78402
rect 137560 78338 137612 78344
rect 137572 77625 137600 78338
rect 137664 78198 137692 79784
rect 137802 79744 137830 80036
rect 137894 79937 137922 80036
rect 137986 79966 138014 80036
rect 137974 79960 138026 79966
rect 137880 79928 137936 79937
rect 137974 79902 138026 79908
rect 137880 79863 137936 79872
rect 138078 79801 138106 80036
rect 138170 79830 138198 80036
rect 138262 79971 138290 80036
rect 138248 79962 138304 79971
rect 138354 79966 138382 80036
rect 138248 79897 138304 79906
rect 138342 79960 138394 79966
rect 138446 79937 138474 80036
rect 138342 79902 138394 79908
rect 138432 79928 138488 79937
rect 138432 79863 138434 79872
rect 138486 79863 138488 79872
rect 138434 79834 138486 79840
rect 138158 79824 138210 79830
rect 137756 79716 137830 79744
rect 137926 79792 137982 79801
rect 137926 79727 137982 79736
rect 138064 79792 138120 79801
rect 138538 79778 138566 80036
rect 138158 79766 138210 79772
rect 138064 79727 138120 79736
rect 138308 79750 138566 79778
rect 137756 78674 137784 79716
rect 137836 79620 137888 79626
rect 137836 79562 137888 79568
rect 137744 78668 137796 78674
rect 137744 78610 137796 78616
rect 137848 78606 137876 79562
rect 137836 78600 137888 78606
rect 137836 78542 137888 78548
rect 137744 78532 137796 78538
rect 137744 78474 137796 78480
rect 137652 78192 137704 78198
rect 137652 78134 137704 78140
rect 137558 77616 137614 77625
rect 137558 77551 137614 77560
rect 137558 77480 137614 77489
rect 137558 77415 137614 77424
rect 137468 77036 137520 77042
rect 137468 76978 137520 76984
rect 137572 64874 137600 77415
rect 137756 72554 137784 78474
rect 137834 78296 137890 78305
rect 137834 78231 137890 78240
rect 137848 77926 137876 78231
rect 137836 77920 137888 77926
rect 137836 77862 137888 77868
rect 137940 74186 137968 79727
rect 138020 79688 138072 79694
rect 138020 79630 138072 79636
rect 138032 78577 138060 79630
rect 138204 79552 138256 79558
rect 138204 79494 138256 79500
rect 138018 78568 138074 78577
rect 138018 78503 138074 78512
rect 138110 78432 138166 78441
rect 138110 78367 138166 78376
rect 138124 78334 138152 78367
rect 138112 78328 138164 78334
rect 138112 78270 138164 78276
rect 138110 77888 138166 77897
rect 138110 77823 138166 77832
rect 137928 74180 137980 74186
rect 137928 74122 137980 74128
rect 137744 72548 137796 72554
rect 137744 72490 137796 72496
rect 138020 71188 138072 71194
rect 138020 71130 138072 71136
rect 137388 64846 137600 64874
rect 137388 58682 137416 64846
rect 137376 58676 137428 58682
rect 137376 58618 137428 58624
rect 138032 6186 138060 71130
rect 138124 69834 138152 77823
rect 138216 70038 138244 79494
rect 138308 77353 138336 79750
rect 138388 79688 138440 79694
rect 138630 79676 138658 80036
rect 138722 79778 138750 80036
rect 138814 79966 138842 80036
rect 138906 79966 138934 80036
rect 138802 79960 138854 79966
rect 138802 79902 138854 79908
rect 138894 79960 138946 79966
rect 138998 79937 139026 80036
rect 138894 79902 138946 79908
rect 138984 79928 139040 79937
rect 138984 79863 139040 79872
rect 138940 79824 138992 79830
rect 138846 79792 138902 79801
rect 138722 79750 138846 79778
rect 139090 79801 139118 80036
rect 139182 79898 139210 80036
rect 139274 79966 139302 80036
rect 139262 79960 139314 79966
rect 139262 79902 139314 79908
rect 139366 79898 139394 80036
rect 139170 79892 139222 79898
rect 139170 79834 139222 79840
rect 139354 79892 139406 79898
rect 139354 79834 139406 79840
rect 138940 79766 138992 79772
rect 139076 79792 139132 79801
rect 138846 79727 138902 79736
rect 138388 79630 138440 79636
rect 138584 79648 138658 79676
rect 138294 77344 138350 77353
rect 138294 77279 138350 77288
rect 138308 73846 138336 77279
rect 138296 73840 138348 73846
rect 138296 73782 138348 73788
rect 138204 70032 138256 70038
rect 138204 69974 138256 69980
rect 138112 69828 138164 69834
rect 138112 69770 138164 69776
rect 138216 40730 138244 69974
rect 138400 64874 138428 79630
rect 138480 79620 138532 79626
rect 138480 79562 138532 79568
rect 138308 64846 138428 64874
rect 138204 40724 138256 40730
rect 138204 40666 138256 40672
rect 138308 39370 138336 64846
rect 138492 64802 138520 79562
rect 138584 78305 138612 79648
rect 138756 78328 138808 78334
rect 138570 78296 138626 78305
rect 138570 78231 138626 78240
rect 138754 78296 138756 78305
rect 138808 78296 138810 78305
rect 138754 78231 138810 78240
rect 138860 75914 138888 79727
rect 138952 77489 138980 79766
rect 139076 79727 139132 79736
rect 139306 79792 139362 79801
rect 139458 79744 139486 80036
rect 139550 79937 139578 80036
rect 139536 79928 139592 79937
rect 139536 79863 139592 79872
rect 139642 79778 139670 80036
rect 139734 79937 139762 80036
rect 139720 79928 139776 79937
rect 139720 79863 139776 79872
rect 139826 79830 139854 80036
rect 139814 79824 139866 79830
rect 139306 79727 139362 79736
rect 139032 79688 139084 79694
rect 139032 79630 139084 79636
rect 138938 77480 138994 77489
rect 138938 77415 138994 77424
rect 139044 75914 139072 79630
rect 139124 79620 139176 79626
rect 139124 79562 139176 79568
rect 138768 75886 138888 75914
rect 138952 75886 139072 75914
rect 138768 75274 138796 75886
rect 138756 75268 138808 75274
rect 138756 75210 138808 75216
rect 138952 70530 138980 75886
rect 139136 71194 139164 79562
rect 139216 79552 139268 79558
rect 139216 79494 139268 79500
rect 139228 78985 139256 79494
rect 139214 78976 139270 78985
rect 139214 78911 139270 78920
rect 139124 71188 139176 71194
rect 139124 71130 139176 71136
rect 138676 70502 138980 70530
rect 138676 68882 138704 70502
rect 139228 70394 139256 78911
rect 139320 72962 139348 79727
rect 139412 79716 139486 79744
rect 139550 79750 139670 79778
rect 139812 79792 139814 79801
rect 139866 79792 139868 79801
rect 139412 77897 139440 79716
rect 139550 79676 139578 79750
rect 139812 79727 139868 79736
rect 139504 79648 139578 79676
rect 139768 79688 139820 79694
rect 139398 77888 139454 77897
rect 139398 77823 139454 77832
rect 139504 75818 139532 79648
rect 139918 79676 139946 80036
rect 139768 79630 139820 79636
rect 139872 79648 139946 79676
rect 140010 79676 140038 80036
rect 140102 79937 140130 80036
rect 140194 79966 140222 80036
rect 140182 79960 140234 79966
rect 140088 79928 140144 79937
rect 140182 79902 140234 79908
rect 140088 79863 140144 79872
rect 140102 79778 140130 79863
rect 140102 79750 140176 79778
rect 140010 79648 140084 79676
rect 139676 79620 139728 79626
rect 139676 79562 139728 79568
rect 139584 79552 139636 79558
rect 139584 79494 139636 79500
rect 139596 79354 139624 79494
rect 139584 79348 139636 79354
rect 139584 79290 139636 79296
rect 139582 78976 139638 78985
rect 139582 78911 139638 78920
rect 139596 76294 139624 78911
rect 139584 76288 139636 76294
rect 139584 76230 139636 76236
rect 139492 75812 139544 75818
rect 139492 75754 139544 75760
rect 139308 72956 139360 72962
rect 139308 72898 139360 72904
rect 139688 70394 139716 79562
rect 138768 70366 139256 70394
rect 139596 70366 139716 70394
rect 138664 68876 138716 68882
rect 138664 68818 138716 68824
rect 138480 64796 138532 64802
rect 138480 64738 138532 64744
rect 138768 55962 138796 70366
rect 139596 70242 139624 70366
rect 139584 70236 139636 70242
rect 139584 70178 139636 70184
rect 139400 62348 139452 62354
rect 139400 62290 139452 62296
rect 138756 55956 138808 55962
rect 138756 55898 138808 55904
rect 138664 53848 138716 53854
rect 138664 53790 138716 53796
rect 138296 39364 138348 39370
rect 138296 39306 138348 39312
rect 138020 6180 138072 6186
rect 138020 6122 138072 6128
rect 137284 3664 137336 3670
rect 137284 3606 137336 3612
rect 138676 3534 138704 53790
rect 139412 16574 139440 62290
rect 139780 53174 139808 79630
rect 139872 78198 139900 79648
rect 139952 79348 140004 79354
rect 139952 79290 140004 79296
rect 139860 78192 139912 78198
rect 139860 78134 139912 78140
rect 139964 70394 139992 79290
rect 140056 77897 140084 79648
rect 140148 79234 140176 79750
rect 140286 79744 140314 80036
rect 140378 79937 140406 80036
rect 140364 79928 140420 79937
rect 140470 79898 140498 80036
rect 140364 79863 140420 79872
rect 140458 79892 140510 79898
rect 140458 79834 140510 79840
rect 140240 79716 140314 79744
rect 140410 79792 140466 79801
rect 140562 79744 140590 80036
rect 140654 79937 140682 80036
rect 140746 79966 140774 80036
rect 140838 79966 140866 80036
rect 140930 79966 140958 80036
rect 140734 79960 140786 79966
rect 140640 79928 140696 79937
rect 140734 79902 140786 79908
rect 140826 79960 140878 79966
rect 140826 79902 140878 79908
rect 140918 79960 140970 79966
rect 140918 79902 140970 79908
rect 140640 79863 140696 79872
rect 141022 79812 141050 80036
rect 140700 79801 141050 79812
rect 140410 79727 140466 79736
rect 140240 79354 140268 79716
rect 140228 79348 140280 79354
rect 140228 79290 140280 79296
rect 140148 79206 140360 79234
rect 140136 78328 140188 78334
rect 140136 78270 140188 78276
rect 140042 77888 140098 77897
rect 140042 77823 140098 77832
rect 140044 77716 140096 77722
rect 140044 77658 140096 77664
rect 140056 77489 140084 77658
rect 140042 77480 140098 77489
rect 140042 77415 140098 77424
rect 139872 70366 139992 70394
rect 139872 64870 139900 70366
rect 139860 64864 139912 64870
rect 139860 64806 139912 64812
rect 140044 63572 140096 63578
rect 140044 63514 140096 63520
rect 139768 53168 139820 53174
rect 139768 53110 139820 53116
rect 139412 16546 139624 16574
rect 138848 4888 138900 4894
rect 138848 4830 138900 4836
rect 137652 3528 137704 3534
rect 137652 3470 137704 3476
rect 138664 3528 138716 3534
rect 138664 3470 138716 3476
rect 136456 3256 136508 3262
rect 136456 3198 136508 3204
rect 136468 480 136496 3198
rect 137664 480 137692 3470
rect 138860 480 138888 4830
rect 134126 354 134238 480
rect 133892 326 134238 354
rect 134126 -960 134238 326
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 139596 354 139624 16546
rect 140056 3262 140084 63514
rect 140148 55214 140176 78270
rect 140228 78192 140280 78198
rect 140228 78134 140280 78140
rect 140240 75342 140268 78134
rect 140228 75336 140280 75342
rect 140228 75278 140280 75284
rect 140332 73914 140360 79206
rect 140320 73908 140372 73914
rect 140320 73850 140372 73856
rect 140136 55208 140188 55214
rect 140136 55150 140188 55156
rect 140424 36582 140452 79727
rect 140516 79716 140590 79744
rect 140686 79792 141050 79801
rect 140742 79784 141050 79792
rect 141114 79744 141142 80036
rect 141206 79937 141234 80036
rect 141192 79928 141248 79937
rect 141192 79863 141194 79872
rect 141246 79863 141248 79872
rect 141194 79834 141246 79840
rect 141206 79803 141234 79834
rect 141298 79744 141326 80036
rect 140686 79727 140742 79736
rect 141068 79716 141142 79744
rect 141252 79716 141326 79744
rect 140516 78334 140544 79716
rect 140872 79688 140924 79694
rect 140872 79630 140924 79636
rect 140964 79688 141016 79694
rect 140964 79630 141016 79636
rect 140596 79620 140648 79626
rect 140596 79562 140648 79568
rect 140504 78328 140556 78334
rect 140504 78270 140556 78276
rect 140502 77752 140558 77761
rect 140502 77687 140558 77696
rect 140516 77314 140544 77687
rect 140504 77308 140556 77314
rect 140504 77250 140556 77256
rect 140608 72894 140636 79562
rect 140780 77444 140832 77450
rect 140780 77386 140832 77392
rect 140596 72888 140648 72894
rect 140596 72830 140648 72836
rect 140792 72622 140820 77386
rect 140884 76809 140912 79630
rect 140870 76800 140926 76809
rect 140870 76735 140926 76744
rect 140780 72616 140832 72622
rect 140780 72558 140832 72564
rect 140780 68876 140832 68882
rect 140780 68818 140832 68824
rect 140412 36576 140464 36582
rect 140412 36518 140464 36524
rect 140792 16574 140820 68818
rect 140976 68338 141004 79630
rect 141068 76430 141096 79716
rect 141148 79620 141200 79626
rect 141148 79562 141200 79568
rect 141160 78985 141188 79562
rect 141252 79354 141280 79716
rect 141390 79676 141418 80036
rect 141482 79830 141510 80036
rect 141470 79824 141522 79830
rect 141470 79766 141522 79772
rect 141574 79744 141602 80036
rect 141666 79812 141694 80036
rect 141758 79937 141786 80036
rect 141850 79966 141878 80036
rect 141942 79966 141970 80036
rect 141838 79960 141890 79966
rect 141744 79928 141800 79937
rect 141838 79902 141890 79908
rect 141930 79960 141982 79966
rect 141930 79902 141982 79908
rect 142034 79898 142062 80036
rect 142126 79966 142154 80036
rect 142114 79960 142166 79966
rect 142114 79902 142166 79908
rect 142218 79898 142246 80036
rect 142310 79966 142338 80036
rect 142402 79966 142430 80036
rect 142298 79960 142350 79966
rect 142298 79902 142350 79908
rect 142390 79960 142442 79966
rect 142390 79902 142442 79908
rect 141744 79863 141800 79872
rect 142022 79892 142074 79898
rect 142022 79834 142074 79840
rect 142206 79892 142258 79898
rect 142206 79834 142258 79840
rect 141838 79824 141890 79830
rect 141666 79784 141740 79812
rect 141574 79716 141648 79744
rect 141344 79648 141418 79676
rect 141240 79348 141292 79354
rect 141240 79290 141292 79296
rect 141146 78976 141202 78985
rect 141146 78911 141202 78920
rect 141056 76424 141108 76430
rect 141056 76366 141108 76372
rect 141160 68406 141188 78911
rect 141240 78668 141292 78674
rect 141240 78610 141292 78616
rect 141252 78577 141280 78610
rect 141238 78568 141294 78577
rect 141238 78503 141294 78512
rect 141252 77450 141280 78503
rect 141344 77897 141372 79648
rect 141516 79620 141568 79626
rect 141516 79562 141568 79568
rect 141424 79348 141476 79354
rect 141424 79290 141476 79296
rect 141330 77888 141386 77897
rect 141330 77823 141386 77832
rect 141240 77444 141292 77450
rect 141240 77386 141292 77392
rect 141436 75206 141464 79290
rect 141528 78674 141556 79562
rect 141516 78668 141568 78674
rect 141516 78610 141568 78616
rect 141516 78532 141568 78538
rect 141516 78474 141568 78480
rect 141528 75449 141556 78474
rect 141620 76498 141648 79716
rect 141712 78538 141740 79784
rect 141838 79766 141890 79772
rect 141930 79824 141982 79830
rect 142114 79824 142166 79830
rect 141982 79772 142016 79778
rect 141930 79766 142016 79772
rect 141850 79676 141878 79766
rect 141942 79750 142016 79766
rect 141804 79648 141878 79676
rect 141700 78532 141752 78538
rect 141700 78474 141752 78480
rect 141698 78432 141754 78441
rect 141698 78367 141754 78376
rect 141608 76492 141660 76498
rect 141608 76434 141660 76440
rect 141514 75440 141570 75449
rect 141514 75375 141570 75384
rect 141424 75200 141476 75206
rect 141424 75142 141476 75148
rect 141424 71528 141476 71534
rect 141424 71470 141476 71476
rect 141148 68400 141200 68406
rect 141148 68342 141200 68348
rect 140964 68332 141016 68338
rect 140964 68274 141016 68280
rect 140792 16546 141280 16574
rect 140044 3256 140096 3262
rect 140044 3198 140096 3204
rect 141252 480 141280 16546
rect 141436 3330 141464 71470
rect 141712 70394 141740 78367
rect 141804 76226 141832 79648
rect 141988 78690 142016 79750
rect 142080 79772 142114 79778
rect 142298 79824 142350 79830
rect 142080 79766 142166 79772
rect 142264 79772 142298 79778
rect 142264 79766 142350 79772
rect 142080 79750 142154 79766
rect 142264 79750 142338 79766
rect 142080 78742 142108 79750
rect 142160 79688 142212 79694
rect 142160 79630 142212 79636
rect 142172 78878 142200 79630
rect 142160 78872 142212 78878
rect 142160 78814 142212 78820
rect 141896 78662 142016 78690
rect 142068 78736 142120 78742
rect 142068 78678 142120 78684
rect 141896 76673 141924 78662
rect 141976 78600 142028 78606
rect 141976 78542 142028 78548
rect 141988 77858 142016 78542
rect 141976 77852 142028 77858
rect 141976 77794 142028 77800
rect 142264 77586 142292 79750
rect 142344 79688 142396 79694
rect 142494 79676 142522 80036
rect 142586 79971 142614 80036
rect 142572 79962 142628 79971
rect 142572 79897 142628 79906
rect 142678 79898 142706 80036
rect 142770 79966 142798 80036
rect 142862 79971 142890 80036
rect 142758 79960 142810 79966
rect 142758 79902 142810 79908
rect 142848 79962 142904 79971
rect 142666 79892 142718 79898
rect 142848 79897 142904 79906
rect 142954 79898 142982 80036
rect 143046 79971 143074 80036
rect 143032 79962 143088 79971
rect 142666 79834 142718 79840
rect 142942 79892 142994 79898
rect 143032 79897 143088 79906
rect 143138 79898 143166 80036
rect 142942 79834 142994 79840
rect 143126 79892 143178 79898
rect 143126 79834 143178 79840
rect 142710 79792 142766 79801
rect 142710 79727 142766 79736
rect 142894 79792 142950 79801
rect 142894 79727 142950 79736
rect 143078 79792 143134 79801
rect 143230 79744 143258 80036
rect 143078 79727 143134 79736
rect 142620 79688 142672 79694
rect 142494 79648 142568 79676
rect 142344 79630 142396 79636
rect 142356 77761 142384 79630
rect 142434 78976 142490 78985
rect 142434 78911 142490 78920
rect 142448 78674 142476 78911
rect 142436 78668 142488 78674
rect 142436 78610 142488 78616
rect 142540 78520 142568 79648
rect 142620 79630 142672 79636
rect 142448 78492 142568 78520
rect 142448 78130 142476 78492
rect 142526 78432 142582 78441
rect 142632 78402 142660 79630
rect 142724 78606 142752 79727
rect 142804 79620 142856 79626
rect 142804 79562 142856 79568
rect 142712 78600 142764 78606
rect 142712 78542 142764 78548
rect 142526 78367 142582 78376
rect 142620 78396 142672 78402
rect 142436 78124 142488 78130
rect 142436 78066 142488 78072
rect 142342 77752 142398 77761
rect 142342 77687 142398 77696
rect 142252 77580 142304 77586
rect 142252 77522 142304 77528
rect 141882 76664 141938 76673
rect 141882 76599 141938 76608
rect 141792 76220 141844 76226
rect 141792 76162 141844 76168
rect 142436 71460 142488 71466
rect 142436 71402 142488 71408
rect 142160 71324 142212 71330
rect 142160 71266 142212 71272
rect 141620 70366 141740 70394
rect 141620 68474 141648 70366
rect 142172 68882 142200 71266
rect 142160 68876 142212 68882
rect 142160 68818 142212 68824
rect 142252 68808 142304 68814
rect 142252 68750 142304 68756
rect 141608 68468 141660 68474
rect 141608 68410 141660 68416
rect 142264 4894 142292 68750
rect 142344 68672 142396 68678
rect 142344 68614 142396 68620
rect 142356 45626 142384 68614
rect 142448 53854 142476 71402
rect 142436 53848 142488 53854
rect 142436 53790 142488 53796
rect 142344 45620 142396 45626
rect 142344 45562 142396 45568
rect 142540 6914 142568 78367
rect 142620 78338 142672 78344
rect 142712 77716 142764 77722
rect 142712 77658 142764 77664
rect 142724 68814 142752 77658
rect 142816 72826 142844 79562
rect 142804 72820 142856 72826
rect 142804 72762 142856 72768
rect 142816 71534 142844 72762
rect 142804 71528 142856 71534
rect 142804 71470 142856 71476
rect 142804 71392 142856 71398
rect 142804 71334 142856 71340
rect 142712 68808 142764 68814
rect 142712 68750 142764 68756
rect 142816 62354 142844 71334
rect 142908 68678 142936 79727
rect 142988 79688 143040 79694
rect 142988 79630 143040 79636
rect 143000 77466 143028 79630
rect 143092 77586 143120 79727
rect 143184 79716 143258 79744
rect 143322 79744 143350 80036
rect 143414 79971 143442 80036
rect 143400 79962 143456 79971
rect 143506 79966 143534 80036
rect 143598 79966 143626 80036
rect 143400 79897 143456 79906
rect 143494 79960 143546 79966
rect 143494 79902 143546 79908
rect 143586 79960 143638 79966
rect 143586 79902 143638 79908
rect 143690 79812 143718 80036
rect 143782 79966 143810 80036
rect 143770 79960 143822 79966
rect 143770 79902 143822 79908
rect 143874 79812 143902 80036
rect 143966 79937 143994 80036
rect 143952 79928 144008 79937
rect 143952 79863 144008 79872
rect 143644 79784 143718 79812
rect 143828 79784 143902 79812
rect 143644 79778 143672 79784
rect 143460 79750 143672 79778
rect 143322 79716 143396 79744
rect 143080 77580 143132 77586
rect 143080 77522 143132 77528
rect 143000 77438 143120 77466
rect 142988 77308 143040 77314
rect 142988 77250 143040 77256
rect 143000 71194 143028 77250
rect 143092 72758 143120 77438
rect 143184 74254 143212 79716
rect 143264 79620 143316 79626
rect 143264 79562 143316 79568
rect 143276 77722 143304 79562
rect 143264 77716 143316 77722
rect 143264 77658 143316 77664
rect 143264 77580 143316 77586
rect 143264 77522 143316 77528
rect 143172 74248 143224 74254
rect 143172 74190 143224 74196
rect 143080 72752 143132 72758
rect 143080 72694 143132 72700
rect 142988 71188 143040 71194
rect 142988 71130 143040 71136
rect 143092 70394 143120 72694
rect 143184 71398 143212 74190
rect 143276 71466 143304 77522
rect 143368 77330 143396 79716
rect 143460 78169 143488 79750
rect 143632 79552 143684 79558
rect 143632 79494 143684 79500
rect 143724 79552 143776 79558
rect 143724 79494 143776 79500
rect 143540 79484 143592 79490
rect 143540 79426 143592 79432
rect 143552 79354 143580 79426
rect 143540 79348 143592 79354
rect 143540 79290 143592 79296
rect 143538 78704 143594 78713
rect 143538 78639 143594 78648
rect 143446 78160 143502 78169
rect 143446 78095 143502 78104
rect 143460 77586 143488 78095
rect 143448 77580 143500 77586
rect 143448 77522 143500 77528
rect 143368 77302 143488 77330
rect 143356 76220 143408 76226
rect 143356 76162 143408 76168
rect 143264 71460 143316 71466
rect 143264 71402 143316 71408
rect 143172 71392 143224 71398
rect 143172 71334 143224 71340
rect 143000 70366 143120 70394
rect 142896 68672 142948 68678
rect 142896 68614 142948 68620
rect 143000 63578 143028 70366
rect 143368 68513 143396 76162
rect 143460 71330 143488 77302
rect 143448 71324 143500 71330
rect 143448 71266 143500 71272
rect 143448 71188 143500 71194
rect 143448 71130 143500 71136
rect 143354 68504 143410 68513
rect 143354 68439 143410 68448
rect 142988 63572 143040 63578
rect 142988 63514 143040 63520
rect 142804 62348 142856 62354
rect 142804 62290 142856 62296
rect 142448 6886 142568 6914
rect 142252 4888 142304 4894
rect 142252 4830 142304 4836
rect 141424 3324 141476 3330
rect 141424 3266 141476 3272
rect 142448 480 142476 6886
rect 143460 3534 143488 71130
rect 143552 6186 143580 78639
rect 143644 77314 143672 79494
rect 143736 77314 143764 79494
rect 143828 78577 143856 79784
rect 144058 79744 144086 80036
rect 144150 79898 144178 80036
rect 144138 79892 144190 79898
rect 144138 79834 144190 79840
rect 144242 79812 144270 80036
rect 144334 79966 144362 80036
rect 144322 79960 144374 79966
rect 144322 79902 144374 79908
rect 144242 79784 144316 79812
rect 144288 79744 144316 79784
rect 144426 79744 144454 80036
rect 144012 79716 144086 79744
rect 144196 79716 144316 79744
rect 144380 79716 144454 79744
rect 143908 79416 143960 79422
rect 143908 79358 143960 79364
rect 143920 78674 143948 79358
rect 143908 78668 143960 78674
rect 143908 78610 143960 78616
rect 143814 78568 143870 78577
rect 143814 78503 143870 78512
rect 143632 77308 143684 77314
rect 143632 77250 143684 77256
rect 143724 77308 143776 77314
rect 143724 77250 143776 77256
rect 143828 67634 143856 78503
rect 143908 77308 143960 77314
rect 143908 77250 143960 77256
rect 143920 74526 143948 77250
rect 143908 74520 143960 74526
rect 143908 74462 143960 74468
rect 143906 74352 143962 74361
rect 143906 74287 143962 74296
rect 143920 73098 143948 74287
rect 144012 74050 144040 79716
rect 144092 79620 144144 79626
rect 144092 79562 144144 79568
rect 144104 78985 144132 79562
rect 144196 79354 144224 79716
rect 144276 79620 144328 79626
rect 144276 79562 144328 79568
rect 144184 79348 144236 79354
rect 144184 79290 144236 79296
rect 144090 78976 144146 78985
rect 144090 78911 144146 78920
rect 144000 74044 144052 74050
rect 144000 73986 144052 73992
rect 143908 73092 143960 73098
rect 143908 73034 143960 73040
rect 144012 69630 144040 73986
rect 144104 73982 144132 78911
rect 144196 78470 144224 79290
rect 144184 78464 144236 78470
rect 144184 78406 144236 78412
rect 144184 77580 144236 77586
rect 144184 77522 144236 77528
rect 144092 73976 144144 73982
rect 144092 73918 144144 73924
rect 144000 69624 144052 69630
rect 144000 69566 144052 69572
rect 143644 67606 143856 67634
rect 143644 53446 143672 67606
rect 143632 53440 143684 53446
rect 143632 53382 143684 53388
rect 144196 23526 144224 77522
rect 144288 74338 144316 79562
rect 144380 78713 144408 79716
rect 144518 79676 144546 80036
rect 144610 79966 144638 80036
rect 144702 79966 144730 80036
rect 144794 79966 144822 80036
rect 144598 79960 144650 79966
rect 144598 79902 144650 79908
rect 144690 79960 144742 79966
rect 144690 79902 144742 79908
rect 144782 79960 144834 79966
rect 144782 79902 144834 79908
rect 144886 79812 144914 80036
rect 144840 79801 144914 79812
rect 144826 79792 144914 79801
rect 144736 79756 144788 79762
rect 144882 79784 144914 79792
rect 144978 79744 145006 80036
rect 144826 79727 144882 79736
rect 144736 79698 144788 79704
rect 144932 79716 145006 79744
rect 144472 79648 144546 79676
rect 144366 78704 144422 78713
rect 144366 78639 144422 78648
rect 144472 74610 144500 79648
rect 144644 79620 144696 79626
rect 144644 79562 144696 79568
rect 144472 74582 144592 74610
rect 144460 74520 144512 74526
rect 144460 74462 144512 74468
rect 144288 74310 144408 74338
rect 144276 74044 144328 74050
rect 144276 73986 144328 73992
rect 144288 58682 144316 73986
rect 144380 72690 144408 74310
rect 144472 73778 144500 74462
rect 144460 73772 144512 73778
rect 144460 73714 144512 73720
rect 144368 72684 144420 72690
rect 144368 72626 144420 72632
rect 144380 63102 144408 72626
rect 144472 69018 144500 73714
rect 144460 69012 144512 69018
rect 144460 68954 144512 68960
rect 144564 68785 144592 74582
rect 144656 74458 144684 79562
rect 144748 76226 144776 79698
rect 144828 79688 144880 79694
rect 144828 79630 144880 79636
rect 144736 76220 144788 76226
rect 144736 76162 144788 76168
rect 144644 74452 144696 74458
rect 144644 74394 144696 74400
rect 144656 74050 144684 74394
rect 144644 74044 144696 74050
rect 144644 73986 144696 73992
rect 144840 70553 144868 79630
rect 144932 78810 144960 79716
rect 145070 79676 145098 80036
rect 145162 79898 145190 80036
rect 145150 79892 145202 79898
rect 145150 79834 145202 79840
rect 145254 79778 145282 80036
rect 145024 79648 145098 79676
rect 145208 79750 145282 79778
rect 145346 79778 145374 80036
rect 145438 79898 145466 80036
rect 145426 79892 145478 79898
rect 145426 79834 145478 79840
rect 145346 79750 145466 79778
rect 144920 78804 144972 78810
rect 144920 78746 144972 78752
rect 145024 77314 145052 79648
rect 145104 79552 145156 79558
rect 145104 79494 145156 79500
rect 145012 77308 145064 77314
rect 145012 77250 145064 77256
rect 145116 75886 145144 79494
rect 145104 75880 145156 75886
rect 145104 75822 145156 75828
rect 145208 73914 145236 79750
rect 145438 79642 145466 79750
rect 145530 79744 145558 80036
rect 145622 79898 145650 80036
rect 145714 79966 145742 80036
rect 145702 79960 145754 79966
rect 145702 79902 145754 79908
rect 145806 79898 145834 80036
rect 145898 79971 145926 80036
rect 145884 79962 145940 79971
rect 145610 79892 145662 79898
rect 145610 79834 145662 79840
rect 145794 79892 145846 79898
rect 145884 79897 145940 79906
rect 145794 79834 145846 79840
rect 145990 79830 146018 80036
rect 145978 79824 146030 79830
rect 145838 79792 145894 79801
rect 145530 79716 145604 79744
rect 145978 79766 146030 79772
rect 146082 79778 146110 80036
rect 146174 79898 146202 80036
rect 146266 79898 146294 80036
rect 146358 79966 146386 80036
rect 146450 79966 146478 80036
rect 146346 79960 146398 79966
rect 146346 79902 146398 79908
rect 146438 79960 146490 79966
rect 146438 79902 146490 79908
rect 146162 79892 146214 79898
rect 146162 79834 146214 79840
rect 146254 79892 146306 79898
rect 146254 79834 146306 79840
rect 146358 79812 146386 79902
rect 146358 79784 146432 79812
rect 146082 79750 146248 79778
rect 145838 79727 145894 79736
rect 146220 79744 146248 79750
rect 145300 79614 145466 79642
rect 145300 79257 145328 79614
rect 145380 79552 145432 79558
rect 145380 79494 145432 79500
rect 145286 79248 145342 79257
rect 145286 79183 145342 79192
rect 145196 73908 145248 73914
rect 145196 73850 145248 73856
rect 145208 73506 145236 73850
rect 145196 73500 145248 73506
rect 145196 73442 145248 73448
rect 144826 70544 144882 70553
rect 144826 70479 144882 70488
rect 145300 70394 145328 79183
rect 145392 77625 145420 79494
rect 145472 79484 145524 79490
rect 145472 79426 145524 79432
rect 145378 77616 145434 77625
rect 145378 77551 145434 77560
rect 145392 76090 145420 77551
rect 145380 76084 145432 76090
rect 145380 76026 145432 76032
rect 145484 75410 145512 79426
rect 145472 75404 145524 75410
rect 145472 75346 145524 75352
rect 145024 70366 145328 70394
rect 145484 70394 145512 75346
rect 145576 74526 145604 79716
rect 145656 79688 145708 79694
rect 145656 79630 145708 79636
rect 145748 79688 145800 79694
rect 145748 79630 145800 79636
rect 145668 75682 145696 79630
rect 145760 78305 145788 79630
rect 145852 79490 145880 79727
rect 146220 79716 146340 79744
rect 146024 79688 146076 79694
rect 146024 79630 146076 79636
rect 146116 79688 146168 79694
rect 146116 79630 146168 79636
rect 145840 79484 145892 79490
rect 145840 79426 145892 79432
rect 145746 78296 145802 78305
rect 145746 78231 145802 78240
rect 145656 75676 145708 75682
rect 145656 75618 145708 75624
rect 145668 74866 145696 75618
rect 145656 74860 145708 74866
rect 145656 74802 145708 74808
rect 145564 74520 145616 74526
rect 145564 74462 145616 74468
rect 145656 73500 145708 73506
rect 145656 73442 145708 73448
rect 145484 70366 145604 70394
rect 144550 68776 144606 68785
rect 144550 68711 144606 68720
rect 145024 64874 145052 70366
rect 144932 64846 145052 64874
rect 144368 63096 144420 63102
rect 144368 63038 144420 63044
rect 144276 58676 144328 58682
rect 144276 58618 144328 58624
rect 144932 46238 144960 64846
rect 144920 46232 144972 46238
rect 144920 46174 144972 46180
rect 145576 24138 145604 70366
rect 145668 35222 145696 73442
rect 145656 35216 145708 35222
rect 145656 35158 145708 35164
rect 145760 25566 145788 78231
rect 146036 76702 146064 79630
rect 146128 77761 146156 79630
rect 146208 79620 146260 79626
rect 146208 79562 146260 79568
rect 146220 79354 146248 79562
rect 146208 79348 146260 79354
rect 146208 79290 146260 79296
rect 146114 77752 146170 77761
rect 146114 77687 146170 77696
rect 146116 77308 146168 77314
rect 146116 77250 146168 77256
rect 146024 76696 146076 76702
rect 146024 76638 146076 76644
rect 146024 76084 146076 76090
rect 146024 76026 146076 76032
rect 145932 74860 145984 74866
rect 145932 74802 145984 74808
rect 145840 74520 145892 74526
rect 145840 74462 145892 74468
rect 145852 74118 145880 74462
rect 145840 74112 145892 74118
rect 145840 74054 145892 74060
rect 145852 51746 145880 74054
rect 145944 60042 145972 74802
rect 146036 67590 146064 76026
rect 146128 74322 146156 77250
rect 146312 76945 146340 79716
rect 146298 76936 146354 76945
rect 146298 76871 146354 76880
rect 146116 74316 146168 74322
rect 146116 74258 146168 74264
rect 146024 67584 146076 67590
rect 146024 67526 146076 67532
rect 146128 63578 146156 74258
rect 146404 69562 146432 79784
rect 146542 79744 146570 80036
rect 146634 79812 146662 80036
rect 146726 79966 146754 80036
rect 146818 79966 146846 80036
rect 146714 79960 146766 79966
rect 146712 79928 146714 79937
rect 146806 79960 146858 79966
rect 146766 79928 146768 79937
rect 146806 79902 146858 79908
rect 146712 79863 146768 79872
rect 146634 79784 146800 79812
rect 146910 79801 146938 80036
rect 146542 79716 146616 79744
rect 146484 79620 146536 79626
rect 146484 79562 146536 79568
rect 146496 75682 146524 79562
rect 146588 78334 146616 79716
rect 146668 79552 146720 79558
rect 146668 79494 146720 79500
rect 146576 78328 146628 78334
rect 146576 78270 146628 78276
rect 146680 75750 146708 79494
rect 146772 77926 146800 79784
rect 146896 79792 146952 79801
rect 146896 79727 146952 79736
rect 146910 79676 146938 79727
rect 146864 79648 146938 79676
rect 147002 79676 147030 80036
rect 147094 79812 147122 80036
rect 147186 79966 147214 80036
rect 147174 79960 147226 79966
rect 147174 79902 147226 79908
rect 147278 79898 147306 80036
rect 147266 79892 147318 79898
rect 147266 79834 147318 79840
rect 147094 79784 147168 79812
rect 147140 79744 147168 79784
rect 147370 79744 147398 80036
rect 147462 79801 147490 80036
rect 147554 79898 147582 80036
rect 147646 79971 147674 80036
rect 147632 79962 147688 79971
rect 147542 79892 147594 79898
rect 147632 79897 147688 79906
rect 147542 79834 147594 79840
rect 147738 79812 147766 80036
rect 147140 79716 147260 79744
rect 147002 79648 147076 79676
rect 146760 77920 146812 77926
rect 146760 77862 146812 77868
rect 146772 77518 146800 77862
rect 146760 77512 146812 77518
rect 146760 77454 146812 77460
rect 146668 75744 146720 75750
rect 146668 75686 146720 75692
rect 146484 75676 146536 75682
rect 146484 75618 146536 75624
rect 146496 75002 146524 75618
rect 146484 74996 146536 75002
rect 146484 74938 146536 74944
rect 146680 72826 146708 75686
rect 146668 72820 146720 72826
rect 146668 72762 146720 72768
rect 146864 70394 146892 79648
rect 146944 79552 146996 79558
rect 146942 79520 146944 79529
rect 146996 79520 146998 79529
rect 146942 79455 146998 79464
rect 146956 77790 146984 79455
rect 147048 79064 147076 79648
rect 147128 79620 147180 79626
rect 147128 79562 147180 79568
rect 147140 79529 147168 79562
rect 147126 79520 147182 79529
rect 147126 79455 147182 79464
rect 147048 79036 147168 79064
rect 146944 77784 146996 77790
rect 146944 77726 146996 77732
rect 146942 76936 146998 76945
rect 146942 76871 146998 76880
rect 146680 70366 146892 70394
rect 146392 69556 146444 69562
rect 146392 69498 146444 69504
rect 146300 69012 146352 69018
rect 146300 68954 146352 68960
rect 146116 63572 146168 63578
rect 146116 63514 146168 63520
rect 145932 60036 145984 60042
rect 145932 59978 145984 59984
rect 145840 51740 145892 51746
rect 145840 51682 145892 51688
rect 145748 25560 145800 25566
rect 145748 25502 145800 25508
rect 145564 24132 145616 24138
rect 145564 24074 145616 24080
rect 144184 23520 144236 23526
rect 144184 23462 144236 23468
rect 144920 23520 144972 23526
rect 144920 23462 144972 23468
rect 144932 16574 144960 23462
rect 146312 16574 146340 68954
rect 146680 64874 146708 70366
rect 146404 64846 146708 64874
rect 146404 58818 146432 64846
rect 146392 58812 146444 58818
rect 146392 58754 146444 58760
rect 144932 16546 145512 16574
rect 146312 16546 146892 16574
rect 143540 6180 143592 6186
rect 143540 6122 143592 6128
rect 143540 3732 143592 3738
rect 143540 3674 143592 3680
rect 143448 3528 143500 3534
rect 143448 3470 143500 3476
rect 143552 480 143580 3674
rect 144736 3528 144788 3534
rect 144736 3470 144788 3476
rect 144748 480 144776 3470
rect 140014 354 140126 480
rect 139596 326 140126 354
rect 140014 -960 140126 326
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145484 354 145512 16546
rect 146864 3482 146892 16546
rect 146956 4146 146984 76871
rect 147140 75478 147168 79036
rect 147128 75472 147180 75478
rect 147128 75414 147180 75420
rect 147232 75138 147260 79716
rect 147324 79716 147398 79744
rect 147448 79792 147504 79801
rect 147692 79784 147766 79812
rect 147692 79744 147720 79784
rect 147448 79727 147504 79736
rect 147600 79716 147720 79744
rect 147324 77897 147352 79716
rect 147496 79620 147548 79626
rect 147496 79562 147548 79568
rect 147404 79552 147456 79558
rect 147402 79520 147404 79529
rect 147456 79520 147458 79529
rect 147402 79455 147458 79464
rect 147508 79132 147536 79562
rect 147600 79286 147628 79716
rect 147830 79676 147858 80036
rect 147922 79898 147950 80036
rect 147910 79892 147962 79898
rect 147910 79834 147962 79840
rect 148014 79801 148042 80036
rect 148106 79898 148134 80036
rect 148094 79892 148146 79898
rect 148094 79834 148146 79840
rect 148000 79792 148056 79801
rect 148000 79727 148056 79736
rect 147692 79648 147858 79676
rect 147956 79688 148008 79694
rect 147692 79529 147720 79648
rect 148198 79676 148226 80036
rect 148290 79778 148318 80036
rect 148382 79966 148410 80036
rect 148474 79966 148502 80036
rect 148566 79966 148594 80036
rect 148370 79960 148422 79966
rect 148370 79902 148422 79908
rect 148462 79960 148514 79966
rect 148554 79960 148606 79966
rect 148462 79902 148514 79908
rect 148552 79928 148554 79937
rect 148606 79928 148608 79937
rect 148552 79863 148608 79872
rect 148566 79837 148594 79863
rect 148506 79792 148562 79801
rect 148290 79750 148364 79778
rect 148198 79648 148272 79676
rect 147956 79630 148008 79636
rect 147678 79520 147734 79529
rect 147678 79455 147734 79464
rect 147588 79280 147640 79286
rect 147588 79222 147640 79228
rect 147508 79104 147628 79132
rect 147310 77888 147366 77897
rect 147310 77823 147366 77832
rect 147404 77784 147456 77790
rect 147404 77726 147456 77732
rect 147312 77512 147364 77518
rect 147312 77454 147364 77460
rect 147220 75132 147272 75138
rect 147220 75074 147272 75080
rect 147036 73092 147088 73098
rect 147036 73034 147088 73040
rect 146944 4140 146996 4146
rect 146944 4082 146996 4088
rect 147048 3670 147076 73034
rect 147232 70394 147260 75074
rect 147140 70366 147260 70394
rect 147140 69766 147168 70366
rect 147128 69760 147180 69766
rect 147128 69702 147180 69708
rect 147128 69624 147180 69630
rect 147128 69566 147180 69572
rect 147140 3942 147168 69566
rect 147324 64190 147352 77454
rect 147312 64184 147364 64190
rect 147312 64126 147364 64132
rect 147220 63572 147272 63578
rect 147220 63514 147272 63520
rect 147128 3936 147180 3942
rect 147128 3878 147180 3884
rect 147232 3874 147260 63514
rect 147416 62830 147444 77726
rect 147404 62824 147456 62830
rect 147404 62766 147456 62772
rect 147312 60036 147364 60042
rect 147312 59978 147364 59984
rect 147220 3868 147272 3874
rect 147220 3810 147272 3816
rect 147036 3664 147088 3670
rect 147036 3606 147088 3612
rect 147324 3602 147352 59978
rect 147600 50454 147628 79104
rect 147692 75546 147720 79455
rect 147864 79280 147916 79286
rect 147864 79222 147916 79228
rect 147772 77648 147824 77654
rect 147772 77590 147824 77596
rect 147680 75540 147732 75546
rect 147680 75482 147732 75488
rect 147680 53440 147732 53446
rect 147680 53382 147732 53388
rect 147588 50448 147640 50454
rect 147588 50390 147640 50396
rect 147692 16574 147720 53382
rect 147784 36922 147812 77590
rect 147876 53242 147904 79222
rect 147968 78878 147996 79630
rect 148048 79552 148100 79558
rect 148140 79552 148192 79558
rect 148048 79494 148100 79500
rect 148138 79520 148140 79529
rect 148192 79520 148194 79529
rect 147956 78872 148008 78878
rect 147956 78814 148008 78820
rect 148060 75614 148088 79494
rect 148138 79455 148194 79464
rect 148140 78940 148192 78946
rect 148140 78882 148192 78888
rect 148152 78402 148180 78882
rect 148140 78396 148192 78402
rect 148140 78338 148192 78344
rect 148048 75608 148100 75614
rect 148048 75550 148100 75556
rect 147864 53236 147916 53242
rect 147864 53178 147916 53184
rect 148152 51814 148180 78338
rect 148244 77042 148272 79648
rect 148336 78266 148364 79750
rect 148506 79727 148562 79736
rect 148658 79744 148686 80036
rect 148750 79937 148778 80036
rect 148736 79928 148792 79937
rect 148736 79863 148792 79872
rect 148842 79744 148870 80036
rect 148934 79898 148962 80036
rect 148922 79892 148974 79898
rect 148922 79834 148974 79840
rect 149026 79830 149054 80036
rect 149014 79824 149066 79830
rect 149014 79766 149066 79772
rect 148416 79688 148468 79694
rect 148416 79630 148468 79636
rect 148324 78260 148376 78266
rect 148324 78202 148376 78208
rect 148336 77586 148364 78202
rect 148428 77994 148456 79630
rect 148416 77988 148468 77994
rect 148416 77930 148468 77936
rect 148324 77580 148376 77586
rect 148324 77522 148376 77528
rect 148232 77036 148284 77042
rect 148232 76978 148284 76984
rect 148244 69698 148272 76978
rect 148428 75914 148456 77930
rect 148520 77654 148548 79727
rect 148658 79716 148732 79744
rect 148842 79716 148916 79744
rect 148600 79620 148652 79626
rect 148600 79562 148652 79568
rect 148612 78033 148640 79562
rect 148704 78305 148732 79716
rect 148784 79620 148836 79626
rect 148784 79562 148836 79568
rect 148690 78296 148746 78305
rect 148690 78231 148746 78240
rect 148598 78024 148654 78033
rect 148598 77959 148600 77968
rect 148652 77959 148654 77968
rect 148600 77930 148652 77936
rect 148612 77899 148640 77930
rect 148690 77888 148746 77897
rect 148690 77823 148746 77832
rect 148508 77648 148560 77654
rect 148508 77590 148560 77596
rect 148600 77580 148652 77586
rect 148600 77522 148652 77528
rect 148428 75886 148548 75914
rect 148324 75880 148376 75886
rect 148324 75822 148376 75828
rect 148232 69692 148284 69698
rect 148232 69634 148284 69640
rect 148140 51808 148192 51814
rect 148140 51750 148192 51756
rect 147772 36916 147824 36922
rect 147772 36858 147824 36864
rect 147692 16546 147904 16574
rect 147404 4140 147456 4146
rect 147404 4082 147456 4088
rect 147312 3596 147364 3602
rect 147312 3538 147364 3544
rect 146864 3454 147168 3482
rect 147140 480 147168 3454
rect 147416 3330 147444 4082
rect 147404 3324 147456 3330
rect 147404 3266 147456 3272
rect 145902 354 146014 480
rect 145484 326 146014 354
rect 145902 -960 146014 326
rect 147098 -960 147210 480
rect 147876 354 147904 16546
rect 148336 3806 148364 75822
rect 148416 67584 148468 67590
rect 148416 67526 148468 67532
rect 148324 3800 148376 3806
rect 148324 3742 148376 3748
rect 148428 3738 148456 67526
rect 148520 32706 148548 75886
rect 148612 46306 148640 77522
rect 148704 49298 148732 77823
rect 148796 76974 148824 79562
rect 148888 78402 148916 79716
rect 148968 79688 149020 79694
rect 149118 79676 149146 80036
rect 149210 79778 149238 80036
rect 149302 79971 149330 80036
rect 149288 79962 149344 79971
rect 149288 79897 149344 79906
rect 149394 79898 149422 80036
rect 149486 79898 149514 80036
rect 149578 79898 149606 80036
rect 149382 79892 149434 79898
rect 149382 79834 149434 79840
rect 149474 79892 149526 79898
rect 149474 79834 149526 79840
rect 149566 79892 149618 79898
rect 149566 79834 149618 79840
rect 149334 79792 149390 79801
rect 149210 79750 149284 79778
rect 149118 79648 149192 79676
rect 148968 79630 149020 79636
rect 148876 78396 148928 78402
rect 148876 78338 148928 78344
rect 148876 77988 148928 77994
rect 148876 77930 148928 77936
rect 148784 76968 148836 76974
rect 148784 76910 148836 76916
rect 148796 65618 148824 76910
rect 148888 75410 148916 77930
rect 148980 77489 149008 79630
rect 149060 79144 149112 79150
rect 149060 79086 149112 79092
rect 148966 77480 149022 77489
rect 148966 77415 149022 77424
rect 148876 75404 148928 75410
rect 148876 75346 148928 75352
rect 148784 65612 148836 65618
rect 148784 65554 148836 65560
rect 148692 49292 148744 49298
rect 148692 49234 148744 49240
rect 148600 46300 148652 46306
rect 148600 46242 148652 46248
rect 149072 36854 149100 79086
rect 149164 73642 149192 79648
rect 149256 78849 149284 79750
rect 149670 79744 149698 80036
rect 149334 79727 149390 79736
rect 149242 78840 149298 78849
rect 149242 78775 149298 78784
rect 149152 73636 149204 73642
rect 149152 73578 149204 73584
rect 149256 64874 149284 78775
rect 149348 78266 149376 79727
rect 149624 79716 149698 79744
rect 149762 79744 149790 80036
rect 149854 79898 149882 80036
rect 149842 79892 149894 79898
rect 149842 79834 149894 79840
rect 149946 79744 149974 80036
rect 150038 79971 150066 80036
rect 150024 79962 150080 79971
rect 150024 79897 150080 79906
rect 150130 79898 150158 80036
rect 150118 79892 150170 79898
rect 150118 79834 150170 79840
rect 150222 79778 150250 80036
rect 150314 79937 150342 80036
rect 150300 79928 150356 79937
rect 150300 79863 150356 79872
rect 150222 79750 150296 79778
rect 149762 79716 149836 79744
rect 149946 79716 150112 79744
rect 149428 79688 149480 79694
rect 149480 79648 149560 79676
rect 149428 79630 149480 79636
rect 149428 79484 149480 79490
rect 149428 79426 149480 79432
rect 149336 78260 149388 78266
rect 149336 78202 149388 78208
rect 149440 75274 149468 79426
rect 149532 78742 149560 79648
rect 149624 79642 149652 79716
rect 149808 79642 149836 79716
rect 149624 79614 149744 79642
rect 149808 79614 150020 79642
rect 149612 79552 149664 79558
rect 149612 79494 149664 79500
rect 149520 78736 149572 78742
rect 149520 78678 149572 78684
rect 149624 78305 149652 79494
rect 149716 79150 149744 79614
rect 149796 79552 149848 79558
rect 149796 79494 149848 79500
rect 149704 79144 149756 79150
rect 149704 79086 149756 79092
rect 149610 78296 149666 78305
rect 149610 78231 149666 78240
rect 149808 76362 149836 79494
rect 149888 79280 149940 79286
rect 149888 79222 149940 79228
rect 149900 77761 149928 79222
rect 149886 77752 149942 77761
rect 149886 77687 149942 77696
rect 149796 76356 149848 76362
rect 149796 76298 149848 76304
rect 149428 75268 149480 75274
rect 149428 75210 149480 75216
rect 149704 73976 149756 73982
rect 149704 73918 149756 73924
rect 149164 64846 149284 64874
rect 149164 43654 149192 64846
rect 149152 43648 149204 43654
rect 149152 43590 149204 43596
rect 149060 36848 149112 36854
rect 149060 36790 149112 36796
rect 148508 32700 148560 32706
rect 148508 32642 148560 32648
rect 149716 4146 149744 73918
rect 149808 64326 149836 76298
rect 149992 74254 150020 79614
rect 150084 78674 150112 79716
rect 150164 79688 150216 79694
rect 150164 79630 150216 79636
rect 150176 79132 150204 79630
rect 150268 79234 150296 79750
rect 150406 79676 150434 80036
rect 150498 79744 150526 80036
rect 150590 79898 150618 80036
rect 150682 79966 150710 80036
rect 150774 79966 150802 80036
rect 150866 79971 150894 80036
rect 150670 79960 150722 79966
rect 150670 79902 150722 79908
rect 150762 79960 150814 79966
rect 150762 79902 150814 79908
rect 150852 79962 150908 79971
rect 150578 79892 150630 79898
rect 150852 79897 150908 79906
rect 150578 79834 150630 79840
rect 150716 79824 150768 79830
rect 150716 79766 150768 79772
rect 150624 79756 150676 79762
rect 150498 79716 150572 79744
rect 150360 79648 150434 79676
rect 150360 79422 150388 79648
rect 150544 79558 150572 79716
rect 150624 79698 150676 79704
rect 150532 79552 150584 79558
rect 150532 79494 150584 79500
rect 150348 79416 150400 79422
rect 150348 79358 150400 79364
rect 150268 79206 150480 79234
rect 150176 79121 150296 79132
rect 150162 79112 150296 79121
rect 150218 79104 150296 79112
rect 150162 79047 150218 79056
rect 150164 78736 150216 78742
rect 150164 78678 150216 78684
rect 150072 78668 150124 78674
rect 150072 78610 150124 78616
rect 150084 76566 150112 78610
rect 150176 78062 150204 78678
rect 150164 78056 150216 78062
rect 150164 77998 150216 78004
rect 150072 76560 150124 76566
rect 150072 76502 150124 76508
rect 150072 75268 150124 75274
rect 150072 75210 150124 75216
rect 149980 74248 150032 74254
rect 149980 74190 150032 74196
rect 149980 73636 150032 73642
rect 149980 73578 150032 73584
rect 149796 64320 149848 64326
rect 149796 64262 149848 64268
rect 149796 63096 149848 63102
rect 149796 63038 149848 63044
rect 149704 4140 149756 4146
rect 149704 4082 149756 4088
rect 148416 3732 148468 3738
rect 148416 3674 148468 3680
rect 149520 3664 149572 3670
rect 149520 3606 149572 3612
rect 149532 480 149560 3606
rect 149808 2922 149836 63038
rect 149992 57458 150020 73578
rect 149980 57452 150032 57458
rect 149980 57394 150032 57400
rect 150084 49094 150112 75210
rect 150072 49088 150124 49094
rect 150072 49030 150124 49036
rect 150176 23050 150204 77998
rect 150268 62898 150296 79104
rect 150346 78976 150402 78985
rect 150346 78911 150402 78920
rect 150256 62892 150308 62898
rect 150256 62834 150308 62840
rect 150164 23044 150216 23050
rect 150164 22986 150216 22992
rect 150360 7886 150388 78911
rect 150452 77897 150480 79206
rect 150438 77888 150494 77897
rect 150438 77823 150494 77832
rect 150544 42362 150572 79494
rect 150636 69018 150664 79698
rect 150728 79393 150756 79766
rect 150958 79744 150986 80036
rect 151050 79966 151078 80036
rect 151142 79971 151170 80036
rect 151038 79960 151090 79966
rect 151038 79902 151090 79908
rect 151128 79962 151184 79971
rect 151128 79897 151184 79906
rect 151084 79824 151136 79830
rect 151084 79766 151136 79772
rect 151234 79778 151262 80036
rect 151326 79966 151354 80036
rect 151418 79971 151446 80036
rect 151314 79960 151366 79966
rect 151314 79902 151366 79908
rect 151404 79962 151460 79971
rect 151404 79897 151460 79906
rect 150958 79716 151032 79744
rect 150714 79384 150770 79393
rect 150714 79319 150770 79328
rect 150728 76634 150756 79319
rect 150806 79112 150862 79121
rect 151004 79082 151032 79716
rect 151096 79150 151124 79766
rect 151234 79750 151308 79778
rect 151176 79688 151228 79694
rect 151176 79630 151228 79636
rect 151084 79144 151136 79150
rect 151084 79086 151136 79092
rect 150806 79047 150862 79056
rect 150992 79076 151044 79082
rect 150716 76628 150768 76634
rect 150716 76570 150768 76576
rect 150624 69012 150676 69018
rect 150624 68954 150676 68960
rect 150636 68882 150664 68954
rect 150624 68876 150676 68882
rect 150624 68818 150676 68824
rect 150532 42356 150584 42362
rect 150532 42298 150584 42304
rect 150820 9246 150848 79047
rect 150992 79018 151044 79024
rect 151096 76906 151124 79086
rect 151084 76900 151136 76906
rect 151084 76842 151136 76848
rect 151084 76696 151136 76702
rect 151084 76638 151136 76644
rect 150900 76628 150952 76634
rect 150900 76570 150952 76576
rect 150912 32638 150940 76570
rect 150900 32632 150952 32638
rect 150900 32574 150952 32580
rect 150808 9240 150860 9246
rect 150808 9182 150860 9188
rect 150348 7880 150400 7886
rect 150348 7822 150400 7828
rect 150624 3936 150676 3942
rect 150624 3878 150676 3884
rect 149796 2916 149848 2922
rect 149796 2858 149848 2864
rect 150636 480 150664 3878
rect 151096 3534 151124 76638
rect 151188 71670 151216 79630
rect 151280 78713 151308 79750
rect 151418 79676 151446 79897
rect 151510 79812 151538 80036
rect 151602 79966 151630 80036
rect 151590 79960 151642 79966
rect 151694 79937 151722 80036
rect 151590 79902 151642 79908
rect 151680 79928 151736 79937
rect 151680 79863 151736 79872
rect 151694 79812 151722 79863
rect 151510 79801 151584 79812
rect 151510 79792 151598 79801
rect 151510 79784 151542 79792
rect 151542 79727 151598 79736
rect 151648 79784 151722 79812
rect 151418 79648 151492 79676
rect 151358 79112 151414 79121
rect 151358 79047 151414 79056
rect 151266 78704 151322 78713
rect 151266 78639 151322 78648
rect 151268 77240 151320 77246
rect 151268 77182 151320 77188
rect 151280 76770 151308 77182
rect 151268 76764 151320 76770
rect 151268 76706 151320 76712
rect 151176 71664 151228 71670
rect 151176 71606 151228 71612
rect 151188 70394 151216 71606
rect 151372 70394 151400 79047
rect 151464 77194 151492 79648
rect 151544 79552 151596 79558
rect 151544 79494 151596 79500
rect 151556 79014 151584 79494
rect 151544 79008 151596 79014
rect 151544 78950 151596 78956
rect 151648 77294 151676 79784
rect 151786 79744 151814 80036
rect 151878 79778 151906 80036
rect 151970 79898 151998 80036
rect 151958 79892 152010 79898
rect 151958 79834 152010 79840
rect 152062 79801 152090 80036
rect 152154 79966 152182 80036
rect 152142 79960 152194 79966
rect 152246 79937 152274 80036
rect 152142 79902 152194 79908
rect 152232 79928 152288 79937
rect 152232 79863 152234 79872
rect 152286 79863 152288 79872
rect 152234 79834 152286 79840
rect 152048 79792 152104 79801
rect 151878 79750 151952 79778
rect 151740 79716 151814 79744
rect 151740 78577 151768 79716
rect 151820 79620 151872 79626
rect 151820 79562 151872 79568
rect 151726 78568 151782 78577
rect 151726 78503 151782 78512
rect 151832 77314 151860 79562
rect 151820 77308 151872 77314
rect 151648 77266 151768 77294
rect 151464 77166 151676 77194
rect 151188 70366 151308 70394
rect 151372 70366 151584 70394
rect 151176 69012 151228 69018
rect 151176 68954 151228 68960
rect 151188 17542 151216 68954
rect 151280 29918 151308 70366
rect 151556 53174 151584 70366
rect 151544 53168 151596 53174
rect 151544 53110 151596 53116
rect 151268 29912 151320 29918
rect 151268 29854 151320 29860
rect 151176 17536 151228 17542
rect 151176 17478 151228 17484
rect 151648 10606 151676 77166
rect 151740 73846 151768 77266
rect 151820 77250 151872 77256
rect 151728 73840 151780 73846
rect 151728 73782 151780 73788
rect 151924 71738 151952 79750
rect 152338 79778 152366 80036
rect 152430 79966 152458 80036
rect 152418 79960 152470 79966
rect 152418 79902 152470 79908
rect 152522 79830 152550 80036
rect 152048 79727 152104 79736
rect 152188 79756 152240 79762
rect 152188 79698 152240 79704
rect 152292 79750 152366 79778
rect 152510 79824 152562 79830
rect 152510 79766 152562 79772
rect 152004 79688 152056 79694
rect 152004 79630 152056 79636
rect 152094 79656 152150 79665
rect 152016 78130 152044 79630
rect 152094 79591 152150 79600
rect 152108 79490 152136 79591
rect 152096 79484 152148 79490
rect 152096 79426 152148 79432
rect 152004 78124 152056 78130
rect 152004 78066 152056 78072
rect 151912 71732 151964 71738
rect 151912 71674 151964 71680
rect 152108 71618 152136 79426
rect 151924 71590 152136 71618
rect 151924 60178 151952 71590
rect 152200 70394 152228 79698
rect 152292 73166 152320 79750
rect 152614 79744 152642 80036
rect 152706 79966 152734 80036
rect 152798 79966 152826 80036
rect 152890 79966 152918 80036
rect 152694 79960 152746 79966
rect 152786 79960 152838 79966
rect 152694 79902 152746 79908
rect 152784 79928 152786 79937
rect 152878 79960 152930 79966
rect 152838 79928 152840 79937
rect 152982 79937 153010 80036
rect 152878 79902 152930 79908
rect 152968 79928 153024 79937
rect 152784 79863 152840 79872
rect 152968 79863 153024 79872
rect 153074 79830 153102 80036
rect 153166 79898 153194 80036
rect 153258 79966 153286 80036
rect 153246 79960 153298 79966
rect 153246 79902 153298 79908
rect 153154 79892 153206 79898
rect 153154 79834 153206 79840
rect 152924 79824 152976 79830
rect 152924 79766 152976 79772
rect 153062 79824 153114 79830
rect 153350 79812 153378 80036
rect 153442 79966 153470 80036
rect 153430 79960 153482 79966
rect 153430 79902 153482 79908
rect 153350 79784 153424 79812
rect 153062 79766 153114 79772
rect 152614 79716 152688 79744
rect 152464 79688 152516 79694
rect 152464 79630 152516 79636
rect 152372 78464 152424 78470
rect 152372 78406 152424 78412
rect 152280 73160 152332 73166
rect 152280 73102 152332 73108
rect 152292 72146 152320 73102
rect 152280 72140 152332 72146
rect 152280 72082 152332 72088
rect 152016 70366 152228 70394
rect 151912 60172 151964 60178
rect 151912 60114 151964 60120
rect 152016 57390 152044 70366
rect 152004 57384 152056 57390
rect 152004 57326 152056 57332
rect 151636 10600 151688 10606
rect 151636 10542 151688 10548
rect 152384 6914 152412 78406
rect 152476 71602 152504 79630
rect 152556 78124 152608 78130
rect 152556 78066 152608 78072
rect 152464 71596 152516 71602
rect 152464 71538 152516 71544
rect 152476 13326 152504 71538
rect 152568 68950 152596 78066
rect 152660 73817 152688 79716
rect 152832 79688 152884 79694
rect 152752 79648 152832 79676
rect 152752 74186 152780 79648
rect 152832 79630 152884 79636
rect 152832 79552 152884 79558
rect 152832 79494 152884 79500
rect 152844 79393 152872 79494
rect 152830 79384 152886 79393
rect 152830 79319 152886 79328
rect 152740 74180 152792 74186
rect 152740 74122 152792 74128
rect 152646 73808 152702 73817
rect 152646 73743 152702 73752
rect 152740 72140 152792 72146
rect 152740 72082 152792 72088
rect 152648 71732 152700 71738
rect 152648 71674 152700 71680
rect 152556 68944 152608 68950
rect 152556 68886 152608 68892
rect 152464 13320 152516 13326
rect 152464 13262 152516 13268
rect 152568 11966 152596 68886
rect 152660 39642 152688 71674
rect 152752 47734 152780 72082
rect 152740 47728 152792 47734
rect 152740 47670 152792 47676
rect 152648 39636 152700 39642
rect 152648 39578 152700 39584
rect 152844 16114 152872 79319
rect 152936 73545 152964 79766
rect 153200 79756 153252 79762
rect 153200 79698 153252 79704
rect 153016 79688 153068 79694
rect 153014 79656 153016 79665
rect 153068 79656 153070 79665
rect 153014 79591 153070 79600
rect 152922 73536 152978 73545
rect 152922 73471 152978 73480
rect 153028 18902 153056 79591
rect 153108 79008 153160 79014
rect 153108 78950 153160 78956
rect 153120 76702 153148 78950
rect 153212 77602 153240 79698
rect 153396 79540 153424 79784
rect 153534 79778 153562 80036
rect 153626 79937 153654 80036
rect 153612 79928 153668 79937
rect 153612 79863 153668 79872
rect 153488 79750 153562 79778
rect 153488 79608 153516 79750
rect 153718 79744 153746 80036
rect 153810 79966 153838 80036
rect 153798 79960 153850 79966
rect 153902 79937 153930 80036
rect 153798 79902 153850 79908
rect 153888 79928 153944 79937
rect 153888 79863 153944 79872
rect 153994 79812 154022 80036
rect 154086 79966 154114 80036
rect 154178 79966 154206 80036
rect 154074 79960 154126 79966
rect 154074 79902 154126 79908
rect 154166 79960 154218 79966
rect 154166 79902 154218 79908
rect 154270 79898 154298 80036
rect 154362 79971 154390 80036
rect 154348 79962 154404 79971
rect 154454 79966 154482 80036
rect 154258 79892 154310 79898
rect 154348 79897 154404 79906
rect 154442 79960 154494 79966
rect 154442 79902 154494 79908
rect 154546 79898 154574 80036
rect 154638 79898 154666 80036
rect 154730 79966 154758 80036
rect 154822 79966 154850 80036
rect 154914 79966 154942 80036
rect 154718 79960 154770 79966
rect 154718 79902 154770 79908
rect 154810 79960 154862 79966
rect 154810 79902 154862 79908
rect 154902 79960 154954 79966
rect 155006 79937 155034 80036
rect 154902 79902 154954 79908
rect 154992 79928 155048 79937
rect 154258 79834 154310 79840
rect 154534 79892 154586 79898
rect 154534 79834 154586 79840
rect 154626 79892 154678 79898
rect 154992 79863 155048 79872
rect 154626 79834 154678 79840
rect 155098 79830 155126 80036
rect 153948 79784 154022 79812
rect 154764 79824 154816 79830
rect 154118 79792 154174 79801
rect 153718 79716 153792 79744
rect 153488 79580 153608 79608
rect 153396 79512 153516 79540
rect 153212 77574 153424 77602
rect 153290 77480 153346 77489
rect 153290 77415 153346 77424
rect 153108 76696 153160 76702
rect 153108 76638 153160 76644
rect 153200 73772 153252 73778
rect 153200 73714 153252 73720
rect 153212 27198 153240 73714
rect 153304 35494 153332 77415
rect 153396 74390 153424 77574
rect 153488 77178 153516 79512
rect 153476 77172 153528 77178
rect 153476 77114 153528 77120
rect 153384 74384 153436 74390
rect 153384 74326 153436 74332
rect 153488 73914 153516 77114
rect 153476 73908 153528 73914
rect 153476 73850 153528 73856
rect 153580 71641 153608 79580
rect 153658 79520 153714 79529
rect 153658 79455 153714 79464
rect 153672 79354 153700 79455
rect 153660 79348 153712 79354
rect 153660 79290 153712 79296
rect 153566 71632 153622 71641
rect 153566 71567 153622 71576
rect 153580 67634 153608 71567
rect 153764 69426 153792 79716
rect 153948 79694 153976 79784
rect 154764 79766 154816 79772
rect 155086 79824 155138 79830
rect 155086 79766 155138 79772
rect 155190 79778 155218 80036
rect 155282 79966 155310 80036
rect 155374 79971 155402 80036
rect 155270 79960 155322 79966
rect 155270 79902 155322 79908
rect 155360 79962 155416 79971
rect 155466 79966 155494 80036
rect 155558 79966 155586 80036
rect 155650 79971 155678 80036
rect 155360 79897 155416 79906
rect 155454 79960 155506 79966
rect 155454 79902 155506 79908
rect 155546 79960 155598 79966
rect 155546 79902 155598 79908
rect 155636 79962 155692 79971
rect 155636 79897 155692 79906
rect 155454 79824 155506 79830
rect 154118 79727 154174 79736
rect 154396 79756 154448 79762
rect 153844 79688 153896 79694
rect 153844 79630 153896 79636
rect 153936 79688 153988 79694
rect 153936 79630 153988 79636
rect 154028 79688 154080 79694
rect 154028 79630 154080 79636
rect 153856 79540 153884 79630
rect 153856 79512 153976 79540
rect 153844 79416 153896 79422
rect 153842 79384 153844 79393
rect 153896 79384 153898 79393
rect 153842 79319 153898 79328
rect 153948 74497 153976 79512
rect 154040 74633 154068 79630
rect 154026 74624 154082 74633
rect 154026 74559 154082 74568
rect 154028 74520 154080 74526
rect 153934 74488 153990 74497
rect 154028 74462 154080 74468
rect 153934 74423 153990 74432
rect 153752 69420 153804 69426
rect 153752 69362 153804 69368
rect 153580 67606 153884 67634
rect 153292 35488 153344 35494
rect 153292 35430 153344 35436
rect 153200 27192 153252 27198
rect 153200 27134 153252 27140
rect 153016 18896 153068 18902
rect 153016 18838 153068 18844
rect 152832 16108 152884 16114
rect 152832 16050 152884 16056
rect 152556 11960 152608 11966
rect 152556 11902 152608 11908
rect 152384 6886 153056 6914
rect 151820 4140 151872 4146
rect 151820 4082 151872 4088
rect 151084 3528 151136 3534
rect 151084 3470 151136 3476
rect 151832 480 151860 4082
rect 153028 480 153056 6886
rect 153856 6458 153884 67606
rect 153948 14754 153976 74423
rect 154040 73137 154068 74462
rect 154026 73128 154082 73137
rect 154026 73063 154082 73072
rect 154040 58750 154068 73063
rect 154028 58744 154080 58750
rect 154028 58686 154080 58692
rect 153936 14748 153988 14754
rect 153936 14690 153988 14696
rect 153844 6452 153896 6458
rect 153844 6394 153896 6400
rect 154132 5098 154160 79727
rect 154396 79698 154448 79704
rect 154672 79756 154724 79762
rect 154672 79698 154724 79704
rect 154212 79688 154264 79694
rect 154212 79630 154264 79636
rect 154302 79656 154358 79665
rect 154224 74526 154252 79630
rect 154302 79591 154358 79600
rect 154212 74520 154264 74526
rect 154212 74462 154264 74468
rect 154212 74384 154264 74390
rect 154212 74326 154264 74332
rect 154224 38214 154252 74326
rect 154316 73778 154344 79591
rect 154408 79529 154436 79698
rect 154488 79688 154540 79694
rect 154488 79630 154540 79636
rect 154394 79520 154450 79529
rect 154394 79455 154450 79464
rect 154396 79416 154448 79422
rect 154396 79358 154448 79364
rect 154304 73772 154356 73778
rect 154304 73714 154356 73720
rect 154212 38208 154264 38214
rect 154212 38150 154264 38156
rect 154408 20262 154436 79358
rect 154500 77353 154528 79630
rect 154578 79520 154634 79529
rect 154578 79455 154634 79464
rect 154486 77344 154542 77353
rect 154486 77279 154542 77288
rect 154592 74534 154620 79455
rect 154684 79014 154712 79698
rect 154672 79008 154724 79014
rect 154672 78950 154724 78956
rect 154500 74506 154620 74534
rect 154500 74118 154528 74506
rect 154488 74112 154540 74118
rect 154488 74054 154540 74060
rect 154776 68921 154804 79766
rect 154856 79756 154908 79762
rect 155190 79750 155356 79778
rect 155742 79812 155770 80036
rect 155604 79784 155770 79812
rect 155506 79772 155540 79778
rect 155454 79766 155540 79772
rect 155466 79750 155540 79766
rect 154856 79698 154908 79704
rect 154868 76974 154896 79698
rect 155040 79688 155092 79694
rect 155040 79630 155092 79636
rect 154948 79620 155000 79626
rect 154948 79562 155000 79568
rect 154856 76968 154908 76974
rect 154856 76910 154908 76916
rect 154762 68912 154818 68921
rect 154762 68847 154818 68856
rect 154776 61266 154804 68847
rect 154960 61985 154988 79562
rect 155052 63345 155080 79630
rect 155132 79620 155184 79626
rect 155132 79562 155184 79568
rect 155144 79529 155172 79562
rect 155130 79520 155186 79529
rect 155130 79455 155186 79464
rect 155328 79370 155356 79750
rect 155406 79656 155462 79665
rect 155406 79591 155408 79600
rect 155460 79591 155462 79600
rect 155408 79562 155460 79568
rect 155408 79416 155460 79422
rect 155236 79342 155356 79370
rect 155406 79384 155408 79393
rect 155460 79384 155462 79393
rect 155130 78160 155186 78169
rect 155130 78095 155186 78104
rect 155144 67590 155172 78095
rect 155236 73030 155264 79342
rect 155406 79319 155462 79328
rect 155420 79268 155448 79319
rect 155328 79240 155448 79268
rect 155328 76922 155356 79240
rect 155512 79200 155540 79750
rect 155420 79172 155540 79200
rect 155420 77110 155448 79172
rect 155604 77217 155632 79784
rect 155834 79778 155862 80036
rect 155926 79937 155954 80036
rect 155912 79928 155968 79937
rect 156018 79898 156046 80036
rect 155912 79863 155968 79872
rect 156006 79892 156058 79898
rect 156006 79834 156058 79840
rect 155834 79750 155908 79778
rect 155774 79656 155830 79665
rect 155774 79591 155830 79600
rect 155684 79484 155736 79490
rect 155684 79426 155736 79432
rect 155696 79393 155724 79426
rect 155682 79384 155738 79393
rect 155682 79319 155738 79328
rect 155590 77208 155646 77217
rect 155590 77143 155646 77152
rect 155408 77104 155460 77110
rect 155408 77046 155460 77052
rect 155328 76894 155540 76922
rect 155224 73024 155276 73030
rect 155224 72966 155276 72972
rect 155408 73024 155460 73030
rect 155408 72966 155460 72972
rect 155132 67584 155184 67590
rect 155132 67526 155184 67532
rect 155038 63336 155094 63345
rect 155038 63271 155094 63280
rect 154946 61976 155002 61985
rect 154946 61911 155002 61920
rect 154764 61260 154816 61266
rect 154764 61202 154816 61208
rect 155224 61260 155276 61266
rect 155224 61202 155276 61208
rect 154396 20256 154448 20262
rect 154396 20198 154448 20204
rect 155236 20194 155264 61202
rect 155420 42294 155448 72966
rect 155408 42288 155460 42294
rect 155408 42230 155460 42236
rect 155512 41002 155540 76894
rect 155500 40996 155552 41002
rect 155500 40938 155552 40944
rect 155604 34066 155632 77143
rect 155592 34060 155644 34066
rect 155592 34002 155644 34008
rect 155224 20188 155276 20194
rect 155224 20130 155276 20136
rect 155696 20126 155724 79319
rect 155788 79150 155816 79591
rect 155880 79422 155908 79750
rect 156110 79744 156138 80036
rect 156202 79966 156230 80036
rect 156190 79960 156242 79966
rect 156190 79902 156242 79908
rect 156294 79812 156322 80036
rect 156386 79966 156414 80036
rect 156374 79960 156426 79966
rect 156374 79902 156426 79908
rect 156478 79812 156506 80036
rect 156248 79784 156322 79812
rect 156432 79784 156506 79812
rect 156110 79716 156184 79744
rect 156052 79620 156104 79626
rect 156052 79562 156104 79568
rect 155960 79552 156012 79558
rect 155960 79494 156012 79500
rect 155868 79416 155920 79422
rect 155868 79358 155920 79364
rect 155868 79280 155920 79286
rect 155868 79222 155920 79228
rect 155776 79144 155828 79150
rect 155776 79086 155828 79092
rect 155774 78976 155830 78985
rect 155774 78911 155830 78920
rect 155684 20120 155736 20126
rect 155684 20062 155736 20068
rect 155788 19990 155816 78911
rect 155880 77081 155908 79222
rect 155866 77072 155922 77081
rect 155866 77007 155922 77016
rect 155868 74996 155920 75002
rect 155868 74938 155920 74944
rect 155776 19984 155828 19990
rect 155776 19926 155828 19932
rect 155408 6180 155460 6186
rect 155408 6122 155460 6128
rect 154120 5092 154172 5098
rect 154120 5034 154172 5040
rect 154212 2916 154264 2922
rect 154212 2858 154264 2864
rect 154224 480 154252 2858
rect 155420 480 155448 6122
rect 155880 3942 155908 74938
rect 155972 74050 156000 79494
rect 156064 74361 156092 79562
rect 156156 78713 156184 79716
rect 156142 78704 156198 78713
rect 156142 78639 156198 78648
rect 156144 78124 156196 78130
rect 156144 78066 156196 78072
rect 156156 77625 156184 78066
rect 156142 77616 156198 77625
rect 156142 77551 156198 77560
rect 156050 74352 156106 74361
rect 156050 74287 156106 74296
rect 155960 74044 156012 74050
rect 155960 73986 156012 73992
rect 156248 73137 156276 79784
rect 156432 79778 156460 79784
rect 156386 79750 156460 79778
rect 156386 79744 156414 79750
rect 156570 79744 156598 80036
rect 156662 79937 156690 80036
rect 156648 79928 156704 79937
rect 156648 79863 156704 79872
rect 156340 79716 156414 79744
rect 156524 79716 156598 79744
rect 156340 75750 156368 79716
rect 156420 79620 156472 79626
rect 156420 79562 156472 79568
rect 156328 75744 156380 75750
rect 156328 75686 156380 75692
rect 156234 73128 156290 73137
rect 156234 73063 156290 73072
rect 156248 70394 156276 73063
rect 156432 72282 156460 79562
rect 156524 73001 156552 79716
rect 156754 79676 156782 80036
rect 156846 79830 156874 80036
rect 156834 79824 156886 79830
rect 156834 79766 156886 79772
rect 156938 79778 156966 80036
rect 157030 79937 157058 80036
rect 157122 79966 157150 80036
rect 157110 79960 157162 79966
rect 157016 79928 157072 79937
rect 157110 79902 157162 79908
rect 157016 79863 157072 79872
rect 157214 79830 157242 80036
rect 157202 79824 157254 79830
rect 156938 79750 157012 79778
rect 157306 79812 157334 80036
rect 157398 79966 157426 80036
rect 157386 79960 157438 79966
rect 157490 79937 157518 80036
rect 157386 79902 157438 79908
rect 157476 79928 157532 79937
rect 157476 79863 157532 79872
rect 157306 79801 157380 79812
rect 157306 79792 157394 79801
rect 157306 79784 157338 79792
rect 157202 79766 157254 79772
rect 156602 79656 156658 79665
rect 156754 79648 156828 79676
rect 156984 79665 157012 79750
rect 157582 79744 157610 80036
rect 157674 79830 157702 80036
rect 157766 79966 157794 80036
rect 157754 79960 157806 79966
rect 157754 79902 157806 79908
rect 157662 79824 157714 79830
rect 157754 79824 157806 79830
rect 157662 79766 157714 79772
rect 157752 79792 157754 79801
rect 157806 79792 157808 79801
rect 157338 79727 157394 79736
rect 157536 79716 157610 79744
rect 157752 79727 157808 79736
rect 157156 79688 157208 79694
rect 156602 79591 156658 79600
rect 156510 72992 156566 73001
rect 156510 72927 156566 72936
rect 156524 72321 156552 72927
rect 156616 72758 156644 79591
rect 156696 79552 156748 79558
rect 156696 79494 156748 79500
rect 156708 75834 156736 79494
rect 156800 77625 156828 79648
rect 156970 79656 157026 79665
rect 157156 79630 157208 79636
rect 156970 79591 157026 79600
rect 157064 79620 157116 79626
rect 156880 79416 156932 79422
rect 156880 79358 156932 79364
rect 156786 77616 156842 77625
rect 156786 77551 156842 77560
rect 156708 75806 156828 75834
rect 156696 75744 156748 75750
rect 156696 75686 156748 75692
rect 156604 72752 156656 72758
rect 156604 72694 156656 72700
rect 156510 72312 156566 72321
rect 156420 72276 156472 72282
rect 156510 72247 156566 72256
rect 156420 72218 156472 72224
rect 156248 70366 156552 70394
rect 155958 26888 156014 26897
rect 155958 26823 156014 26832
rect 155972 16574 156000 26823
rect 155972 16546 156184 16574
rect 155868 3936 155920 3942
rect 155868 3878 155920 3884
rect 148294 354 148406 480
rect 147876 326 148406 354
rect 148294 -960 148406 326
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156156 354 156184 16546
rect 156524 13258 156552 70366
rect 156604 58676 156656 58682
rect 156604 58618 156656 58624
rect 156512 13252 156564 13258
rect 156512 13194 156564 13200
rect 156616 3398 156644 58618
rect 156708 40934 156736 75686
rect 156800 75002 156828 75806
rect 156788 74996 156840 75002
rect 156788 74938 156840 74944
rect 156786 74352 156842 74361
rect 156786 74287 156842 74296
rect 156696 40928 156748 40934
rect 156696 40870 156748 40876
rect 156800 36786 156828 74287
rect 156892 72865 156920 79358
rect 156984 76838 157012 79591
rect 157064 79562 157116 79568
rect 157076 79393 157104 79562
rect 157062 79384 157118 79393
rect 157062 79319 157118 79328
rect 157076 77790 157104 79319
rect 157064 77784 157116 77790
rect 157064 77726 157116 77732
rect 157168 76922 157196 79630
rect 157248 79620 157300 79626
rect 157248 79562 157300 79568
rect 157432 79620 157484 79626
rect 157432 79562 157484 79568
rect 157260 78577 157288 79562
rect 157340 79416 157392 79422
rect 157340 79358 157392 79364
rect 157246 78568 157302 78577
rect 157246 78503 157302 78512
rect 157076 76894 157196 76922
rect 156972 76832 157024 76838
rect 156972 76774 157024 76780
rect 156970 73128 157026 73137
rect 156970 73063 157026 73072
rect 156878 72856 156934 72865
rect 156878 72791 156934 72800
rect 156984 72729 157012 73063
rect 156970 72720 157026 72729
rect 156970 72655 157026 72664
rect 157076 72593 157104 76894
rect 157156 76832 157208 76838
rect 157156 76774 157208 76780
rect 157062 72584 157118 72593
rect 156892 72542 157062 72570
rect 156788 36780 156840 36786
rect 156788 36722 156840 36728
rect 156892 31278 156920 72542
rect 157062 72519 157118 72528
rect 157062 72448 157118 72457
rect 157062 72383 157118 72392
rect 156970 72312 157026 72321
rect 156970 72247 157026 72256
rect 156880 31272 156932 31278
rect 156880 31214 156932 31220
rect 156984 25838 157012 72247
rect 156972 25832 157024 25838
rect 156972 25774 157024 25780
rect 157076 24410 157104 72383
rect 157064 24404 157116 24410
rect 157064 24346 157116 24352
rect 157168 22982 157196 76774
rect 157260 72690 157288 78503
rect 157248 72684 157300 72690
rect 157248 72626 157300 72632
rect 157352 66230 157380 79358
rect 157444 78402 157472 79562
rect 157536 79422 157564 79716
rect 157858 79676 157886 80036
rect 157614 79656 157670 79665
rect 157614 79591 157670 79600
rect 157720 79648 157886 79676
rect 157524 79416 157576 79422
rect 157524 79358 157576 79364
rect 157522 78976 157578 78985
rect 157522 78911 157578 78920
rect 157432 78396 157484 78402
rect 157432 78338 157484 78344
rect 157432 77784 157484 77790
rect 157432 77726 157484 77732
rect 157340 66224 157392 66230
rect 157340 66166 157392 66172
rect 157156 22976 157208 22982
rect 157156 22918 157208 22924
rect 157444 21690 157472 77726
rect 157432 21684 157484 21690
rect 157432 21626 157484 21632
rect 157536 21622 157564 78911
rect 157628 78538 157656 79591
rect 157720 78577 157748 79648
rect 157950 79608 157978 80036
rect 158042 79966 158070 80036
rect 158134 79966 158162 80036
rect 158030 79960 158082 79966
rect 158030 79902 158082 79908
rect 158122 79960 158174 79966
rect 158122 79902 158174 79908
rect 158076 79824 158128 79830
rect 158076 79766 158128 79772
rect 157904 79580 157978 79608
rect 157800 79552 157852 79558
rect 157800 79494 157852 79500
rect 157706 78568 157762 78577
rect 157616 78532 157668 78538
rect 157706 78503 157762 78512
rect 157616 78474 157668 78480
rect 157708 78396 157760 78402
rect 157708 78338 157760 78344
rect 157720 71738 157748 78338
rect 157812 72622 157840 79494
rect 157904 74526 157932 79580
rect 157984 79484 158036 79490
rect 157984 79426 158036 79432
rect 157996 78674 158024 79426
rect 157984 78668 158036 78674
rect 157984 78610 158036 78616
rect 158088 75993 158116 79766
rect 158226 79676 158254 80036
rect 158180 79648 158254 79676
rect 158074 75984 158130 75993
rect 158074 75919 158130 75928
rect 157982 75848 158038 75857
rect 158180 75834 158208 79648
rect 158318 79608 158346 80036
rect 158410 79966 158438 80036
rect 158502 79966 158530 80036
rect 158398 79960 158450 79966
rect 158398 79902 158450 79908
rect 158490 79960 158542 79966
rect 158594 79937 158622 80036
rect 158490 79902 158542 79908
rect 158580 79928 158636 79937
rect 158580 79863 158636 79872
rect 158398 79824 158450 79830
rect 158396 79792 158398 79801
rect 158450 79792 158452 79801
rect 158686 79778 158714 80036
rect 158778 79966 158806 80036
rect 158766 79960 158818 79966
rect 158870 79937 158898 80036
rect 158766 79902 158818 79908
rect 158856 79928 158912 79937
rect 158962 79898 158990 80036
rect 158856 79863 158912 79872
rect 158950 79892 159002 79898
rect 158950 79834 159002 79840
rect 158810 79792 158866 79801
rect 158686 79750 158760 79778
rect 158396 79727 158452 79736
rect 158626 79656 158682 79665
rect 158272 79580 158346 79608
rect 158444 79620 158496 79626
rect 158272 79393 158300 79580
rect 158626 79591 158682 79600
rect 158444 79562 158496 79568
rect 158258 79384 158314 79393
rect 158258 79319 158314 79328
rect 158038 75806 158208 75834
rect 157982 75783 158038 75792
rect 157892 74520 157944 74526
rect 157892 74462 157944 74468
rect 157800 72616 157852 72622
rect 157800 72558 157852 72564
rect 157708 71732 157760 71738
rect 157708 71674 157760 71680
rect 157996 29850 158024 75783
rect 158168 74520 158220 74526
rect 158168 74462 158220 74468
rect 158076 71732 158128 71738
rect 158076 71674 158128 71680
rect 158088 70854 158116 71674
rect 158076 70848 158128 70854
rect 158076 70790 158128 70796
rect 158088 35426 158116 70790
rect 158180 42226 158208 74462
rect 158272 72554 158300 79319
rect 158456 78792 158484 79562
rect 158364 78764 158484 78792
rect 158260 72548 158312 72554
rect 158260 72490 158312 72496
rect 158364 71738 158392 78764
rect 158444 78668 158496 78674
rect 158444 78610 158496 78616
rect 158352 71732 158404 71738
rect 158352 71674 158404 71680
rect 158456 71126 158484 78610
rect 158640 78282 158668 79591
rect 158732 78849 158760 79750
rect 158810 79727 158866 79736
rect 158904 79756 158956 79762
rect 158824 79150 158852 79727
rect 158904 79698 158956 79704
rect 158812 79144 158864 79150
rect 158812 79086 158864 79092
rect 158718 78840 158774 78849
rect 158718 78775 158774 78784
rect 158640 78254 158760 78282
rect 158628 71732 158680 71738
rect 158628 71674 158680 71680
rect 158640 71194 158668 71674
rect 158628 71188 158680 71194
rect 158628 71130 158680 71136
rect 158444 71120 158496 71126
rect 158444 71062 158496 71068
rect 158456 70394 158484 71062
rect 158456 70366 158576 70394
rect 158168 42220 158220 42226
rect 158168 42162 158220 42168
rect 158076 35420 158128 35426
rect 158076 35362 158128 35368
rect 157984 29844 158036 29850
rect 157984 29786 158036 29792
rect 157524 21616 157576 21622
rect 157524 21558 157576 21564
rect 158548 14686 158576 70366
rect 158536 14680 158588 14686
rect 158536 14622 158588 14628
rect 158640 6390 158668 71130
rect 158732 21554 158760 78254
rect 158916 75914 158944 79698
rect 159054 79676 159082 80036
rect 159146 79937 159174 80036
rect 159238 79966 159266 80036
rect 159330 79966 159358 80036
rect 159226 79960 159278 79966
rect 159132 79928 159188 79937
rect 159226 79902 159278 79908
rect 159318 79960 159370 79966
rect 159318 79902 159370 79908
rect 159422 79898 159450 80036
rect 159514 79966 159542 80036
rect 159502 79960 159554 79966
rect 159502 79902 159554 79908
rect 159132 79863 159188 79872
rect 159410 79892 159462 79898
rect 159410 79834 159462 79840
rect 159180 79824 159232 79830
rect 159178 79792 159180 79801
rect 159232 79792 159234 79801
rect 159178 79727 159234 79736
rect 159456 79756 159508 79762
rect 159054 79648 159128 79676
rect 158916 75886 159036 75914
rect 159008 71262 159036 75886
rect 159100 71738 159128 79648
rect 159192 73982 159220 79727
rect 159606 79744 159634 80036
rect 159698 79971 159726 80036
rect 159684 79962 159740 79971
rect 159790 79966 159818 80036
rect 159882 79971 159910 80036
rect 159684 79897 159740 79906
rect 159778 79960 159830 79966
rect 159778 79902 159830 79908
rect 159868 79962 159924 79971
rect 159868 79897 159924 79906
rect 159974 79898 160002 80036
rect 159962 79892 160014 79898
rect 159962 79834 160014 79840
rect 159732 79824 159784 79830
rect 159732 79766 159784 79772
rect 159914 79792 159970 79801
rect 159456 79698 159508 79704
rect 159560 79716 159634 79744
rect 159364 79688 159416 79694
rect 159364 79630 159416 79636
rect 159272 79620 159324 79626
rect 159272 79562 159324 79568
rect 159180 73976 159232 73982
rect 159180 73918 159232 73924
rect 159088 71732 159140 71738
rect 159088 71674 159140 71680
rect 158996 71256 159048 71262
rect 158996 71198 159048 71204
rect 159284 57866 159312 79562
rect 159376 66162 159404 79630
rect 159364 66156 159416 66162
rect 159364 66098 159416 66104
rect 159468 63510 159496 79698
rect 159560 79676 159588 79716
rect 159560 79648 159680 79676
rect 159548 79552 159600 79558
rect 159548 79494 159600 79500
rect 159560 71670 159588 79494
rect 159652 72894 159680 79648
rect 159640 72888 159692 72894
rect 159640 72830 159692 72836
rect 159548 71664 159600 71670
rect 159548 71606 159600 71612
rect 159560 70394 159588 71606
rect 159652 70514 159680 72830
rect 159744 71913 159772 79766
rect 159824 79756 159876 79762
rect 160066 79744 160094 80036
rect 160158 79801 160186 80036
rect 160250 79966 160278 80036
rect 160238 79960 160290 79966
rect 160342 79937 160370 80036
rect 160434 79966 160462 80036
rect 160422 79960 160474 79966
rect 160238 79902 160290 79908
rect 160328 79928 160384 79937
rect 160422 79902 160474 79908
rect 160328 79863 160384 79872
rect 160526 79812 160554 80036
rect 160618 79966 160646 80036
rect 160606 79960 160658 79966
rect 160606 79902 160658 79908
rect 160710 79898 160738 80036
rect 160698 79892 160750 79898
rect 159914 79727 159970 79736
rect 159824 79698 159876 79704
rect 159836 79665 159864 79698
rect 159822 79656 159878 79665
rect 159822 79591 159878 79600
rect 159836 78198 159864 79591
rect 159824 78192 159876 78198
rect 159824 78134 159876 78140
rect 159928 78044 159956 79727
rect 159836 78016 159956 78044
rect 160020 79716 160094 79744
rect 160144 79792 160200 79801
rect 160388 79784 160554 79812
rect 160604 79826 160660 79835
rect 160698 79834 160750 79840
rect 160144 79727 160200 79736
rect 160284 79756 160336 79762
rect 159730 71904 159786 71913
rect 159730 71839 159786 71848
rect 159640 70508 159692 70514
rect 159640 70450 159692 70456
rect 159560 70366 159772 70394
rect 159456 63504 159508 63510
rect 159456 63446 159508 63452
rect 159272 57860 159324 57866
rect 159272 57802 159324 57808
rect 159744 28490 159772 70366
rect 159732 28484 159784 28490
rect 159732 28426 159784 28432
rect 158720 21548 158772 21554
rect 158720 21490 158772 21496
rect 159836 21486 159864 78016
rect 160020 75041 160048 79716
rect 160284 79698 160336 79704
rect 160192 79688 160244 79694
rect 160098 79656 160154 79665
rect 160192 79630 160244 79636
rect 160098 79591 160154 79600
rect 160112 78062 160140 79591
rect 160204 78742 160232 79630
rect 160296 79354 160324 79698
rect 160284 79348 160336 79354
rect 160284 79290 160336 79296
rect 160192 78736 160244 78742
rect 160192 78678 160244 78684
rect 160100 78056 160152 78062
rect 160100 77998 160152 78004
rect 160204 77908 160232 78678
rect 160112 77880 160232 77908
rect 160006 75032 160062 75041
rect 160006 74967 160062 74976
rect 159916 71732 159968 71738
rect 159916 71674 159968 71680
rect 159928 71466 159956 71674
rect 159916 71460 159968 71466
rect 159916 71402 159968 71408
rect 159824 21480 159876 21486
rect 159824 21422 159876 21428
rect 158902 11656 158958 11665
rect 158902 11591 158958 11600
rect 158628 6384 158680 6390
rect 158628 6326 158680 6332
rect 156604 3392 156656 3398
rect 156604 3334 156656 3340
rect 157800 3392 157852 3398
rect 157800 3334 157852 3340
rect 157812 480 157840 3334
rect 158916 480 158944 11591
rect 159928 10538 159956 71402
rect 160008 70508 160060 70514
rect 160008 70450 160060 70456
rect 160020 11898 160048 70450
rect 160112 16046 160140 77880
rect 160192 72072 160244 72078
rect 160192 72014 160244 72020
rect 160100 16040 160152 16046
rect 160100 15982 160152 15988
rect 160204 15978 160232 72014
rect 160296 18834 160324 79290
rect 160388 79121 160416 79784
rect 160802 79778 160830 80036
rect 160894 79966 160922 80036
rect 160986 79966 161014 80036
rect 161078 79966 161106 80036
rect 161170 79966 161198 80036
rect 160882 79960 160934 79966
rect 160882 79902 160934 79908
rect 160974 79960 161026 79966
rect 160974 79902 161026 79908
rect 161066 79960 161118 79966
rect 161066 79902 161118 79908
rect 161158 79960 161210 79966
rect 161158 79902 161210 79908
rect 161262 79830 161290 80036
rect 161354 79971 161382 80036
rect 161340 79962 161396 79971
rect 161446 79966 161474 80036
rect 161340 79897 161396 79906
rect 161434 79960 161486 79966
rect 161434 79902 161486 79908
rect 160604 79761 160660 79770
rect 160756 79750 160830 79778
rect 160882 79824 160934 79830
rect 161158 79824 161210 79830
rect 161032 79784 161158 79812
rect 160934 79772 160968 79778
rect 160882 79766 160968 79772
rect 160894 79750 160968 79766
rect 160560 79620 160612 79626
rect 160560 79562 160612 79568
rect 160466 79520 160522 79529
rect 160466 79455 160522 79464
rect 160374 79112 160430 79121
rect 160374 79047 160430 79056
rect 160388 71534 160416 79047
rect 160376 71528 160428 71534
rect 160376 71470 160428 71476
rect 160480 64870 160508 79455
rect 160572 72078 160600 79562
rect 160756 79529 160784 79750
rect 160836 79620 160888 79626
rect 160836 79562 160888 79568
rect 160742 79520 160798 79529
rect 160742 79455 160798 79464
rect 160756 74322 160784 79455
rect 160744 74316 160796 74322
rect 160744 74258 160796 74264
rect 160560 72072 160612 72078
rect 160560 72014 160612 72020
rect 160848 71058 160876 79562
rect 160836 71052 160888 71058
rect 160836 70994 160888 71000
rect 160940 67697 160968 79750
rect 160926 67688 160982 67697
rect 160926 67623 160982 67632
rect 161032 67561 161060 79784
rect 161158 79766 161210 79772
rect 161250 79824 161302 79830
rect 161250 79766 161302 79772
rect 161538 79744 161566 80036
rect 161630 79937 161658 80036
rect 161722 79966 161750 80036
rect 161814 79966 161842 80036
rect 161710 79960 161762 79966
rect 161616 79928 161672 79937
rect 161710 79902 161762 79908
rect 161802 79960 161854 79966
rect 161802 79902 161854 79908
rect 161906 79898 161934 80036
rect 161998 79971 162026 80036
rect 161984 79962 162040 79971
rect 162090 79966 162118 80036
rect 161616 79863 161672 79872
rect 161894 79892 161946 79898
rect 161984 79897 162040 79906
rect 162078 79960 162130 79966
rect 162078 79902 162130 79908
rect 161894 79834 161946 79840
rect 161664 79824 161716 79830
rect 161664 79766 161716 79772
rect 161492 79716 161566 79744
rect 161296 79688 161348 79694
rect 161202 79656 161258 79665
rect 161112 79620 161164 79626
rect 161492 79676 161520 79716
rect 161492 79648 161612 79676
rect 161296 79630 161348 79636
rect 161202 79591 161258 79600
rect 161112 79562 161164 79568
rect 161124 78577 161152 79562
rect 161216 79558 161244 79591
rect 161204 79552 161256 79558
rect 161204 79494 161256 79500
rect 161110 78568 161166 78577
rect 161110 78503 161166 78512
rect 161112 78056 161164 78062
rect 161112 77998 161164 78004
rect 161124 71602 161152 77998
rect 161216 74458 161244 79494
rect 161308 79132 161336 79630
rect 161308 79104 161428 79132
rect 161400 75818 161428 79104
rect 161388 75812 161440 75818
rect 161388 75754 161440 75760
rect 161204 74452 161256 74458
rect 161204 74394 161256 74400
rect 161296 74316 161348 74322
rect 161296 74258 161348 74264
rect 161202 74216 161258 74225
rect 161202 74151 161258 74160
rect 161112 71596 161164 71602
rect 161112 71538 161164 71544
rect 161018 67552 161074 67561
rect 161018 67487 161074 67496
rect 160468 64864 160520 64870
rect 160468 64806 160520 64812
rect 160374 33824 160430 33833
rect 160374 33759 160430 33768
rect 160284 18828 160336 18834
rect 160284 18770 160336 18776
rect 160192 15972 160244 15978
rect 160192 15914 160244 15920
rect 160008 11892 160060 11898
rect 160008 11834 160060 11840
rect 159916 10532 159968 10538
rect 159916 10474 159968 10480
rect 160388 6914 160416 33759
rect 161124 32570 161152 71538
rect 161216 38146 161244 74151
rect 161204 38140 161256 38146
rect 161204 38082 161256 38088
rect 161112 32564 161164 32570
rect 161112 32506 161164 32512
rect 161308 29782 161336 74258
rect 161296 29776 161348 29782
rect 161296 29718 161348 29724
rect 161294 15872 161350 15881
rect 161294 15807 161350 15816
rect 160112 6886 160416 6914
rect 160112 480 160140 6886
rect 161308 480 161336 15807
rect 161400 9178 161428 75754
rect 161584 71398 161612 79648
rect 161676 78878 161704 79766
rect 161756 79756 161808 79762
rect 162182 79744 162210 80036
rect 162274 79966 162302 80036
rect 162262 79960 162314 79966
rect 162262 79902 162314 79908
rect 162366 79801 162394 80036
rect 162458 79830 162486 80036
rect 162446 79824 162498 79830
rect 161756 79698 161808 79704
rect 162136 79716 162210 79744
rect 162352 79792 162408 79801
rect 162550 79812 162578 80036
rect 162642 79966 162670 80036
rect 162734 79966 162762 80036
rect 162630 79960 162682 79966
rect 162722 79960 162774 79966
rect 162630 79902 162682 79908
rect 162720 79928 162722 79937
rect 162774 79928 162776 79937
rect 162720 79863 162776 79872
rect 162676 79824 162728 79830
rect 162550 79784 162676 79812
rect 162446 79766 162498 79772
rect 162826 79812 162854 80036
rect 162918 79971 162946 80036
rect 162904 79962 162960 79971
rect 162904 79897 162960 79906
rect 163010 79830 163038 80036
rect 163102 79898 163130 80036
rect 163194 79966 163222 80036
rect 163182 79960 163234 79966
rect 163286 79937 163314 80036
rect 163378 79966 163406 80036
rect 163366 79960 163418 79966
rect 163182 79902 163234 79908
rect 163272 79928 163328 79937
rect 163090 79892 163142 79898
rect 163366 79902 163418 79908
rect 163272 79863 163328 79872
rect 163090 79834 163142 79840
rect 162676 79766 162728 79772
rect 162780 79784 162854 79812
rect 162998 79824 163050 79830
rect 162352 79727 162408 79736
rect 161664 78872 161716 78878
rect 161664 78814 161716 78820
rect 161664 78532 161716 78538
rect 161664 78474 161716 78480
rect 161676 72418 161704 78474
rect 161664 72412 161716 72418
rect 161664 72354 161716 72360
rect 161768 71670 161796 79698
rect 162032 79688 162084 79694
rect 161846 79656 161902 79665
rect 162032 79630 162084 79636
rect 161846 79591 161848 79600
rect 161900 79591 161902 79600
rect 161848 79562 161900 79568
rect 161756 71664 161808 71670
rect 161756 71606 161808 71612
rect 161572 71392 161624 71398
rect 161572 71334 161624 71340
rect 161584 68882 161612 71334
rect 161768 68950 161796 71606
rect 161756 68944 161808 68950
rect 161756 68886 161808 68892
rect 161572 68876 161624 68882
rect 161572 68818 161624 68824
rect 161860 55214 161888 79562
rect 161938 79520 161994 79529
rect 161938 79455 161994 79464
rect 161952 77858 161980 79455
rect 162044 78674 162072 79630
rect 162136 79393 162164 79716
rect 162214 79656 162270 79665
rect 162582 79656 162638 79665
rect 162214 79591 162270 79600
rect 162400 79620 162452 79626
rect 162122 79384 162178 79393
rect 162122 79319 162178 79328
rect 162124 79280 162176 79286
rect 162124 79222 162176 79228
rect 162032 78668 162084 78674
rect 162032 78610 162084 78616
rect 162136 78282 162164 79222
rect 162044 78254 162164 78282
rect 161940 77852 161992 77858
rect 161940 77794 161992 77800
rect 161860 55186 161980 55214
rect 161952 20058 161980 55186
rect 161940 20052 161992 20058
rect 161940 19994 161992 20000
rect 161388 9172 161440 9178
rect 161388 9114 161440 9120
rect 162044 7750 162072 78254
rect 162228 77194 162256 79591
rect 162582 79591 162584 79600
rect 162400 79562 162452 79568
rect 162636 79591 162638 79600
rect 162584 79562 162636 79568
rect 162308 79552 162360 79558
rect 162412 79529 162440 79562
rect 162492 79552 162544 79558
rect 162308 79494 162360 79500
rect 162398 79520 162454 79529
rect 162320 77314 162348 79494
rect 162492 79494 162544 79500
rect 162398 79455 162454 79464
rect 162400 78668 162452 78674
rect 162400 78610 162452 78616
rect 162308 77308 162360 77314
rect 162308 77250 162360 77256
rect 162228 77178 162348 77194
rect 162228 77172 162360 77178
rect 162228 77166 162308 77172
rect 162308 77114 162360 77120
rect 162124 71528 162176 71534
rect 162124 71470 162176 71476
rect 162136 43586 162164 71470
rect 162124 43580 162176 43586
rect 162124 43522 162176 43528
rect 162320 33998 162348 77114
rect 162412 71380 162440 78610
rect 162504 71777 162532 79494
rect 162596 76566 162624 79562
rect 162674 79520 162730 79529
rect 162674 79455 162730 79464
rect 162584 76560 162636 76566
rect 162584 76502 162636 76508
rect 162490 71768 162546 71777
rect 162490 71703 162546 71712
rect 162584 71664 162636 71670
rect 162584 71606 162636 71612
rect 162596 71534 162624 71606
rect 162584 71528 162636 71534
rect 162584 71470 162636 71476
rect 162412 71352 162624 71380
rect 162596 70922 162624 71352
rect 162584 70916 162636 70922
rect 162584 70858 162636 70864
rect 162492 68944 162544 68950
rect 162492 68886 162544 68892
rect 162400 68876 162452 68882
rect 162400 68818 162452 68824
rect 162308 33992 162360 33998
rect 162308 33934 162360 33940
rect 162412 27130 162440 68818
rect 162400 27124 162452 27130
rect 162400 27066 162452 27072
rect 162504 7818 162532 68886
rect 162492 7812 162544 7818
rect 162492 7754 162544 7760
rect 162032 7744 162084 7750
rect 162032 7686 162084 7692
rect 162596 5030 162624 70858
rect 162688 10470 162716 79455
rect 162780 78577 162808 79784
rect 162998 79766 163050 79772
rect 163320 79824 163372 79830
rect 163320 79766 163372 79772
rect 162860 79688 162912 79694
rect 162860 79630 162912 79636
rect 162950 79656 163006 79665
rect 162766 78568 162822 78577
rect 162766 78503 162822 78512
rect 162872 56574 162900 79630
rect 162950 79591 163006 79600
rect 163044 79620 163096 79626
rect 162964 78606 162992 79591
rect 163044 79562 163096 79568
rect 162952 78600 163004 78606
rect 162952 78542 163004 78548
rect 163056 78130 163084 79562
rect 163332 78690 163360 79766
rect 163470 79744 163498 80036
rect 163562 79966 163590 80036
rect 163550 79960 163602 79966
rect 163654 79937 163682 80036
rect 163550 79902 163602 79908
rect 163640 79928 163696 79937
rect 163640 79863 163696 79872
rect 163596 79824 163648 79830
rect 163746 79812 163774 80036
rect 163838 79898 163866 80036
rect 163826 79892 163878 79898
rect 163826 79834 163878 79840
rect 163596 79766 163648 79772
rect 163700 79784 163774 79812
rect 163148 78662 163360 78690
rect 163424 79716 163498 79744
rect 163044 78124 163096 78130
rect 163044 78066 163096 78072
rect 163148 75936 163176 78662
rect 163228 78600 163280 78606
rect 163228 78542 163280 78548
rect 163240 77294 163268 78542
rect 163240 77266 163360 77294
rect 162964 75908 163176 75936
rect 162964 60654 162992 75908
rect 163044 75268 163096 75274
rect 163044 75210 163096 75216
rect 163056 68678 163084 75210
rect 163136 75200 163188 75206
rect 163136 75142 163188 75148
rect 163148 69902 163176 75142
rect 163332 73166 163360 77266
rect 163320 73160 163372 73166
rect 163320 73102 163372 73108
rect 163424 70394 163452 79716
rect 163608 79529 163636 79766
rect 163594 79520 163650 79529
rect 163594 79455 163650 79464
rect 163504 79144 163556 79150
rect 163504 79086 163556 79092
rect 163240 70366 163452 70394
rect 163136 69896 163188 69902
rect 163136 69838 163188 69844
rect 163240 69834 163268 70366
rect 163228 69828 163280 69834
rect 163228 69770 163280 69776
rect 163044 68672 163096 68678
rect 163044 68614 163096 68620
rect 162952 60648 163004 60654
rect 162952 60590 163004 60596
rect 162860 56568 162912 56574
rect 162860 56510 162912 56516
rect 163516 39574 163544 79086
rect 163596 77308 163648 77314
rect 163596 77250 163648 77256
rect 163608 61713 163636 77250
rect 163700 75274 163728 79784
rect 163930 79744 163958 80036
rect 164022 79812 164050 80036
rect 164114 79966 164142 80036
rect 164102 79960 164154 79966
rect 164100 79928 164102 79937
rect 164154 79928 164156 79937
rect 164100 79863 164156 79872
rect 164022 79784 164096 79812
rect 163884 79716 163958 79744
rect 163780 79688 163832 79694
rect 163778 79656 163780 79665
rect 163832 79656 163834 79665
rect 163778 79591 163834 79600
rect 163792 78282 163820 79591
rect 163884 78713 163912 79716
rect 163964 79620 164016 79626
rect 163964 79562 164016 79568
rect 163870 78704 163926 78713
rect 163870 78639 163926 78648
rect 163976 78402 164004 79562
rect 163964 78396 164016 78402
rect 163964 78338 164016 78344
rect 163792 78254 164004 78282
rect 163870 78160 163926 78169
rect 163870 78095 163926 78104
rect 163688 75268 163740 75274
rect 163688 75210 163740 75216
rect 163688 73160 163740 73166
rect 163688 73102 163740 73108
rect 163700 72962 163728 73102
rect 163688 72956 163740 72962
rect 163688 72898 163740 72904
rect 163700 70394 163728 72898
rect 163700 70366 163820 70394
rect 163594 61704 163650 61713
rect 163594 61639 163650 61648
rect 163504 39568 163556 39574
rect 163504 39510 163556 39516
rect 163792 25770 163820 70366
rect 163884 28422 163912 78095
rect 163976 70394 164004 78254
rect 164068 75206 164096 79784
rect 164206 79778 164234 80036
rect 164160 79750 164234 79778
rect 164298 79778 164326 80036
rect 164390 79937 164418 80036
rect 164376 79928 164432 79937
rect 164482 79898 164510 80036
rect 164574 79898 164602 80036
rect 164376 79863 164432 79872
rect 164470 79892 164522 79898
rect 164470 79834 164522 79840
rect 164562 79892 164614 79898
rect 164562 79834 164614 79840
rect 164666 79778 164694 80036
rect 164298 79750 164372 79778
rect 164160 77625 164188 79750
rect 164344 79694 164372 79750
rect 164436 79750 164694 79778
rect 164758 79778 164786 80036
rect 164850 79898 164878 80036
rect 164942 79937 164970 80036
rect 164928 79928 164984 79937
rect 164838 79892 164890 79898
rect 165034 79898 165062 80036
rect 165126 79966 165154 80036
rect 165218 79966 165246 80036
rect 165114 79960 165166 79966
rect 165114 79902 165166 79908
rect 165206 79960 165258 79966
rect 165206 79902 165258 79908
rect 164928 79863 164984 79872
rect 165022 79892 165074 79898
rect 164838 79834 164890 79840
rect 165022 79834 165074 79840
rect 165126 79778 165154 79902
rect 165310 79812 165338 80036
rect 165402 79898 165430 80036
rect 165494 79937 165522 80036
rect 165480 79928 165536 79937
rect 165390 79892 165442 79898
rect 165480 79863 165536 79872
rect 165390 79834 165442 79840
rect 164758 79750 164832 79778
rect 164240 79688 164292 79694
rect 164240 79630 164292 79636
rect 164332 79688 164384 79694
rect 164332 79630 164384 79636
rect 164252 79257 164280 79630
rect 164238 79248 164294 79257
rect 164238 79183 164294 79192
rect 164436 78606 164464 79750
rect 164516 79688 164568 79694
rect 164516 79630 164568 79636
rect 164608 79688 164660 79694
rect 164608 79630 164660 79636
rect 164700 79688 164752 79694
rect 164700 79630 164752 79636
rect 164424 78600 164476 78606
rect 164424 78542 164476 78548
rect 164240 78532 164292 78538
rect 164240 78474 164292 78480
rect 164146 77616 164202 77625
rect 164146 77551 164202 77560
rect 164056 75200 164108 75206
rect 164056 75142 164108 75148
rect 163976 70366 164188 70394
rect 164056 70100 164108 70106
rect 164056 70042 164108 70048
rect 163964 69896 164016 69902
rect 163964 69838 164016 69844
rect 163872 28416 163924 28422
rect 163872 28358 163924 28364
rect 163780 25764 163832 25770
rect 163780 25706 163832 25712
rect 163976 14550 164004 69838
rect 164068 69834 164096 70042
rect 164056 69828 164108 69834
rect 164056 69770 164108 69776
rect 163964 14544 164016 14550
rect 163964 14486 164016 14492
rect 164068 13190 164096 69770
rect 164056 13184 164108 13190
rect 164056 13126 164108 13132
rect 162676 10464 162728 10470
rect 162676 10406 162728 10412
rect 164160 9110 164188 70366
rect 164252 22914 164280 78474
rect 164424 76288 164476 76294
rect 164424 76230 164476 76236
rect 164332 73228 164384 73234
rect 164332 73170 164384 73176
rect 164344 31210 164372 73170
rect 164436 43518 164464 76230
rect 164528 69970 164556 79630
rect 164620 70038 164648 79630
rect 164608 70032 164660 70038
rect 164608 69974 164660 69980
rect 164516 69964 164568 69970
rect 164516 69906 164568 69912
rect 164712 69902 164740 79630
rect 164804 77489 164832 79750
rect 164988 79750 165154 79778
rect 165264 79784 165338 79812
rect 165434 79792 165490 79801
rect 164884 79688 164936 79694
rect 164884 79630 164936 79636
rect 164896 78538 164924 79630
rect 164884 78532 164936 78538
rect 164884 78474 164936 78480
rect 164790 77480 164846 77489
rect 164790 77415 164846 77424
rect 164884 74452 164936 74458
rect 164884 74394 164936 74400
rect 164700 69896 164752 69902
rect 164700 69838 164752 69844
rect 164896 55214 164924 74394
rect 164988 73234 165016 79750
rect 165160 79688 165212 79694
rect 165066 79656 165122 79665
rect 165160 79630 165212 79636
rect 165066 79591 165068 79600
rect 165120 79591 165122 79600
rect 165068 79562 165120 79568
rect 165080 74662 165108 79562
rect 165172 79354 165200 79630
rect 165160 79348 165212 79354
rect 165160 79290 165212 79296
rect 165158 79248 165214 79257
rect 165158 79183 165214 79192
rect 165068 74656 165120 74662
rect 165068 74598 165120 74604
rect 164976 73228 165028 73234
rect 164976 73170 165028 73176
rect 164896 55186 165016 55214
rect 164988 50386 165016 55186
rect 164976 50380 165028 50386
rect 164976 50322 165028 50328
rect 164424 43512 164476 43518
rect 164424 43454 164476 43460
rect 165172 35358 165200 79183
rect 165264 77761 165292 79784
rect 165356 79736 165434 79744
rect 165586 79744 165614 80036
rect 165356 79727 165490 79736
rect 165356 79716 165476 79727
rect 165540 79716 165614 79744
rect 165678 79744 165706 80036
rect 165770 79971 165798 80036
rect 165756 79962 165812 79971
rect 165756 79897 165812 79906
rect 165862 79812 165890 80036
rect 165954 79971 165982 80036
rect 165940 79962 165996 79971
rect 165940 79897 165996 79906
rect 166046 79830 166074 80036
rect 166138 79898 166166 80036
rect 166126 79892 166178 79898
rect 166126 79834 166178 79840
rect 166230 79830 166258 80036
rect 166322 79966 166350 80036
rect 166310 79960 166362 79966
rect 166310 79902 166362 79908
rect 166034 79824 166086 79830
rect 165862 79784 165982 79812
rect 165678 79716 165752 79744
rect 165250 77752 165306 77761
rect 165250 77687 165306 77696
rect 165250 77616 165306 77625
rect 165250 77551 165306 77560
rect 165264 76158 165292 77551
rect 165252 76152 165304 76158
rect 165252 76094 165304 76100
rect 165252 70304 165304 70310
rect 165252 70246 165304 70252
rect 165264 69970 165292 70246
rect 165252 69964 165304 69970
rect 165252 69906 165304 69912
rect 165160 35352 165212 35358
rect 165160 35294 165212 35300
rect 164332 31204 164384 31210
rect 164332 31146 164384 31152
rect 165264 24342 165292 69906
rect 165356 27062 165384 79716
rect 165540 79608 165568 79716
rect 165448 79580 165568 79608
rect 165620 79620 165672 79626
rect 165448 77722 165476 79580
rect 165620 79562 165672 79568
rect 165528 79348 165580 79354
rect 165528 79290 165580 79296
rect 165540 79257 165568 79290
rect 165526 79248 165582 79257
rect 165526 79183 165582 79192
rect 165632 79121 165660 79562
rect 165618 79112 165674 79121
rect 165618 79047 165674 79056
rect 165618 78704 165674 78713
rect 165618 78639 165674 78648
rect 165528 78600 165580 78606
rect 165528 78542 165580 78548
rect 165540 78441 165568 78542
rect 165526 78432 165582 78441
rect 165526 78367 165582 78376
rect 165436 77716 165488 77722
rect 165436 77658 165488 77664
rect 165448 76294 165476 77658
rect 165540 77518 165568 78367
rect 165528 77512 165580 77518
rect 165528 77454 165580 77460
rect 165436 76288 165488 76294
rect 165436 76230 165488 76236
rect 165436 76152 165488 76158
rect 165436 76094 165488 76100
rect 165344 27056 165396 27062
rect 165344 26998 165396 27004
rect 165252 24336 165304 24342
rect 165252 24278 165304 24284
rect 164884 24132 164936 24138
rect 164884 24074 164936 24080
rect 164240 22908 164292 22914
rect 164240 22850 164292 22856
rect 164148 9104 164200 9110
rect 164148 9046 164200 9052
rect 162584 5024 162636 5030
rect 162584 4966 162636 4972
rect 164896 4010 164924 24074
rect 165448 6322 165476 76094
rect 165528 70168 165580 70174
rect 165528 70110 165580 70116
rect 165540 69902 165568 70110
rect 165528 69896 165580 69902
rect 165528 69838 165580 69844
rect 165436 6316 165488 6322
rect 165436 6258 165488 6264
rect 165540 6254 165568 69838
rect 165632 36718 165660 78639
rect 165724 70242 165752 79716
rect 165804 79688 165856 79694
rect 165954 79676 165982 79784
rect 166032 79792 166034 79801
rect 166218 79824 166270 79830
rect 166086 79792 166088 79801
rect 166218 79766 166270 79772
rect 166414 79744 166442 80036
rect 166506 79830 166534 80036
rect 166494 79824 166546 79830
rect 166598 79801 166626 80036
rect 166690 79966 166718 80036
rect 166782 79966 166810 80036
rect 166678 79960 166730 79966
rect 166678 79902 166730 79908
rect 166770 79960 166822 79966
rect 166874 79937 166902 80036
rect 166966 79966 166994 80036
rect 166954 79960 167006 79966
rect 166770 79902 166822 79908
rect 166860 79928 166916 79937
rect 166954 79902 167006 79908
rect 167058 79898 167086 80036
rect 167150 79966 167178 80036
rect 167242 79966 167270 80036
rect 167334 79966 167362 80036
rect 167138 79960 167190 79966
rect 167138 79902 167190 79908
rect 167230 79960 167282 79966
rect 167230 79902 167282 79908
rect 167322 79960 167374 79966
rect 167426 79937 167454 80036
rect 167322 79902 167374 79908
rect 167412 79928 167468 79937
rect 166860 79863 166916 79872
rect 167046 79892 167098 79898
rect 166494 79766 166546 79772
rect 166584 79792 166640 79801
rect 166032 79727 166088 79736
rect 166368 79716 166442 79744
rect 166874 79778 166902 79863
rect 167518 79898 167546 80036
rect 167610 79966 167638 80036
rect 167702 79966 167730 80036
rect 167598 79960 167650 79966
rect 167598 79902 167650 79908
rect 167690 79960 167742 79966
rect 167690 79902 167742 79908
rect 167412 79863 167468 79872
rect 167506 79892 167558 79898
rect 167046 79834 167098 79840
rect 167506 79834 167558 79840
rect 166584 79727 166640 79736
rect 166736 79750 166902 79778
rect 167184 79756 167236 79762
rect 165954 79648 166028 79676
rect 165804 79630 165856 79636
rect 165816 79257 165844 79630
rect 165896 79552 165948 79558
rect 165896 79494 165948 79500
rect 165802 79248 165858 79257
rect 165802 79183 165858 79192
rect 165816 77790 165844 79183
rect 165804 77784 165856 77790
rect 165804 77726 165856 77732
rect 165712 70236 165764 70242
rect 165712 70178 165764 70184
rect 165908 67153 165936 79494
rect 166000 67561 166028 79648
rect 166264 79620 166316 79626
rect 166264 79562 166316 79568
rect 166172 79144 166224 79150
rect 166172 79086 166224 79092
rect 166184 78878 166212 79086
rect 166172 78872 166224 78878
rect 166172 78814 166224 78820
rect 166276 78810 166304 79562
rect 166264 78804 166316 78810
rect 166264 78746 166316 78752
rect 166264 78464 166316 78470
rect 166264 78406 166316 78412
rect 166172 78396 166224 78402
rect 166172 78338 166224 78344
rect 165986 67552 166042 67561
rect 165986 67487 166042 67496
rect 165894 67144 165950 67153
rect 165894 67079 165950 67088
rect 166184 60722 166212 78338
rect 166172 60716 166224 60722
rect 166172 60658 166224 60664
rect 166276 47666 166304 78406
rect 166368 73574 166396 79716
rect 166632 79688 166684 79694
rect 166632 79630 166684 79636
rect 166448 79620 166500 79626
rect 166500 79580 166580 79608
rect 166448 79562 166500 79568
rect 166448 79484 166500 79490
rect 166448 79426 166500 79432
rect 166460 77654 166488 79426
rect 166448 77648 166500 77654
rect 166448 77590 166500 77596
rect 166356 73568 166408 73574
rect 166356 73510 166408 73516
rect 166552 70360 166580 79580
rect 166644 73681 166672 79630
rect 166736 77926 166764 79750
rect 167184 79698 167236 79704
rect 166816 79688 166868 79694
rect 166814 79656 166816 79665
rect 166868 79656 166870 79665
rect 166998 79656 167054 79665
rect 166814 79591 166870 79600
rect 166920 79600 166998 79608
rect 166920 79591 167054 79600
rect 166920 79580 167040 79591
rect 166816 79552 166868 79558
rect 166816 79494 166868 79500
rect 166724 77920 166776 77926
rect 166724 77862 166776 77868
rect 166630 73672 166686 73681
rect 166630 73607 166686 73616
rect 166724 70372 166776 70378
rect 166552 70332 166724 70360
rect 166724 70314 166776 70320
rect 166446 70272 166502 70281
rect 166356 70236 166408 70242
rect 166446 70207 166502 70216
rect 166356 70178 166408 70184
rect 166264 47660 166316 47666
rect 166264 47602 166316 47608
rect 166368 40866 166396 70178
rect 166356 40860 166408 40866
rect 166356 40802 166408 40808
rect 165620 36712 165672 36718
rect 165620 36654 165672 36660
rect 165620 35216 165672 35222
rect 165620 35158 165672 35164
rect 165632 16574 165660 35158
rect 166460 29714 166488 70207
rect 166630 70136 166686 70145
rect 166630 70071 166686 70080
rect 166448 29708 166500 29714
rect 166448 29650 166500 29656
rect 165632 16546 166120 16574
rect 165528 6248 165580 6254
rect 165528 6190 165580 6196
rect 164884 4004 164936 4010
rect 164884 3946 164936 3952
rect 163688 3868 163740 3874
rect 163688 3810 163740 3816
rect 162492 3596 162544 3602
rect 162492 3538 162544 3544
rect 162504 480 162532 3538
rect 163700 480 163728 3810
rect 164884 3800 164936 3806
rect 164884 3742 164936 3748
rect 164896 480 164924 3742
rect 166092 480 166120 16546
rect 166644 15910 166672 70071
rect 166632 15904 166684 15910
rect 166632 15846 166684 15852
rect 166736 11830 166764 70314
rect 166828 18766 166856 79494
rect 166920 70281 166948 79580
rect 167000 78804 167052 78810
rect 167000 78746 167052 78752
rect 167012 74458 167040 78746
rect 167000 74452 167052 74458
rect 167000 74394 167052 74400
rect 166906 70272 166962 70281
rect 166906 70207 166962 70216
rect 167012 60734 167040 74394
rect 167196 73166 167224 79698
rect 167368 79688 167420 79694
rect 167368 79630 167420 79636
rect 167460 79688 167512 79694
rect 167460 79630 167512 79636
rect 167552 79688 167604 79694
rect 167794 79676 167822 80036
rect 167886 79778 167914 80036
rect 167978 79966 168006 80036
rect 168070 79966 168098 80036
rect 168162 79966 168190 80036
rect 168254 79971 168282 80036
rect 167966 79960 168018 79966
rect 167966 79902 168018 79908
rect 168058 79960 168110 79966
rect 168058 79902 168110 79908
rect 168150 79960 168202 79966
rect 168150 79902 168202 79908
rect 168240 79962 168296 79971
rect 168240 79897 168296 79906
rect 168104 79824 168156 79830
rect 168102 79792 168104 79801
rect 168156 79792 168158 79801
rect 167886 79750 168052 79778
rect 167552 79630 167604 79636
rect 167748 79648 167822 79676
rect 167918 79656 167974 79665
rect 167276 79620 167328 79626
rect 167276 79562 167328 79568
rect 167288 79257 167316 79562
rect 167274 79248 167330 79257
rect 167274 79183 167330 79192
rect 167276 78192 167328 78198
rect 167276 78134 167328 78140
rect 167184 73160 167236 73166
rect 167184 73102 167236 73108
rect 167092 72480 167144 72486
rect 167092 72422 167144 72428
rect 166920 60706 167040 60734
rect 166816 18760 166868 18766
rect 166816 18702 166868 18708
rect 166724 11824 166776 11830
rect 166724 11766 166776 11772
rect 166920 10402 166948 60706
rect 167000 46232 167052 46238
rect 167000 46174 167052 46180
rect 167012 16574 167040 46174
rect 167104 40798 167132 72422
rect 167288 69834 167316 78134
rect 167276 69828 167328 69834
rect 167276 69770 167328 69776
rect 167380 69018 167408 79630
rect 167472 73817 167500 79630
rect 167458 73808 167514 73817
rect 167458 73743 167514 73752
rect 167564 73409 167592 79630
rect 167644 79484 167696 79490
rect 167644 79426 167696 79432
rect 167656 78470 167684 79426
rect 167644 78464 167696 78470
rect 167644 78406 167696 78412
rect 167748 78169 167776 79648
rect 168024 79642 168052 79750
rect 168346 79778 168374 80036
rect 168438 79937 168466 80036
rect 168530 79966 168558 80036
rect 168622 79971 168650 80036
rect 168518 79960 168570 79966
rect 168424 79928 168480 79937
rect 168518 79902 168570 79908
rect 168608 79962 168664 79971
rect 168608 79897 168664 79906
rect 168424 79863 168480 79872
rect 168472 79824 168524 79830
rect 168346 79750 168420 79778
rect 168714 79812 168742 80036
rect 168806 79966 168834 80036
rect 168794 79960 168846 79966
rect 168794 79902 168846 79908
rect 168898 79812 168926 80036
rect 168990 79966 169018 80036
rect 169082 79966 169110 80036
rect 169174 79966 169202 80036
rect 168978 79960 169030 79966
rect 169070 79960 169122 79966
rect 168978 79902 169030 79908
rect 169068 79928 169070 79937
rect 169162 79960 169214 79966
rect 169122 79928 169124 79937
rect 169162 79902 169214 79908
rect 169266 79898 169294 80036
rect 169358 79898 169386 80036
rect 169068 79863 169124 79872
rect 169254 79892 169306 79898
rect 169254 79834 169306 79840
rect 169346 79892 169398 79898
rect 169346 79834 169398 79840
rect 169450 79830 169478 80036
rect 169438 79824 169490 79830
rect 168714 79784 168788 79812
rect 168898 79784 169064 79812
rect 168472 79766 168524 79772
rect 168102 79727 168158 79736
rect 168024 79614 168328 79642
rect 167918 79591 167974 79600
rect 167828 79484 167880 79490
rect 167828 79426 167880 79432
rect 167734 78160 167790 78169
rect 167734 78095 167790 78104
rect 167840 75138 167868 79426
rect 167828 75132 167880 75138
rect 167828 75074 167880 75080
rect 167550 73400 167606 73409
rect 167550 73335 167606 73344
rect 167368 69012 167420 69018
rect 167368 68954 167420 68960
rect 167840 45014 167868 75074
rect 167932 46238 167960 79591
rect 168104 79552 168156 79558
rect 168104 79494 168156 79500
rect 168116 73098 168144 79494
rect 168194 79248 168250 79257
rect 168194 79183 168250 79192
rect 168104 73092 168156 73098
rect 168104 73034 168156 73040
rect 168012 69012 168064 69018
rect 168012 68954 168064 68960
rect 167920 46232 167972 46238
rect 167920 46174 167972 46180
rect 167828 45008 167880 45014
rect 167828 44950 167880 44956
rect 167092 40792 167144 40798
rect 167092 40734 167144 40740
rect 168024 17338 168052 68954
rect 168116 17406 168144 73034
rect 168208 22846 168236 79183
rect 168300 78402 168328 79614
rect 168392 79121 168420 79750
rect 168378 79112 168434 79121
rect 168378 79047 168434 79056
rect 168288 78396 168340 78402
rect 168288 78338 168340 78344
rect 168196 22840 168248 22846
rect 168196 22782 168248 22788
rect 168104 17400 168156 17406
rect 168104 17342 168156 17348
rect 168012 17332 168064 17338
rect 168012 17274 168064 17280
rect 167012 16546 167224 16574
rect 166908 10396 166960 10402
rect 166908 10338 166960 10344
rect 167196 480 167224 16546
rect 168300 9042 168328 78338
rect 168392 72486 168420 79047
rect 168484 78538 168512 79766
rect 168564 79620 168616 79626
rect 168564 79562 168616 79568
rect 168472 78532 168524 78538
rect 168472 78474 168524 78480
rect 168472 73636 168524 73642
rect 168472 73578 168524 73584
rect 168380 72480 168432 72486
rect 168380 72422 168432 72428
rect 168380 70440 168432 70446
rect 168380 70382 168432 70388
rect 168392 55214 168420 70382
rect 168484 57934 168512 73578
rect 168576 61441 168604 79562
rect 168656 77852 168708 77858
rect 168656 77794 168708 77800
rect 168668 72486 168696 77794
rect 168656 72480 168708 72486
rect 168656 72422 168708 72428
rect 168760 69630 168788 79784
rect 168932 79688 168984 79694
rect 168932 79630 168984 79636
rect 169036 79642 169064 79784
rect 169542 79812 169570 80036
rect 169634 79966 169662 80036
rect 169726 79971 169754 80036
rect 169622 79960 169674 79966
rect 169622 79902 169674 79908
rect 169712 79962 169768 79971
rect 169712 79897 169768 79906
rect 169542 79784 169616 79812
rect 169438 79766 169490 79772
rect 169392 79688 169444 79694
rect 169298 79656 169354 79665
rect 168840 75880 168892 75886
rect 168840 75822 168892 75828
rect 168748 69624 168800 69630
rect 168748 69566 168800 69572
rect 168852 68950 168880 75822
rect 168944 69902 168972 79630
rect 169036 79614 169156 79642
rect 169024 79552 169076 79558
rect 169024 79494 169076 79500
rect 168932 69896 168984 69902
rect 168932 69838 168984 69844
rect 168840 68944 168892 68950
rect 168840 68886 168892 68892
rect 169036 64802 169064 79494
rect 169128 70446 169156 79614
rect 169208 79620 169260 79626
rect 169392 79630 169444 79636
rect 169482 79656 169538 79665
rect 169298 79591 169354 79600
rect 169208 79562 169260 79568
rect 169220 73642 169248 79562
rect 169312 79490 169340 79591
rect 169300 79484 169352 79490
rect 169300 79426 169352 79432
rect 169208 73636 169260 73642
rect 169208 73578 169260 73584
rect 169116 70440 169168 70446
rect 169116 70382 169168 70388
rect 169024 64796 169076 64802
rect 169024 64738 169076 64744
rect 168562 61432 168618 61441
rect 168562 61367 168618 61376
rect 169312 58682 169340 79426
rect 169404 75993 169432 79630
rect 169482 79591 169484 79600
rect 169536 79591 169538 79600
rect 169484 79562 169536 79568
rect 169390 75984 169446 75993
rect 169390 75919 169446 75928
rect 169496 70394 169524 79562
rect 169588 75886 169616 79784
rect 169668 79756 169720 79762
rect 169818 79744 169846 80036
rect 169910 79898 169938 80036
rect 169898 79892 169950 79898
rect 169898 79834 169950 79840
rect 170002 79744 170030 80036
rect 170094 79801 170122 80036
rect 169668 79698 169720 79704
rect 169772 79716 169846 79744
rect 169956 79716 170030 79744
rect 170080 79792 170136 79801
rect 170080 79727 170136 79736
rect 170186 79744 170214 80036
rect 170278 79966 170306 80036
rect 170266 79960 170318 79966
rect 170266 79902 170318 79908
rect 170370 79898 170398 80036
rect 170462 79937 170490 80036
rect 170448 79928 170504 79937
rect 170358 79892 170410 79898
rect 170554 79898 170582 80036
rect 170448 79863 170504 79872
rect 170542 79892 170594 79898
rect 170358 79834 170410 79840
rect 170542 79834 170594 79840
rect 170404 79756 170456 79762
rect 170186 79716 170260 79744
rect 169680 79257 169708 79698
rect 169666 79248 169722 79257
rect 169666 79183 169722 79192
rect 169680 77994 169708 79183
rect 169668 77988 169720 77994
rect 169668 77930 169720 77936
rect 169772 77178 169800 79716
rect 169852 79620 169904 79626
rect 169852 79562 169904 79568
rect 169864 78849 169892 79562
rect 169850 78840 169906 78849
rect 169850 78775 169906 78784
rect 169760 77172 169812 77178
rect 169760 77114 169812 77120
rect 169772 76362 169800 77114
rect 169760 76356 169812 76362
rect 169760 76298 169812 76304
rect 169576 75880 169628 75886
rect 169576 75822 169628 75828
rect 169496 70366 169708 70394
rect 169392 69896 169444 69902
rect 169392 69838 169444 69844
rect 169404 68814 169432 69838
rect 169484 69624 169536 69630
rect 169484 69566 169536 69572
rect 169496 68882 169524 69566
rect 169576 68944 169628 68950
rect 169576 68886 169628 68892
rect 169484 68876 169536 68882
rect 169484 68818 169536 68824
rect 169392 68808 169444 68814
rect 169392 68750 169444 68756
rect 169300 58676 169352 58682
rect 169300 58618 169352 58624
rect 168472 57928 168524 57934
rect 168472 57870 168524 57876
rect 168380 55208 168432 55214
rect 168380 55150 168432 55156
rect 168472 51740 168524 51746
rect 168472 51682 168524 51688
rect 168484 16574 168512 51682
rect 169404 39506 169432 68750
rect 169392 39500 169444 39506
rect 169392 39442 169444 39448
rect 169496 31142 169524 68818
rect 169484 31136 169536 31142
rect 169484 31078 169536 31084
rect 169588 28354 169616 68886
rect 169680 33930 169708 70366
rect 169864 64874 169892 78775
rect 169956 78305 169984 79716
rect 170232 79665 170260 79716
rect 170646 79744 170674 80036
rect 170738 79937 170766 80036
rect 170830 79966 170858 80036
rect 170818 79960 170870 79966
rect 170724 79928 170780 79937
rect 170818 79902 170870 79908
rect 170724 79863 170780 79872
rect 170922 79830 170950 80036
rect 171014 79971 171042 80036
rect 171000 79962 171056 79971
rect 171000 79897 171056 79906
rect 170772 79824 170824 79830
rect 170772 79766 170824 79772
rect 170910 79824 170962 79830
rect 170910 79766 170962 79772
rect 170646 79716 170720 79744
rect 170404 79698 170456 79704
rect 170312 79688 170364 79694
rect 170218 79656 170274 79665
rect 170036 79620 170088 79626
rect 170312 79630 170364 79636
rect 170218 79591 170274 79600
rect 170036 79562 170088 79568
rect 169942 78296 169998 78305
rect 169942 78231 169998 78240
rect 170048 78198 170076 79562
rect 170036 78192 170088 78198
rect 170036 78134 170088 78140
rect 170232 70394 170260 79591
rect 170324 75449 170352 79630
rect 170416 76786 170444 79698
rect 170496 79620 170548 79626
rect 170496 79562 170548 79568
rect 170508 77353 170536 79562
rect 170494 77344 170550 77353
rect 170494 77279 170550 77288
rect 170586 76936 170642 76945
rect 170586 76871 170642 76880
rect 170692 76888 170720 79716
rect 170784 79642 170812 79766
rect 171106 79744 171134 80036
rect 171198 79778 171226 80036
rect 171290 79966 171318 80036
rect 171382 79971 171410 80036
rect 171278 79960 171330 79966
rect 171278 79902 171330 79908
rect 171368 79962 171424 79971
rect 171368 79897 171424 79906
rect 171474 79898 171502 80036
rect 171566 79937 171594 80036
rect 171658 79966 171686 80036
rect 171750 79966 171778 80036
rect 171842 79966 171870 80036
rect 171934 79966 171962 80036
rect 172026 79971 172054 80036
rect 171646 79960 171698 79966
rect 171552 79928 171608 79937
rect 171462 79892 171514 79898
rect 171646 79902 171698 79908
rect 171738 79960 171790 79966
rect 171738 79902 171790 79908
rect 171830 79960 171882 79966
rect 171830 79902 171882 79908
rect 171922 79960 171974 79966
rect 171922 79902 171974 79908
rect 172012 79962 172068 79971
rect 172118 79966 172146 80036
rect 172012 79897 172068 79906
rect 172106 79960 172158 79966
rect 172106 79902 172158 79908
rect 171552 79863 171608 79872
rect 171462 79834 171514 79840
rect 171692 79824 171744 79830
rect 171198 79750 171364 79778
rect 171692 79766 171744 79772
rect 171782 79792 171838 79801
rect 171060 79716 171134 79744
rect 170954 79656 171010 79665
rect 170784 79614 170904 79642
rect 170772 79552 170824 79558
rect 170772 79494 170824 79500
rect 170784 77353 170812 79494
rect 170876 77489 170904 79614
rect 170954 79591 171010 79600
rect 170862 77480 170918 77489
rect 170862 77415 170918 77424
rect 170770 77344 170826 77353
rect 170770 77279 170826 77288
rect 170864 77308 170916 77314
rect 170864 77250 170916 77256
rect 170600 76786 170628 76871
rect 170692 76860 170812 76888
rect 170416 76758 170720 76786
rect 170588 76356 170640 76362
rect 170588 76298 170640 76304
rect 170310 75440 170366 75449
rect 170310 75375 170366 75384
rect 170232 70366 170352 70394
rect 169772 64846 169892 64874
rect 169668 33924 169720 33930
rect 169668 33866 169720 33872
rect 169576 28348 169628 28354
rect 169576 28290 169628 28296
rect 168484 16546 169616 16574
rect 168288 9036 168340 9042
rect 168288 8978 168340 8984
rect 168380 4004 168432 4010
rect 168380 3946 168432 3952
rect 168392 480 168420 3946
rect 169588 480 169616 16546
rect 169772 7682 169800 64846
rect 169760 7676 169812 7682
rect 169760 7618 169812 7624
rect 170324 4894 170352 70366
rect 170600 39438 170628 76298
rect 170588 39432 170640 39438
rect 170588 39374 170640 39380
rect 170692 38078 170720 76758
rect 170784 76537 170812 76860
rect 170770 76528 170826 76537
rect 170770 76463 170826 76472
rect 170680 38072 170732 38078
rect 170680 38014 170732 38020
rect 170402 37904 170458 37913
rect 170402 37839 170458 37848
rect 170312 4888 170364 4894
rect 170312 4830 170364 4836
rect 170416 3806 170444 37839
rect 170784 35290 170812 76463
rect 170772 35284 170824 35290
rect 170772 35226 170824 35232
rect 170876 33862 170904 77250
rect 170864 33856 170916 33862
rect 170864 33798 170916 33804
rect 170968 13122 170996 79591
rect 171060 69902 171088 79716
rect 171140 79620 171192 79626
rect 171140 79562 171192 79568
rect 171152 79082 171180 79562
rect 171140 79076 171192 79082
rect 171140 79018 171192 79024
rect 171230 78840 171286 78849
rect 171230 78775 171286 78784
rect 171138 78160 171194 78169
rect 171138 78095 171194 78104
rect 171152 77314 171180 78095
rect 171140 77308 171192 77314
rect 171140 77250 171192 77256
rect 171048 69896 171100 69902
rect 171048 69838 171100 69844
rect 171244 28286 171272 78775
rect 171336 74322 171364 79750
rect 171416 79756 171468 79762
rect 171416 79698 171468 79704
rect 171428 78985 171456 79698
rect 171508 79688 171560 79694
rect 171508 79630 171560 79636
rect 171414 78976 171470 78985
rect 171414 78911 171470 78920
rect 171324 74316 171376 74322
rect 171324 74258 171376 74264
rect 171324 73772 171376 73778
rect 171324 73714 171376 73720
rect 171336 29646 171364 73714
rect 171428 49026 171456 78911
rect 171520 76809 171548 79630
rect 171600 79416 171652 79422
rect 171600 79358 171652 79364
rect 171612 78946 171640 79358
rect 171600 78940 171652 78946
rect 171600 78882 171652 78888
rect 171704 78577 171732 79766
rect 172058 79792 172114 79801
rect 171782 79727 171784 79736
rect 171836 79727 171838 79736
rect 171968 79756 172020 79762
rect 171784 79698 171836 79704
rect 172210 79778 172238 80036
rect 172302 79971 172330 80036
rect 172288 79962 172344 79971
rect 172394 79966 172422 80036
rect 172288 79897 172344 79906
rect 172382 79960 172434 79966
rect 172382 79902 172434 79908
rect 172486 79898 172514 80036
rect 172578 79898 172606 80036
rect 172474 79892 172526 79898
rect 172474 79834 172526 79840
rect 172566 79892 172618 79898
rect 172566 79834 172618 79840
rect 172210 79750 172284 79778
rect 172058 79727 172060 79736
rect 171968 79698 172020 79704
rect 172112 79727 172114 79736
rect 172060 79698 172112 79704
rect 171784 79620 171836 79626
rect 171784 79562 171836 79568
rect 171690 78568 171746 78577
rect 171690 78503 171746 78512
rect 171598 77888 171654 77897
rect 171598 77823 171654 77832
rect 171612 77042 171640 77823
rect 171600 77036 171652 77042
rect 171600 76978 171652 76984
rect 171506 76800 171562 76809
rect 171506 76735 171562 76744
rect 171520 72350 171548 76735
rect 171704 73778 171732 78503
rect 171692 73772 171744 73778
rect 171692 73714 171744 73720
rect 171508 72344 171560 72350
rect 171508 72286 171560 72292
rect 171796 68921 171824 79562
rect 171980 79393 172008 79698
rect 171966 79384 172022 79393
rect 171966 79319 172022 79328
rect 171966 79248 172022 79257
rect 171966 79183 172022 79192
rect 171876 78328 171928 78334
rect 171876 78270 171928 78276
rect 171888 77858 171916 78270
rect 171876 77852 171928 77858
rect 171876 77794 171928 77800
rect 171874 77752 171930 77761
rect 171874 77687 171930 77696
rect 171782 68912 171838 68921
rect 171782 68847 171838 68856
rect 171416 49020 171468 49026
rect 171416 48962 171468 48968
rect 171324 29640 171376 29646
rect 171324 29582 171376 29588
rect 171232 28280 171284 28286
rect 171232 28222 171284 28228
rect 171888 26994 171916 77687
rect 171876 26988 171928 26994
rect 171876 26930 171928 26936
rect 171784 25560 171836 25566
rect 171784 25502 171836 25508
rect 170956 13116 171008 13122
rect 170956 13058 171008 13064
rect 170404 3800 170456 3806
rect 170404 3742 170456 3748
rect 170772 3732 170824 3738
rect 170772 3674 170824 3680
rect 170784 480 170812 3674
rect 171796 3534 171824 25502
rect 171980 17270 172008 79183
rect 171968 17264 172020 17270
rect 171874 17232 171930 17241
rect 171968 17206 172020 17212
rect 171874 17167 171930 17176
rect 171888 3602 171916 17167
rect 172072 14482 172100 79698
rect 172152 79620 172204 79626
rect 172152 79562 172204 79568
rect 172164 76129 172192 79562
rect 172150 76120 172206 76129
rect 172150 76055 172206 76064
rect 172256 75993 172284 79750
rect 172336 79756 172388 79762
rect 172670 79744 172698 80036
rect 172762 79937 172790 80036
rect 172854 79966 172882 80036
rect 172842 79960 172894 79966
rect 172748 79928 172804 79937
rect 172842 79902 172894 79908
rect 172748 79863 172804 79872
rect 172946 79830 172974 80036
rect 173038 79966 173066 80036
rect 173130 79966 173158 80036
rect 173026 79960 173078 79966
rect 173026 79902 173078 79908
rect 173118 79960 173170 79966
rect 173118 79902 173170 79908
rect 172934 79824 172986 79830
rect 173222 79801 173250 80036
rect 173314 79966 173342 80036
rect 173302 79960 173354 79966
rect 173302 79902 173354 79908
rect 173208 79792 173264 79801
rect 172934 79766 172986 79772
rect 172336 79698 172388 79704
rect 172624 79716 172698 79744
rect 173084 79750 173208 79778
rect 172348 79393 172376 79698
rect 172428 79688 172480 79694
rect 172428 79630 172480 79636
rect 172334 79384 172390 79393
rect 172334 79319 172390 79328
rect 172242 75984 172298 75993
rect 172242 75919 172298 75928
rect 172348 75206 172376 79319
rect 172440 78198 172468 79630
rect 172428 78192 172480 78198
rect 172428 78134 172480 78140
rect 172520 76900 172572 76906
rect 172520 76842 172572 76848
rect 172336 75200 172388 75206
rect 172336 75142 172388 75148
rect 172152 74316 172204 74322
rect 172152 74258 172204 74264
rect 172164 73710 172192 74258
rect 172152 73704 172204 73710
rect 172152 73646 172204 73652
rect 172164 42158 172192 73646
rect 172244 72344 172296 72350
rect 172244 72286 172296 72292
rect 172256 43450 172284 72286
rect 172426 71360 172482 71369
rect 172426 71295 172428 71304
rect 172480 71295 172482 71304
rect 172428 71266 172480 71272
rect 172244 43444 172296 43450
rect 172244 43386 172296 43392
rect 172152 42152 172204 42158
rect 172152 42094 172204 42100
rect 172532 24206 172560 76842
rect 172624 75993 172652 79716
rect 172888 79688 172940 79694
rect 172940 79648 173020 79676
rect 172888 79630 172940 79636
rect 172796 79620 172848 79626
rect 172796 79562 172848 79568
rect 172808 78985 172836 79562
rect 172888 79484 172940 79490
rect 172888 79426 172940 79432
rect 172794 78976 172850 78985
rect 172794 78911 172850 78920
rect 172610 75984 172666 75993
rect 172610 75919 172666 75928
rect 172808 67634 172836 78911
rect 172900 75274 172928 79426
rect 172992 79393 173020 79648
rect 172978 79384 173034 79393
rect 172978 79319 173034 79328
rect 172992 75313 173020 79319
rect 173084 76022 173112 79750
rect 173208 79727 173264 79736
rect 173406 79744 173434 80036
rect 173498 79812 173526 80036
rect 173590 79966 173618 80036
rect 173682 79966 173710 80036
rect 173774 79966 173802 80036
rect 173578 79960 173630 79966
rect 173578 79902 173630 79908
rect 173670 79960 173722 79966
rect 173670 79902 173722 79908
rect 173762 79960 173814 79966
rect 173762 79902 173814 79908
rect 173716 79824 173768 79830
rect 173498 79784 173664 79812
rect 173406 79716 173480 79744
rect 173164 79688 173216 79694
rect 173164 79630 173216 79636
rect 173072 76016 173124 76022
rect 173072 75958 173124 75964
rect 172978 75304 173034 75313
rect 172888 75268 172940 75274
rect 172978 75239 173034 75248
rect 172888 75210 172940 75216
rect 173176 73817 173204 79630
rect 173256 79620 173308 79626
rect 173256 79562 173308 79568
rect 173268 79257 173296 79562
rect 173348 79552 173400 79558
rect 173348 79494 173400 79500
rect 173254 79248 173310 79257
rect 173254 79183 173310 79192
rect 173256 79076 173308 79082
rect 173256 79018 173308 79024
rect 173268 75342 173296 79018
rect 173360 76362 173388 79494
rect 173452 79404 173480 79716
rect 173452 79376 173572 79404
rect 173440 79280 173492 79286
rect 173440 79222 173492 79228
rect 173452 78985 173480 79222
rect 173544 79218 173572 79376
rect 173532 79212 173584 79218
rect 173532 79154 173584 79160
rect 173438 78976 173494 78985
rect 173438 78911 173494 78920
rect 173348 76356 173400 76362
rect 173348 76298 173400 76304
rect 173256 75336 173308 75342
rect 173256 75278 173308 75284
rect 173162 73808 173218 73817
rect 173162 73743 173218 73752
rect 172624 67606 172836 67634
rect 173360 67634 173388 76298
rect 173452 76294 173480 78911
rect 173544 76906 173572 79154
rect 173636 78849 173664 79784
rect 173866 79778 173894 80036
rect 173958 79966 173986 80036
rect 173946 79960 173998 79966
rect 173944 79928 173946 79937
rect 173998 79928 174000 79937
rect 174050 79898 174078 80036
rect 174142 79937 174170 80036
rect 174128 79928 174184 79937
rect 173944 79863 174000 79872
rect 174038 79892 174090 79898
rect 174128 79863 174184 79872
rect 174038 79834 174090 79840
rect 173716 79766 173768 79772
rect 173622 78840 173678 78849
rect 173622 78775 173678 78784
rect 173532 76900 173584 76906
rect 173532 76842 173584 76848
rect 173440 76288 173492 76294
rect 173440 76230 173492 76236
rect 173360 67606 173572 67634
rect 172624 25634 172652 67606
rect 173544 40730 173572 67606
rect 173532 40724 173584 40730
rect 173532 40666 173584 40672
rect 173636 38010 173664 78775
rect 173728 76401 173756 79766
rect 173820 79750 173894 79778
rect 174082 79792 174138 79801
rect 173992 79756 174044 79762
rect 173714 76392 173770 76401
rect 173714 76327 173770 76336
rect 173716 76288 173768 76294
rect 173716 76230 173768 76236
rect 173624 38004 173676 38010
rect 173624 37946 173676 37952
rect 173728 32502 173756 76230
rect 173820 76129 173848 79750
rect 174082 79727 174138 79736
rect 174234 79744 174262 80036
rect 174326 79898 174354 80036
rect 174418 79898 174446 80036
rect 174510 79966 174538 80036
rect 174498 79960 174550 79966
rect 174602 79937 174630 80036
rect 174694 79966 174722 80036
rect 174682 79960 174734 79966
rect 174498 79902 174550 79908
rect 174588 79928 174644 79937
rect 174314 79892 174366 79898
rect 174314 79834 174366 79840
rect 174406 79892 174458 79898
rect 174682 79902 174734 79908
rect 174588 79863 174644 79872
rect 174406 79834 174458 79840
rect 174498 79824 174550 79830
rect 174358 79792 174414 79801
rect 173992 79698 174044 79704
rect 173900 79688 173952 79694
rect 173900 79630 173952 79636
rect 173912 79354 173940 79630
rect 173900 79348 173952 79354
rect 173900 79290 173952 79296
rect 173806 76120 173862 76129
rect 173806 76055 173862 76064
rect 173808 76016 173860 76022
rect 173808 75958 173860 75964
rect 173716 32496 173768 32502
rect 173716 32438 173768 32444
rect 172612 25628 172664 25634
rect 172612 25570 172664 25576
rect 172520 24200 172572 24206
rect 172520 24142 172572 24148
rect 172060 14476 172112 14482
rect 172060 14418 172112 14424
rect 173820 6186 173848 75958
rect 173900 75948 173952 75954
rect 173900 75890 173952 75896
rect 173912 7614 173940 75890
rect 174004 74934 174032 79698
rect 174096 78606 174124 79727
rect 174234 79716 174308 79744
rect 174358 79727 174414 79736
rect 174496 79792 174498 79801
rect 174602 79812 174630 79863
rect 174550 79792 174552 79801
rect 174602 79784 174676 79812
rect 174496 79727 174552 79736
rect 174176 79620 174228 79626
rect 174176 79562 174228 79568
rect 174084 78600 174136 78606
rect 174084 78542 174136 78548
rect 173992 74928 174044 74934
rect 173992 74870 174044 74876
rect 173992 74792 174044 74798
rect 173992 74734 174044 74740
rect 174004 22778 174032 74734
rect 174188 71774 174216 79562
rect 174280 78985 174308 79716
rect 174266 78976 174322 78985
rect 174266 78911 174322 78920
rect 174280 74798 174308 78911
rect 174372 76022 174400 79727
rect 174544 79688 174596 79694
rect 174544 79630 174596 79636
rect 174452 79620 174504 79626
rect 174452 79562 174504 79568
rect 174464 79393 174492 79562
rect 174450 79384 174506 79393
rect 174450 79319 174506 79328
rect 174556 79200 174584 79630
rect 174464 79172 174584 79200
rect 174360 76016 174412 76022
rect 174360 75958 174412 75964
rect 174464 75857 174492 79172
rect 174544 79076 174596 79082
rect 174544 79018 174596 79024
rect 174556 75954 174584 79018
rect 174544 75948 174596 75954
rect 174544 75890 174596 75896
rect 174450 75848 174506 75857
rect 174450 75783 174506 75792
rect 174268 74792 174320 74798
rect 174268 74734 174320 74740
rect 174096 71746 174216 71774
rect 174096 39370 174124 71746
rect 174648 67634 174676 79784
rect 174786 79778 174814 80036
rect 174878 79937 174906 80036
rect 174864 79928 174920 79937
rect 174970 79898 174998 80036
rect 174864 79863 174920 79872
rect 174958 79892 175010 79898
rect 174958 79834 175010 79840
rect 174910 79792 174966 79801
rect 174786 79750 174860 79778
rect 174728 79484 174780 79490
rect 174728 79426 174780 79432
rect 174740 74225 174768 79426
rect 174832 79082 174860 79750
rect 175062 79778 175090 80036
rect 174910 79727 174966 79736
rect 175016 79750 175090 79778
rect 174924 79370 174952 79727
rect 175016 79490 175044 79750
rect 175154 79642 175182 80036
rect 175246 79937 175274 80036
rect 175232 79928 175288 79937
rect 175232 79863 175288 79872
rect 175338 79778 175366 80036
rect 175430 79937 175458 80036
rect 175522 79966 175550 80036
rect 175510 79960 175562 79966
rect 175416 79928 175472 79937
rect 175510 79902 175562 79908
rect 175416 79863 175472 79872
rect 175464 79824 175516 79830
rect 175338 79750 175412 79778
rect 175614 79778 175642 80036
rect 175706 79898 175734 80036
rect 175694 79892 175746 79898
rect 175694 79834 175746 79840
rect 175464 79766 175516 79772
rect 175108 79614 175182 79642
rect 175280 79620 175332 79626
rect 175004 79484 175056 79490
rect 175004 79426 175056 79432
rect 174924 79342 175044 79370
rect 174820 79076 174872 79082
rect 174820 79018 174872 79024
rect 174818 78840 174874 78849
rect 174818 78775 174874 78784
rect 174726 74216 174782 74225
rect 174726 74151 174782 74160
rect 174648 67606 174768 67634
rect 174740 47598 174768 67606
rect 174728 47592 174780 47598
rect 174728 47534 174780 47540
rect 174832 42090 174860 78775
rect 174910 77616 174966 77625
rect 174910 77551 174966 77560
rect 174924 75177 174952 77551
rect 174910 75168 174966 75177
rect 174910 75103 174966 75112
rect 174912 74928 174964 74934
rect 174912 74870 174964 74876
rect 174924 70990 174952 74870
rect 174912 70984 174964 70990
rect 174912 70926 174964 70932
rect 174820 42084 174872 42090
rect 174820 42026 174872 42032
rect 174084 39364 174136 39370
rect 174084 39306 174136 39312
rect 174924 26926 174952 70926
rect 174912 26920 174964 26926
rect 174912 26862 174964 26868
rect 175016 25566 175044 79342
rect 175108 77625 175136 79614
rect 175280 79562 175332 79568
rect 175188 79348 175240 79354
rect 175188 79290 175240 79296
rect 175200 78674 175228 79290
rect 175292 78849 175320 79562
rect 175278 78840 175334 78849
rect 175278 78775 175334 78784
rect 175278 78704 175334 78713
rect 175188 78668 175240 78674
rect 175278 78639 175334 78648
rect 175188 78610 175240 78616
rect 175094 77616 175150 77625
rect 175094 77551 175150 77560
rect 175188 76016 175240 76022
rect 175188 75958 175240 75964
rect 175200 75585 175228 75958
rect 175186 75576 175242 75585
rect 175186 75511 175242 75520
rect 175094 74216 175150 74225
rect 175094 74151 175150 74160
rect 175004 25560 175056 25566
rect 175004 25502 175056 25508
rect 173992 22772 174044 22778
rect 173992 22714 174044 22720
rect 175108 11762 175136 74151
rect 175096 11756 175148 11762
rect 175096 11698 175148 11704
rect 173900 7608 173952 7614
rect 173900 7550 173952 7556
rect 173808 6180 173860 6186
rect 173808 6122 173860 6128
rect 175200 4826 175228 75511
rect 175292 44946 175320 78639
rect 175384 74322 175412 79750
rect 175372 74316 175424 74322
rect 175372 74258 175424 74264
rect 175476 71777 175504 79766
rect 175568 79750 175642 79778
rect 175568 73778 175596 79750
rect 175798 79744 175826 80036
rect 175890 79898 175918 80036
rect 175982 79937 176010 80036
rect 175968 79928 176024 79937
rect 175878 79892 175930 79898
rect 175968 79863 176024 79872
rect 175878 79834 175930 79840
rect 175752 79716 175826 79744
rect 175922 79792 175978 79801
rect 176074 79744 176102 80036
rect 176166 79801 176194 80036
rect 176258 79966 176286 80036
rect 176350 79966 176378 80036
rect 176246 79960 176298 79966
rect 176246 79902 176298 79908
rect 176338 79960 176390 79966
rect 176338 79902 176390 79908
rect 176292 79824 176344 79830
rect 175922 79727 175924 79736
rect 175648 79620 175700 79626
rect 175648 79562 175700 79568
rect 175660 79257 175688 79562
rect 175752 79393 175780 79716
rect 175976 79727 175978 79736
rect 175924 79698 175976 79704
rect 176028 79716 176102 79744
rect 176152 79792 176208 79801
rect 176152 79727 176208 79736
rect 176290 79792 176292 79801
rect 176442 79812 176470 80036
rect 176534 79937 176562 80036
rect 176520 79928 176576 79937
rect 176520 79863 176576 79872
rect 176534 79830 176562 79863
rect 176344 79792 176346 79801
rect 176290 79727 176346 79736
rect 176396 79784 176470 79812
rect 176522 79824 176574 79830
rect 175936 79472 175964 79698
rect 176028 79540 176056 79716
rect 176106 79656 176162 79665
rect 176162 79614 176240 79642
rect 176106 79591 176162 79600
rect 176028 79512 176148 79540
rect 175936 79444 176056 79472
rect 175738 79384 175794 79393
rect 175738 79319 175794 79328
rect 175832 79280 175884 79286
rect 175646 79248 175702 79257
rect 175832 79222 175884 79228
rect 175922 79248 175978 79257
rect 175646 79183 175702 79192
rect 175844 79082 175872 79222
rect 175922 79183 175978 79192
rect 175832 79076 175884 79082
rect 175832 79018 175884 79024
rect 175738 78840 175794 78849
rect 175738 78775 175794 78784
rect 175556 73772 175608 73778
rect 175556 73714 175608 73720
rect 175462 71768 175518 71777
rect 175462 71703 175518 71712
rect 175752 70394 175780 78775
rect 175752 70366 175872 70394
rect 175280 44940 175332 44946
rect 175280 44882 175332 44888
rect 175844 36650 175872 70366
rect 175832 36644 175884 36650
rect 175832 36586 175884 36592
rect 175936 33794 175964 79183
rect 176028 53106 176056 79444
rect 176120 70145 176148 79512
rect 176212 78810 176240 79614
rect 176200 78804 176252 78810
rect 176200 78746 176252 78752
rect 176200 74316 176252 74322
rect 176200 74258 176252 74264
rect 176106 70136 176162 70145
rect 176106 70071 176162 70080
rect 176016 53100 176068 53106
rect 176016 53042 176068 53048
rect 176212 37942 176240 74258
rect 176200 37936 176252 37942
rect 176200 37878 176252 37884
rect 175924 33788 175976 33794
rect 175924 33730 175976 33736
rect 176304 24138 176332 79727
rect 176396 78713 176424 79784
rect 176522 79766 176574 79772
rect 176476 79688 176528 79694
rect 176626 79676 176654 80036
rect 176718 79971 176746 80036
rect 176704 79962 176760 79971
rect 176704 79897 176760 79906
rect 176810 79744 176838 80036
rect 176476 79630 176528 79636
rect 176580 79648 176654 79676
rect 176764 79716 176838 79744
rect 176382 78704 176438 78713
rect 176382 78639 176438 78648
rect 176488 77294 176516 79630
rect 176580 77897 176608 79648
rect 176658 79384 176714 79393
rect 176658 79319 176714 79328
rect 176566 77888 176622 77897
rect 176566 77823 176622 77832
rect 176396 77266 176516 77294
rect 176292 24132 176344 24138
rect 176292 24074 176344 24080
rect 176396 18698 176424 77266
rect 176566 75712 176622 75721
rect 176566 75647 176622 75656
rect 176476 73772 176528 73778
rect 176476 73714 176528 73720
rect 176384 18692 176436 18698
rect 176384 18634 176436 18640
rect 176488 8974 176516 73714
rect 176580 10334 176608 75647
rect 176672 32434 176700 79319
rect 176764 79082 176792 79716
rect 176902 79642 176930 80036
rect 176856 79614 176930 79642
rect 176994 79642 177022 80036
rect 177086 79898 177114 80036
rect 177074 79892 177126 79898
rect 177074 79834 177126 79840
rect 177178 79778 177206 80036
rect 177270 79830 177298 80036
rect 177362 79971 177390 80036
rect 177348 79962 177404 79971
rect 177348 79897 177404 79906
rect 177132 79750 177206 79778
rect 177258 79824 177310 79830
rect 177258 79766 177310 79772
rect 176994 79614 177068 79642
rect 176752 79076 176804 79082
rect 176752 79018 176804 79024
rect 176856 70394 176884 79614
rect 176936 79484 176988 79490
rect 176936 79426 176988 79432
rect 176764 70366 176884 70394
rect 176764 68542 176792 70366
rect 176948 69630 176976 79426
rect 177040 78674 177068 79614
rect 177028 78668 177080 78674
rect 177028 78610 177080 78616
rect 177040 77314 177068 78610
rect 177028 77308 177080 77314
rect 177028 77250 177080 77256
rect 176936 69624 176988 69630
rect 176936 69566 176988 69572
rect 176752 68536 176804 68542
rect 176752 68478 176804 68484
rect 177132 66094 177160 79750
rect 177362 79744 177390 79897
rect 177454 79880 177482 80036
rect 177546 79948 177574 80036
rect 177546 79937 177620 79948
rect 177868 79937 177896 80038
rect 177948 80028 178000 80034
rect 177948 79970 178000 79976
rect 178040 80028 178092 80034
rect 178040 79970 178092 79976
rect 177546 79928 177634 79937
rect 177546 79920 177578 79928
rect 177454 79852 177528 79880
rect 177854 79928 177910 79937
rect 177634 79886 177712 79914
rect 177578 79863 177634 79872
rect 177500 79801 177528 79852
rect 177486 79792 177542 79801
rect 177362 79716 177436 79744
rect 177542 79750 177620 79778
rect 177486 79727 177542 79736
rect 177408 79676 177436 79716
rect 177302 79656 177358 79665
rect 177408 79648 177528 79676
rect 177302 79591 177358 79600
rect 177212 79076 177264 79082
rect 177212 79018 177264 79024
rect 177224 76430 177252 79018
rect 177212 76424 177264 76430
rect 177212 76366 177264 76372
rect 177224 75954 177252 76366
rect 177212 75948 177264 75954
rect 177212 75890 177264 75896
rect 177316 67634 177344 79591
rect 177396 79416 177448 79422
rect 177396 79358 177448 79364
rect 177408 78470 177436 79358
rect 177396 78464 177448 78470
rect 177396 78406 177448 78412
rect 177316 67606 177436 67634
rect 177120 66088 177172 66094
rect 177120 66030 177172 66036
rect 177408 64874 177436 67606
rect 177316 64846 177436 64874
rect 176660 32428 176712 32434
rect 176660 32370 176712 32376
rect 177316 31074 177344 64846
rect 177500 51746 177528 79648
rect 177592 76673 177620 79750
rect 177684 77625 177712 79886
rect 177764 79892 177816 79898
rect 177854 79863 177910 79872
rect 177764 79834 177816 79840
rect 177670 77616 177726 77625
rect 177670 77551 177726 77560
rect 177776 77353 177804 79834
rect 177856 79824 177908 79830
rect 177856 79766 177908 79772
rect 177868 78169 177896 79766
rect 177960 78849 177988 79970
rect 178052 79354 178080 79970
rect 178144 79626 178172 80106
rect 178222 79792 178278 79801
rect 178222 79727 178278 79736
rect 178132 79620 178184 79626
rect 178132 79562 178184 79568
rect 178236 79490 178264 79727
rect 178328 79558 178356 80174
rect 178316 79552 178368 79558
rect 178316 79494 178368 79500
rect 178224 79484 178276 79490
rect 178224 79426 178276 79432
rect 178040 79348 178092 79354
rect 178040 79290 178092 79296
rect 178420 79150 178448 80679
rect 183704 80702 183836 80708
rect 183652 80650 183704 80656
rect 183836 80650 183888 80656
rect 186424 80510 186452 80854
rect 186412 80504 186464 80510
rect 186412 80446 186464 80452
rect 183742 80336 183798 80345
rect 183742 80271 183798 80280
rect 178684 79960 178736 79966
rect 178684 79902 178736 79908
rect 180890 79928 180946 79937
rect 178696 79257 178724 79902
rect 180890 79863 180946 79872
rect 180062 79656 180118 79665
rect 180062 79591 180118 79600
rect 178682 79248 178738 79257
rect 178682 79183 178738 79192
rect 178408 79144 178460 79150
rect 178408 79086 178460 79092
rect 178040 78940 178092 78946
rect 178040 78882 178092 78888
rect 179328 78940 179380 78946
rect 179328 78882 179380 78888
rect 177946 78840 178002 78849
rect 177946 78775 178002 78784
rect 177854 78160 177910 78169
rect 177854 78095 177910 78104
rect 177762 77344 177818 77353
rect 177672 77308 177724 77314
rect 177762 77279 177818 77288
rect 177672 77250 177724 77256
rect 177578 76664 177634 76673
rect 177578 76599 177634 76608
rect 177684 76514 177712 77250
rect 177592 76486 177712 76514
rect 177488 51740 177540 51746
rect 177488 51682 177540 51688
rect 177592 44878 177620 76486
rect 177672 75948 177724 75954
rect 177672 75890 177724 75896
rect 177580 44872 177632 44878
rect 177580 44814 177632 44820
rect 177684 36582 177712 75890
rect 177868 64874 177896 78095
rect 177946 77344 178002 77353
rect 177946 77279 178002 77288
rect 177776 64846 177896 64874
rect 177672 36576 177724 36582
rect 177672 36518 177724 36524
rect 177776 35222 177804 64846
rect 177764 35216 177816 35222
rect 177764 35158 177816 35164
rect 177304 31068 177356 31074
rect 177304 31010 177356 31016
rect 177960 18630 177988 77279
rect 177948 18624 178000 18630
rect 177948 18566 178000 18572
rect 178052 16574 178080 78882
rect 178684 78804 178736 78810
rect 178684 78746 178736 78752
rect 178406 72448 178462 72457
rect 178406 72383 178462 72392
rect 178420 72350 178448 72383
rect 178408 72344 178460 72350
rect 178408 72286 178460 72292
rect 178052 16546 178632 16574
rect 176568 10328 176620 10334
rect 176568 10270 176620 10276
rect 176476 8968 176528 8974
rect 176476 8910 176528 8916
rect 175188 4820 175240 4826
rect 175188 4762 175240 4768
rect 174268 3800 174320 3806
rect 174268 3742 174320 3748
rect 171968 3664 172020 3670
rect 171968 3606 172020 3612
rect 171876 3596 171928 3602
rect 171876 3538 171928 3544
rect 171784 3528 171836 3534
rect 171784 3470 171836 3476
rect 171980 480 172008 3606
rect 173164 3528 173216 3534
rect 173164 3470 173216 3476
rect 173176 480 173204 3470
rect 174280 480 174308 3742
rect 177856 3596 177908 3602
rect 177856 3538 177908 3544
rect 175464 3460 175516 3466
rect 175464 3402 175516 3408
rect 175476 480 175504 3402
rect 176660 3392 176712 3398
rect 176660 3334 176712 3340
rect 176672 480 176700 3334
rect 177868 480 177896 3538
rect 156574 354 156686 480
rect 156156 326 156686 354
rect 156574 -960 156686 326
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 178604 354 178632 16546
rect 178696 3874 178724 78746
rect 179340 78606 179368 78882
rect 179972 78872 180024 78878
rect 179972 78814 180024 78820
rect 180076 78826 180104 79591
rect 180904 79393 180932 79863
rect 180890 79384 180946 79393
rect 180890 79319 180946 79328
rect 181904 79348 181956 79354
rect 181904 79290 181956 79296
rect 180156 79144 180208 79150
rect 180156 79086 180208 79092
rect 180168 79014 180196 79086
rect 180156 79008 180208 79014
rect 180156 78950 180208 78956
rect 178960 78600 179012 78606
rect 178960 78542 179012 78548
rect 179328 78600 179380 78606
rect 179328 78542 179380 78548
rect 178776 77648 178828 77654
rect 178776 77590 178828 77596
rect 178788 14618 178816 77590
rect 178972 77489 179000 78542
rect 179984 78470 180012 78814
rect 180076 78798 180196 78826
rect 179972 78464 180024 78470
rect 179972 78406 180024 78412
rect 178958 77480 179014 77489
rect 178958 77415 179014 77424
rect 180062 76664 180118 76673
rect 180062 76599 180118 76608
rect 179326 76392 179382 76401
rect 179326 76327 179382 76336
rect 179234 75440 179290 75449
rect 179234 75375 179290 75384
rect 178868 74656 178920 74662
rect 178868 74598 178920 74604
rect 178880 21418 178908 74598
rect 178868 21412 178920 21418
rect 178868 21354 178920 21360
rect 178776 14612 178828 14618
rect 178776 14554 178828 14560
rect 178684 3868 178736 3874
rect 178684 3810 178736 3816
rect 179248 3738 179276 75375
rect 179236 3732 179288 3738
rect 179236 3674 179288 3680
rect 179340 3534 179368 76327
rect 179694 73128 179750 73137
rect 179694 73063 179750 73072
rect 179708 72418 179736 73063
rect 179696 72412 179748 72418
rect 179696 72354 179748 72360
rect 179420 69556 179472 69562
rect 179420 69498 179472 69504
rect 179432 16574 179460 69498
rect 179432 16546 180012 16574
rect 179328 3528 179380 3534
rect 179328 3470 179380 3476
rect 179984 3482 180012 16546
rect 180076 3618 180104 76599
rect 180168 4962 180196 78798
rect 180708 77852 180760 77858
rect 180708 77794 180760 77800
rect 180430 77752 180486 77761
rect 180430 77687 180486 77696
rect 180340 77512 180392 77518
rect 180340 77454 180392 77460
rect 180246 73536 180302 73545
rect 180246 73471 180302 73480
rect 180156 4956 180208 4962
rect 180156 4898 180208 4904
rect 180260 3738 180288 73471
rect 180352 73154 180380 77454
rect 180444 77353 180472 77687
rect 180430 77344 180486 77353
rect 180430 77279 180486 77288
rect 180352 73126 180472 73154
rect 180340 72820 180392 72826
rect 180340 72762 180392 72768
rect 180352 4078 180380 72762
rect 180444 17474 180472 73126
rect 180616 72412 180668 72418
rect 180616 72354 180668 72360
rect 180628 71806 180656 72354
rect 180616 71800 180668 71806
rect 180616 71742 180668 71748
rect 180720 68610 180748 77794
rect 181628 77784 181680 77790
rect 181628 77726 181680 77732
rect 181352 76628 181404 76634
rect 181352 76570 181404 76576
rect 180800 75676 180852 75682
rect 180800 75618 180852 75624
rect 180708 68604 180760 68610
rect 180708 68546 180760 68552
rect 180432 17468 180484 17474
rect 180432 17410 180484 17416
rect 180812 16574 180840 75618
rect 181258 73128 181314 73137
rect 181258 73063 181314 73072
rect 181272 72282 181300 73063
rect 181260 72276 181312 72282
rect 181260 72218 181312 72224
rect 181272 71874 181300 72218
rect 181260 71868 181312 71874
rect 181260 71810 181312 71816
rect 181364 70394 181392 76570
rect 181536 75608 181588 75614
rect 181536 75550 181588 75556
rect 181364 70366 181484 70394
rect 181168 69420 181220 69426
rect 181168 69362 181220 69368
rect 181180 66201 181208 69362
rect 181166 66192 181222 66201
rect 181166 66127 181222 66136
rect 180812 16546 181024 16574
rect 180340 4072 180392 4078
rect 180340 4014 180392 4020
rect 180248 3732 180300 3738
rect 180248 3674 180300 3680
rect 180076 3590 180380 3618
rect 179984 3454 180288 3482
rect 180260 480 180288 3454
rect 180352 3398 180380 3590
rect 180340 3392 180392 3398
rect 180340 3334 180392 3340
rect 179022 354 179134 480
rect 178604 326 179134 354
rect 179022 -960 179134 326
rect 180218 -960 180330 480
rect 180996 354 181024 16546
rect 181456 4010 181484 70366
rect 181444 4004 181496 4010
rect 181444 3946 181496 3952
rect 181548 3194 181576 75550
rect 181640 25702 181668 77726
rect 181916 77722 181944 79290
rect 183756 79150 183784 80271
rect 186516 80102 186544 80951
rect 187160 80374 187188 80951
rect 187148 80368 187200 80374
rect 187148 80310 187200 80316
rect 186504 80096 186556 80102
rect 186504 80038 186556 80044
rect 183744 79144 183796 79150
rect 183744 79086 183796 79092
rect 187436 78713 187464 80951
rect 188172 80850 188200 81194
rect 188160 80844 188212 80850
rect 188160 80786 188212 80792
rect 188264 80782 188292 194890
rect 188356 143410 188384 201719
rect 188448 193186 188476 259655
rect 189172 195016 189224 195022
rect 189172 194958 189224 194964
rect 189080 194880 189132 194886
rect 189080 194822 189132 194828
rect 188436 193180 188488 193186
rect 188436 193122 188488 193128
rect 188436 178084 188488 178090
rect 188436 178026 188488 178032
rect 188448 144226 188476 178026
rect 188528 145988 188580 145994
rect 188528 145930 188580 145936
rect 188436 144220 188488 144226
rect 188436 144162 188488 144168
rect 188344 143404 188396 143410
rect 188344 143346 188396 143352
rect 188252 80776 188304 80782
rect 188252 80718 188304 80724
rect 187422 78704 187478 78713
rect 187422 78639 187478 78648
rect 184478 78568 184534 78577
rect 184478 78503 184534 78512
rect 186410 78568 186466 78577
rect 186410 78503 186466 78512
rect 187422 78568 187478 78577
rect 187422 78503 187478 78512
rect 183468 78464 183520 78470
rect 183468 78406 183520 78412
rect 183008 78328 183060 78334
rect 183008 78270 183060 78276
rect 182824 77920 182876 77926
rect 182824 77862 182876 77868
rect 181904 77716 181956 77722
rect 181904 77658 181956 77664
rect 181996 72820 182048 72826
rect 181996 72762 182048 72768
rect 182008 72350 182036 72762
rect 181996 72344 182048 72350
rect 181996 72286 182048 72292
rect 182008 64874 182036 72286
rect 182180 68604 182232 68610
rect 182180 68546 182232 68552
rect 182008 64846 182128 64874
rect 181628 25696 181680 25702
rect 181628 25638 181680 25644
rect 182100 3670 182128 64846
rect 182088 3664 182140 3670
rect 182088 3606 182140 3612
rect 181536 3188 181588 3194
rect 181536 3130 181588 3136
rect 181414 354 181526 480
rect 180996 326 181526 354
rect 182192 354 182220 68546
rect 182836 24274 182864 77862
rect 183020 77858 183048 78270
rect 183008 77852 183060 77858
rect 183008 77794 183060 77800
rect 183282 77072 183338 77081
rect 183282 77007 183338 77016
rect 183296 76673 183324 77007
rect 183282 76664 183338 76673
rect 183282 76599 183338 76608
rect 182824 24268 182876 24274
rect 182824 24210 182876 24216
rect 183480 3806 183508 78406
rect 183560 78260 183612 78266
rect 183560 78202 183612 78208
rect 183572 71738 183600 78202
rect 184492 76974 184520 78503
rect 184480 76968 184532 76974
rect 184480 76910 184532 76916
rect 184204 76900 184256 76906
rect 184204 76842 184256 76848
rect 184216 76362 184244 76842
rect 184204 76356 184256 76362
rect 184204 76298 184256 76304
rect 184492 76022 184520 76910
rect 184480 76016 184532 76022
rect 184480 75958 184532 75964
rect 183744 73568 183796 73574
rect 183744 73510 183796 73516
rect 183560 71732 183612 71738
rect 183560 71674 183612 71680
rect 183560 64184 183612 64190
rect 183560 64126 183612 64132
rect 183572 16574 183600 64126
rect 183756 61577 183784 73510
rect 186424 70922 186452 78503
rect 187436 77110 187464 78503
rect 187424 77104 187476 77110
rect 187424 77046 187476 77052
rect 187700 75472 187752 75478
rect 187700 75414 187752 75420
rect 186412 70916 186464 70922
rect 186412 70858 186464 70864
rect 185584 69760 185636 69766
rect 185584 69702 185636 69708
rect 183834 69048 183890 69057
rect 183834 68983 183890 68992
rect 183848 68746 183876 68983
rect 183836 68740 183888 68746
rect 183836 68682 183888 68688
rect 183742 61568 183798 61577
rect 183742 61503 183798 61512
rect 183572 16546 183784 16574
rect 183468 3800 183520 3806
rect 183468 3742 183520 3748
rect 183756 480 183784 16546
rect 185596 3398 185624 69702
rect 186320 58812 186372 58818
rect 186320 58754 186372 58760
rect 186332 16574 186360 58754
rect 187712 16574 187740 75414
rect 188540 74390 188568 145930
rect 188804 77104 188856 77110
rect 188804 77046 188856 77052
rect 188816 75954 188844 77046
rect 188804 75948 188856 75954
rect 188804 75890 188856 75896
rect 188528 74384 188580 74390
rect 188528 74326 188580 74332
rect 188250 68776 188306 68785
rect 188250 68711 188306 68720
rect 188264 68678 188292 68711
rect 188252 68672 188304 68678
rect 188252 68614 188304 68620
rect 188264 67726 188292 68614
rect 188252 67720 188304 67726
rect 188252 67662 188304 67668
rect 188066 66192 188122 66201
rect 188066 66127 188068 66136
rect 188120 66127 188122 66136
rect 188068 66098 188120 66104
rect 188618 65104 188674 65113
rect 188618 65039 188674 65048
rect 188632 65006 188660 65039
rect 188620 65000 188672 65006
rect 188620 64942 188672 64948
rect 189092 63345 189120 194822
rect 189184 67590 189212 194958
rect 189276 143138 189304 263638
rect 189632 262880 189684 262886
rect 189632 262822 189684 262828
rect 189540 260500 189592 260506
rect 189540 260442 189592 260448
rect 189354 260264 189410 260273
rect 189354 260199 189410 260208
rect 189448 260228 189500 260234
rect 189264 143132 189316 143138
rect 189264 143074 189316 143080
rect 189368 141438 189396 260199
rect 189448 260170 189500 260176
rect 189460 141642 189488 260170
rect 189552 143206 189580 260442
rect 189644 145518 189672 262822
rect 189816 260024 189868 260030
rect 189816 259966 189868 259972
rect 189724 196512 189776 196518
rect 189724 196454 189776 196460
rect 189632 145512 189684 145518
rect 189632 145454 189684 145460
rect 189632 143472 189684 143478
rect 189632 143414 189684 143420
rect 189540 143200 189592 143206
rect 189540 143142 189592 143148
rect 189448 141636 189500 141642
rect 189448 141578 189500 141584
rect 189356 141432 189408 141438
rect 189356 141374 189408 141380
rect 189356 140412 189408 140418
rect 189356 140354 189408 140360
rect 189262 139360 189318 139369
rect 189262 139295 189318 139304
rect 189172 67584 189224 67590
rect 189172 67526 189224 67532
rect 189184 66910 189212 67526
rect 189172 66904 189224 66910
rect 189172 66846 189224 66852
rect 189078 63336 189134 63345
rect 189078 63271 189134 63280
rect 189276 56273 189304 139295
rect 189368 60654 189396 140354
rect 189446 139088 189502 139097
rect 189446 139023 189502 139032
rect 189356 60648 189408 60654
rect 189460 60625 189488 139023
rect 189644 74497 189672 143414
rect 189736 80714 189764 196454
rect 189828 144838 189856 259966
rect 189908 259616 189960 259622
rect 189908 259558 189960 259564
rect 189920 145382 189948 259558
rect 190000 145648 190052 145654
rect 190000 145590 190052 145596
rect 189908 145376 189960 145382
rect 189908 145318 189960 145324
rect 189816 144832 189868 144838
rect 189816 144774 189868 144780
rect 189816 140344 189868 140350
rect 189816 140286 189868 140292
rect 189724 80708 189776 80714
rect 189724 80650 189776 80656
rect 189630 74488 189686 74497
rect 189630 74423 189686 74432
rect 189644 73817 189672 74423
rect 189630 73808 189686 73817
rect 189630 73743 189686 73752
rect 189828 72894 189856 140286
rect 189908 140208 189960 140214
rect 189908 140150 189960 140156
rect 189920 79422 189948 140150
rect 189908 79416 189960 79422
rect 189908 79358 189960 79364
rect 190012 73030 190040 145590
rect 190472 144430 190500 264998
rect 190920 263764 190972 263770
rect 190920 263706 190972 263712
rect 190828 262608 190880 262614
rect 190828 262550 190880 262556
rect 190552 197192 190604 197198
rect 190552 197134 190604 197140
rect 190460 144424 190512 144430
rect 190460 144366 190512 144372
rect 190000 73024 190052 73030
rect 190000 72966 190052 72972
rect 189816 72888 189868 72894
rect 189816 72830 189868 72836
rect 189722 68232 189778 68241
rect 189722 68167 189778 68176
rect 189356 60590 189408 60596
rect 189446 60616 189502 60625
rect 189368 60042 189396 60590
rect 189446 60551 189502 60560
rect 189630 60616 189686 60625
rect 189630 60551 189686 60560
rect 189644 60217 189672 60551
rect 189630 60208 189686 60217
rect 189630 60143 189686 60152
rect 189356 60036 189408 60042
rect 189356 59978 189408 59984
rect 189262 56264 189318 56273
rect 189262 56199 189318 56208
rect 189736 16574 189764 68167
rect 190460 62824 190512 62830
rect 190460 62766 190512 62772
rect 186332 16546 186912 16574
rect 187712 16546 188568 16574
rect 189736 16546 189856 16574
rect 186136 4072 186188 4078
rect 186136 4014 186188 4020
rect 185584 3392 185636 3398
rect 185584 3334 185636 3340
rect 184940 3188 184992 3194
rect 184940 3130 184992 3136
rect 184952 480 184980 3130
rect 186148 480 186176 4014
rect 182518 354 182630 480
rect 182192 326 182630 354
rect 181414 -960 181526 326
rect 182518 -960 182630 326
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 186884 354 186912 16546
rect 188540 480 188568 16546
rect 189828 4078 189856 16546
rect 189816 4072 189868 4078
rect 189816 4014 189868 4020
rect 189724 3392 189776 3398
rect 189724 3334 189776 3340
rect 189736 480 189764 3334
rect 187302 354 187414 480
rect 186884 326 187414 354
rect 187302 -960 187414 326
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190472 354 190500 62766
rect 190564 57905 190592 197134
rect 190736 195900 190788 195906
rect 190736 195842 190788 195848
rect 190644 195424 190696 195430
rect 190644 195366 190696 195372
rect 190656 75750 190684 195366
rect 190644 75744 190696 75750
rect 190644 75686 190696 75692
rect 190748 75002 190776 195842
rect 190840 144566 190868 262550
rect 190932 145450 190960 263706
rect 191748 262880 191800 262886
rect 191748 262822 191800 262828
rect 191760 262614 191788 262822
rect 191748 262608 191800 262614
rect 191748 262550 191800 262556
rect 192208 262472 192260 262478
rect 192208 262414 192260 262420
rect 191104 260432 191156 260438
rect 191104 260374 191156 260380
rect 191012 259684 191064 259690
rect 191012 259626 191064 259632
rect 190920 145444 190972 145450
rect 190920 145386 190972 145392
rect 191024 144634 191052 259626
rect 191012 144628 191064 144634
rect 191012 144570 191064 144576
rect 190828 144560 190880 144566
rect 190828 144502 190880 144508
rect 191116 144498 191144 260374
rect 191932 196988 191984 196994
rect 191932 196930 191984 196936
rect 191840 195356 191892 195362
rect 191840 195298 191892 195304
rect 191194 180840 191250 180849
rect 191194 180775 191250 180784
rect 191104 144492 191156 144498
rect 191104 144434 191156 144440
rect 190918 138816 190974 138825
rect 190918 138751 190974 138760
rect 190736 74996 190788 75002
rect 190736 74938 190788 74944
rect 190932 60489 190960 138751
rect 191102 138544 191158 138553
rect 191102 138479 191158 138488
rect 191116 71126 191144 138479
rect 191208 114481 191236 180775
rect 191286 146160 191342 146169
rect 191286 146095 191342 146104
rect 191300 140865 191328 146095
rect 191470 145752 191526 145761
rect 191470 145687 191526 145696
rect 191380 144900 191432 144906
rect 191380 144842 191432 144848
rect 191286 140856 191342 140865
rect 191286 140791 191342 140800
rect 191288 140276 191340 140282
rect 191288 140218 191340 140224
rect 191194 114472 191250 114481
rect 191194 114407 191250 114416
rect 191194 81968 191250 81977
rect 191194 81903 191250 81912
rect 191208 71194 191236 81903
rect 191300 79354 191328 140218
rect 191288 79348 191340 79354
rect 191288 79290 191340 79296
rect 191196 71188 191248 71194
rect 191196 71130 191248 71136
rect 191104 71120 191156 71126
rect 191104 71062 191156 71068
rect 191392 61849 191420 144842
rect 191484 77042 191512 145687
rect 191562 144800 191618 144809
rect 191562 144735 191618 144744
rect 191472 77036 191524 77042
rect 191472 76978 191524 76984
rect 191378 61840 191434 61849
rect 191378 61775 191434 61784
rect 190918 60480 190974 60489
rect 190918 60415 190974 60424
rect 190550 57896 190606 57905
rect 190550 57831 190606 57840
rect 191576 52193 191604 144735
rect 191748 77036 191800 77042
rect 191748 76978 191800 76984
rect 191760 76634 191788 76978
rect 191748 76628 191800 76634
rect 191748 76570 191800 76576
rect 191746 60480 191802 60489
rect 191746 60415 191802 60424
rect 191760 60081 191788 60415
rect 191746 60072 191802 60081
rect 191746 60007 191802 60016
rect 191746 57896 191802 57905
rect 191746 57831 191802 57840
rect 191760 57497 191788 57831
rect 191746 57488 191802 57497
rect 191746 57423 191802 57432
rect 191852 55049 191880 195298
rect 191944 69698 191972 196930
rect 192116 196648 192168 196654
rect 192116 196590 192168 196596
rect 192024 195288 192076 195294
rect 192024 195230 192076 195236
rect 191932 69692 191984 69698
rect 191932 69634 191984 69640
rect 192036 63481 192064 195230
rect 192128 70446 192156 196590
rect 192220 141846 192248 262414
rect 192312 146266 192340 265610
rect 196440 265600 196492 265606
rect 196440 265542 196492 265548
rect 193864 265532 193916 265538
rect 193864 265474 193916 265480
rect 193588 265328 193640 265334
rect 193588 265270 193640 265276
rect 193220 265124 193272 265130
rect 193220 265066 193272 265072
rect 192484 262744 192536 262750
rect 192484 262686 192536 262692
rect 192392 260364 192444 260370
rect 192392 260306 192444 260312
rect 192300 146260 192352 146266
rect 192300 146202 192352 146208
rect 192300 145784 192352 145790
rect 192300 145726 192352 145732
rect 192208 141840 192260 141846
rect 192208 141782 192260 141788
rect 192208 140344 192260 140350
rect 192208 140286 192260 140292
rect 192116 70440 192168 70446
rect 192116 70382 192168 70388
rect 192116 69692 192168 69698
rect 192116 69634 192168 69640
rect 192022 63472 192078 63481
rect 192022 63407 192078 63416
rect 192128 59129 192156 69634
rect 192114 59120 192170 59129
rect 192114 59055 192170 59064
rect 191838 55040 191894 55049
rect 191838 54975 191894 54984
rect 191852 54777 191880 54975
rect 191838 54768 191894 54777
rect 191838 54703 191894 54712
rect 191562 52184 191618 52193
rect 191562 52119 191618 52128
rect 192220 50561 192248 140286
rect 192312 74526 192340 145726
rect 192404 142050 192432 260306
rect 192496 144770 192524 262686
rect 192668 261384 192720 261390
rect 192668 261326 192720 261332
rect 192576 261248 192628 261254
rect 192576 261190 192628 261196
rect 192588 146130 192616 261190
rect 192680 149598 192708 261326
rect 192668 149592 192720 149598
rect 192668 149534 192720 149540
rect 192852 148232 192904 148238
rect 192852 148174 192904 148180
rect 192576 146124 192628 146130
rect 192576 146066 192628 146072
rect 192760 145852 192812 145858
rect 192760 145794 192812 145800
rect 192484 144764 192536 144770
rect 192484 144706 192536 144712
rect 192392 142044 192444 142050
rect 192392 141986 192444 141992
rect 192668 140140 192720 140146
rect 192668 140082 192720 140088
rect 192576 140072 192628 140078
rect 192576 140014 192628 140020
rect 192300 74520 192352 74526
rect 192300 74462 192352 74468
rect 192588 71058 192616 140014
rect 192680 75138 192708 140082
rect 192668 75132 192720 75138
rect 192668 75074 192720 75080
rect 192576 71052 192628 71058
rect 192576 70994 192628 71000
rect 192772 70854 192800 145794
rect 192760 70848 192812 70854
rect 192760 70790 192812 70796
rect 192300 70440 192352 70446
rect 192300 70382 192352 70388
rect 192312 66230 192340 70382
rect 192300 66224 192352 66230
rect 192300 66166 192352 66172
rect 192864 53417 192892 148174
rect 193232 145625 193260 265066
rect 193404 196784 193456 196790
rect 193404 196726 193456 196732
rect 193312 195492 193364 195498
rect 193312 195434 193364 195440
rect 193218 145616 193274 145625
rect 193218 145551 193274 145560
rect 193220 140684 193272 140690
rect 193220 140626 193272 140632
rect 193232 140593 193260 140626
rect 193218 140584 193274 140593
rect 193218 140519 193274 140528
rect 193128 66224 193180 66230
rect 193128 66166 193180 66172
rect 193140 65550 193168 66166
rect 193128 65544 193180 65550
rect 193128 65486 193180 65492
rect 193126 63472 193182 63481
rect 193126 63407 193182 63416
rect 193140 63209 193168 63407
rect 193126 63200 193182 63209
rect 193126 63135 193182 63144
rect 193126 59120 193182 59129
rect 193126 59055 193182 59064
rect 193140 58857 193168 59055
rect 193126 58848 193182 58857
rect 193126 58783 193182 58792
rect 192850 53408 192906 53417
rect 192850 53343 192906 53352
rect 193324 50969 193352 195434
rect 193416 63510 193444 196726
rect 193496 196580 193548 196586
rect 193496 196522 193548 196528
rect 193508 71262 193536 196522
rect 193600 139738 193628 265270
rect 193772 264988 193824 264994
rect 193772 264930 193824 264936
rect 193680 262676 193732 262682
rect 193680 262618 193732 262624
rect 193692 141506 193720 262618
rect 193784 144294 193812 264930
rect 193876 144702 193904 265474
rect 196256 265464 196308 265470
rect 196256 265406 196308 265412
rect 195152 265192 195204 265198
rect 195152 265134 195204 265140
rect 195060 259480 195112 259486
rect 195060 259422 195112 259428
rect 194692 197056 194744 197062
rect 194692 196998 194744 197004
rect 194140 195764 194192 195770
rect 194140 195706 194192 195712
rect 193956 147076 194008 147082
rect 193956 147018 194008 147024
rect 193864 144696 193916 144702
rect 193864 144638 193916 144644
rect 193772 144288 193824 144294
rect 193772 144230 193824 144236
rect 193864 142112 193916 142118
rect 193864 142054 193916 142060
rect 193680 141500 193732 141506
rect 193680 141442 193732 141448
rect 193680 140752 193732 140758
rect 193678 140720 193680 140729
rect 193732 140720 193734 140729
rect 193678 140655 193734 140664
rect 193588 139732 193640 139738
rect 193588 139674 193640 139680
rect 193678 138952 193734 138961
rect 193678 138887 193734 138896
rect 193586 78568 193642 78577
rect 193586 78503 193588 78512
rect 193640 78503 193642 78512
rect 193588 78474 193640 78480
rect 193496 71256 193548 71262
rect 193496 71198 193548 71204
rect 193404 63504 193456 63510
rect 193404 63446 193456 63452
rect 193416 62830 193444 63446
rect 193404 62824 193456 62830
rect 193404 62766 193456 62772
rect 193692 61577 193720 138887
rect 193876 71466 193904 142054
rect 193968 79558 193996 147018
rect 194046 139360 194102 139369
rect 194046 139295 194102 139304
rect 194060 80442 194088 139295
rect 194048 80436 194100 80442
rect 194048 80378 194100 80384
rect 193956 79552 194008 79558
rect 193956 79494 194008 79500
rect 193864 71460 193916 71466
rect 193864 71402 193916 71408
rect 193862 66872 193918 66881
rect 193862 66807 193918 66816
rect 193678 61568 193734 61577
rect 193678 61503 193734 61512
rect 193402 59936 193458 59945
rect 193402 59871 193458 59880
rect 193310 50960 193366 50969
rect 193310 50895 193366 50904
rect 192206 50552 192262 50561
rect 192206 50487 192262 50496
rect 191840 50448 191892 50454
rect 191840 50390 191892 50396
rect 191852 16574 191880 50390
rect 193416 16574 193444 59871
rect 191852 16546 192064 16574
rect 193416 16546 193812 16574
rect 192036 480 192064 16546
rect 193220 4072 193272 4078
rect 193220 4014 193272 4020
rect 193232 480 193260 4014
rect 193784 3482 193812 16546
rect 193876 4078 193904 66807
rect 194152 57866 194180 195706
rect 194600 195560 194652 195566
rect 194600 195502 194652 195508
rect 194324 145716 194376 145722
rect 194324 145658 194376 145664
rect 194232 141976 194284 141982
rect 194232 141918 194284 141924
rect 194140 57860 194192 57866
rect 194140 57802 194192 57808
rect 194244 52057 194272 141918
rect 194336 71670 194364 145658
rect 194508 79552 194560 79558
rect 194508 79494 194560 79500
rect 194520 79354 194548 79494
rect 194508 79348 194560 79354
rect 194508 79290 194560 79296
rect 194508 78532 194560 78538
rect 194508 78474 194560 78480
rect 194520 77314 194548 78474
rect 194508 77308 194560 77314
rect 194508 77250 194560 77256
rect 194324 71664 194376 71670
rect 194324 71606 194376 71612
rect 194508 57860 194560 57866
rect 194508 57802 194560 57808
rect 194520 57322 194548 57802
rect 194508 57316 194560 57322
rect 194508 57258 194560 57264
rect 194612 55185 194640 195502
rect 194704 59265 194732 196998
rect 194876 196852 194928 196858
rect 194876 196794 194928 196800
rect 194784 193044 194836 193050
rect 194784 192986 194836 192992
rect 194690 59256 194746 59265
rect 194690 59191 194746 59200
rect 194796 57769 194824 192986
rect 194888 64870 194916 196794
rect 194968 147552 195020 147558
rect 194968 147494 195020 147500
rect 194980 73710 195008 147494
rect 195072 143342 195100 259422
rect 195164 146033 195192 265134
rect 195612 199300 195664 199306
rect 195612 199242 195664 199248
rect 195244 186720 195296 186726
rect 195244 186662 195296 186668
rect 195150 146024 195206 146033
rect 195150 145959 195206 145968
rect 195060 143336 195112 143342
rect 195060 143278 195112 143284
rect 195152 141908 195204 141914
rect 195152 141850 195204 141856
rect 194968 73704 195020 73710
rect 194968 73646 195020 73652
rect 195164 71602 195192 141850
rect 195256 78946 195284 186662
rect 195336 147484 195388 147490
rect 195336 147426 195388 147432
rect 195348 81297 195376 147426
rect 195520 145920 195572 145926
rect 195520 145862 195572 145868
rect 195428 140480 195480 140486
rect 195428 140422 195480 140428
rect 195334 81288 195390 81297
rect 195334 81223 195390 81232
rect 195244 78940 195296 78946
rect 195244 78882 195296 78888
rect 195256 78441 195284 78882
rect 195440 78742 195468 140422
rect 195428 78736 195480 78742
rect 195428 78678 195480 78684
rect 195242 78432 195298 78441
rect 195242 78367 195298 78376
rect 195532 75818 195560 145862
rect 195624 139505 195652 199242
rect 196072 197124 196124 197130
rect 196072 197066 196124 197072
rect 195980 192500 196032 192506
rect 195980 192442 196032 192448
rect 195610 139496 195666 139505
rect 195610 139431 195666 139440
rect 195520 75812 195572 75818
rect 195520 75754 195572 75760
rect 195152 71596 195204 71602
rect 195152 71538 195204 71544
rect 195150 70408 195206 70417
rect 195150 70343 195206 70352
rect 195164 69562 195192 70343
rect 195152 69556 195204 69562
rect 195152 69498 195204 69504
rect 195164 69086 195192 69498
rect 195152 69080 195204 69086
rect 195152 69022 195204 69028
rect 194876 64864 194928 64870
rect 194876 64806 194928 64812
rect 194888 64258 194916 64806
rect 194876 64252 194928 64258
rect 194876 64194 194928 64200
rect 195058 59256 195114 59265
rect 195058 59191 195114 59200
rect 195072 58721 195100 59191
rect 195058 58712 195114 58721
rect 195058 58647 195114 58656
rect 194782 57760 194838 57769
rect 194782 57695 194838 57704
rect 195058 57760 195114 57769
rect 195058 57695 195114 57704
rect 195072 57361 195100 57695
rect 195058 57352 195114 57361
rect 195058 57287 195114 57296
rect 194598 55176 194654 55185
rect 194598 55111 194654 55120
rect 194612 54641 194640 55111
rect 194598 54632 194654 54641
rect 194598 54567 194654 54576
rect 195992 53689 196020 192442
rect 196084 61713 196112 197066
rect 196164 196716 196216 196722
rect 196164 196658 196216 196664
rect 196176 66065 196204 196658
rect 196268 139806 196296 265406
rect 196348 260908 196400 260914
rect 196348 260850 196400 260856
rect 196360 141778 196388 260850
rect 196452 146878 196480 265542
rect 197728 265396 197780 265402
rect 197728 265338 197780 265344
rect 197636 265260 197688 265266
rect 197636 265202 197688 265208
rect 196532 262404 196584 262410
rect 196532 262346 196584 262352
rect 196440 146872 196492 146878
rect 196440 146814 196492 146820
rect 196544 146198 196572 262346
rect 196624 261044 196676 261050
rect 196624 260986 196676 260992
rect 196532 146192 196584 146198
rect 196532 146134 196584 146140
rect 196636 146062 196664 260986
rect 196716 260976 196768 260982
rect 196716 260918 196768 260924
rect 196728 147626 196756 260918
rect 197544 197328 197596 197334
rect 197544 197270 197596 197276
rect 197452 196920 197504 196926
rect 197452 196862 197504 196868
rect 197360 192568 197412 192574
rect 197360 192510 197412 192516
rect 196808 184068 196860 184074
rect 196808 184010 196860 184016
rect 196820 147801 196848 184010
rect 196900 148776 196952 148782
rect 196900 148718 196952 148724
rect 196806 147792 196862 147801
rect 196806 147727 196862 147736
rect 196716 147620 196768 147626
rect 196716 147562 196768 147568
rect 196624 146056 196676 146062
rect 196624 145998 196676 146004
rect 196808 143268 196860 143274
rect 196808 143210 196860 143216
rect 196348 141772 196400 141778
rect 196348 141714 196400 141720
rect 196716 140004 196768 140010
rect 196716 139946 196768 139952
rect 196256 139800 196308 139806
rect 196256 139742 196308 139748
rect 196530 138680 196586 138689
rect 196530 138615 196586 138624
rect 196544 69970 196572 138615
rect 196728 77246 196756 139946
rect 196716 77240 196768 77246
rect 196716 77182 196768 77188
rect 196820 71534 196848 143210
rect 196808 71528 196860 71534
rect 196808 71470 196860 71476
rect 196912 71398 196940 148718
rect 196992 147416 197044 147422
rect 196992 147358 197044 147364
rect 197004 81161 197032 147358
rect 197084 147348 197136 147354
rect 197084 147290 197136 147296
rect 196990 81152 197046 81161
rect 196990 81087 197046 81096
rect 196900 71392 196952 71398
rect 196900 71334 196952 71340
rect 196532 69964 196584 69970
rect 196532 69906 196584 69912
rect 196624 69624 196676 69630
rect 196624 69566 196676 69572
rect 196162 66056 196218 66065
rect 196162 65991 196218 66000
rect 196438 66056 196494 66065
rect 196438 65991 196494 66000
rect 196452 65521 196480 65991
rect 196438 65512 196494 65521
rect 196438 65447 196494 65456
rect 196070 61704 196126 61713
rect 196070 61639 196126 61648
rect 195978 53680 196034 53689
rect 195978 53615 196034 53624
rect 195992 53281 196020 53615
rect 195978 53272 196034 53281
rect 195978 53207 196034 53216
rect 194230 52048 194286 52057
rect 194230 51983 194286 51992
rect 194598 47560 194654 47569
rect 194598 47495 194654 47504
rect 194612 16574 194640 47495
rect 194612 16546 195192 16574
rect 193864 4072 193916 4078
rect 193864 4014 193916 4020
rect 193784 3454 194456 3482
rect 194428 480 194456 3454
rect 190798 354 190910 480
rect 190472 326 190910 354
rect 190798 -960 190910 326
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195164 354 195192 16546
rect 196636 4146 196664 69566
rect 197096 46753 197124 147290
rect 197082 46744 197138 46753
rect 197082 46679 197138 46688
rect 197372 45529 197400 192510
rect 197464 60874 197492 196862
rect 197556 74534 197584 197270
rect 197648 139670 197676 265202
rect 197740 141574 197768 265338
rect 218072 262886 218100 703582
rect 218808 703474 218836 703582
rect 218950 703520 219062 704960
rect 234632 703582 235028 703610
rect 218992 703474 219020 703520
rect 218808 703446 219020 703474
rect 234632 273970 234660 703582
rect 235000 703474 235028 703582
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 299492 703582 299980 703610
rect 235184 703474 235212 703520
rect 235000 703446 235212 703474
rect 267660 699718 267688 703520
rect 283852 700534 283880 703520
rect 283840 700528 283892 700534
rect 283840 700470 283892 700476
rect 265624 699712 265676 699718
rect 265624 699654 265676 699660
rect 267648 699712 267700 699718
rect 267648 699654 267700 699660
rect 265636 276729 265664 699654
rect 265622 276720 265678 276729
rect 265622 276655 265678 276664
rect 234620 273964 234672 273970
rect 234620 273906 234672 273912
rect 299492 264246 299520 703582
rect 299952 703474 299980 703582
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 412652 703582 413508 703610
rect 300136 703474 300164 703520
rect 299952 703446 300164 703474
rect 332520 700398 332548 703520
rect 348804 702434 348832 703520
rect 364996 702434 365024 703520
rect 347792 702406 348832 702434
rect 364352 702406 365024 702434
rect 332508 700392 332560 700398
rect 332508 700334 332560 700340
rect 299480 264240 299532 264246
rect 299480 264182 299532 264188
rect 347792 263498 347820 702406
rect 364352 275330 364380 702406
rect 397472 699718 397500 703520
rect 396724 699712 396776 699718
rect 396724 699654 396776 699660
rect 397460 699712 397512 699718
rect 397460 699654 397512 699660
rect 396736 280838 396764 699654
rect 396724 280832 396776 280838
rect 396724 280774 396776 280780
rect 364340 275324 364392 275330
rect 364340 275266 364392 275272
rect 347780 263492 347832 263498
rect 347780 263434 347832 263440
rect 412652 262993 412680 703582
rect 413480 703474 413508 703582
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494072 703582 494652 703610
rect 413664 703474 413692 703520
rect 413480 703446 413692 703474
rect 429856 699718 429884 703520
rect 428464 699712 428516 699718
rect 428464 699654 428516 699660
rect 429844 699712 429896 699718
rect 429844 699654 429896 699660
rect 428476 271153 428504 699654
rect 462332 279478 462360 703520
rect 478524 702434 478552 703520
rect 477512 702406 478552 702434
rect 462320 279472 462372 279478
rect 462320 279414 462372 279420
rect 428462 271144 428518 271153
rect 428462 271079 428518 271088
rect 412638 262984 412694 262993
rect 412638 262919 412694 262928
rect 218060 262880 218112 262886
rect 477512 262857 477540 702406
rect 494072 269822 494100 703582
rect 494624 703474 494652 703582
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 494808 703474 494836 703520
rect 494624 703446 494836 703474
rect 525064 700392 525116 700398
rect 525064 700334 525116 700340
rect 494060 269816 494112 269822
rect 494060 269758 494112 269764
rect 525076 268394 525104 700334
rect 527192 278050 527220 703520
rect 543476 700330 543504 703520
rect 559668 700398 559696 703520
rect 559656 700392 559708 700398
rect 559656 700334 559708 700340
rect 543464 700324 543516 700330
rect 543464 700266 543516 700272
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683194 580212 683839
rect 580172 683188 580224 683194
rect 580172 683130 580224 683136
rect 580172 670744 580224 670750
rect 580170 670712 580172 670721
rect 580224 670712 580226 670721
rect 580170 670647 580226 670656
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580184 643142 580212 643991
rect 580172 643136 580224 643142
rect 580172 643078 580224 643084
rect 580170 630864 580226 630873
rect 580170 630799 580226 630808
rect 580184 630698 580212 630799
rect 580172 630692 580224 630698
rect 580172 630634 580224 630640
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580184 616894 580212 617471
rect 580172 616888 580224 616894
rect 580172 616830 580224 616836
rect 579802 591016 579858 591025
rect 579802 590951 579858 590960
rect 579816 590714 579844 590951
rect 579804 590708 579856 590714
rect 579804 590650 579856 590656
rect 580170 577688 580226 577697
rect 580170 577623 580226 577632
rect 580184 576910 580212 577623
rect 580172 576904 580224 576910
rect 580172 576846 580224 576852
rect 579802 564360 579858 564369
rect 579802 564295 579858 564304
rect 579816 563106 579844 564295
rect 579804 563100 579856 563106
rect 579804 563042 579856 563048
rect 580170 537840 580226 537849
rect 580170 537775 580226 537784
rect 580184 536858 580212 537775
rect 580172 536852 580224 536858
rect 580172 536794 580224 536800
rect 580170 524512 580226 524521
rect 580170 524447 580172 524456
rect 580224 524447 580226 524456
rect 580172 524418 580224 524424
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 580184 510678 580212 511255
rect 580172 510672 580224 510678
rect 580172 510614 580224 510620
rect 580170 484664 580226 484673
rect 580170 484599 580226 484608
rect 580184 484430 580212 484599
rect 580172 484424 580224 484430
rect 580172 484366 580224 484372
rect 579986 471472 580042 471481
rect 579986 471407 580042 471416
rect 580000 470626 580028 471407
rect 579988 470620 580040 470626
rect 579988 470562 580040 470568
rect 580170 458144 580226 458153
rect 580170 458079 580226 458088
rect 580184 456822 580212 458079
rect 580172 456816 580224 456822
rect 580172 456758 580224 456764
rect 580170 431624 580226 431633
rect 580170 431559 580226 431568
rect 580184 430642 580212 431559
rect 580172 430636 580224 430642
rect 580172 430578 580224 430584
rect 580170 418296 580226 418305
rect 580170 418231 580226 418240
rect 580184 418198 580212 418231
rect 580172 418192 580224 418198
rect 580172 418134 580224 418140
rect 580170 404968 580226 404977
rect 580170 404903 580226 404912
rect 580184 404394 580212 404903
rect 580172 404388 580224 404394
rect 580172 404330 580224 404336
rect 580170 378448 580226 378457
rect 580170 378383 580226 378392
rect 580184 378214 580212 378383
rect 580172 378208 580224 378214
rect 580172 378150 580224 378156
rect 580262 365120 580318 365129
rect 580262 365055 580318 365064
rect 580172 351960 580224 351966
rect 580170 351928 580172 351937
rect 580224 351928 580226 351937
rect 580170 351863 580226 351872
rect 580170 325272 580226 325281
rect 580170 325207 580226 325216
rect 580184 324358 580212 325207
rect 580172 324352 580224 324358
rect 580172 324294 580224 324300
rect 579986 312080 580042 312089
rect 579986 312015 580042 312024
rect 580000 311914 580028 312015
rect 579988 311908 580040 311914
rect 579988 311850 580040 311856
rect 580170 298752 580226 298761
rect 580170 298687 580226 298696
rect 580184 298178 580212 298687
rect 580172 298172 580224 298178
rect 580172 298114 580224 298120
rect 527180 278044 527232 278050
rect 527180 277986 527232 277992
rect 580170 272232 580226 272241
rect 580170 272167 580226 272176
rect 580184 271930 580212 272167
rect 580172 271924 580224 271930
rect 580172 271866 580224 271872
rect 525064 268388 525116 268394
rect 525064 268330 525116 268336
rect 580276 263566 580304 365055
rect 580264 263560 580316 263566
rect 580264 263502 580316 263508
rect 580356 263084 580408 263090
rect 580356 263026 580408 263032
rect 218060 262822 218112 262828
rect 477498 262848 477554 262857
rect 477498 262783 477554 262792
rect 472624 261316 472676 261322
rect 472624 261258 472676 261264
rect 471244 260296 471296 260302
rect 471244 260238 471296 260244
rect 199290 210352 199346 210361
rect 199290 210287 199346 210296
rect 198922 200288 198978 200297
rect 198922 200223 198978 200232
rect 198004 198212 198056 198218
rect 198004 198154 198056 198160
rect 197912 148912 197964 148918
rect 197912 148854 197964 148860
rect 197820 148844 197872 148850
rect 197820 148786 197872 148792
rect 197728 141568 197780 141574
rect 197728 141510 197780 141516
rect 197636 139664 197688 139670
rect 197636 139606 197688 139612
rect 197726 137456 197782 137465
rect 197726 137391 197782 137400
rect 197634 79928 197690 79937
rect 197634 79863 197690 79872
rect 197648 79626 197676 79863
rect 197636 79620 197688 79626
rect 197636 79562 197688 79568
rect 197648 78810 197676 79562
rect 197636 78804 197688 78810
rect 197636 78746 197688 78752
rect 197556 74506 197676 74534
rect 197544 66088 197596 66094
rect 197544 66030 197596 66036
rect 197556 65113 197584 66030
rect 197542 65104 197598 65113
rect 197542 65039 197598 65048
rect 197556 64938 197584 65039
rect 197544 64932 197596 64938
rect 197544 64874 197596 64880
rect 197464 60846 197584 60874
rect 197452 60716 197504 60722
rect 197452 60658 197504 60664
rect 197464 60110 197492 60658
rect 197452 60104 197504 60110
rect 197452 60046 197504 60052
rect 197450 56536 197506 56545
rect 197556 56522 197584 60846
rect 197648 56574 197676 74506
rect 197740 70106 197768 137391
rect 197728 70100 197780 70106
rect 197728 70042 197780 70048
rect 197832 60722 197860 148786
rect 197924 67153 197952 148854
rect 198016 80458 198044 198154
rect 198832 198076 198884 198082
rect 198832 198018 198884 198024
rect 198740 186448 198792 186454
rect 198740 186390 198792 186396
rect 198188 152856 198240 152862
rect 198188 152798 198240 152804
rect 198096 147280 198148 147286
rect 198096 147222 198148 147228
rect 198108 81025 198136 147222
rect 198094 81016 198150 81025
rect 198094 80951 198150 80960
rect 198016 80430 198136 80458
rect 198002 80064 198058 80073
rect 198002 79999 198058 80008
rect 198016 79762 198044 79999
rect 198004 79756 198056 79762
rect 198004 79698 198056 79704
rect 198016 78878 198044 79698
rect 198108 79014 198136 80430
rect 198096 79008 198148 79014
rect 198096 78950 198148 78956
rect 198004 78872 198056 78878
rect 198004 78814 198056 78820
rect 198108 78305 198136 78950
rect 198094 78296 198150 78305
rect 198094 78231 198150 78240
rect 198200 72962 198228 152798
rect 198752 147801 198780 186390
rect 198738 147792 198794 147801
rect 198738 147727 198794 147736
rect 198740 75540 198792 75546
rect 198740 75482 198792 75488
rect 198188 72956 198240 72962
rect 198188 72898 198240 72904
rect 197910 67144 197966 67153
rect 197910 67079 197966 67088
rect 197820 60716 197872 60722
rect 197820 60658 197872 60664
rect 197506 56494 197584 56522
rect 197636 56568 197688 56574
rect 197636 56510 197688 56516
rect 197450 56471 197506 56480
rect 197464 56137 197492 56471
rect 197450 56128 197506 56137
rect 197450 56063 197506 56072
rect 197648 55894 197676 56510
rect 197636 55888 197688 55894
rect 197636 55830 197688 55836
rect 197452 53236 197504 53242
rect 197452 53178 197504 53184
rect 197358 45520 197414 45529
rect 197358 45455 197414 45464
rect 197372 44849 197400 45455
rect 197358 44840 197414 44849
rect 197358 44775 197414 44784
rect 197464 16574 197492 53178
rect 197464 16546 197952 16574
rect 196624 4140 196676 4146
rect 196624 4082 196676 4088
rect 196808 4072 196860 4078
rect 196808 4014 196860 4020
rect 196820 480 196848 4014
rect 197924 480 197952 16546
rect 195582 354 195694 480
rect 195164 326 195694 354
rect 195582 -960 195694 326
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 198752 354 198780 75482
rect 198844 55865 198872 198018
rect 198936 63073 198964 200223
rect 199108 192432 199160 192438
rect 199108 192374 199160 192380
rect 199016 186652 199068 186658
rect 199016 186594 199068 186600
rect 199028 70530 199056 186594
rect 199120 74474 199148 192374
rect 199200 186516 199252 186522
rect 199200 186458 199252 186464
rect 199212 78033 199240 186458
rect 199304 148306 199332 210287
rect 471256 206990 471284 260238
rect 472636 245614 472664 261258
rect 580172 259412 580224 259418
rect 580172 259354 580224 259360
rect 580184 258913 580212 259354
rect 580170 258904 580226 258913
rect 580170 258839 580226 258848
rect 472624 245608 472676 245614
rect 580172 245608 580224 245614
rect 472624 245550 472676 245556
rect 580170 245576 580172 245585
rect 580224 245576 580226 245585
rect 580170 245511 580226 245520
rect 580368 219065 580396 263026
rect 580448 262812 580500 262818
rect 580448 262754 580500 262760
rect 580460 232393 580488 262754
rect 580446 232384 580502 232393
rect 580446 232319 580502 232328
rect 580354 219056 580410 219065
rect 580354 218991 580410 219000
rect 471244 206984 471296 206990
rect 471244 206926 471296 206932
rect 579804 206984 579856 206990
rect 579804 206926 579856 206932
rect 579816 205737 579844 206926
rect 579802 205728 579858 205737
rect 579802 205663 579858 205672
rect 200302 200424 200358 200433
rect 200302 200359 200358 200368
rect 199660 198144 199712 198150
rect 199660 198086 199712 198092
rect 199384 152720 199436 152726
rect 199384 152662 199436 152668
rect 199292 148300 199344 148306
rect 199292 148242 199344 148248
rect 199198 78024 199254 78033
rect 199198 77959 199254 77968
rect 199120 74446 199332 74474
rect 199028 70502 199240 70530
rect 199016 70032 199068 70038
rect 199016 69974 199068 69980
rect 199028 69766 199056 69974
rect 199108 69896 199160 69902
rect 199108 69838 199160 69844
rect 199016 69760 199068 69766
rect 199016 69702 199068 69708
rect 199120 69698 199148 69838
rect 199108 69692 199160 69698
rect 199108 69634 199160 69640
rect 199212 68921 199240 70502
rect 199304 69766 199332 74446
rect 199396 70310 199424 152662
rect 199476 148572 199528 148578
rect 199476 148514 199528 148520
rect 199488 79830 199516 148514
rect 199568 148368 199620 148374
rect 199568 148310 199620 148316
rect 199580 80918 199608 148310
rect 199568 80912 199620 80918
rect 199568 80854 199620 80860
rect 199476 79824 199528 79830
rect 199476 79766 199528 79772
rect 199384 70304 199436 70310
rect 199384 70246 199436 70252
rect 199292 69760 199344 69766
rect 199292 69702 199344 69708
rect 199672 69698 199700 198086
rect 200120 193860 200172 193866
rect 200120 193802 200172 193808
rect 199752 152788 199804 152794
rect 199752 152730 199804 152736
rect 199764 70174 199792 152730
rect 199752 70168 199804 70174
rect 199752 70110 199804 70116
rect 199660 69692 199712 69698
rect 199660 69634 199712 69640
rect 199198 68912 199254 68921
rect 199198 68847 199254 68856
rect 199212 68241 199240 68847
rect 199198 68232 199254 68241
rect 199198 68167 199254 68176
rect 198922 63064 198978 63073
rect 198922 62999 198978 63008
rect 198830 55856 198886 55865
rect 198830 55791 198886 55800
rect 200132 50833 200160 193802
rect 200212 192364 200264 192370
rect 200212 192306 200264 192312
rect 200224 53825 200252 192306
rect 200316 67561 200344 200359
rect 204258 200152 204314 200161
rect 204258 200087 204314 200096
rect 201500 199504 201552 199510
rect 201500 199446 201552 199452
rect 200764 194200 200816 194206
rect 200764 194142 200816 194148
rect 200396 155712 200448 155718
rect 200396 155654 200448 155660
rect 200408 71330 200436 155654
rect 200580 155508 200632 155514
rect 200580 155450 200632 155456
rect 200486 152416 200542 152425
rect 200486 152351 200542 152360
rect 200396 71324 200448 71330
rect 200396 71266 200448 71272
rect 200500 70242 200528 152351
rect 200592 74458 200620 155450
rect 200672 148640 200724 148646
rect 200672 148582 200724 148588
rect 200580 74452 200632 74458
rect 200580 74394 200632 74400
rect 200684 70378 200712 148582
rect 200776 78742 200804 194142
rect 201512 173505 201540 199446
rect 202420 199028 202472 199034
rect 202420 198970 202472 198976
rect 201776 192772 201828 192778
rect 201776 192714 201828 192720
rect 201684 185700 201736 185706
rect 201684 185642 201736 185648
rect 201498 173496 201554 173505
rect 201498 173431 201554 173440
rect 200948 147212 201000 147218
rect 200948 147154 201000 147160
rect 200856 147144 200908 147150
rect 200856 147086 200908 147092
rect 200764 78736 200816 78742
rect 200764 78678 200816 78684
rect 200868 76906 200896 147086
rect 200960 80753 200988 147154
rect 200946 80744 201002 80753
rect 200946 80679 201002 80688
rect 201408 78736 201460 78742
rect 201408 78678 201460 78684
rect 201420 77489 201448 78678
rect 201406 77480 201462 77489
rect 201406 77415 201462 77424
rect 200856 76900 200908 76906
rect 200856 76842 200908 76848
rect 201500 75404 201552 75410
rect 201500 75346 201552 75352
rect 200762 71088 200818 71097
rect 200762 71023 200818 71032
rect 200672 70372 200724 70378
rect 200672 70314 200724 70320
rect 200488 70236 200540 70242
rect 200488 70178 200540 70184
rect 200302 67552 200358 67561
rect 200302 67487 200358 67496
rect 200210 53816 200266 53825
rect 200210 53751 200266 53760
rect 200118 50824 200174 50833
rect 200118 50759 200174 50768
rect 200776 3806 200804 71023
rect 201406 68912 201462 68921
rect 201406 68847 201462 68856
rect 201420 68610 201448 68847
rect 201408 68604 201460 68610
rect 201408 68546 201460 68552
rect 201420 67658 201448 68546
rect 201408 67652 201460 67658
rect 201408 67594 201460 67600
rect 201406 67552 201462 67561
rect 201406 67487 201462 67496
rect 201420 67017 201448 67487
rect 201406 67008 201462 67017
rect 201406 66943 201462 66952
rect 201406 53816 201462 53825
rect 201406 53751 201462 53760
rect 201420 53145 201448 53751
rect 201406 53136 201462 53145
rect 201406 53071 201462 53080
rect 201406 50824 201462 50833
rect 201406 50759 201462 50768
rect 201420 50425 201448 50759
rect 201406 50416 201462 50425
rect 201406 50351 201462 50360
rect 201512 11694 201540 75346
rect 201696 58993 201724 185642
rect 201682 58984 201738 58993
rect 201682 58919 201738 58928
rect 201788 56001 201816 192714
rect 201868 155644 201920 155650
rect 201868 155586 201920 155592
rect 201774 55992 201830 56001
rect 201774 55927 201830 55936
rect 201592 49292 201644 49298
rect 201592 49234 201644 49240
rect 201500 11688 201552 11694
rect 201500 11630 201552 11636
rect 201604 6914 201632 49234
rect 201880 45554 201908 155586
rect 201960 155576 202012 155582
rect 201960 155518 202012 155524
rect 201972 69018 202000 155518
rect 202144 155236 202196 155242
rect 202144 155178 202196 155184
rect 202052 148708 202104 148714
rect 202052 148650 202104 148656
rect 201960 69012 202012 69018
rect 201960 68954 202012 68960
rect 202064 61441 202092 148650
rect 202156 73098 202184 155178
rect 202328 150272 202380 150278
rect 202328 150214 202380 150220
rect 202236 148504 202288 148510
rect 202236 148446 202288 148452
rect 202248 78402 202276 148446
rect 202340 79286 202368 150214
rect 202328 79280 202380 79286
rect 202328 79222 202380 79228
rect 202236 78396 202288 78402
rect 202236 78338 202288 78344
rect 202144 73092 202196 73098
rect 202144 73034 202196 73040
rect 202432 71777 202460 198970
rect 203156 198008 203208 198014
rect 203156 197950 203208 197956
rect 202880 193996 202932 194002
rect 202880 193938 202932 193944
rect 202512 193928 202564 193934
rect 202512 193870 202564 193876
rect 202418 71768 202474 71777
rect 202418 71703 202474 71712
rect 202050 61432 202106 61441
rect 202050 61367 202106 61376
rect 202524 49609 202552 193870
rect 202786 71768 202842 71777
rect 202786 71703 202842 71712
rect 202800 71097 202828 71703
rect 202786 71088 202842 71097
rect 202786 71023 202842 71032
rect 202786 58984 202842 58993
rect 202786 58919 202842 58928
rect 202800 58585 202828 58919
rect 202786 58576 202842 58585
rect 202786 58511 202842 58520
rect 202892 55214 202920 193938
rect 203064 192840 203116 192846
rect 203064 192782 203116 192788
rect 202972 192704 203024 192710
rect 202972 192646 203024 192652
rect 202984 64802 203012 192646
rect 203076 68746 203104 192782
rect 203168 77178 203196 197950
rect 203340 155440 203392 155446
rect 203340 155382 203392 155388
rect 203248 151088 203300 151094
rect 203248 151030 203300 151036
rect 203156 77172 203208 77178
rect 203156 77114 203208 77120
rect 203064 68740 203116 68746
rect 203064 68682 203116 68688
rect 202972 64796 203024 64802
rect 202972 64738 203024 64744
rect 202984 64190 203012 64738
rect 202972 64184 203024 64190
rect 202972 64126 203024 64132
rect 202880 55208 202932 55214
rect 202880 55150 202932 55156
rect 202892 54534 202920 55150
rect 202880 54528 202932 54534
rect 202880 54470 202932 54476
rect 202510 49600 202566 49609
rect 202510 49535 202566 49544
rect 203260 46889 203288 151030
rect 203352 57934 203380 155382
rect 203524 155372 203576 155378
rect 203524 155314 203576 155320
rect 203432 155304 203484 155310
rect 203432 155246 203484 155252
rect 203444 68882 203472 155246
rect 203432 68876 203484 68882
rect 203432 68818 203484 68824
rect 203536 68814 203564 155314
rect 203708 149864 203760 149870
rect 203708 149806 203760 149812
rect 203616 148436 203668 148442
rect 203616 148378 203668 148384
rect 203628 68950 203656 148378
rect 203720 79218 203748 149806
rect 203708 79212 203760 79218
rect 203708 79154 203760 79160
rect 203708 74248 203760 74254
rect 203708 74190 203760 74196
rect 203616 68944 203668 68950
rect 203616 68886 203668 68892
rect 203524 68808 203576 68814
rect 203524 68750 203576 68756
rect 203340 57928 203392 57934
rect 203340 57870 203392 57876
rect 203246 46880 203302 46889
rect 203246 46815 203302 46824
rect 201788 45526 201908 45554
rect 201788 44169 201816 45526
rect 201774 44160 201830 44169
rect 201774 44095 201830 44104
rect 202786 44160 202842 44169
rect 202786 44095 202842 44104
rect 202800 43489 202828 44095
rect 202786 43480 202842 43489
rect 202786 43415 202842 43424
rect 202696 11688 202748 11694
rect 202696 11630 202748 11636
rect 201512 6886 201632 6914
rect 200304 3800 200356 3806
rect 200304 3742 200356 3748
rect 200764 3800 200816 3806
rect 200764 3742 200816 3748
rect 200316 480 200344 3742
rect 201512 480 201540 6886
rect 202708 480 202736 11630
rect 203720 4078 203748 74190
rect 204272 72826 204300 200087
rect 208584 199232 208636 199238
rect 208584 199174 208636 199180
rect 208492 198892 208544 198898
rect 208492 198834 208544 198840
rect 208400 198824 208452 198830
rect 208400 198766 208452 198772
rect 207020 194064 207072 194070
rect 207020 194006 207072 194012
rect 205640 193112 205692 193118
rect 205640 193054 205692 193060
rect 204352 192976 204404 192982
rect 204352 192918 204404 192924
rect 204260 72820 204312 72826
rect 204260 72762 204312 72768
rect 204364 70990 204392 192918
rect 204720 152652 204772 152658
rect 204720 152594 204772 152600
rect 204444 150204 204496 150210
rect 204444 150146 204496 150152
rect 204352 70984 204404 70990
rect 204352 70926 204404 70932
rect 204168 68740 204220 68746
rect 204168 68682 204220 68688
rect 204180 68338 204208 68682
rect 204168 68332 204220 68338
rect 204168 68274 204220 68280
rect 204168 57928 204220 57934
rect 204168 57870 204220 57876
rect 204180 57254 204208 57870
rect 204168 57248 204220 57254
rect 204168 57190 204220 57196
rect 204456 49337 204484 150146
rect 204536 147008 204588 147014
rect 204536 146950 204588 146956
rect 204442 49328 204498 49337
rect 204442 49263 204498 49272
rect 204548 48113 204576 146950
rect 204628 146940 204680 146946
rect 204628 146882 204680 146888
rect 204640 52465 204668 146882
rect 204732 71738 204760 152594
rect 204812 152584 204864 152590
rect 204812 152526 204864 152532
rect 204824 78334 204852 152526
rect 204904 150340 204956 150346
rect 204904 150282 204956 150288
rect 204812 78328 204864 78334
rect 204812 78270 204864 78276
rect 204916 78169 204944 150282
rect 204902 78160 204958 78169
rect 204902 78095 204958 78104
rect 204720 71732 204772 71738
rect 204720 71674 204772 71680
rect 204732 71194 204760 71674
rect 204720 71188 204772 71194
rect 204720 71130 204772 71136
rect 204626 52456 204682 52465
rect 204626 52391 204682 52400
rect 204640 51785 204668 52391
rect 204626 51776 204682 51785
rect 204626 51711 204682 51720
rect 204718 49328 204774 49337
rect 204718 49263 204774 49272
rect 204732 48929 204760 49263
rect 204718 48920 204774 48929
rect 204718 48855 204774 48864
rect 204534 48104 204590 48113
rect 204534 48039 204590 48048
rect 204810 48104 204866 48113
rect 204810 48039 204866 48048
rect 204824 47569 204852 48039
rect 204810 47560 204866 47569
rect 204810 47495 204866 47504
rect 204260 46300 204312 46306
rect 204260 46242 204312 46248
rect 204272 16574 204300 46242
rect 205652 42809 205680 193054
rect 205732 186380 205784 186386
rect 205732 186322 205784 186328
rect 205744 75857 205772 186322
rect 206192 152516 206244 152522
rect 206192 152458 206244 152464
rect 205824 150408 205876 150414
rect 205824 150350 205876 150356
rect 205730 75848 205786 75857
rect 205730 75783 205786 75792
rect 205836 50289 205864 150350
rect 205916 150068 205968 150074
rect 205916 150010 205968 150016
rect 205928 74322 205956 150010
rect 206100 150000 206152 150006
rect 206100 149942 206152 149948
rect 206008 149932 206060 149938
rect 206008 149874 206060 149880
rect 205916 74316 205968 74322
rect 205916 74258 205968 74264
rect 206020 73778 206048 149874
rect 206112 75721 206140 149942
rect 206204 78470 206232 152458
rect 206284 150136 206336 150142
rect 206284 150078 206336 150084
rect 206296 78674 206324 150078
rect 206376 149796 206428 149802
rect 206376 149738 206428 149744
rect 206388 78849 206416 149738
rect 206468 145580 206520 145586
rect 206468 145522 206520 145528
rect 206374 78840 206430 78849
rect 206374 78775 206430 78784
rect 206284 78668 206336 78674
rect 206284 78610 206336 78616
rect 206480 78606 206508 145522
rect 206468 78600 206520 78606
rect 206468 78542 206520 78548
rect 206192 78464 206244 78470
rect 206192 78406 206244 78412
rect 207032 77761 207060 194006
rect 207112 192908 207164 192914
rect 207112 192850 207164 192856
rect 207018 77752 207074 77761
rect 207018 77687 207074 77696
rect 207124 76430 207152 192850
rect 207112 76424 207164 76430
rect 207112 76366 207164 76372
rect 206098 75712 206154 75721
rect 206098 75647 206154 75656
rect 206008 73772 206060 73778
rect 206008 73714 206060 73720
rect 207020 65612 207072 65618
rect 207020 65554 207072 65560
rect 205822 50280 205878 50289
rect 205822 50215 205878 50224
rect 205638 42800 205694 42809
rect 205638 42735 205694 42744
rect 205652 42129 205680 42735
rect 205638 42120 205694 42129
rect 205638 42055 205694 42064
rect 205640 32700 205692 32706
rect 205640 32642 205692 32648
rect 205652 16574 205680 32642
rect 204272 16546 205128 16574
rect 205652 16546 206232 16574
rect 203892 4140 203944 4146
rect 203892 4082 203944 4088
rect 203708 4072 203760 4078
rect 203708 4014 203760 4020
rect 203904 480 203932 4082
rect 205100 480 205128 16546
rect 206204 480 206232 16546
rect 199078 354 199190 480
rect 198752 326 199190 354
rect 199078 -960 199190 326
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207032 354 207060 65554
rect 208412 64841 208440 198766
rect 208504 73166 208532 198834
rect 208596 80850 208624 199174
rect 580172 193180 580224 193186
rect 580172 193122 580224 193128
rect 208674 192672 208730 192681
rect 208674 192607 208730 192616
rect 208584 80844 208636 80850
rect 208584 80786 208636 80792
rect 208688 76265 208716 192607
rect 580184 192545 580212 193122
rect 580170 192536 580226 192545
rect 580170 192471 580226 192480
rect 580170 179208 580226 179217
rect 580170 179143 580226 179152
rect 580184 178090 580212 179143
rect 580172 178084 580224 178090
rect 580172 178026 580224 178032
rect 580172 166320 580224 166326
rect 580172 166262 580224 166268
rect 580184 165889 580212 166262
rect 580170 165880 580226 165889
rect 580170 165815 580226 165824
rect 580262 152688 580318 152697
rect 580262 152623 580318 152632
rect 580276 143546 580304 152623
rect 580356 146328 580408 146334
rect 580356 146270 580408 146276
rect 580264 143540 580316 143546
rect 580264 143482 580316 143488
rect 549904 140956 549956 140962
rect 549904 140898 549956 140904
rect 286322 139768 286378 139777
rect 286322 139703 286378 139712
rect 234620 80844 234672 80850
rect 234620 80786 234672 80792
rect 224224 76832 224276 76838
rect 224224 76774 224276 76780
rect 208674 76256 208730 76265
rect 208674 76191 208730 76200
rect 208492 73160 208544 73166
rect 208492 73102 208544 73108
rect 220084 72820 220136 72826
rect 220084 72762 220136 72768
rect 217324 71188 217376 71194
rect 217324 71130 217376 71136
rect 213918 67280 213974 67289
rect 213918 67215 213974 67224
rect 208398 64832 208454 64841
rect 208398 64767 208454 64776
rect 208412 64433 208440 64767
rect 208398 64424 208454 64433
rect 208398 64359 208454 64368
rect 209870 54904 209926 54913
rect 209870 54839 209926 54848
rect 208400 36916 208452 36922
rect 208400 36858 208452 36864
rect 208412 16574 208440 36858
rect 208412 16546 208624 16574
rect 208596 480 208624 16546
rect 209884 6914 209912 54839
rect 211160 51808 211212 51814
rect 211160 51750 211212 51756
rect 211172 16574 211200 51750
rect 212538 45112 212594 45121
rect 212538 45047 212594 45056
rect 212552 16574 212580 45047
rect 213932 16574 213960 67215
rect 215300 57452 215352 57458
rect 215300 57394 215352 57400
rect 211172 16546 211752 16574
rect 212552 16546 213408 16574
rect 213932 16546 214512 16574
rect 209792 6886 209912 6914
rect 209792 480 209820 6886
rect 210976 3800 211028 3806
rect 210976 3742 211028 3748
rect 210988 480 211016 3742
rect 207358 354 207470 480
rect 207032 326 207470 354
rect 207358 -960 207470 326
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 211724 354 211752 16546
rect 213380 480 213408 16546
rect 214484 480 214512 16546
rect 212142 354 212254 480
rect 211724 326 212254 354
rect 212142 -960 212254 326
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215312 354 215340 57394
rect 216680 43648 216732 43654
rect 216680 43590 216732 43596
rect 216692 16574 216720 43590
rect 216692 16546 216904 16574
rect 216876 480 216904 16546
rect 217336 3398 217364 71130
rect 218152 49088 218204 49094
rect 218152 49030 218204 49036
rect 218164 16574 218192 49030
rect 219440 23044 219492 23050
rect 219440 22986 219492 22992
rect 219452 16574 219480 22986
rect 218164 16546 219296 16574
rect 219452 16546 220032 16574
rect 217324 3392 217376 3398
rect 217324 3334 217376 3340
rect 218060 3392 218112 3398
rect 218060 3334 218112 3340
rect 218072 480 218100 3334
rect 219268 480 219296 16546
rect 215638 354 215750 480
rect 215312 326 215750 354
rect 215638 -960 215750 326
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220004 354 220032 16546
rect 220096 3806 220124 72762
rect 220818 68368 220874 68377
rect 220818 68303 220874 68312
rect 220832 16574 220860 68303
rect 222200 36848 222252 36854
rect 222200 36790 222252 36796
rect 222212 16574 222240 36790
rect 220832 16546 221136 16574
rect 222212 16546 222792 16574
rect 220084 3800 220136 3806
rect 220084 3742 220136 3748
rect 220422 354 220534 480
rect 220004 326 220534 354
rect 221108 354 221136 16546
rect 222764 480 222792 16546
rect 224236 4078 224264 76774
rect 229742 73944 229798 73953
rect 229742 73879 229798 73888
rect 224960 64320 225012 64326
rect 224960 64262 225012 64268
rect 224972 16574 225000 64262
rect 227720 62892 227772 62898
rect 227720 62834 227772 62840
rect 227732 16574 227760 62834
rect 229098 30968 229154 30977
rect 229098 30903 229154 30912
rect 229112 16574 229140 30903
rect 224972 16546 225184 16574
rect 227732 16546 228312 16574
rect 229112 16546 229416 16574
rect 223948 4072 224000 4078
rect 223948 4014 224000 4020
rect 224224 4072 224276 4078
rect 224224 4014 224276 4020
rect 223960 480 223988 4014
rect 225156 480 225184 16546
rect 227536 7880 227588 7886
rect 227536 7822 227588 7828
rect 226340 4004 226392 4010
rect 226340 3946 226392 3952
rect 226352 480 226380 3946
rect 227548 480 227576 7822
rect 221526 354 221638 480
rect 221108 326 221638 354
rect 220422 -960 220534 326
rect 221526 -960 221638 326
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228284 354 228312 16546
rect 228702 354 228814 480
rect 228284 326 228814 354
rect 229388 354 229416 16546
rect 229756 3398 229784 73879
rect 231858 56400 231914 56409
rect 231858 56335 231914 56344
rect 229744 3392 229796 3398
rect 229744 3334 229796 3340
rect 231032 3392 231084 3398
rect 231032 3334 231084 3340
rect 231044 480 231072 3334
rect 229806 354 229918 480
rect 229388 326 229918 354
rect 228702 -960 228814 326
rect 229806 -960 229918 326
rect 231002 -960 231114 480
rect 231872 354 231900 56335
rect 233240 42356 233292 42362
rect 233240 42298 233292 42304
rect 233252 16574 233280 42298
rect 233252 16546 233464 16574
rect 233436 480 233464 16546
rect 234632 11694 234660 80786
rect 270500 80776 270552 80782
rect 270500 80718 270552 80724
rect 252560 80164 252612 80170
rect 252560 80106 252612 80112
rect 238760 79484 238812 79490
rect 238760 79426 238812 79432
rect 237380 53168 237432 53174
rect 237380 53110 237432 53116
rect 236000 32632 236052 32638
rect 236000 32574 236052 32580
rect 234712 17536 234764 17542
rect 234712 17478 234764 17484
rect 234620 11688 234672 11694
rect 234620 11630 234672 11636
rect 234724 6914 234752 17478
rect 236012 16574 236040 32574
rect 237392 16574 237420 53110
rect 238772 16574 238800 79426
rect 247040 76764 247092 76770
rect 247040 76706 247092 76712
rect 242898 67416 242954 67425
rect 242898 67351 242954 67360
rect 236012 16546 236592 16574
rect 237392 16546 237696 16574
rect 238772 16546 239352 16574
rect 235816 11688 235868 11694
rect 235816 11630 235868 11636
rect 234632 6886 234752 6914
rect 234632 480 234660 6886
rect 235828 480 235856 11630
rect 232198 354 232310 480
rect 231872 326 232310 354
rect 232198 -960 232310 326
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236564 354 236592 16546
rect 236982 354 237094 480
rect 236564 326 237094 354
rect 237668 354 237696 16546
rect 239324 480 239352 16546
rect 241704 9240 241756 9246
rect 241704 9182 241756 9188
rect 240508 4072 240560 4078
rect 240508 4014 240560 4020
rect 240520 480 240548 4014
rect 241716 480 241744 9182
rect 242912 480 242940 67351
rect 245658 61296 245714 61305
rect 245658 61231 245714 61240
rect 242992 29912 243044 29918
rect 242992 29854 243044 29860
rect 243004 16574 243032 29854
rect 245672 16574 245700 61231
rect 247052 16574 247080 76706
rect 248420 73840 248472 73846
rect 248420 73782 248472 73788
rect 243004 16546 244136 16574
rect 245672 16546 245976 16574
rect 247052 16546 247632 16574
rect 244108 480 244136 16546
rect 245200 10600 245252 10606
rect 245200 10542 245252 10548
rect 245212 480 245240 10542
rect 238086 354 238198 480
rect 237668 326 238198 354
rect 236982 -960 237094 326
rect 238086 -960 238198 326
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 245948 354 245976 16546
rect 247604 480 247632 16546
rect 246366 354 246478 480
rect 245948 326 246478 354
rect 246366 -960 246478 326
rect 247562 -960 247674 480
rect 248432 354 248460 73782
rect 249798 62112 249854 62121
rect 249798 62047 249854 62056
rect 249812 16574 249840 62047
rect 251180 39636 251232 39642
rect 251180 39578 251232 39584
rect 249812 16546 250024 16574
rect 249996 480 250024 16546
rect 251192 480 251220 39578
rect 252572 16574 252600 80106
rect 255964 78192 256016 78198
rect 255964 78134 256016 78140
rect 253940 76696 253992 76702
rect 253940 76638 253992 76644
rect 253952 16574 253980 76638
rect 255976 73846 256004 78134
rect 269764 77308 269816 77314
rect 269764 77250 269816 77256
rect 260838 76664 260894 76673
rect 260838 76599 260894 76608
rect 255964 73840 256016 73846
rect 255964 73782 256016 73788
rect 259458 64424 259514 64433
rect 259458 64359 259514 64368
rect 255320 57384 255372 57390
rect 255320 57326 255372 57332
rect 255332 16574 255360 57326
rect 256700 47728 256752 47734
rect 256700 47670 256752 47676
rect 252572 16546 253520 16574
rect 253952 16546 254256 16574
rect 255332 16546 255912 16574
rect 252376 11960 252428 11966
rect 252376 11902 252428 11908
rect 252388 480 252416 11902
rect 253492 480 253520 16546
rect 248758 354 248870 480
rect 248432 326 248870 354
rect 248758 -960 248870 326
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254228 354 254256 16546
rect 255884 480 255912 16546
rect 254646 354 254758 480
rect 254228 326 254758 354
rect 254646 -960 254758 326
rect 255842 -960 255954 480
rect 256712 354 256740 47670
rect 258264 13320 258316 13326
rect 258264 13262 258316 13268
rect 258276 480 258304 13262
rect 259472 11694 259500 64359
rect 260852 16574 260880 76599
rect 262220 74180 262272 74186
rect 262220 74122 262272 74128
rect 262232 16574 262260 74122
rect 269776 73914 269804 77250
rect 269120 73908 269172 73914
rect 269120 73850 269172 73856
rect 269764 73908 269816 73914
rect 269764 73850 269816 73856
rect 263600 60172 263652 60178
rect 263600 60114 263652 60120
rect 263612 16574 263640 60114
rect 267738 44976 267794 44985
rect 267738 44911 267794 44920
rect 264978 28248 265034 28257
rect 264978 28183 265034 28192
rect 260852 16546 261800 16574
rect 262232 16546 262536 16574
rect 263612 16546 264192 16574
rect 259552 16108 259604 16114
rect 259552 16050 259604 16056
rect 259460 11688 259512 11694
rect 259460 11630 259512 11636
rect 259564 6914 259592 16050
rect 260656 11688 260708 11694
rect 260656 11630 260708 11636
rect 259472 6886 259592 6914
rect 259472 480 259500 6886
rect 260668 480 260696 11630
rect 261772 480 261800 16546
rect 257038 354 257150 480
rect 256712 326 257150 354
rect 257038 -960 257150 326
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262508 354 262536 16546
rect 264164 480 264192 16546
rect 262926 354 263038 480
rect 262508 326 263038 354
rect 262926 -960 263038 326
rect 264122 -960 264234 480
rect 264992 354 265020 28183
rect 266360 18896 266412 18902
rect 266360 18838 266412 18844
rect 266372 16574 266400 18838
rect 266372 16546 266584 16574
rect 266556 480 266584 16546
rect 267752 480 267780 44911
rect 267832 38208 267884 38214
rect 267832 38150 267884 38156
rect 267844 16574 267872 38150
rect 269132 16574 269160 73850
rect 270512 16574 270540 80718
rect 285680 79144 285732 79150
rect 285680 79086 285732 79092
rect 284300 74112 284352 74118
rect 284300 74054 284352 74060
rect 274638 65648 274694 65657
rect 274638 65583 274694 65592
rect 274652 16574 274680 65583
rect 277398 61976 277454 61985
rect 277398 61911 277454 61920
rect 276020 35488 276072 35494
rect 276020 35430 276072 35436
rect 267844 16546 268424 16574
rect 269132 16546 270080 16574
rect 270512 16546 270816 16574
rect 274652 16546 274864 16574
rect 265318 354 265430 480
rect 264992 326 265430 354
rect 265318 -960 265430 326
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268396 354 268424 16546
rect 270052 480 270080 16546
rect 268814 354 268926 480
rect 268396 326 268926 354
rect 268814 -960 268926 326
rect 270010 -960 270122 480
rect 270788 354 270816 16546
rect 272432 6452 272484 6458
rect 272432 6394 272484 6400
rect 272444 480 272472 6394
rect 273628 5092 273680 5098
rect 273628 5034 273680 5040
rect 273640 480 273668 5034
rect 274836 480 274864 16546
rect 276032 4010 276060 35430
rect 277412 16574 277440 61911
rect 281540 58744 281592 58750
rect 281540 58686 281592 58692
rect 278778 53544 278834 53553
rect 278778 53479 278834 53488
rect 278792 16574 278820 53479
rect 280160 20256 280212 20262
rect 280160 20198 280212 20204
rect 280172 16574 280200 20198
rect 277412 16546 278360 16574
rect 278792 16546 279096 16574
rect 280172 16546 280752 16574
rect 276112 14748 276164 14754
rect 276112 14690 276164 14696
rect 276020 4004 276072 4010
rect 276020 3946 276072 3952
rect 276124 3482 276152 14690
rect 276756 4004 276808 4010
rect 276756 3946 276808 3952
rect 276032 3454 276152 3482
rect 276032 480 276060 3454
rect 271206 354 271318 480
rect 270788 326 271318 354
rect 271206 -960 271318 326
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 276768 354 276796 3946
rect 278332 480 278360 16546
rect 277094 354 277206 480
rect 276768 326 277206 354
rect 277094 -960 277206 326
rect 278290 -960 278402 480
rect 279068 354 279096 16546
rect 280724 480 280752 16546
rect 279486 354 279598 480
rect 279068 326 279598 354
rect 279486 -960 279598 326
rect 280682 -960 280794 480
rect 281552 354 281580 58686
rect 282920 27192 282972 27198
rect 282920 27134 282972 27140
rect 282932 16574 282960 27134
rect 282932 16546 283144 16574
rect 283116 480 283144 16546
rect 284312 480 284340 74054
rect 284390 43616 284446 43625
rect 284390 43551 284446 43560
rect 284404 16574 284432 43551
rect 285692 16574 285720 79086
rect 286336 20670 286364 139703
rect 327722 139632 327778 139641
rect 327722 139567 327778 139576
rect 288440 80708 288492 80714
rect 288440 80650 288492 80656
rect 286324 20664 286376 20670
rect 286324 20606 286376 20612
rect 287060 20188 287112 20194
rect 287060 20130 287112 20136
rect 287072 16574 287100 20130
rect 288452 16574 288480 80650
rect 302240 80096 302292 80102
rect 302240 80038 302292 80044
rect 291842 77888 291898 77897
rect 291842 77823 291898 77832
rect 289820 76016 289872 76022
rect 289820 75958 289872 75964
rect 284404 16546 284984 16574
rect 285692 16546 286640 16574
rect 287072 16546 287376 16574
rect 288452 16546 289032 16574
rect 281878 354 281990 480
rect 281552 326 281990 354
rect 281878 -960 281990 326
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 284956 354 284984 16546
rect 286612 480 286640 16546
rect 285374 354 285486 480
rect 284956 326 285486 354
rect 285374 -960 285486 326
rect 286570 -960 286682 480
rect 287348 354 287376 16546
rect 289004 480 289032 16546
rect 287766 354 287878 480
rect 287348 326 287878 354
rect 287766 -960 287878 326
rect 288962 -960 289074 480
rect 289832 354 289860 75958
rect 291856 19990 291884 77823
rect 296720 75948 296772 75954
rect 296720 75890 296772 75896
rect 295340 66904 295392 66910
rect 295340 66846 295392 66852
rect 292578 63336 292634 63345
rect 292578 63271 292634 63280
rect 291200 19984 291252 19990
rect 291200 19926 291252 19932
rect 291844 19984 291896 19990
rect 291844 19926 291896 19932
rect 291212 16574 291240 19926
rect 291212 16546 291424 16574
rect 291396 480 291424 16546
rect 292592 480 292620 63271
rect 292672 42288 292724 42294
rect 292672 42230 292724 42236
rect 292684 16574 292712 42230
rect 293960 20120 294012 20126
rect 293960 20062 294012 20068
rect 293972 16574 294000 20062
rect 295352 16574 295380 66846
rect 296732 16574 296760 75890
rect 297364 74044 297416 74050
rect 297364 73986 297416 73992
rect 292684 16546 293264 16574
rect 293972 16546 294920 16574
rect 295352 16546 295656 16574
rect 296732 16546 297312 16574
rect 290158 354 290270 480
rect 289832 326 290270 354
rect 290158 -960 290270 326
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293236 354 293264 16546
rect 294892 480 294920 16546
rect 293654 354 293766 480
rect 293236 326 293766 354
rect 293654 -960 293766 326
rect 294850 -960 294962 480
rect 295628 354 295656 16546
rect 297284 480 297312 16546
rect 297376 3058 297404 73986
rect 299478 60208 299534 60217
rect 299478 60143 299534 60152
rect 299492 3482 299520 60143
rect 300860 40996 300912 41002
rect 300860 40938 300912 40944
rect 299572 34060 299624 34066
rect 299572 34002 299624 34008
rect 299584 4010 299612 34002
rect 300872 16574 300900 40938
rect 302252 16574 302280 80038
rect 304998 73808 305054 73817
rect 304998 73743 305054 73752
rect 304264 71868 304316 71874
rect 304264 71810 304316 71816
rect 303620 36780 303672 36786
rect 303620 36722 303672 36728
rect 303632 16574 303660 36722
rect 300872 16546 301544 16574
rect 302252 16546 303200 16574
rect 303632 16546 303936 16574
rect 299572 4004 299624 4010
rect 299572 3946 299624 3952
rect 300768 4004 300820 4010
rect 300768 3946 300820 3952
rect 299492 3454 299704 3482
rect 297364 3052 297416 3058
rect 297364 2994 297416 3000
rect 298468 3052 298520 3058
rect 298468 2994 298520 3000
rect 298480 480 298508 2994
rect 299676 480 299704 3454
rect 300780 480 300808 3946
rect 296046 354 296158 480
rect 295628 326 296158 354
rect 296046 -960 296158 326
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301516 354 301544 16546
rect 303172 480 303200 16546
rect 301934 354 302046 480
rect 301516 326 302046 354
rect 301934 -960 302046 326
rect 303130 -960 303242 480
rect 303908 354 303936 16546
rect 304276 4146 304304 71810
rect 305012 16574 305040 73743
rect 327736 73166 327764 139567
rect 549916 86970 549944 140898
rect 576122 140176 576178 140185
rect 576122 140111 576178 140120
rect 549904 86964 549956 86970
rect 549904 86906 549956 86912
rect 382278 79520 382334 79529
rect 382278 79455 382334 79464
rect 376760 79076 376812 79082
rect 376760 79018 376812 79024
rect 337384 78124 337436 78130
rect 337384 78066 337436 78072
rect 327724 73160 327776 73166
rect 327724 73102 327776 73108
rect 311164 72752 311216 72758
rect 311164 72694 311216 72700
rect 309140 40928 309192 40934
rect 309140 40870 309192 40876
rect 309152 16574 309180 40870
rect 310520 25832 310572 25838
rect 310520 25774 310572 25780
rect 310532 16574 310560 25774
rect 305012 16546 305592 16574
rect 309152 16546 309824 16574
rect 310532 16546 311112 16574
rect 304264 4140 304316 4146
rect 304264 4082 304316 4088
rect 305564 480 305592 16546
rect 307944 13252 307996 13258
rect 307944 13194 307996 13200
rect 306748 3936 306800 3942
rect 306748 3878 306800 3884
rect 306760 480 306788 3878
rect 307956 480 307984 13194
rect 309048 4140 309100 4146
rect 309048 4082 309100 4088
rect 309060 480 309088 4082
rect 304326 354 304438 480
rect 303908 326 304438 354
rect 304326 -960 304438 326
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 309796 354 309824 16546
rect 311084 3482 311112 16546
rect 311176 3942 311204 72694
rect 318800 72684 318852 72690
rect 318800 72626 318852 72632
rect 313278 57488 313334 57497
rect 313278 57423 313334 57432
rect 313292 16574 313320 57423
rect 315302 56264 315358 56273
rect 315302 56199 315358 56208
rect 314660 24404 314712 24410
rect 314660 24346 314712 24352
rect 313292 16546 313872 16574
rect 311164 3936 311216 3942
rect 311164 3878 311216 3884
rect 312636 3936 312688 3942
rect 312636 3878 312688 3884
rect 311084 3454 311480 3482
rect 311452 480 311480 3454
rect 312648 480 312676 3878
rect 313844 480 313872 16546
rect 310214 354 310326 480
rect 309796 326 310326 354
rect 310214 -960 310326 326
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314672 354 314700 24346
rect 315316 3330 315344 56199
rect 317420 31272 317472 31278
rect 317420 31214 317472 31220
rect 316132 22976 316184 22982
rect 316132 22918 316184 22924
rect 316144 16574 316172 22918
rect 317432 16574 317460 31214
rect 318812 16574 318840 72626
rect 324964 72616 325016 72622
rect 324964 72558 325016 72564
rect 322940 71800 322992 71806
rect 322940 71742 322992 71748
rect 320178 61840 320234 61849
rect 320178 61775 320234 61784
rect 320192 16574 320220 61775
rect 321560 35420 321612 35426
rect 321560 35362 321612 35368
rect 321572 16574 321600 35362
rect 316144 16546 316264 16574
rect 317432 16546 318104 16574
rect 318812 16546 319760 16574
rect 320192 16546 320496 16574
rect 321572 16546 322152 16574
rect 315304 3324 315356 3330
rect 315304 3266 315356 3272
rect 316236 480 316264 16546
rect 317328 3324 317380 3330
rect 317328 3266 317380 3272
rect 317340 480 317368 3266
rect 314998 354 315110 480
rect 314672 326 315110 354
rect 314998 -960 315110 326
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318076 354 318104 16546
rect 319732 480 319760 16546
rect 318494 354 318606 480
rect 318076 326 318606 354
rect 318494 -960 318606 326
rect 319690 -960 319802 480
rect 320468 354 320496 16546
rect 322124 480 322152 16546
rect 320886 354 320998 480
rect 320468 326 320998 354
rect 320886 -960 320998 326
rect 322082 -960 322194 480
rect 322952 354 322980 71742
rect 324320 65544 324372 65550
rect 324320 65486 324372 65492
rect 324332 3210 324360 65486
rect 324412 14680 324464 14686
rect 324412 14622 324464 14628
rect 324424 3398 324452 14622
rect 324412 3392 324464 3398
rect 324412 3334 324464 3340
rect 324332 3182 324452 3210
rect 324976 3194 325004 72558
rect 332600 72548 332652 72554
rect 332600 72490 332652 72496
rect 331218 63200 331274 63209
rect 331218 63135 331274 63144
rect 327078 58848 327134 58857
rect 327078 58783 327134 58792
rect 327092 16574 327120 58783
rect 328460 42220 328512 42226
rect 328460 42162 328512 42168
rect 328472 16574 328500 42162
rect 329840 21684 329892 21690
rect 329840 21626 329892 21632
rect 329852 16574 329880 21626
rect 327092 16546 328040 16574
rect 328472 16546 328776 16574
rect 329852 16546 330432 16574
rect 325608 3392 325660 3398
rect 325608 3334 325660 3340
rect 324424 480 324452 3182
rect 324964 3188 325016 3194
rect 324964 3130 325016 3136
rect 325620 480 325648 3334
rect 326804 3188 326856 3194
rect 326804 3130 326856 3136
rect 326816 480 326844 3130
rect 328012 480 328040 16546
rect 323278 354 323390 480
rect 322952 326 323390 354
rect 323278 -960 323390 326
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 328748 354 328776 16546
rect 330404 480 330432 16546
rect 329166 354 329278 480
rect 328748 326 329278 354
rect 329166 -960 329278 326
rect 330362 -960 330474 480
rect 331232 354 331260 63135
rect 332612 3398 332640 72490
rect 336004 71120 336056 71126
rect 336004 71062 336056 71068
rect 333978 54768 334034 54777
rect 333978 54703 334034 54712
rect 332692 29844 332744 29850
rect 332692 29786 332744 29792
rect 332600 3392 332652 3398
rect 332600 3334 332652 3340
rect 332704 480 332732 29786
rect 333992 16574 334020 54703
rect 333992 16546 334664 16574
rect 333888 3392 333940 3398
rect 333888 3334 333940 3340
rect 333900 480 333928 3334
rect 331558 354 331670 480
rect 331232 326 331670 354
rect 331558 -960 331670 326
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 334636 354 334664 16546
rect 336016 3194 336044 71062
rect 337396 21622 337424 78066
rect 353300 76628 353352 76634
rect 353300 76570 353352 76576
rect 347780 73976 347832 73982
rect 347780 73918 347832 73924
rect 346400 65000 346452 65006
rect 346400 64942 346452 64948
rect 338118 60072 338174 60081
rect 338118 60007 338174 60016
rect 336740 21616 336792 21622
rect 336740 21558 336792 21564
rect 337384 21616 337436 21622
rect 337384 21558 337436 21564
rect 336752 16574 336780 21558
rect 338132 16574 338160 60007
rect 345020 57316 345072 57322
rect 345020 57258 345072 57264
rect 340972 39568 341024 39574
rect 340972 39510 341024 39516
rect 339500 28484 339552 28490
rect 339500 28426 339552 28432
rect 336752 16546 337056 16574
rect 338132 16546 338712 16574
rect 336280 6384 336332 6390
rect 336280 6326 336332 6332
rect 336004 3188 336056 3194
rect 336004 3130 336056 3136
rect 336292 480 336320 6326
rect 335054 354 335166 480
rect 334636 326 335166 354
rect 335054 -960 335166 326
rect 336250 -960 336362 480
rect 337028 354 337056 16546
rect 338684 480 338712 16546
rect 337446 354 337558 480
rect 337028 326 337558 354
rect 337446 -960 337558 326
rect 338642 -960 338754 480
rect 339512 354 339540 28426
rect 340984 480 341012 39510
rect 343640 21548 343692 21554
rect 343640 21490 343692 21496
rect 343652 16574 343680 21490
rect 345032 16574 345060 57258
rect 346412 16574 346440 64942
rect 347792 16574 347820 73918
rect 349160 62824 349212 62830
rect 349160 62766 349212 62772
rect 343652 16546 344600 16574
rect 345032 16546 345336 16574
rect 346412 16546 346992 16574
rect 347792 16546 348096 16574
rect 342904 10532 342956 10538
rect 342904 10474 342956 10480
rect 342168 3188 342220 3194
rect 342168 3130 342220 3136
rect 342180 480 342208 3130
rect 339838 354 339950 480
rect 339512 326 339950 354
rect 339838 -960 339950 326
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 342916 354 342944 10474
rect 344572 480 344600 16546
rect 343334 354 343446 480
rect 342916 326 343446 354
rect 343334 -960 343446 326
rect 344530 -960 344642 480
rect 345308 354 345336 16546
rect 346964 480 346992 16546
rect 348068 480 348096 16546
rect 349172 3210 349200 62766
rect 351918 53408 351974 53417
rect 351918 53343 351974 53352
rect 350540 21480 350592 21486
rect 350540 21422 350592 21428
rect 350552 16574 350580 21422
rect 351932 16574 351960 53343
rect 353312 16574 353340 76570
rect 375380 72480 375432 72486
rect 375380 72422 375432 72428
rect 367100 71052 367152 71058
rect 367100 70994 367152 71000
rect 354680 69828 354732 69834
rect 354680 69770 354732 69776
rect 354692 16574 354720 69770
rect 358820 64252 358872 64258
rect 358820 64194 358872 64200
rect 356058 50688 356114 50697
rect 356058 50623 356114 50632
rect 356072 16574 356100 50623
rect 357440 32564 357492 32570
rect 357440 32506 357492 32512
rect 350552 16546 351224 16574
rect 351932 16546 352880 16574
rect 353312 16546 353616 16574
rect 354692 16546 355272 16574
rect 356072 16546 356376 16574
rect 349252 11892 349304 11898
rect 349252 11834 349304 11840
rect 349264 3398 349292 11834
rect 349252 3392 349304 3398
rect 349252 3334 349304 3340
rect 350448 3392 350500 3398
rect 350448 3334 350500 3340
rect 349172 3182 349292 3210
rect 349264 480 349292 3182
rect 350460 480 350488 3334
rect 345726 354 345838 480
rect 345308 326 345838 354
rect 345726 -960 345838 326
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351196 354 351224 16546
rect 352852 480 352880 16546
rect 351614 354 351726 480
rect 351196 326 351726 354
rect 351614 -960 351726 326
rect 352810 -960 352922 480
rect 353588 354 353616 16546
rect 355244 480 355272 16546
rect 356348 480 356376 16546
rect 357452 3210 357480 32506
rect 357532 18828 357584 18834
rect 357532 18770 357584 18776
rect 357544 3398 357572 18770
rect 358832 16574 358860 64194
rect 362958 58712 363014 58721
rect 362958 58647 363014 58656
rect 361580 43580 361632 43586
rect 361580 43522 361632 43528
rect 361592 16574 361620 43522
rect 362972 16574 363000 58647
rect 364982 54632 365038 54641
rect 364982 54567 365038 54576
rect 358832 16546 359504 16574
rect 361592 16546 361896 16574
rect 362972 16546 363552 16574
rect 357532 3392 357584 3398
rect 357532 3334 357584 3340
rect 358728 3392 358780 3398
rect 358728 3334 358780 3340
rect 357452 3182 357572 3210
rect 357544 480 357572 3182
rect 358740 480 358768 3334
rect 354006 354 354118 480
rect 353588 326 354118 354
rect 354006 -960 354118 326
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359476 354 359504 16546
rect 361120 16040 361172 16046
rect 361120 15982 361172 15988
rect 361132 480 361160 15982
rect 359894 354 360006 480
rect 359476 326 360006 354
rect 359894 -960 360006 326
rect 361090 -960 361202 480
rect 361868 354 361896 16546
rect 363524 480 363552 16546
rect 364616 15972 364668 15978
rect 364616 15914 364668 15920
rect 364628 480 364656 15914
rect 364996 3398 365024 54567
rect 365812 29776 365864 29782
rect 365812 29718 365864 29724
rect 364984 3392 365036 3398
rect 364984 3334 365036 3340
rect 365824 480 365852 29718
rect 367112 16574 367140 70994
rect 369858 52184 369914 52193
rect 369858 52119 369914 52128
rect 368480 50380 368532 50386
rect 368480 50322 368532 50328
rect 368492 16574 368520 50322
rect 369872 16574 369900 52119
rect 373998 52048 374054 52057
rect 373998 51983 374054 51992
rect 372620 38140 372672 38146
rect 372620 38082 372672 38088
rect 372632 16574 372660 38082
rect 367112 16546 367784 16574
rect 368492 16546 369440 16574
rect 369872 16546 370176 16574
rect 372632 16546 372936 16574
rect 367008 3392 367060 3398
rect 367008 3334 367060 3340
rect 367020 480 367048 3334
rect 362286 354 362398 480
rect 361868 326 362398 354
rect 362286 -960 362398 326
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 367756 354 367784 16546
rect 369412 480 369440 16546
rect 368174 354 368286 480
rect 367756 326 368286 354
rect 368174 -960 368286 326
rect 369370 -960 369482 480
rect 370148 354 370176 16546
rect 371700 9172 371752 9178
rect 371700 9114 371752 9120
rect 371712 480 371740 9114
rect 372908 480 372936 16546
rect 374012 1170 374040 51983
rect 374092 27124 374144 27130
rect 374092 27066 374144 27072
rect 374104 3398 374132 27066
rect 375392 16574 375420 72422
rect 376772 16574 376800 79018
rect 380898 65512 380954 65521
rect 380898 65447 380954 65456
rect 379520 20052 379572 20058
rect 379520 19994 379572 20000
rect 375392 16546 376064 16574
rect 376772 16546 377720 16574
rect 374092 3392 374144 3398
rect 374092 3334 374144 3340
rect 375288 3392 375340 3398
rect 375288 3334 375340 3340
rect 374012 1142 374132 1170
rect 374104 480 374132 1142
rect 375300 480 375328 3334
rect 370566 354 370678 480
rect 370148 326 370678 354
rect 370566 -960 370678 326
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376036 354 376064 16546
rect 377692 480 377720 16546
rect 378876 7812 378928 7818
rect 378876 7754 378928 7760
rect 378888 480 378916 7754
rect 376454 354 376566 480
rect 376036 326 376566 354
rect 376454 -960 376566 326
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379532 354 379560 19994
rect 380912 16574 380940 65447
rect 380912 16546 381216 16574
rect 381188 480 381216 16546
rect 382292 3398 382320 79455
rect 448520 79348 448572 79354
rect 448520 79290 448572 79296
rect 393320 78056 393372 78062
rect 393320 77998 393372 78004
rect 389180 76560 389232 76566
rect 389180 76502 389232 76508
rect 382922 61704 382978 61713
rect 382922 61639 382978 61648
rect 382372 5024 382424 5030
rect 382372 4966 382424 4972
rect 382280 3392 382332 3398
rect 382280 3334 382332 3340
rect 382384 480 382412 4966
rect 382936 3194 382964 61639
rect 387798 53272 387854 53281
rect 387798 53207 387854 53216
rect 385040 33992 385092 33998
rect 385040 33934 385092 33940
rect 385052 16574 385080 33934
rect 385052 16546 386000 16574
rect 383568 3392 383620 3398
rect 383568 3334 383620 3340
rect 382924 3188 382976 3194
rect 382924 3130 382976 3136
rect 383580 480 383608 3334
rect 384764 3188 384816 3194
rect 384764 3130 384816 3136
rect 384776 480 384804 3130
rect 385972 480 386000 16546
rect 386696 10464 386748 10470
rect 386696 10406 386748 10412
rect 379950 354 380062 480
rect 379532 326 380062 354
rect 379950 -960 380062 326
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 386708 354 386736 10406
rect 387126 354 387238 480
rect 386708 326 387238 354
rect 387812 354 387840 53207
rect 389192 16574 389220 76502
rect 390558 47696 390614 47705
rect 390558 47631 390614 47640
rect 389192 16546 389496 16574
rect 389468 480 389496 16546
rect 390572 3398 390600 47631
rect 391940 25764 391992 25770
rect 391940 25706 391992 25712
rect 391952 16574 391980 25706
rect 393332 16574 393360 77998
rect 400864 77988 400916 77994
rect 400864 77930 400916 77936
rect 396080 60104 396132 60110
rect 396080 60046 396132 60052
rect 394700 55888 394752 55894
rect 394700 55830 394752 55836
rect 394712 16574 394740 55830
rect 391952 16546 392624 16574
rect 393332 16546 394280 16574
rect 394712 16546 395384 16574
rect 390652 7744 390704 7750
rect 390652 7686 390704 7692
rect 390560 3392 390612 3398
rect 390560 3334 390612 3340
rect 390664 480 390692 7686
rect 391848 3392 391900 3398
rect 391848 3334 391900 3340
rect 391860 480 391888 3334
rect 388230 354 388342 480
rect 387812 326 388342 354
rect 387126 -960 387238 326
rect 388230 -960 388342 326
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 392596 354 392624 16546
rect 394252 480 394280 16546
rect 395356 480 395384 16546
rect 393014 354 393126 480
rect 392596 326 393126 354
rect 393014 -960 393126 326
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396092 354 396120 60046
rect 398840 60036 398892 60042
rect 398840 59978 398892 59984
rect 397460 28416 397512 28422
rect 397460 28358 397512 28364
rect 397472 16574 397500 28358
rect 397472 16546 397776 16574
rect 397748 480 397776 16546
rect 398852 3210 398880 59978
rect 400876 15978 400904 77930
rect 412640 69760 412692 69766
rect 412640 69702 412692 69708
rect 402980 67720 403032 67726
rect 402980 67662 403032 67668
rect 400954 56128 401010 56137
rect 400954 56063 401010 56072
rect 400864 15972 400916 15978
rect 400864 15914 400916 15920
rect 398932 13184 398984 13190
rect 398932 13126 398984 13132
rect 398944 3398 398972 13126
rect 400968 3398 400996 56063
rect 402992 16574 403020 67662
rect 405738 50552 405794 50561
rect 405738 50487 405794 50496
rect 405752 16574 405780 50487
rect 408498 44840 408554 44849
rect 408498 44775 408554 44784
rect 408512 16574 408540 44775
rect 409880 24336 409932 24342
rect 409880 24278 409932 24284
rect 409892 16574 409920 24278
rect 402992 16546 403664 16574
rect 405752 16546 406056 16574
rect 408512 16546 409184 16574
rect 409892 16546 410840 16574
rect 401324 3868 401376 3874
rect 401324 3810 401376 3816
rect 398932 3392 398984 3398
rect 398932 3334 398984 3340
rect 400128 3392 400180 3398
rect 400128 3334 400180 3340
rect 400956 3392 401008 3398
rect 400956 3334 401008 3340
rect 398852 3182 398972 3210
rect 398944 480 398972 3182
rect 400140 480 400168 3334
rect 401336 480 401364 3810
rect 402520 3392 402572 3398
rect 402520 3334 402572 3340
rect 402532 480 402560 3334
rect 403636 480 403664 16546
rect 404820 9104 404872 9110
rect 404820 9046 404872 9052
rect 404832 480 404860 9046
rect 406028 480 406056 16546
rect 407212 14612 407264 14618
rect 407212 14554 407264 14560
rect 407120 14544 407172 14550
rect 407120 14486 407172 14492
rect 407132 3210 407160 14486
rect 407224 3398 407252 14554
rect 407212 3392 407264 3398
rect 407212 3334 407264 3340
rect 408408 3392 408460 3398
rect 408408 3334 408460 3340
rect 407132 3182 407252 3210
rect 407224 480 407252 3182
rect 408420 480 408448 3334
rect 396510 354 396622 480
rect 396092 326 396622 354
rect 396510 -960 396622 326
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409156 354 409184 16546
rect 410812 480 410840 16546
rect 411904 6316 411956 6322
rect 411904 6258 411956 6264
rect 411916 480 411944 6258
rect 409574 354 409686 480
rect 409156 326 409686 354
rect 409574 -960 409686 326
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 412652 354 412680 69702
rect 423678 67144 423734 67153
rect 423678 67079 423734 67088
rect 414662 63064 414718 63073
rect 414662 62999 414718 63008
rect 414296 6248 414348 6254
rect 414296 6190 414348 6196
rect 414308 480 414336 6190
rect 414676 3398 414704 62999
rect 418802 57352 418858 57361
rect 418802 57287 418858 57296
rect 418160 35352 418212 35358
rect 418160 35294 418212 35300
rect 416780 22908 416832 22914
rect 416780 22850 416832 22856
rect 415492 17468 415544 17474
rect 415492 17410 415544 17416
rect 414664 3392 414716 3398
rect 414664 3334 414716 3340
rect 415504 480 415532 17410
rect 416792 16574 416820 22850
rect 418172 16574 418200 35294
rect 416792 16546 417464 16574
rect 418172 16546 418568 16574
rect 416688 3392 416740 3398
rect 416688 3334 416740 3340
rect 416700 480 416728 3334
rect 413070 354 413182 480
rect 412652 326 413182 354
rect 413070 -960 413182 326
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417436 354 417464 16546
rect 417854 354 417966 480
rect 417436 326 417966 354
rect 418540 354 418568 16546
rect 418816 3398 418844 57287
rect 420920 31204 420972 31210
rect 420920 31146 420972 31152
rect 418804 3392 418856 3398
rect 418804 3334 418856 3340
rect 420184 3392 420236 3398
rect 420184 3334 420236 3340
rect 420196 480 420224 3334
rect 418958 354 419070 480
rect 418540 326 419070 354
rect 417854 -960 417966 326
rect 418958 -960 419070 326
rect 420154 -960 420266 480
rect 420932 354 420960 31146
rect 422300 21412 422352 21418
rect 422300 21354 422352 21360
rect 422312 16574 422340 21354
rect 422312 16546 422616 16574
rect 422588 480 422616 16546
rect 423692 3398 423720 67079
rect 430578 67008 430634 67017
rect 430578 66943 430634 66952
rect 423770 54496 423826 54505
rect 423770 54431 423826 54440
rect 423680 3392 423732 3398
rect 423680 3334 423732 3340
rect 423784 480 423812 54431
rect 426440 43512 426492 43518
rect 426440 43454 426492 43460
rect 425060 27056 425112 27062
rect 425060 26998 425112 27004
rect 425072 16574 425100 26998
rect 426452 16574 426480 43454
rect 427820 40860 427872 40866
rect 427820 40802 427872 40808
rect 427832 16574 427860 40802
rect 430592 16574 430620 66943
rect 437478 61568 437534 61577
rect 437478 61503 437534 61512
rect 432602 53136 432658 53145
rect 432602 53071 432658 53080
rect 431960 18760 432012 18766
rect 431960 18702 432012 18708
rect 425072 16546 425744 16574
rect 426452 16546 426848 16574
rect 427832 16546 428504 16574
rect 430592 16546 430896 16574
rect 424968 3392 425020 3398
rect 424968 3334 425020 3340
rect 424980 480 425008 3334
rect 421350 354 421462 480
rect 420932 326 421462 354
rect 421350 -960 421462 326
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 425716 354 425744 16546
rect 426134 354 426246 480
rect 425716 326 426246 354
rect 426820 354 426848 16546
rect 428476 480 428504 16546
rect 429660 4956 429712 4962
rect 429660 4898 429712 4904
rect 429672 480 429700 4898
rect 430868 480 430896 16546
rect 431972 3330 432000 18702
rect 432052 15904 432104 15910
rect 432052 15846 432104 15852
rect 431960 3324 432012 3330
rect 431960 3266 432012 3272
rect 432064 480 432092 15846
rect 432616 3398 432644 53071
rect 436100 25696 436152 25702
rect 436100 25638 436152 25644
rect 436112 16574 436140 25638
rect 436112 16546 436784 16574
rect 435088 10396 435140 10402
rect 435088 10338 435140 10344
rect 432604 3392 432656 3398
rect 432604 3334 432656 3340
rect 434444 3392 434496 3398
rect 434444 3334 434496 3340
rect 433248 3324 433300 3330
rect 433248 3266 433300 3272
rect 433260 480 433288 3266
rect 434456 480 434484 3334
rect 427238 354 427350 480
rect 426820 326 427350 354
rect 426134 -960 426246 326
rect 427238 -960 427350 326
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435100 354 435128 10338
rect 436756 480 436784 16546
rect 435518 354 435630 480
rect 435100 326 435630 354
rect 435518 -960 435630 326
rect 436714 -960 436826 480
rect 437492 354 437520 61503
rect 440238 50416 440294 50425
rect 440238 50351 440294 50360
rect 439136 11824 439188 11830
rect 439136 11766 439188 11772
rect 439148 480 439176 11766
rect 440252 3398 440280 50351
rect 444380 47660 444432 47666
rect 444380 47602 444432 47608
rect 440332 36712 440384 36718
rect 440332 36654 440384 36660
rect 440240 3392 440292 3398
rect 440240 3334 440292 3340
rect 440344 480 440372 36654
rect 441620 29708 441672 29714
rect 441620 29650 441672 29656
rect 441632 16574 441660 29650
rect 443000 24268 443052 24274
rect 443000 24210 443052 24216
rect 443012 16574 443040 24210
rect 444392 16574 444420 47602
rect 445760 17400 445812 17406
rect 445760 17342 445812 17348
rect 441632 16546 442672 16574
rect 443012 16546 443408 16574
rect 444392 16546 445064 16574
rect 441528 3392 441580 3398
rect 441528 3334 441580 3340
rect 441540 480 441568 3334
rect 442644 480 442672 16546
rect 437910 354 438022 480
rect 437492 326 438022 354
rect 437910 -960 438022 326
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443380 354 443408 16546
rect 445036 480 445064 16546
rect 443798 354 443910 480
rect 443380 326 443910 354
rect 443798 -960 443910 326
rect 444994 -960 445106 480
rect 445772 354 445800 17342
rect 447416 3800 447468 3806
rect 447416 3742 447468 3748
rect 447428 480 447456 3742
rect 448532 3210 448560 79290
rect 483020 79008 483072 79014
rect 483020 78950 483072 78956
rect 468574 77616 468630 77625
rect 468574 77551 468630 77560
rect 453304 75336 453356 75342
rect 453304 75278 453356 75284
rect 450542 55992 450598 56001
rect 450542 55927 450598 55936
rect 449900 46232 449952 46238
rect 449900 46174 449952 46180
rect 448612 17332 448664 17338
rect 448612 17274 448664 17280
rect 448624 3398 448652 17274
rect 449912 16574 449940 46174
rect 449912 16546 450492 16574
rect 450464 3482 450492 16546
rect 450556 4146 450584 55927
rect 452658 43480 452714 43489
rect 452658 43415 452714 43424
rect 452672 6914 452700 43415
rect 453316 16574 453344 75278
rect 465172 73908 465224 73914
rect 465172 73850 465224 73856
rect 456800 73840 456852 73846
rect 456800 73782 456852 73788
rect 454682 49192 454738 49201
rect 454682 49127 454738 49136
rect 453316 16546 453436 16574
rect 452672 6886 453344 6914
rect 450544 4140 450596 4146
rect 450544 4082 450596 4088
rect 451004 4140 451056 4146
rect 451004 4082 451056 4088
rect 450464 3454 450952 3482
rect 448612 3392 448664 3398
rect 448612 3334 448664 3340
rect 449808 3392 449860 3398
rect 449808 3334 449860 3340
rect 448532 3182 448652 3210
rect 448624 480 448652 3182
rect 449820 480 449848 3334
rect 450924 480 450952 3454
rect 451016 3194 451044 4082
rect 451004 3188 451056 3194
rect 451004 3130 451056 3136
rect 452108 3188 452160 3194
rect 452108 3130 452160 3136
rect 452120 480 452148 3130
rect 453316 480 453344 6886
rect 453408 3806 453436 16546
rect 453396 3800 453448 3806
rect 453396 3742 453448 3748
rect 454500 3732 454552 3738
rect 454500 3674 454552 3680
rect 454512 480 454540 3674
rect 454696 2922 454724 49127
rect 456812 3398 456840 73782
rect 464344 68332 464396 68338
rect 464344 68274 464396 68280
rect 459558 61432 459614 61441
rect 459558 61367 459614 61376
rect 458180 45008 458232 45014
rect 458180 44950 458232 44956
rect 458192 16574 458220 44950
rect 459572 16574 459600 61367
rect 463698 46336 463754 46345
rect 463698 46271 463754 46280
rect 462320 40792 462372 40798
rect 462320 40734 462372 40740
rect 460940 22840 460992 22846
rect 460940 22782 460992 22788
rect 460952 16574 460980 22782
rect 458192 16546 459232 16574
rect 459572 16546 459968 16574
rect 460952 16546 461624 16574
rect 456892 9036 456944 9042
rect 456892 8978 456944 8984
rect 456800 3392 456852 3398
rect 456800 3334 456852 3340
rect 454684 2916 454736 2922
rect 454684 2858 454736 2864
rect 455696 2916 455748 2922
rect 455696 2858 455748 2864
rect 455708 480 455736 2858
rect 456904 480 456932 8978
rect 458088 3392 458140 3398
rect 458088 3334 458140 3340
rect 458100 480 458128 3334
rect 459204 480 459232 16546
rect 446190 354 446302 480
rect 445772 326 446302 354
rect 446190 -960 446302 326
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 459940 354 459968 16546
rect 461596 480 461624 16546
rect 460358 354 460470 480
rect 459940 326 460470 354
rect 460358 -960 460470 326
rect 461554 -960 461666 480
rect 462332 354 462360 40734
rect 463712 16574 463740 46271
rect 463712 16546 464016 16574
rect 463988 480 464016 16546
rect 464356 3398 464384 68274
rect 464344 3392 464396 3398
rect 464344 3334 464396 3340
rect 465184 480 465212 73850
rect 467840 58676 467892 58682
rect 467840 58618 467892 58624
rect 466460 31136 466512 31142
rect 466460 31078 466512 31084
rect 466472 16574 466500 31078
rect 467852 16574 467880 58618
rect 468588 54534 468616 77551
rect 472624 64184 472676 64190
rect 472624 64126 472676 64132
rect 468484 54528 468536 54534
rect 468484 54470 468536 54476
rect 468576 54528 468628 54534
rect 468576 54470 468628 54476
rect 466472 16546 467512 16574
rect 467852 16546 468248 16574
rect 466276 3392 466328 3398
rect 466276 3334 466328 3340
rect 466288 480 466316 3334
rect 467484 480 467512 16546
rect 462750 354 462862 480
rect 462332 326 462862 354
rect 462750 -960 462862 326
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468220 354 468248 16546
rect 468496 3398 468524 54470
rect 470600 39500 470652 39506
rect 470600 39442 470652 39448
rect 468484 3392 468536 3398
rect 468484 3334 468536 3340
rect 469864 3392 469916 3398
rect 469864 3334 469916 3340
rect 469876 480 469904 3334
rect 468638 354 468750 480
rect 468220 326 468750 354
rect 468638 -960 468750 326
rect 469834 -960 469946 480
rect 470612 354 470640 39442
rect 471980 21616 472032 21622
rect 471980 21558 472032 21564
rect 471992 16574 472020 21558
rect 471992 16546 472296 16574
rect 472268 480 472296 16546
rect 472636 3398 472664 64126
rect 473452 57248 473504 57254
rect 473452 57190 473504 57196
rect 473464 16574 473492 57190
rect 476118 51912 476174 51921
rect 476118 51847 476174 51856
rect 474740 33924 474792 33930
rect 474740 33866 474792 33872
rect 474752 16574 474780 33866
rect 476132 16574 476160 51847
rect 481640 39432 481692 39438
rect 481640 39374 481692 39380
rect 477500 28348 477552 28354
rect 477500 28290 477552 28296
rect 477512 16574 477540 28290
rect 481652 16574 481680 39374
rect 483032 16574 483060 78950
rect 500960 78940 501012 78946
rect 500960 78882 501012 78888
rect 486422 75440 486478 75449
rect 486422 75375 486478 75384
rect 484398 51776 484454 51785
rect 484398 51711 484454 51720
rect 484412 16574 484440 51711
rect 486436 16574 486464 75375
rect 498200 69692 498252 69698
rect 498200 69634 498252 69640
rect 489918 55856 489974 55865
rect 489918 55791 489974 55800
rect 488540 38072 488592 38078
rect 488540 38014 488592 38020
rect 488552 16574 488580 38014
rect 473464 16546 474136 16574
rect 474752 16546 475792 16574
rect 476132 16546 476528 16574
rect 477512 16546 478184 16574
rect 481652 16546 481772 16574
rect 483032 16546 484072 16574
rect 484412 16546 484808 16574
rect 486436 16546 486556 16574
rect 488552 16546 488856 16574
rect 472624 3392 472676 3398
rect 472624 3334 472676 3340
rect 473452 3392 473504 3398
rect 473452 3334 473504 3340
rect 473464 480 473492 3334
rect 471030 354 471142 480
rect 470612 326 471142 354
rect 471030 -960 471142 326
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474108 354 474136 16546
rect 475764 480 475792 16546
rect 474526 354 474638 480
rect 474108 326 474638 354
rect 474526 -960 474638 326
rect 475722 -960 475834 480
rect 476500 354 476528 16546
rect 478156 480 478184 16546
rect 478880 15972 478932 15978
rect 478880 15914 478932 15920
rect 476918 354 477030 480
rect 476500 326 477030 354
rect 476918 -960 477030 326
rect 478114 -960 478226 480
rect 478892 354 478920 15914
rect 480536 3664 480588 3670
rect 480536 3606 480588 3612
rect 480548 480 480576 3606
rect 481744 480 481772 16546
rect 482836 7676 482888 7682
rect 482836 7618 482888 7624
rect 482848 480 482876 7618
rect 484044 480 484072 16546
rect 479310 354 479422 480
rect 478892 326 479422 354
rect 479310 -960 479422 326
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 484780 354 484808 16546
rect 486424 4888 486476 4894
rect 486424 4830 486476 4836
rect 486436 480 486464 4830
rect 486528 3670 486556 16546
rect 486516 3664 486568 3670
rect 486516 3606 486568 3612
rect 487620 3596 487672 3602
rect 487620 3538 487672 3544
rect 487632 480 487660 3538
rect 488828 480 488856 16546
rect 489932 3602 489960 55791
rect 494058 49056 494114 49065
rect 494058 48991 494114 49000
rect 491300 35284 491352 35290
rect 491300 35226 491352 35232
rect 490012 33856 490064 33862
rect 490012 33798 490064 33804
rect 489920 3596 489972 3602
rect 489920 3538 489972 3544
rect 490024 3482 490052 33798
rect 491312 16574 491340 35226
rect 494072 16574 494100 48991
rect 495438 46200 495494 46209
rect 495438 46135 495494 46144
rect 491312 16546 492352 16574
rect 494072 16546 494744 16574
rect 490748 3596 490800 3602
rect 490748 3538 490800 3544
rect 489932 3454 490052 3482
rect 489932 480 489960 3454
rect 485198 354 485310 480
rect 484780 326 485310 354
rect 485198 -960 485310 326
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 490760 354 490788 3538
rect 492324 480 492352 16546
rect 493048 13116 493100 13122
rect 493048 13058 493100 13064
rect 491086 354 491198 480
rect 490760 326 491198 354
rect 491086 -960 491198 326
rect 492282 -960 492394 480
rect 493060 354 493088 13058
rect 494716 480 494744 16546
rect 493478 354 493590 480
rect 493060 326 493590 354
rect 493478 -960 493590 326
rect 494674 -960 494786 480
rect 495452 354 495480 46135
rect 497096 3800 497148 3806
rect 497096 3742 497148 3748
rect 497108 480 497136 3742
rect 498212 480 498240 69634
rect 499580 49020 499632 49026
rect 499580 48962 499632 48968
rect 498292 42152 498344 42158
rect 498292 42094 498344 42100
rect 498304 16574 498332 42094
rect 499592 16574 499620 48962
rect 500972 16574 501000 78882
rect 523132 78872 523184 78878
rect 523132 78814 523184 78820
rect 521658 75304 521714 75313
rect 506480 75268 506532 75274
rect 521658 75239 521714 75248
rect 506480 75210 506532 75216
rect 504362 68232 504418 68241
rect 504362 68167 504418 68176
rect 502340 43444 502392 43450
rect 502340 43386 502392 43392
rect 502352 16574 502380 43386
rect 503720 17264 503772 17270
rect 503720 17206 503772 17212
rect 498304 16546 498976 16574
rect 499592 16546 500632 16574
rect 500972 16546 501368 16574
rect 502352 16546 503024 16574
rect 495870 354 495982 480
rect 495452 326 495982 354
rect 495870 -960 495982 326
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 498948 354 498976 16546
rect 500604 480 500632 16546
rect 499366 354 499478 480
rect 498948 326 499478 354
rect 499366 -960 499478 326
rect 500562 -960 500674 480
rect 501340 354 501368 16546
rect 502996 480 503024 16546
rect 501758 354 501870 480
rect 501340 326 501870 354
rect 501758 -960 501870 326
rect 502954 -960 503066 480
rect 503732 354 503760 17206
rect 504376 3602 504404 68167
rect 506492 3602 506520 75210
rect 511264 75200 511316 75206
rect 511264 75142 511316 75148
rect 507858 42120 507914 42129
rect 507858 42055 507914 42064
rect 506572 29640 506624 29646
rect 506572 29582 506624 29588
rect 504364 3596 504416 3602
rect 504364 3538 504416 3544
rect 505376 3596 505428 3602
rect 505376 3538 505428 3544
rect 506480 3596 506532 3602
rect 506480 3538 506532 3544
rect 505388 480 505416 3538
rect 506584 3482 506612 29582
rect 507872 16574 507900 42055
rect 509240 28280 509292 28286
rect 509240 28222 509292 28228
rect 509252 16574 509280 28222
rect 511276 16574 511304 75142
rect 511998 64288 512054 64297
rect 511998 64223 512054 64232
rect 507872 16546 508912 16574
rect 509252 16546 509648 16574
rect 511276 16546 511396 16574
rect 507308 3596 507360 3602
rect 507308 3538 507360 3544
rect 506492 3454 506612 3482
rect 506492 480 506520 3454
rect 504150 354 504262 480
rect 503732 326 504262 354
rect 504150 -960 504262 326
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507320 354 507348 3538
rect 508884 480 508912 16546
rect 507646 354 507758 480
rect 507320 326 507758 354
rect 507646 -960 507758 326
rect 508842 -960 508954 480
rect 509620 354 509648 16546
rect 511264 14476 511316 14482
rect 511264 14418 511316 14424
rect 511276 480 511304 14418
rect 511368 3194 511396 16546
rect 511356 3188 511408 3194
rect 511356 3130 511408 3136
rect 510038 354 510150 480
rect 509620 326 510150 354
rect 510038 -960 510150 326
rect 511234 -960 511346 480
rect 512012 354 512040 64223
rect 514022 62928 514078 62937
rect 514022 62863 514078 62872
rect 513380 26988 513432 26994
rect 513380 26930 513432 26936
rect 512430 354 512542 480
rect 512012 326 512542 354
rect 513392 354 513420 26930
rect 514036 3058 514064 62863
rect 520922 47560 520978 47569
rect 520922 47495 520978 47504
rect 516140 40724 516192 40730
rect 516140 40666 516192 40672
rect 516152 16574 516180 40666
rect 520280 25628 520332 25634
rect 520280 25570 520332 25576
rect 518900 19984 518952 19990
rect 518900 19926 518952 19932
rect 518912 16574 518940 19926
rect 516152 16546 517192 16574
rect 518912 16546 519584 16574
rect 514760 3188 514812 3194
rect 514760 3130 514812 3136
rect 514024 3052 514076 3058
rect 514024 2994 514076 3000
rect 514772 480 514800 3130
rect 515956 3052 516008 3058
rect 515956 2994 516008 3000
rect 515968 480 515996 2994
rect 517164 480 517192 16546
rect 518348 3664 518400 3670
rect 518348 3606 518400 3612
rect 518360 480 518388 3606
rect 519556 480 519584 16546
rect 513534 354 513646 480
rect 513392 326 513646 354
rect 512430 -960 512542 326
rect 513534 -960 513646 326
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520292 354 520320 25570
rect 520936 3602 520964 47495
rect 520924 3596 520976 3602
rect 520924 3538 520976 3544
rect 520710 354 520822 480
rect 520292 326 520822 354
rect 521672 354 521700 75239
rect 523144 6914 523172 78814
rect 525800 78804 525852 78810
rect 525800 78746 525852 78752
rect 525062 59936 525118 59945
rect 525062 59871 525118 59880
rect 523052 6886 523172 6914
rect 523052 480 523080 6886
rect 525076 3602 525104 59871
rect 525812 16574 525840 78746
rect 536840 78736 536892 78742
rect 536840 78678 536892 78684
rect 529940 69080 529992 69086
rect 529940 69022 529992 69028
rect 528560 38004 528612 38010
rect 528560 37946 528612 37952
rect 527180 24200 527232 24206
rect 527180 24142 527232 24148
rect 527192 16574 527220 24142
rect 525812 16546 526208 16574
rect 527192 16546 527864 16574
rect 525432 6180 525484 6186
rect 525432 6122 525484 6128
rect 524236 3596 524288 3602
rect 524236 3538 524288 3544
rect 525064 3596 525116 3602
rect 525064 3538 525116 3544
rect 524248 480 524276 3538
rect 525444 480 525472 6122
rect 521814 354 521926 480
rect 521672 326 521926 354
rect 520710 -960 520822 326
rect 521814 -960 521926 326
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526180 354 526208 16546
rect 527836 480 527864 16546
rect 526598 354 526710 480
rect 526180 326 526710 354
rect 526598 -960 526710 326
rect 527794 -960 527906 480
rect 528572 354 528600 37946
rect 528990 354 529102 480
rect 528572 326 529102 354
rect 529952 354 529980 69022
rect 534080 39364 534132 39370
rect 534080 39306 534132 39312
rect 531412 32496 531464 32502
rect 531412 32438 531464 32444
rect 531424 16574 531452 32438
rect 534092 16574 534120 39306
rect 535460 26920 535512 26926
rect 535460 26862 535512 26868
rect 535472 16574 535500 26862
rect 536852 16574 536880 78678
rect 553398 76528 553454 76537
rect 553398 76463 553454 76472
rect 549258 75168 549314 75177
rect 549258 75103 549314 75112
rect 543738 71088 543794 71097
rect 543738 71023 543794 71032
rect 539690 58576 539746 58585
rect 539690 58511 539746 58520
rect 538864 42084 538916 42090
rect 538864 42026 538916 42032
rect 538220 22772 538272 22778
rect 538220 22714 538272 22720
rect 531424 16546 532096 16574
rect 534092 16546 534488 16574
rect 535472 16546 536144 16574
rect 536852 16546 537248 16574
rect 531320 3528 531372 3534
rect 531320 3470 531372 3476
rect 531332 480 531360 3470
rect 530094 354 530206 480
rect 529952 326 530206 354
rect 528990 -960 529102 326
rect 530094 -960 530206 326
rect 531290 -960 531402 480
rect 532068 354 532096 16546
rect 533712 3596 533764 3602
rect 533712 3538 533764 3544
rect 533724 480 533752 3538
rect 532486 354 532598 480
rect 532068 326 532598 354
rect 532486 -960 532598 326
rect 533682 -960 533794 480
rect 534460 354 534488 16546
rect 536116 480 536144 16546
rect 537220 480 537248 16546
rect 534878 354 534990 480
rect 534460 326 534990 354
rect 534878 -960 534990 326
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538232 354 538260 22714
rect 538876 3534 538904 42026
rect 539704 16574 539732 58511
rect 542360 47592 542412 47598
rect 542360 47534 542412 47540
rect 542372 16574 542400 47534
rect 543752 16574 543780 71023
rect 547878 64152 547934 64161
rect 547878 64087 547934 64096
rect 545762 57216 545818 57225
rect 545762 57151 545818 57160
rect 539704 16546 540376 16574
rect 542372 16546 542768 16574
rect 543752 16546 544424 16574
rect 538864 3528 538916 3534
rect 538864 3470 538916 3476
rect 539600 3528 539652 3534
rect 539600 3470 539652 3476
rect 539612 480 539640 3470
rect 538374 354 538486 480
rect 538232 326 538486 354
rect 538374 -960 538486 326
rect 539570 -960 539682 480
rect 540348 354 540376 16546
rect 541992 4820 542044 4826
rect 541992 4762 542044 4768
rect 542004 480 542032 4762
rect 540766 354 540878 480
rect 540348 326 540878 354
rect 540766 -960 540878 326
rect 541962 -960 542074 480
rect 542740 354 542768 16546
rect 544396 480 544424 16546
rect 545488 7608 545540 7614
rect 545488 7550 545540 7556
rect 545500 480 545528 7550
rect 545776 3534 545804 57151
rect 546500 25560 546552 25566
rect 546500 25502 546552 25508
rect 545764 3528 545816 3534
rect 545764 3470 545816 3476
rect 543158 354 543270 480
rect 542740 326 543270 354
rect 543158 -960 543270 326
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546512 354 546540 25502
rect 547892 480 547920 64087
rect 549272 16574 549300 75103
rect 552664 67652 552716 67658
rect 552664 67594 552716 67600
rect 552020 37936 552072 37942
rect 552020 37878 552072 37884
rect 549272 16546 550312 16574
rect 548616 11756 548668 11762
rect 548616 11698 548668 11704
rect 546654 354 546766 480
rect 546512 326 546766 354
rect 546654 -960 546766 326
rect 547850 -960 547962 480
rect 548628 354 548656 11698
rect 550284 480 550312 16546
rect 552032 6914 552060 37878
rect 552676 16574 552704 67594
rect 553412 16574 553440 76463
rect 561678 69592 561734 69601
rect 561678 69527 561734 69536
rect 557538 66872 557594 66881
rect 557538 66807 557594 66816
rect 556160 53100 556212 53106
rect 556160 53042 556212 53048
rect 554780 31068 554832 31074
rect 554780 31010 554832 31016
rect 552676 16546 552796 16574
rect 553412 16546 553808 16574
rect 552032 6886 552704 6914
rect 551468 3528 551520 3534
rect 551468 3470 551520 3476
rect 551480 480 551508 3470
rect 552676 480 552704 6886
rect 552768 3534 552796 16546
rect 552756 3528 552808 3534
rect 552756 3470 552808 3476
rect 553780 480 553808 16546
rect 549046 354 549158 480
rect 548628 326 549158 354
rect 549046 -960 549158 326
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554792 354 554820 31010
rect 556172 16574 556200 53042
rect 557552 16574 557580 66807
rect 560300 44940 560352 44946
rect 560300 44882 560352 44888
rect 558920 36644 558972 36650
rect 558920 36586 558972 36592
rect 558932 16574 558960 36586
rect 560312 16574 560340 44882
rect 561692 16574 561720 69527
rect 574744 64932 574796 64938
rect 574744 64874 574796 64880
rect 567842 62792 567898 62801
rect 567842 62727 567898 62736
rect 565818 48920 565874 48929
rect 565818 48855 565874 48864
rect 563704 33788 563756 33794
rect 563704 33730 563756 33736
rect 556172 16546 556936 16574
rect 557552 16546 558592 16574
rect 558932 16546 559328 16574
rect 560312 16546 560432 16574
rect 561692 16546 562088 16574
rect 556160 8968 556212 8974
rect 556160 8910 556212 8916
rect 556172 480 556200 8910
rect 554934 354 555046 480
rect 554792 326 555046 354
rect 554934 -960 555046 326
rect 556130 -960 556242 480
rect 556908 354 556936 16546
rect 558564 480 558592 16546
rect 557326 354 557438 480
rect 556908 326 557438 354
rect 557326 -960 557438 326
rect 558522 -960 558634 480
rect 559300 354 559328 16546
rect 559718 354 559830 480
rect 559300 326 559830 354
rect 560404 354 560432 16546
rect 562060 480 562088 16546
rect 563060 10328 563112 10334
rect 563060 10270 563112 10276
rect 560822 354 560934 480
rect 560404 326 560934 354
rect 559718 -960 559830 326
rect 560822 -960 560934 326
rect 562018 -960 562130 480
rect 563072 354 563100 10270
rect 563716 3058 563744 33730
rect 564532 24132 564584 24138
rect 564532 24074 564584 24080
rect 564544 6914 564572 24074
rect 565832 16574 565860 48855
rect 567200 18692 567252 18698
rect 567200 18634 567252 18640
rect 567212 16574 567240 18634
rect 565832 16546 566872 16574
rect 567212 16546 567608 16574
rect 564452 6886 564572 6914
rect 563704 3052 563756 3058
rect 563704 2994 563756 3000
rect 564452 480 564480 6886
rect 565636 3052 565688 3058
rect 565636 2994 565688 3000
rect 565648 480 565676 2994
rect 566844 480 566872 16546
rect 563214 354 563326 480
rect 563072 326 563326 354
rect 563214 -960 563326 326
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567580 354 567608 16546
rect 567856 3534 567884 62727
rect 569958 50280 570014 50289
rect 569958 50215 570014 50224
rect 569972 16574 570000 50215
rect 571984 44872 572036 44878
rect 571984 44814 572036 44820
rect 571340 36576 571392 36582
rect 571340 36518 571392 36524
rect 569972 16546 570368 16574
rect 567844 3528 567896 3534
rect 567844 3470 567896 3476
rect 569132 3528 569184 3534
rect 569132 3470 569184 3476
rect 569144 480 569172 3470
rect 570340 480 570368 16546
rect 567998 354 568110 480
rect 567580 326 568110 354
rect 567998 -960 568110 326
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571352 354 571380 36518
rect 571996 3058 572024 44814
rect 574100 18624 574152 18630
rect 574100 18566 574152 18572
rect 574112 16574 574140 18566
rect 574112 16546 574692 16574
rect 572720 3596 572772 3602
rect 572720 3538 572772 3544
rect 571984 3052 572036 3058
rect 571984 2994 572036 3000
rect 572732 480 572760 3538
rect 574664 3482 574692 16546
rect 574756 3602 574784 64874
rect 576136 6866 576164 140111
rect 580368 139369 580396 146270
rect 580540 140888 580592 140894
rect 580540 140830 580592 140836
rect 580448 140820 580500 140826
rect 580448 140762 580500 140768
rect 580354 139360 580410 139369
rect 580354 139295 580410 139304
rect 580264 138712 580316 138718
rect 580264 138654 580316 138660
rect 580172 86964 580224 86970
rect 580172 86906 580224 86912
rect 580184 86193 580212 86906
rect 580170 86184 580226 86193
rect 580170 86119 580226 86128
rect 579988 73160 580040 73166
rect 579988 73102 580040 73108
rect 580000 73001 580028 73102
rect 579986 72992 580042 73001
rect 579986 72927 580042 72936
rect 580276 59673 580304 138654
rect 580354 137320 580410 137329
rect 580354 137255 580410 137264
rect 580368 99521 580396 137255
rect 580460 112849 580488 140762
rect 580552 126041 580580 140830
rect 580538 126032 580594 126041
rect 580538 125967 580594 125976
rect 580446 112840 580502 112849
rect 580446 112775 580502 112784
rect 580354 99512 580410 99521
rect 580354 99447 580410 99456
rect 580262 59664 580318 59673
rect 580262 59599 580318 59608
rect 581092 54528 581144 54534
rect 581092 54470 581144 54476
rect 578240 51740 578292 51746
rect 578240 51682 578292 51688
rect 576860 35216 576912 35222
rect 576860 35158 576912 35164
rect 576872 16574 576900 35158
rect 578252 16574 578280 51682
rect 579988 20664 580040 20670
rect 579988 20606 580040 20612
rect 580000 19825 580028 20606
rect 579986 19816 580042 19825
rect 579986 19751 580042 19760
rect 581104 16574 581132 54470
rect 582380 32428 582432 32434
rect 582380 32370 582432 32376
rect 582392 16574 582420 32370
rect 576872 16546 576992 16574
rect 578252 16546 578648 16574
rect 581104 16546 581776 16574
rect 582392 16546 583432 16574
rect 576124 6860 576176 6866
rect 576124 6802 576176 6808
rect 574744 3596 574796 3602
rect 574744 3538 574796 3544
rect 576308 3596 576360 3602
rect 576308 3538 576360 3544
rect 574664 3454 575152 3482
rect 573916 3052 573968 3058
rect 573916 2994 573968 3000
rect 573928 480 573956 2994
rect 575124 480 575152 3454
rect 576320 480 576348 3538
rect 571494 354 571606 480
rect 571352 326 571606 354
rect 571494 -960 571606 326
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 576964 354 576992 16546
rect 578620 480 578648 16546
rect 580172 6860 580224 6866
rect 580172 6802 580224 6808
rect 580184 6633 580212 6802
rect 580170 6624 580226 6633
rect 580170 6559 580226 6568
rect 581000 3460 581052 3466
rect 581000 3402 581052 3408
rect 581012 480 581040 3402
rect 577382 354 577494 480
rect 576964 326 577494 354
rect 577382 -960 577494 326
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 581748 354 581776 16546
rect 583404 480 583432 16546
rect 582166 354 582278 480
rect 581748 326 582278 354
rect 582166 -960 582278 326
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 3330 671200 3386 671256
rect 3330 579944 3386 580000
rect 3238 566888 3294 566944
rect 3330 553832 3386 553888
rect 2778 527856 2834 527912
rect 3054 501744 3110 501800
rect 3054 475632 3110 475688
rect 3146 449520 3202 449576
rect 2870 410488 2926 410544
rect 3146 358400 3202 358456
rect 3330 345344 3386 345400
rect 3330 319232 3386 319288
rect 3054 267144 3110 267200
rect 3514 658164 3570 658200
rect 3514 658144 3516 658164
rect 3516 658144 3568 658164
rect 3568 658144 3570 658164
rect 3514 632068 3516 632088
rect 3516 632068 3568 632088
rect 3568 632068 3570 632088
rect 3514 632032 3570 632068
rect 3514 619112 3570 619168
rect 3514 606056 3570 606112
rect 3514 514820 3570 514856
rect 3514 514800 3516 514820
rect 3516 514800 3568 514820
rect 3568 514800 3570 514820
rect 3514 462576 3570 462632
rect 3514 423544 3570 423600
rect 3514 397468 3516 397488
rect 3516 397468 3568 397488
rect 3568 397468 3570 397488
rect 3514 397432 3570 397468
rect 3514 371340 3570 371376
rect 3514 371320 3516 371340
rect 3516 371320 3568 371340
rect 3568 371320 3570 371340
rect 3514 306176 3570 306232
rect 3514 293120 3570 293176
rect 2778 214920 2834 214976
rect 3514 254088 3570 254144
rect 3514 241068 3516 241088
rect 3516 241068 3568 241088
rect 3568 241068 3570 241088
rect 3514 241032 3570 241068
rect 3422 201864 3478 201920
rect 109958 200640 110014 200696
rect 107198 200232 107254 200288
rect 105634 200096 105690 200152
rect 103242 199824 103298 199880
rect 3422 188808 3478 188864
rect 3422 162832 3478 162888
rect 3422 149776 3478 149832
rect 3146 110608 3202 110664
rect 3514 136720 3570 136776
rect 4802 76472 4858 76528
rect 3514 71612 3516 71632
rect 3516 71612 3568 71632
rect 3568 71612 3570 71632
rect 3514 71576 3570 71612
rect 3514 58520 3570 58576
rect 3422 6432 3478 6488
rect 7562 75112 7618 75168
rect 31022 139440 31078 139496
rect 11058 72392 11114 72448
rect 8942 68176 8998 68232
rect 7654 65456 7710 65512
rect 17222 33768 17278 33824
rect 21362 73752 21418 73808
rect 24858 66816 24914 66872
rect 27710 51720 27766 51776
rect 39302 48864 39358 48920
rect 44178 47504 44234 47560
rect 46202 64096 46258 64152
rect 49698 46144 49754 46200
rect 54482 73888 54538 73944
rect 56598 54440 56654 54496
rect 75182 62736 75238 62792
rect 77298 57160 77354 57216
rect 80058 66952 80114 67008
rect 84198 59880 84254 59936
rect 93858 65728 93914 65784
rect 93122 65592 93178 65648
rect 92478 62872 92534 62928
rect 100206 74296 100262 74352
rect 97998 58520 98054 58576
rect 100206 73752 100262 73808
rect 100482 148280 100538 148336
rect 100758 52400 100814 52456
rect 101770 52400 101826 52456
rect 100758 51720 100814 51776
rect 100758 49544 100814 49600
rect 100758 48864 100814 48920
rect 102046 49544 102102 49600
rect 100758 48184 100814 48240
rect 101954 48184 102010 48240
rect 100758 47504 100814 47560
rect 102230 64776 102286 64832
rect 102230 64096 102286 64152
rect 102230 46824 102286 46880
rect 102690 46824 102746 46880
rect 102230 46144 102286 46200
rect 104806 195064 104862 195120
rect 104254 192752 104310 192808
rect 103334 64776 103390 64832
rect 103886 60560 103942 60616
rect 103886 59880 103942 59936
rect 104162 76200 104218 76256
rect 104438 186496 104494 186552
rect 104806 60560 104862 60616
rect 103978 55120 104034 55176
rect 103978 54440 104034 54496
rect 104898 54440 104954 54496
rect 106738 192480 106794 192536
rect 108762 198056 108818 198112
rect 107290 74160 107346 74216
rect 107474 185816 107530 185872
rect 107382 67496 107438 67552
rect 105818 57840 105874 57896
rect 106186 57840 106242 57896
rect 105818 57160 105874 57216
rect 108302 186768 108358 186824
rect 107566 59200 107622 59256
rect 107566 58520 107622 58576
rect 108854 66136 108910 66192
rect 110050 68312 110106 68368
rect 108118 63416 108174 63472
rect 110326 63280 110382 63336
rect 108118 62872 108174 62928
rect 110326 62736 110382 62792
rect 111338 68720 111394 68776
rect 111706 198600 111762 198656
rect 111706 71304 111762 71360
rect 111522 65592 111578 65648
rect 112258 76744 112314 76800
rect 112626 77152 112682 77208
rect 112902 190984 112958 191040
rect 112810 71168 112866 71224
rect 112994 75656 113050 75712
rect 113454 75248 113510 75304
rect 114374 199416 114430 199472
rect 113914 70216 113970 70272
rect 114374 77016 114430 77072
rect 112902 68448 112958 68504
rect 112350 66952 112406 67008
rect 113822 54984 113878 55040
rect 113822 54440 113878 54496
rect 115018 139168 115074 139224
rect 115110 138896 115166 138952
rect 114926 71712 114982 71768
rect 115570 193840 115626 193896
rect 116214 146920 116270 146976
rect 116582 76880 116638 76936
rect 116766 138760 116822 138816
rect 117870 140256 117926 140312
rect 117778 80144 117834 80200
rect 118238 259528 118294 259584
rect 116858 74024 116914 74080
rect 118606 198872 118662 198928
rect 118422 75520 118478 75576
rect 119158 142976 119214 143032
rect 119342 142704 119398 142760
rect 120354 198192 120410 198248
rect 119986 196696 120042 196752
rect 119250 138488 119306 138544
rect 120170 194792 120226 194848
rect 120722 199008 120778 199064
rect 120906 142840 120962 142896
rect 127898 262656 127954 262712
rect 126242 262248 126298 262304
rect 133326 262520 133382 262576
rect 133694 262520 133750 262576
rect 140134 264968 140190 265024
rect 138294 260888 138350 260944
rect 138018 260752 138074 260808
rect 138018 260344 138074 260400
rect 138938 260752 138994 260808
rect 141422 262384 141478 262440
rect 142250 260072 142306 260128
rect 143124 260072 143180 260128
rect 143814 260752 143870 260808
rect 144458 260752 144514 260808
rect 143722 260208 143778 260264
rect 144918 260208 144974 260264
rect 144550 259936 144606 259992
rect 145884 260208 145940 260264
rect 146942 263744 146998 263800
rect 125690 259664 125746 259720
rect 148322 262792 148378 262848
rect 151082 263608 151138 263664
rect 149242 260480 149298 260536
rect 150438 262792 150494 262848
rect 151910 270544 151966 270600
rect 151358 262792 151414 262848
rect 153014 262928 153070 262984
rect 154578 275984 154634 276040
rect 160098 260208 160154 260264
rect 160788 260208 160844 260264
rect 163410 264968 163466 265024
rect 162122 262384 162178 262440
rect 163686 262520 163742 262576
rect 163502 260208 163558 260264
rect 164238 259936 164294 259992
rect 166262 265104 166318 265160
rect 166078 263200 166134 263256
rect 166078 262656 166134 262712
rect 165066 259936 165122 259992
rect 167642 265240 167698 265296
rect 166354 263200 166410 263256
rect 167550 263064 167606 263120
rect 167734 263064 167790 263120
rect 171046 260208 171102 260264
rect 171046 259936 171102 259992
rect 180890 260208 180946 260264
rect 162122 259800 162178 259856
rect 160926 259664 160982 259720
rect 130842 259528 130898 259584
rect 180890 259664 180946 259720
rect 185398 259528 185454 259584
rect 186042 259528 186098 259584
rect 123482 199688 123538 199744
rect 120722 79464 120778 79520
rect 120998 75384 121054 75440
rect 119986 72936 120042 72992
rect 119894 72800 119950 72856
rect 115846 68584 115902 68640
rect 115938 68312 115994 68368
rect 121918 139340 121920 139360
rect 121920 139340 121972 139360
rect 121972 139340 121974 139360
rect 121918 139304 121974 139340
rect 122194 139168 122250 139224
rect 131670 199824 131726 199880
rect 131302 199552 131358 199608
rect 123482 140664 123538 140720
rect 123666 148416 123722 148472
rect 122746 139304 122802 139360
rect 122930 139304 122986 139360
rect 124218 141072 124274 141128
rect 125598 143384 125654 143440
rect 125690 142568 125746 142624
rect 125138 140936 125194 140992
rect 131026 198464 131082 198520
rect 126978 145832 127034 145888
rect 126978 142160 127034 142216
rect 128174 142160 128230 142216
rect 130658 141888 130714 141944
rect 130658 141616 130714 141672
rect 131854 145696 131910 145752
rect 132314 197784 132370 197840
rect 132130 185680 132186 185736
rect 132728 199858 132784 199914
rect 132912 199858 132968 199914
rect 132406 185544 132462 185600
rect 132774 197920 132830 197976
rect 132866 186088 132922 186144
rect 132774 185680 132830 185736
rect 132866 185272 132922 185328
rect 133464 199858 133520 199914
rect 133234 185136 133290 185192
rect 133924 199858 133980 199914
rect 134384 199824 134440 199880
rect 133510 197920 133566 197976
rect 133970 199280 134026 199336
rect 133878 198328 133934 198384
rect 133878 185680 133934 185736
rect 133694 185544 133750 185600
rect 134154 197648 134210 197704
rect 134338 198328 134394 198384
rect 134338 197920 134394 197976
rect 134246 197512 134302 197568
rect 134752 199858 134808 199914
rect 134522 197784 134578 197840
rect 134338 186088 134394 186144
rect 134246 185544 134302 185600
rect 135120 199858 135176 199914
rect 135304 199858 135360 199914
rect 135856 199858 135912 199914
rect 134798 197784 134854 197840
rect 134982 198328 135038 198384
rect 134982 185544 135038 185600
rect 136592 199858 136648 199914
rect 137144 199858 137200 199914
rect 137328 199858 137384 199914
rect 135258 199280 135314 199336
rect 135350 197784 135406 197840
rect 135442 192752 135498 192808
rect 135718 186224 135774 186280
rect 135074 185408 135130 185464
rect 136086 198328 136142 198384
rect 135994 197784 136050 197840
rect 135902 183096 135958 183152
rect 136454 199552 136510 199608
rect 136270 197920 136326 197976
rect 136546 199144 136602 199200
rect 136638 186632 136694 186688
rect 137006 186768 137062 186824
rect 137190 186496 137246 186552
rect 137098 185544 137154 185600
rect 132590 148280 132646 148336
rect 137880 199858 137936 199914
rect 138064 199858 138120 199914
rect 138432 199858 138488 199914
rect 138018 199552 138074 199608
rect 138018 192364 138074 192400
rect 138018 192344 138020 192364
rect 138020 192344 138072 192364
rect 138072 192344 138074 192364
rect 138478 190032 138534 190088
rect 138662 196832 138718 196888
rect 138662 195336 138718 195392
rect 139168 199858 139224 199914
rect 139352 199858 139408 199914
rect 138938 199144 138994 199200
rect 138938 198328 138994 198384
rect 138938 189760 138994 189816
rect 138386 177112 138442 177168
rect 139536 199858 139592 199914
rect 139720 199858 139776 199914
rect 139214 186224 139270 186280
rect 139122 185680 139178 185736
rect 140180 199858 140236 199914
rect 139858 198056 139914 198112
rect 139858 195744 139914 195800
rect 140456 199858 140512 199914
rect 140410 199280 140466 199336
rect 140318 198056 140374 198112
rect 140732 199858 140788 199914
rect 140502 189624 140558 189680
rect 139858 186224 139914 186280
rect 140134 186224 140190 186280
rect 139766 179288 139822 179344
rect 139030 174936 139086 174992
rect 137006 147600 137062 147656
rect 132866 143248 132922 143304
rect 141284 199858 141340 199914
rect 140594 185544 140650 185600
rect 141744 199858 141800 199914
rect 141606 192480 141662 192536
rect 141790 198056 141846 198112
rect 142296 199858 142352 199914
rect 142480 199858 142536 199914
rect 142664 199858 142720 199914
rect 141054 185408 141110 185464
rect 140962 185272 141018 185328
rect 141146 144472 141202 144528
rect 138938 143928 138994 143984
rect 139490 139984 139546 140040
rect 141422 141616 141478 141672
rect 141974 185544 142030 185600
rect 142342 198464 142398 198520
rect 142434 198056 142490 198112
rect 142618 199144 142674 199200
rect 143032 199858 143088 199914
rect 143078 199688 143134 199744
rect 142066 170992 142122 171048
rect 142066 161472 142122 161528
rect 142066 161336 142122 161392
rect 142066 151816 142122 151872
rect 142066 151680 142122 151736
rect 141514 141208 141570 141264
rect 142986 185544 143042 185600
rect 143354 192208 143410 192264
rect 143446 192072 143502 192128
rect 143538 191800 143594 191856
rect 143630 191120 143686 191176
rect 144504 199858 144560 199914
rect 144688 199858 144744 199914
rect 143814 190576 143870 190632
rect 144090 190440 144146 190496
rect 144734 190984 144790 191040
rect 144458 190712 144514 190768
rect 145700 199858 145756 199914
rect 145654 192888 145710 192944
rect 145746 190304 145802 190360
rect 146344 199858 146400 199914
rect 146114 198736 146170 198792
rect 145378 185952 145434 186008
rect 146712 199858 146768 199914
rect 146896 199858 146952 199914
rect 147080 199858 147136 199914
rect 146666 191392 146722 191448
rect 147126 189896 147182 189952
rect 147816 199858 147872 199914
rect 147310 181872 147366 181928
rect 147678 191256 147734 191312
rect 147494 186224 147550 186280
rect 146758 179288 146814 179344
rect 142802 144744 142858 144800
rect 142066 142296 142122 142352
rect 144458 144608 144514 144664
rect 143906 141752 143962 141808
rect 145562 144336 145618 144392
rect 145102 142976 145158 143032
rect 146666 143112 146722 143168
rect 148184 199858 148240 199914
rect 148046 190848 148102 190904
rect 148138 187176 148194 187232
rect 149012 199858 149068 199914
rect 149288 199858 149344 199914
rect 147218 144200 147274 144256
rect 147770 144064 147826 144120
rect 148966 199688 149022 199744
rect 148966 199416 149022 199472
rect 148874 186224 148930 186280
rect 149242 193704 149298 193760
rect 149610 197920 149666 197976
rect 149426 194248 149482 194304
rect 150300 199858 150356 199914
rect 149702 193840 149758 193896
rect 149334 191120 149390 191176
rect 149886 185544 149942 185600
rect 150944 199858 151000 199914
rect 151128 199858 151184 199914
rect 150898 186360 150954 186416
rect 148322 142704 148378 142760
rect 149058 141480 149114 141536
rect 149978 142840 150034 142896
rect 151174 199416 151230 199472
rect 151450 185544 151506 185600
rect 151726 199280 151782 199336
rect 152186 195608 152242 195664
rect 150530 141344 150586 141400
rect 150346 140120 150402 140176
rect 152370 198872 152426 198928
rect 152278 185544 152334 185600
rect 152554 185544 152610 185600
rect 153060 199858 153116 199914
rect 152738 186360 152794 186416
rect 152922 199008 152978 199064
rect 153106 196696 153162 196752
rect 153796 199858 153852 199914
rect 153290 186224 153346 186280
rect 152002 146920 152058 146976
rect 152278 142704 152334 142760
rect 153750 196560 153806 196616
rect 154440 199858 154496 199914
rect 154026 196696 154082 196752
rect 153842 186360 153898 186416
rect 153658 186224 153714 186280
rect 153382 149776 153438 149832
rect 153290 145560 153346 145616
rect 152830 141344 152886 141400
rect 153842 142840 153898 142896
rect 154302 197240 154358 197296
rect 154578 196832 154634 196888
rect 154992 199858 155048 199914
rect 155038 193976 155094 194032
rect 154210 185544 154266 185600
rect 153934 140120 153990 140176
rect 155636 199858 155692 199914
rect 155406 185544 155462 185600
rect 154854 149640 154910 149696
rect 155406 142976 155462 143032
rect 154762 140256 154818 140312
rect 156004 199858 156060 199914
rect 156464 199858 156520 199914
rect 155958 199688 156014 199744
rect 156050 186224 156106 186280
rect 124126 139304 124182 139360
rect 126886 139304 126942 139360
rect 129646 139304 129702 139360
rect 131670 139304 131726 139360
rect 132222 139304 132278 139360
rect 138294 139304 138350 139360
rect 151082 139304 151138 139360
rect 152370 139304 152426 139360
rect 155130 139340 155132 139360
rect 155132 139340 155184 139360
rect 155184 139340 155186 139360
rect 155130 139304 155186 139340
rect 156418 192888 156474 192944
rect 156694 199688 156750 199744
rect 157200 199858 157256 199914
rect 157154 199708 157210 199744
rect 157154 199688 157156 199708
rect 157156 199688 157208 199708
rect 157208 199688 157210 199708
rect 158028 199858 158084 199914
rect 157522 193024 157578 193080
rect 156970 185544 157026 185600
rect 156142 152496 156198 152552
rect 156050 150320 156106 150376
rect 156234 150184 156290 150240
rect 157246 147056 157302 147112
rect 158304 199858 158360 199914
rect 158580 199858 158636 199914
rect 158258 186224 158314 186280
rect 158166 185816 158222 185872
rect 157522 152632 157578 152688
rect 159086 192616 159142 192672
rect 158718 185544 158774 185600
rect 159178 179424 159234 179480
rect 159684 199858 159740 199914
rect 160144 199858 160200 199914
rect 158810 145696 158866 145752
rect 157706 144064 157762 144120
rect 157246 143112 157302 143168
rect 157338 142024 157394 142080
rect 160374 199552 160430 199608
rect 160190 186088 160246 186144
rect 160466 186224 160522 186280
rect 160880 199858 160936 199914
rect 161340 199858 161396 199914
rect 160558 178472 160614 178528
rect 161616 199858 161672 199914
rect 161570 199688 161626 199744
rect 161018 185544 161074 185600
rect 160834 181736 160890 181792
rect 160742 177928 160798 177984
rect 161294 171128 161350 171184
rect 161294 170992 161350 171048
rect 161294 161472 161350 161528
rect 161294 161336 161350 161392
rect 161294 151816 161350 151872
rect 161294 151680 161350 151736
rect 160926 145560 160982 145616
rect 162076 199858 162132 199914
rect 162628 199858 162684 199914
rect 161662 193296 161718 193352
rect 162122 199688 162178 199744
rect 162996 199824 163052 199880
rect 163272 199858 163328 199914
rect 163456 199824 163512 199880
rect 163732 199858 163788 199914
rect 162398 199552 162454 199608
rect 162766 198328 162822 198384
rect 162674 186360 162730 186416
rect 162490 186224 162546 186280
rect 162950 198192 163006 198248
rect 162950 198056 163006 198112
rect 162858 192480 162914 192536
rect 162766 179016 162822 179072
rect 163318 198056 163374 198112
rect 163226 186904 163282 186960
rect 163226 186768 163282 186824
rect 163318 186360 163374 186416
rect 163778 199688 163834 199744
rect 164744 199858 164800 199914
rect 165204 199858 165260 199914
rect 163502 186088 163558 186144
rect 164698 199688 164754 199744
rect 164054 186224 164110 186280
rect 163134 148280 163190 148336
rect 162950 145832 163006 145888
rect 162214 143248 162270 143304
rect 161294 142296 161350 142352
rect 162766 144200 162822 144256
rect 163870 143384 163926 143440
rect 164422 183368 164478 183424
rect 164606 198056 164662 198112
rect 164606 186360 164662 186416
rect 164882 186224 164938 186280
rect 165250 192752 165306 192808
rect 165434 199008 165490 199064
rect 165802 190440 165858 190496
rect 166262 199688 166318 199744
rect 165986 185680 166042 185736
rect 165710 185408 165766 185464
rect 165710 185272 165766 185328
rect 165526 178472 165582 178528
rect 166952 199824 167008 199880
rect 166814 199708 166870 199744
rect 166814 199688 166816 199708
rect 166816 199688 166868 199708
rect 166868 199688 166870 199708
rect 166354 180240 166410 180296
rect 166998 198056 167054 198112
rect 166906 185680 166962 185736
rect 166630 185544 166686 185600
rect 167550 199688 167606 199744
rect 167872 199824 167928 199880
rect 168056 199858 168112 199914
rect 168240 199858 168296 199914
rect 168608 199858 168664 199914
rect 168884 199858 168940 199914
rect 169528 199858 169584 199914
rect 168102 199688 168158 199744
rect 167642 198192 167698 198248
rect 167550 185544 167606 185600
rect 167734 197784 167790 197840
rect 167918 198056 167974 198112
rect 167734 185680 167790 185736
rect 168102 198056 168158 198112
rect 168010 185544 168066 185600
rect 168746 199688 168802 199744
rect 169712 199858 169768 199914
rect 169206 185816 169262 185872
rect 169114 179968 169170 180024
rect 165710 148416 165766 148472
rect 169390 193840 169446 193896
rect 169298 185680 169354 185736
rect 169758 199688 169814 199744
rect 170540 199858 170596 199914
rect 170034 199708 170090 199744
rect 170034 199688 170036 199708
rect 170036 199688 170088 199708
rect 170088 199688 170090 199708
rect 171000 199858 171056 199914
rect 171184 199858 171240 199914
rect 171552 199824 171608 199880
rect 169942 196424 169998 196480
rect 169942 195880 169998 195936
rect 169850 186496 169906 186552
rect 169574 185544 169630 185600
rect 164238 145968 164294 146024
rect 164146 144472 164202 144528
rect 167734 144608 167790 144664
rect 166630 144336 166686 144392
rect 166078 141480 166134 141536
rect 169850 147464 169906 147520
rect 170218 198192 170274 198248
rect 170494 199688 170550 199744
rect 170678 199688 170734 199744
rect 170494 198736 170550 198792
rect 170586 186224 170642 186280
rect 170862 199688 170918 199744
rect 170770 198056 170826 198112
rect 171138 199688 171194 199744
rect 171506 199688 171562 199744
rect 170678 184864 170734 184920
rect 171138 147328 171194 147384
rect 171874 185544 171930 185600
rect 172058 185544 172114 185600
rect 172242 185680 172298 185736
rect 172150 185136 172206 185192
rect 173208 199824 173264 199880
rect 173392 199824 173448 199880
rect 172886 186088 172942 186144
rect 173254 199688 173310 199744
rect 173162 185544 173218 185600
rect 173438 198736 173494 198792
rect 173346 185544 173402 185600
rect 173070 185272 173126 185328
rect 173714 185952 173770 186008
rect 174312 199858 174368 199914
rect 174864 199824 174920 199880
rect 174542 186224 174598 186280
rect 175416 199858 175472 199914
rect 175186 199724 175188 199744
rect 175188 199724 175240 199744
rect 175240 199724 175242 199744
rect 175186 199688 175242 199724
rect 175462 199688 175518 199744
rect 175968 199824 176024 199880
rect 176336 199824 176392 199880
rect 176520 199858 176576 199914
rect 174818 198736 174874 198792
rect 176888 199858 176944 199914
rect 174174 150048 174230 150104
rect 174358 149912 174414 149968
rect 175646 185816 175702 185872
rect 175738 185680 175794 185736
rect 176014 185408 176070 185464
rect 176290 186224 176346 186280
rect 176750 197920 176806 197976
rect 176750 197512 176806 197568
rect 176658 186496 176714 186552
rect 173990 147192 174046 147248
rect 173898 146104 173954 146160
rect 174818 140256 174874 140312
rect 177854 186224 177910 186280
rect 177302 176568 177358 176624
rect 176750 141616 176806 141672
rect 176658 141208 176714 141264
rect 178590 140664 178646 140720
rect 180430 198872 180486 198928
rect 180338 147600 180394 147656
rect 174818 139440 174874 139496
rect 180430 139712 180486 139768
rect 179878 139596 179934 139632
rect 179878 139576 179880 139596
rect 179880 139576 179932 139596
rect 179932 139576 179934 139596
rect 180798 140256 180854 140312
rect 182454 144880 182510 144936
rect 181442 140256 181498 140312
rect 182086 140120 182142 140176
rect 182178 139848 182234 139904
rect 183466 144880 183522 144936
rect 183190 139984 183246 140040
rect 184478 141072 184534 141128
rect 184294 140800 184350 140856
rect 184754 139984 184810 140040
rect 184938 140528 184994 140584
rect 185030 140392 185086 140448
rect 185030 140256 185086 140312
rect 185582 143520 185638 143576
rect 185306 139848 185362 139904
rect 186594 262928 186650 262984
rect 186870 259936 186926 259992
rect 187238 202816 187294 202872
rect 186962 149096 187018 149152
rect 186870 143384 186926 143440
rect 186502 142840 186558 142896
rect 186962 142704 187018 142760
rect 186410 141344 186466 141400
rect 186318 140800 186374 140856
rect 185950 140392 186006 140448
rect 155682 139304 155738 139360
rect 159546 139304 159602 139360
rect 160006 139304 160062 139360
rect 163962 139304 164018 139360
rect 179694 139304 179750 139360
rect 180522 139304 180578 139360
rect 122378 138488 122434 138544
rect 186410 139168 186466 139224
rect 187238 174528 187294 174584
rect 187974 262248 188030 262304
rect 187974 260072 188030 260128
rect 187698 143112 187754 143168
rect 187790 142976 187846 143032
rect 188158 259800 188214 259856
rect 188434 259664 188490 259720
rect 188342 201728 188398 201784
rect 188158 143248 188214 143304
rect 187054 138080 187110 138136
rect 122746 137944 122802 138000
rect 122746 128424 122802 128480
rect 122746 122848 122802 122904
rect 122746 122712 122802 122768
rect 122746 113192 122802 113248
rect 122746 113056 122802 113112
rect 122746 103536 122802 103592
rect 122746 103400 122802 103456
rect 122746 93880 122802 93936
rect 122746 93744 122802 93800
rect 122746 89664 122802 89720
rect 122470 81368 122526 81424
rect 186502 80960 186558 81016
rect 187146 80960 187202 81016
rect 187422 80960 187478 81016
rect 122838 80280 122894 80336
rect 177762 80688 177818 80744
rect 178406 80688 178462 80744
rect 132038 80552 132094 80608
rect 131946 80416 132002 80472
rect 131762 80280 131818 80336
rect 124126 79600 124182 79656
rect 125598 76608 125654 76664
rect 129738 75248 129794 75304
rect 130658 79736 130714 79792
rect 130382 78512 130438 78568
rect 130382 75928 130438 75984
rect 130934 79736 130990 79792
rect 130934 75248 130990 75304
rect 131026 72528 131082 72584
rect 131578 75928 131634 75984
rect 177854 80552 177910 80608
rect 131946 78512 132002 78568
rect 132314 79872 132370 79928
rect 132544 79906 132600 79962
rect 133096 79906 133152 79962
rect 133096 79770 133152 79826
rect 133924 79872 133980 79928
rect 132038 77832 132094 77888
rect 132590 76200 132646 76256
rect 133556 79736 133612 79792
rect 133234 77832 133290 77888
rect 133234 72392 133290 72448
rect 133418 77832 133474 77888
rect 134476 79872 134532 79928
rect 134338 79756 134394 79792
rect 134338 79736 134340 79756
rect 134340 79736 134392 79756
rect 134392 79736 134394 79756
rect 133970 77560 134026 77616
rect 133786 74296 133842 74352
rect 133878 66952 133934 67008
rect 134844 79838 134900 79894
rect 134614 79600 134670 79656
rect 134798 79600 134854 79656
rect 134798 78512 134854 78568
rect 135074 73888 135130 73944
rect 135764 79872 135820 79928
rect 135626 79620 135682 79656
rect 135626 79600 135628 79620
rect 135628 79600 135680 79620
rect 135680 79600 135682 79620
rect 135718 77832 135774 77888
rect 135902 79756 135958 79792
rect 135902 79736 135904 79756
rect 135904 79736 135956 79756
rect 135956 79736 135958 79756
rect 136500 79906 136556 79962
rect 135994 77560 136050 77616
rect 135810 76472 135866 76528
rect 136178 78512 136234 78568
rect 136960 79872 137016 79928
rect 136638 79600 136694 79656
rect 137328 79770 137384 79826
rect 136822 79600 136878 79656
rect 136270 74160 136326 74216
rect 136454 73752 136510 73808
rect 136730 78512 136786 78568
rect 136730 77832 136786 77888
rect 136914 78512 136970 78568
rect 137098 79600 137154 79656
rect 137282 79620 137338 79656
rect 137282 79600 137284 79620
rect 137284 79600 137336 79620
rect 137336 79600 137338 79620
rect 137190 78512 137246 78568
rect 137558 78512 137614 78568
rect 137880 79872 137936 79928
rect 138248 79906 138304 79962
rect 138432 79892 138488 79928
rect 138432 79872 138434 79892
rect 138434 79872 138486 79892
rect 138486 79872 138488 79892
rect 137926 79736 137982 79792
rect 138064 79736 138120 79792
rect 137558 77560 137614 77616
rect 137558 77424 137614 77480
rect 137834 78240 137890 78296
rect 138018 78512 138074 78568
rect 138110 78376 138166 78432
rect 138110 77832 138166 77888
rect 138984 79872 139040 79928
rect 138846 79736 138902 79792
rect 138294 77288 138350 77344
rect 138570 78240 138626 78296
rect 138754 78276 138756 78296
rect 138756 78276 138808 78296
rect 138808 78276 138810 78296
rect 138754 78240 138810 78276
rect 139076 79736 139132 79792
rect 139306 79736 139362 79792
rect 139536 79872 139592 79928
rect 139720 79872 139776 79928
rect 138938 77424 138994 77480
rect 139214 78920 139270 78976
rect 139812 79772 139814 79792
rect 139814 79772 139866 79792
rect 139866 79772 139868 79792
rect 139812 79736 139868 79772
rect 139398 77832 139454 77888
rect 140088 79872 140144 79928
rect 139582 78920 139638 78976
rect 140364 79872 140420 79928
rect 140410 79736 140466 79792
rect 140640 79872 140696 79928
rect 140042 77832 140098 77888
rect 140042 77424 140098 77480
rect 140686 79736 140742 79792
rect 141192 79892 141248 79928
rect 141192 79872 141194 79892
rect 141194 79872 141246 79892
rect 141246 79872 141248 79892
rect 140502 77696 140558 77752
rect 140870 76744 140926 76800
rect 141744 79872 141800 79928
rect 141146 78920 141202 78976
rect 141238 78512 141294 78568
rect 141330 77832 141386 77888
rect 141698 78376 141754 78432
rect 141514 75384 141570 75440
rect 142572 79906 142628 79962
rect 142848 79906 142904 79962
rect 143032 79906 143088 79962
rect 142710 79736 142766 79792
rect 142894 79736 142950 79792
rect 143078 79736 143134 79792
rect 142434 78920 142490 78976
rect 142526 78376 142582 78432
rect 142342 77696 142398 77752
rect 141882 76608 141938 76664
rect 143400 79906 143456 79962
rect 143952 79872 144008 79928
rect 143538 78648 143594 78704
rect 143446 78104 143502 78160
rect 143354 68448 143410 68504
rect 143814 78512 143870 78568
rect 143906 74296 143962 74352
rect 144090 78920 144146 78976
rect 144826 79736 144882 79792
rect 144366 78648 144422 78704
rect 145884 79906 145940 79962
rect 145838 79736 145894 79792
rect 145286 79192 145342 79248
rect 144826 70488 144882 70544
rect 145378 77560 145434 77616
rect 145746 78240 145802 78296
rect 144550 68720 144606 68776
rect 146114 77696 146170 77752
rect 146298 76880 146354 76936
rect 146712 79908 146714 79928
rect 146714 79908 146766 79928
rect 146766 79908 146768 79928
rect 146712 79872 146768 79908
rect 146896 79736 146952 79792
rect 147632 79906 147688 79962
rect 146942 79500 146944 79520
rect 146944 79500 146996 79520
rect 146996 79500 146998 79520
rect 146942 79464 146998 79500
rect 147126 79464 147182 79520
rect 146942 76880 146998 76936
rect 147448 79736 147504 79792
rect 147402 79500 147404 79520
rect 147404 79500 147456 79520
rect 147456 79500 147458 79520
rect 147402 79464 147458 79500
rect 148000 79736 148056 79792
rect 148552 79908 148554 79928
rect 148554 79908 148606 79928
rect 148606 79908 148608 79928
rect 148552 79872 148608 79908
rect 147678 79464 147734 79520
rect 147310 77832 147366 77888
rect 148138 79500 148140 79520
rect 148140 79500 148192 79520
rect 148192 79500 148194 79520
rect 148138 79464 148194 79500
rect 148506 79736 148562 79792
rect 148736 79872 148792 79928
rect 148690 78240 148746 78296
rect 148598 77988 148654 78024
rect 148598 77968 148600 77988
rect 148600 77968 148652 77988
rect 148652 77968 148654 77988
rect 148690 77832 148746 77888
rect 149288 79906 149344 79962
rect 148966 77424 149022 77480
rect 149334 79736 149390 79792
rect 149242 78784 149298 78840
rect 150024 79906 150080 79962
rect 150300 79872 150356 79928
rect 149610 78240 149666 78296
rect 149886 77696 149942 77752
rect 150852 79906 150908 79962
rect 150162 79056 150218 79112
rect 150346 78920 150402 78976
rect 150438 77832 150494 77888
rect 151128 79906 151184 79962
rect 151404 79906 151460 79962
rect 150714 79328 150770 79384
rect 150806 79056 150862 79112
rect 151680 79872 151736 79928
rect 151542 79736 151598 79792
rect 151358 79056 151414 79112
rect 151266 78648 151322 78704
rect 152232 79892 152288 79928
rect 152232 79872 152234 79892
rect 152234 79872 152286 79892
rect 152286 79872 152288 79892
rect 151726 78512 151782 78568
rect 152048 79736 152104 79792
rect 152094 79600 152150 79656
rect 152784 79908 152786 79928
rect 152786 79908 152838 79928
rect 152838 79908 152840 79928
rect 152784 79872 152840 79908
rect 152968 79872 153024 79928
rect 152830 79328 152886 79384
rect 152646 73752 152702 73808
rect 153014 79636 153016 79656
rect 153016 79636 153068 79656
rect 153068 79636 153070 79656
rect 153014 79600 153070 79636
rect 152922 73480 152978 73536
rect 153612 79872 153668 79928
rect 153888 79872 153944 79928
rect 154348 79906 154404 79962
rect 154992 79872 155048 79928
rect 153290 77424 153346 77480
rect 153658 79464 153714 79520
rect 153566 71576 153622 71632
rect 154118 79736 154174 79792
rect 155360 79906 155416 79962
rect 155636 79906 155692 79962
rect 153842 79364 153844 79384
rect 153844 79364 153896 79384
rect 153896 79364 153898 79384
rect 153842 79328 153898 79364
rect 154026 74568 154082 74624
rect 153934 74432 153990 74488
rect 154026 73072 154082 73128
rect 154302 79600 154358 79656
rect 154394 79464 154450 79520
rect 154578 79464 154634 79520
rect 154486 77288 154542 77344
rect 154762 68856 154818 68912
rect 155130 79464 155186 79520
rect 155406 79620 155462 79656
rect 155406 79600 155408 79620
rect 155408 79600 155460 79620
rect 155460 79600 155462 79620
rect 155406 79364 155408 79384
rect 155408 79364 155460 79384
rect 155460 79364 155462 79384
rect 155130 78104 155186 78160
rect 155406 79328 155462 79364
rect 155912 79872 155968 79928
rect 155774 79600 155830 79656
rect 155682 79328 155738 79384
rect 155590 77152 155646 77208
rect 155038 63280 155094 63336
rect 154946 61920 155002 61976
rect 155774 78920 155830 78976
rect 155866 77016 155922 77072
rect 156142 78648 156198 78704
rect 156142 77560 156198 77616
rect 156050 74296 156106 74352
rect 156648 79872 156704 79928
rect 156234 73072 156290 73128
rect 157016 79872 157072 79928
rect 157476 79872 157532 79928
rect 156602 79600 156658 79656
rect 157338 79736 157394 79792
rect 157752 79772 157754 79792
rect 157754 79772 157806 79792
rect 157806 79772 157808 79792
rect 157752 79736 157808 79772
rect 156510 72936 156566 72992
rect 156970 79600 157026 79656
rect 156786 77560 156842 77616
rect 156510 72256 156566 72312
rect 155958 26832 156014 26888
rect 156786 74296 156842 74352
rect 157062 79328 157118 79384
rect 157246 78512 157302 78568
rect 156970 73072 157026 73128
rect 156878 72800 156934 72856
rect 156970 72664 157026 72720
rect 157062 72528 157118 72584
rect 157062 72392 157118 72448
rect 156970 72256 157026 72312
rect 157614 79600 157670 79656
rect 157522 78920 157578 78976
rect 157706 78512 157762 78568
rect 158074 75928 158130 75984
rect 157982 75792 158038 75848
rect 158580 79872 158636 79928
rect 158396 79772 158398 79792
rect 158398 79772 158450 79792
rect 158450 79772 158452 79792
rect 158396 79736 158452 79772
rect 158856 79872 158912 79928
rect 158626 79600 158682 79656
rect 158258 79328 158314 79384
rect 158810 79736 158866 79792
rect 158718 78784 158774 78840
rect 159132 79872 159188 79928
rect 159178 79772 159180 79792
rect 159180 79772 159232 79792
rect 159232 79772 159234 79792
rect 159178 79736 159234 79772
rect 159684 79906 159740 79962
rect 159868 79906 159924 79962
rect 159914 79736 159970 79792
rect 160328 79872 160384 79928
rect 159822 79600 159878 79656
rect 160144 79736 160200 79792
rect 160604 79824 160660 79826
rect 159730 71848 159786 71904
rect 160098 79600 160154 79656
rect 160006 74976 160062 75032
rect 158902 11600 158958 11656
rect 160604 79772 160606 79824
rect 160606 79772 160658 79824
rect 160658 79772 160660 79824
rect 161340 79906 161396 79962
rect 160604 79770 160660 79772
rect 160466 79464 160522 79520
rect 160374 79056 160430 79112
rect 160742 79464 160798 79520
rect 160926 67632 160982 67688
rect 161616 79872 161672 79928
rect 161984 79906 162040 79962
rect 161202 79600 161258 79656
rect 161110 78512 161166 78568
rect 161202 74160 161258 74216
rect 161018 67496 161074 67552
rect 160374 33768 160430 33824
rect 161294 15816 161350 15872
rect 162352 79736 162408 79792
rect 162720 79908 162722 79928
rect 162722 79908 162774 79928
rect 162774 79908 162776 79928
rect 162720 79872 162776 79908
rect 162904 79906 162960 79962
rect 163272 79872 163328 79928
rect 161846 79620 161902 79656
rect 161846 79600 161848 79620
rect 161848 79600 161900 79620
rect 161900 79600 161902 79620
rect 161938 79464 161994 79520
rect 162214 79600 162270 79656
rect 162122 79328 162178 79384
rect 162582 79620 162638 79656
rect 162582 79600 162584 79620
rect 162584 79600 162636 79620
rect 162636 79600 162638 79620
rect 162398 79464 162454 79520
rect 162674 79464 162730 79520
rect 162490 71712 162546 71768
rect 162766 78512 162822 78568
rect 162950 79600 163006 79656
rect 163640 79872 163696 79928
rect 163594 79464 163650 79520
rect 164100 79908 164102 79928
rect 164102 79908 164154 79928
rect 164154 79908 164156 79928
rect 164100 79872 164156 79908
rect 163778 79636 163780 79656
rect 163780 79636 163832 79656
rect 163832 79636 163834 79656
rect 163778 79600 163834 79636
rect 163870 78648 163926 78704
rect 163870 78104 163926 78160
rect 163594 61648 163650 61704
rect 164376 79872 164432 79928
rect 164928 79872 164984 79928
rect 165480 79872 165536 79928
rect 164238 79192 164294 79248
rect 164146 77560 164202 77616
rect 164790 77424 164846 77480
rect 165066 79620 165122 79656
rect 165066 79600 165068 79620
rect 165068 79600 165120 79620
rect 165120 79600 165122 79620
rect 165158 79192 165214 79248
rect 165434 79736 165490 79792
rect 165756 79906 165812 79962
rect 165940 79906 165996 79962
rect 165250 77696 165306 77752
rect 165250 77560 165306 77616
rect 165526 79192 165582 79248
rect 165618 79056 165674 79112
rect 165618 78648 165674 78704
rect 165526 78376 165582 78432
rect 166032 79772 166034 79792
rect 166034 79772 166086 79792
rect 166086 79772 166088 79792
rect 166032 79736 166088 79772
rect 166860 79872 166916 79928
rect 166584 79736 166640 79792
rect 167412 79872 167468 79928
rect 165802 79192 165858 79248
rect 165986 67496 166042 67552
rect 165894 67088 165950 67144
rect 166814 79636 166816 79656
rect 166816 79636 166868 79656
rect 166868 79636 166870 79656
rect 166814 79600 166870 79636
rect 166998 79600 167054 79656
rect 166630 73616 166686 73672
rect 166446 70216 166502 70272
rect 166630 70080 166686 70136
rect 166906 70216 166962 70272
rect 168240 79906 168296 79962
rect 167274 79192 167330 79248
rect 167458 73752 167514 73808
rect 167918 79600 167974 79656
rect 168102 79772 168104 79792
rect 168104 79772 168156 79792
rect 168156 79772 168158 79792
rect 168102 79736 168158 79772
rect 168424 79872 168480 79928
rect 168608 79906 168664 79962
rect 169068 79908 169070 79928
rect 169070 79908 169122 79928
rect 169122 79908 169124 79928
rect 169068 79872 169124 79908
rect 167734 78104 167790 78160
rect 167550 73344 167606 73400
rect 168194 79192 168250 79248
rect 168378 79056 168434 79112
rect 169712 79906 169768 79962
rect 169298 79600 169354 79656
rect 168562 61376 168618 61432
rect 169482 79620 169538 79656
rect 169482 79600 169484 79620
rect 169484 79600 169536 79620
rect 169536 79600 169538 79620
rect 169390 75928 169446 75984
rect 170080 79736 170136 79792
rect 170448 79872 170504 79928
rect 169666 79192 169722 79248
rect 169850 78784 169906 78840
rect 170724 79872 170780 79928
rect 171000 79960 171056 79962
rect 171000 79908 171002 79960
rect 171002 79908 171054 79960
rect 171054 79908 171056 79960
rect 171000 79906 171056 79908
rect 170218 79600 170274 79656
rect 169942 78240 169998 78296
rect 170494 77288 170550 77344
rect 170586 76880 170642 76936
rect 171368 79906 171424 79962
rect 171552 79872 171608 79928
rect 172012 79906 172068 79962
rect 170954 79600 171010 79656
rect 170862 77424 170918 77480
rect 170770 77288 170826 77344
rect 170310 75384 170366 75440
rect 170770 76472 170826 76528
rect 170402 37848 170458 37904
rect 171230 78784 171286 78840
rect 171138 78104 171194 78160
rect 171414 78920 171470 78976
rect 171782 79756 171838 79792
rect 171782 79736 171784 79756
rect 171784 79736 171836 79756
rect 171836 79736 171838 79756
rect 172058 79756 172114 79792
rect 172058 79736 172060 79756
rect 172060 79736 172112 79756
rect 172112 79736 172114 79756
rect 172288 79906 172344 79962
rect 171690 78512 171746 78568
rect 171598 77832 171654 77888
rect 171506 76744 171562 76800
rect 171966 79328 172022 79384
rect 171966 79192 172022 79248
rect 171874 77696 171930 77752
rect 171782 68856 171838 68912
rect 171874 17176 171930 17232
rect 172150 76064 172206 76120
rect 172748 79872 172804 79928
rect 172334 79328 172390 79384
rect 172242 75928 172298 75984
rect 172426 71324 172482 71360
rect 172426 71304 172428 71324
rect 172428 71304 172480 71324
rect 172480 71304 172482 71324
rect 172794 78920 172850 78976
rect 172610 75928 172666 75984
rect 172978 79328 173034 79384
rect 173208 79736 173264 79792
rect 172978 75248 173034 75304
rect 173254 79192 173310 79248
rect 173438 78920 173494 78976
rect 173162 73752 173218 73808
rect 173944 79908 173946 79928
rect 173946 79908 173998 79928
rect 173998 79908 174000 79928
rect 173944 79872 174000 79908
rect 174128 79872 174184 79928
rect 173622 78784 173678 78840
rect 173714 76336 173770 76392
rect 174082 79736 174138 79792
rect 174588 79872 174644 79928
rect 173806 76064 173862 76120
rect 174358 79736 174414 79792
rect 174496 79772 174498 79792
rect 174498 79772 174550 79792
rect 174550 79772 174552 79792
rect 174496 79736 174552 79772
rect 174266 78920 174322 78976
rect 174450 79328 174506 79384
rect 174450 75792 174506 75848
rect 174864 79872 174920 79928
rect 174910 79736 174966 79792
rect 175232 79872 175288 79928
rect 175416 79872 175472 79928
rect 174818 78784 174874 78840
rect 174726 74160 174782 74216
rect 174910 77560 174966 77616
rect 174910 75112 174966 75168
rect 175278 78784 175334 78840
rect 175278 78648 175334 78704
rect 175094 77560 175150 77616
rect 175186 75520 175242 75576
rect 175094 74160 175150 74216
rect 175968 79872 176024 79928
rect 175922 79756 175978 79792
rect 175922 79736 175924 79756
rect 175924 79736 175976 79756
rect 175976 79736 175978 79756
rect 176152 79736 176208 79792
rect 176520 79872 176576 79928
rect 176290 79772 176292 79792
rect 176292 79772 176344 79792
rect 176344 79772 176346 79792
rect 176290 79736 176346 79772
rect 176106 79600 176162 79656
rect 175738 79328 175794 79384
rect 175646 79192 175702 79248
rect 175922 79192 175978 79248
rect 175738 78784 175794 78840
rect 175462 71712 175518 71768
rect 176106 70080 176162 70136
rect 176704 79906 176760 79962
rect 176382 78648 176438 78704
rect 176658 79328 176714 79384
rect 176566 77832 176622 77888
rect 176566 75656 176622 75712
rect 177348 79906 177404 79962
rect 177578 79872 177634 79928
rect 177486 79736 177542 79792
rect 177302 79600 177358 79656
rect 177854 79872 177910 79928
rect 177670 77560 177726 77616
rect 178222 79736 178278 79792
rect 183742 80280 183798 80336
rect 180890 79872 180946 79928
rect 180062 79600 180118 79656
rect 178682 79192 178738 79248
rect 177946 78784 178002 78840
rect 177854 78104 177910 78160
rect 177762 77288 177818 77344
rect 177578 76608 177634 76664
rect 177946 77288 178002 77344
rect 178406 72392 178462 72448
rect 180890 79328 180946 79384
rect 178958 77424 179014 77480
rect 180062 76608 180118 76664
rect 179326 76336 179382 76392
rect 179234 75384 179290 75440
rect 179694 73072 179750 73128
rect 180430 77696 180486 77752
rect 180246 73480 180302 73536
rect 180430 77288 180486 77344
rect 181258 73072 181314 73128
rect 181166 66136 181222 66192
rect 187422 78648 187478 78704
rect 184478 78512 184534 78568
rect 186410 78512 186466 78568
rect 187422 78512 187478 78568
rect 183282 77016 183338 77072
rect 183282 76608 183338 76664
rect 183834 68992 183890 69048
rect 183742 61512 183798 61568
rect 188250 68720 188306 68776
rect 188066 66156 188122 66192
rect 188066 66136 188068 66156
rect 188068 66136 188120 66156
rect 188120 66136 188122 66156
rect 188618 65048 188674 65104
rect 189354 260208 189410 260264
rect 189262 139304 189318 139360
rect 189078 63280 189134 63336
rect 189446 139032 189502 139088
rect 189630 74432 189686 74488
rect 189630 73752 189686 73808
rect 189722 68176 189778 68232
rect 189446 60560 189502 60616
rect 189630 60560 189686 60616
rect 189630 60152 189686 60208
rect 189262 56208 189318 56264
rect 191194 180784 191250 180840
rect 190918 138760 190974 138816
rect 191102 138488 191158 138544
rect 191286 146104 191342 146160
rect 191470 145696 191526 145752
rect 191286 140800 191342 140856
rect 191194 114416 191250 114472
rect 191194 81912 191250 81968
rect 191562 144744 191618 144800
rect 191378 61784 191434 61840
rect 190918 60424 190974 60480
rect 190550 57840 190606 57896
rect 191746 60424 191802 60480
rect 191746 60016 191802 60072
rect 191746 57840 191802 57896
rect 191746 57432 191802 57488
rect 192022 63416 192078 63472
rect 192114 59064 192170 59120
rect 191838 54984 191894 55040
rect 191838 54712 191894 54768
rect 191562 52128 191618 52184
rect 193218 145560 193274 145616
rect 193218 140528 193274 140584
rect 193126 63416 193182 63472
rect 193126 63144 193182 63200
rect 193126 59064 193182 59120
rect 193126 58792 193182 58848
rect 192850 53352 192906 53408
rect 193678 140700 193680 140720
rect 193680 140700 193732 140720
rect 193732 140700 193734 140720
rect 193678 140664 193734 140700
rect 193678 138896 193734 138952
rect 193586 78532 193642 78568
rect 193586 78512 193588 78532
rect 193588 78512 193640 78532
rect 193640 78512 193642 78532
rect 194046 139304 194102 139360
rect 193862 66816 193918 66872
rect 193678 61512 193734 61568
rect 193402 59880 193458 59936
rect 193310 50904 193366 50960
rect 192206 50496 192262 50552
rect 194690 59200 194746 59256
rect 195150 145968 195206 146024
rect 195334 81232 195390 81288
rect 195242 78376 195298 78432
rect 195610 139440 195666 139496
rect 195150 70352 195206 70408
rect 195058 59200 195114 59256
rect 195058 58656 195114 58712
rect 194782 57704 194838 57760
rect 195058 57704 195114 57760
rect 195058 57296 195114 57352
rect 194598 55120 194654 55176
rect 194598 54576 194654 54632
rect 196806 147736 196862 147792
rect 196530 138624 196586 138680
rect 196990 81096 197046 81152
rect 196162 66000 196218 66056
rect 196438 66000 196494 66056
rect 196438 65456 196494 65512
rect 196070 61648 196126 61704
rect 195978 53624 196034 53680
rect 195978 53216 196034 53272
rect 194230 51992 194286 52048
rect 194598 47504 194654 47560
rect 197082 46688 197138 46744
rect 265622 276664 265678 276720
rect 428462 271088 428518 271144
rect 412638 262928 412694 262984
rect 580170 697176 580226 697232
rect 580170 683848 580226 683904
rect 580170 670692 580172 670712
rect 580172 670692 580224 670712
rect 580224 670692 580226 670712
rect 580170 670656 580226 670692
rect 580170 644000 580226 644056
rect 580170 630808 580226 630864
rect 580170 617480 580226 617536
rect 579802 590960 579858 591016
rect 580170 577632 580226 577688
rect 579802 564304 579858 564360
rect 580170 537784 580226 537840
rect 580170 524476 580226 524512
rect 580170 524456 580172 524476
rect 580172 524456 580224 524476
rect 580224 524456 580226 524476
rect 580170 511264 580226 511320
rect 580170 484608 580226 484664
rect 579986 471416 580042 471472
rect 580170 458088 580226 458144
rect 580170 431568 580226 431624
rect 580170 418240 580226 418296
rect 580170 404912 580226 404968
rect 580170 378392 580226 378448
rect 580262 365064 580318 365120
rect 580170 351908 580172 351928
rect 580172 351908 580224 351928
rect 580224 351908 580226 351928
rect 580170 351872 580226 351908
rect 580170 325216 580226 325272
rect 579986 312024 580042 312080
rect 580170 298696 580226 298752
rect 580170 272176 580226 272232
rect 477498 262792 477554 262848
rect 199290 210296 199346 210352
rect 198922 200232 198978 200288
rect 197726 137400 197782 137456
rect 197634 79872 197690 79928
rect 197542 65048 197598 65104
rect 197450 56480 197506 56536
rect 198094 80960 198150 81016
rect 198002 80008 198058 80064
rect 198094 78240 198150 78296
rect 198738 147736 198794 147792
rect 197910 67088 197966 67144
rect 197450 56072 197506 56128
rect 197358 45464 197414 45520
rect 197358 44784 197414 44840
rect 580170 258848 580226 258904
rect 580170 245556 580172 245576
rect 580172 245556 580224 245576
rect 580224 245556 580226 245576
rect 580170 245520 580226 245556
rect 580446 232328 580502 232384
rect 580354 219000 580410 219056
rect 579802 205672 579858 205728
rect 200302 200368 200358 200424
rect 199198 77968 199254 78024
rect 199198 68856 199254 68912
rect 199198 68176 199254 68232
rect 198922 63008 198978 63064
rect 198830 55800 198886 55856
rect 204258 200096 204314 200152
rect 200486 152360 200542 152416
rect 201498 173440 201554 173496
rect 200946 80688 201002 80744
rect 201406 77424 201462 77480
rect 200762 71032 200818 71088
rect 200302 67496 200358 67552
rect 200210 53760 200266 53816
rect 200118 50768 200174 50824
rect 201406 68856 201462 68912
rect 201406 67496 201462 67552
rect 201406 66952 201462 67008
rect 201406 53760 201462 53816
rect 201406 53080 201462 53136
rect 201406 50768 201462 50824
rect 201406 50360 201462 50416
rect 201682 58928 201738 58984
rect 201774 55936 201830 55992
rect 202418 71712 202474 71768
rect 202050 61376 202106 61432
rect 202786 71712 202842 71768
rect 202786 71032 202842 71088
rect 202786 58928 202842 58984
rect 202786 58520 202842 58576
rect 202510 49544 202566 49600
rect 203246 46824 203302 46880
rect 201774 44104 201830 44160
rect 202786 44104 202842 44160
rect 202786 43424 202842 43480
rect 204442 49272 204498 49328
rect 204902 78104 204958 78160
rect 204626 52400 204682 52456
rect 204626 51720 204682 51776
rect 204718 49272 204774 49328
rect 204718 48864 204774 48920
rect 204534 48048 204590 48104
rect 204810 48048 204866 48104
rect 204810 47504 204866 47560
rect 205730 75792 205786 75848
rect 206374 78784 206430 78840
rect 207018 77696 207074 77752
rect 206098 75656 206154 75712
rect 205822 50224 205878 50280
rect 205638 42744 205694 42800
rect 205638 42064 205694 42120
rect 208674 192616 208730 192672
rect 580170 192480 580226 192536
rect 580170 179152 580226 179208
rect 580170 165824 580226 165880
rect 580262 152632 580318 152688
rect 286322 139712 286378 139768
rect 208674 76200 208730 76256
rect 213918 67224 213974 67280
rect 208398 64776 208454 64832
rect 208398 64368 208454 64424
rect 209870 54848 209926 54904
rect 212538 45056 212594 45112
rect 220818 68312 220874 68368
rect 229742 73888 229798 73944
rect 229098 30912 229154 30968
rect 231858 56344 231914 56400
rect 242898 67360 242954 67416
rect 245658 61240 245714 61296
rect 249798 62056 249854 62112
rect 260838 76608 260894 76664
rect 259458 64368 259514 64424
rect 267738 44920 267794 44976
rect 264978 28192 265034 28248
rect 274638 65592 274694 65648
rect 277398 61920 277454 61976
rect 278778 53488 278834 53544
rect 284390 43560 284446 43616
rect 327722 139576 327778 139632
rect 291842 77832 291898 77888
rect 292578 63280 292634 63336
rect 299478 60152 299534 60208
rect 304998 73752 305054 73808
rect 576122 140120 576178 140176
rect 382278 79464 382334 79520
rect 313278 57432 313334 57488
rect 315302 56208 315358 56264
rect 320178 61784 320234 61840
rect 331218 63144 331274 63200
rect 327078 58792 327134 58848
rect 333978 54712 334034 54768
rect 338118 60016 338174 60072
rect 351918 53352 351974 53408
rect 356058 50632 356114 50688
rect 362958 58656 363014 58712
rect 364982 54576 365038 54632
rect 369858 52128 369914 52184
rect 373998 51992 374054 52048
rect 380898 65456 380954 65512
rect 382922 61648 382978 61704
rect 387798 53216 387854 53272
rect 390558 47640 390614 47696
rect 400954 56072 401010 56128
rect 405738 50496 405794 50552
rect 408498 44784 408554 44840
rect 423678 67088 423734 67144
rect 414662 63008 414718 63064
rect 418802 57296 418858 57352
rect 430578 66952 430634 67008
rect 423770 54440 423826 54496
rect 437478 61512 437534 61568
rect 432602 53080 432658 53136
rect 440238 50360 440294 50416
rect 468574 77560 468630 77616
rect 450542 55936 450598 55992
rect 452658 43424 452714 43480
rect 454682 49136 454738 49192
rect 459558 61376 459614 61432
rect 463698 46280 463754 46336
rect 476118 51856 476174 51912
rect 486422 75384 486478 75440
rect 484398 51720 484454 51776
rect 489918 55800 489974 55856
rect 494058 49000 494114 49056
rect 495438 46144 495494 46200
rect 521658 75248 521714 75304
rect 504362 68176 504418 68232
rect 507858 42064 507914 42120
rect 511998 64232 512054 64288
rect 514022 62872 514078 62928
rect 520922 47504 520978 47560
rect 525062 59880 525118 59936
rect 553398 76472 553454 76528
rect 549258 75112 549314 75168
rect 543738 71032 543794 71088
rect 539690 58520 539746 58576
rect 547878 64096 547934 64152
rect 545762 57160 545818 57216
rect 561678 69536 561734 69592
rect 557538 66816 557594 66872
rect 567842 62736 567898 62792
rect 565818 48864 565874 48920
rect 569958 50224 570014 50280
rect 580354 139304 580410 139360
rect 580170 86128 580226 86184
rect 579986 72936 580042 72992
rect 580354 137264 580410 137320
rect 580538 125976 580594 126032
rect 580446 112784 580502 112840
rect 580354 99456 580410 99512
rect 580262 59608 580318 59664
rect 579986 19760 580042 19816
rect 580170 6568 580226 6624
<< metal3 >>
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3325 671258 3391 671261
rect -960 671256 3391 671258
rect -960 671200 3330 671256
rect 3386 671200 3391 671256
rect -960 671198 3391 671200
rect -960 671108 480 671198
rect 3325 671195 3391 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3509 658202 3575 658205
rect -960 658200 3575 658202
rect -960 658144 3514 658200
rect 3570 658144 3575 658200
rect -960 658142 3575 658144
rect -960 658052 480 658142
rect 3509 658139 3575 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 3509 632090 3575 632093
rect -960 632088 3575 632090
rect -960 632032 3514 632088
rect 3570 632032 3575 632088
rect -960 632030 3575 632032
rect -960 631940 480 632030
rect 3509 632027 3575 632030
rect 580165 630866 580231 630869
rect 583520 630866 584960 630956
rect 580165 630864 584960 630866
rect 580165 630808 580170 630864
rect 580226 630808 584960 630864
rect 580165 630806 584960 630808
rect 580165 630803 580231 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3509 619170 3575 619173
rect -960 619168 3575 619170
rect -960 619112 3514 619168
rect 3570 619112 3575 619168
rect -960 619110 3575 619112
rect -960 619020 480 619110
rect 3509 619107 3575 619110
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3509 606114 3575 606117
rect -960 606112 3575 606114
rect -960 606056 3514 606112
rect 3570 606056 3575 606112
rect -960 606054 3575 606056
rect -960 605964 480 606054
rect 3509 606051 3575 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 579797 591018 579863 591021
rect 583520 591018 584960 591108
rect 579797 591016 584960 591018
rect 579797 590960 579802 591016
rect 579858 590960 584960 591016
rect 579797 590958 584960 590960
rect 579797 590955 579863 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 3325 580002 3391 580005
rect -960 580000 3391 580002
rect -960 579944 3330 580000
rect 3386 579944 3391 580000
rect -960 579942 3391 579944
rect -960 579852 480 579942
rect 3325 579939 3391 579942
rect 580165 577690 580231 577693
rect 583520 577690 584960 577780
rect 580165 577688 584960 577690
rect 580165 577632 580170 577688
rect 580226 577632 584960 577688
rect 580165 577630 584960 577632
rect 580165 577627 580231 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3233 566946 3299 566949
rect -960 566944 3299 566946
rect -960 566888 3238 566944
rect 3294 566888 3299 566944
rect -960 566886 3299 566888
rect -960 566796 480 566886
rect 3233 566883 3299 566886
rect 579797 564362 579863 564365
rect 583520 564362 584960 564452
rect 579797 564360 584960 564362
rect 579797 564304 579802 564360
rect 579858 564304 584960 564360
rect 579797 564302 584960 564304
rect 579797 564299 579863 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 3325 553890 3391 553893
rect -960 553888 3391 553890
rect -960 553832 3330 553888
rect 3386 553832 3391 553888
rect -960 553830 3391 553832
rect -960 553740 480 553830
rect 3325 553827 3391 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 580165 537842 580231 537845
rect 583520 537842 584960 537932
rect 580165 537840 584960 537842
rect 580165 537784 580170 537840
rect 580226 537784 584960 537840
rect 580165 537782 584960 537784
rect 580165 537779 580231 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 2773 527914 2839 527917
rect -960 527912 2839 527914
rect -960 527856 2778 527912
rect 2834 527856 2839 527912
rect -960 527854 2839 527856
rect -960 527764 480 527854
rect 2773 527851 2839 527854
rect 580165 524514 580231 524517
rect 583520 524514 584960 524604
rect 580165 524512 584960 524514
rect 580165 524456 580170 524512
rect 580226 524456 584960 524512
rect 580165 524454 584960 524456
rect 580165 524451 580231 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 3509 514858 3575 514861
rect -960 514856 3575 514858
rect -960 514800 3514 514856
rect 3570 514800 3575 514856
rect -960 514798 3575 514800
rect -960 514708 480 514798
rect 3509 514795 3575 514798
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 3049 501802 3115 501805
rect -960 501800 3115 501802
rect -960 501744 3054 501800
rect 3110 501744 3115 501800
rect -960 501742 3115 501744
rect -960 501652 480 501742
rect 3049 501739 3115 501742
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 580165 484666 580231 484669
rect 583520 484666 584960 484756
rect 580165 484664 584960 484666
rect 580165 484608 580170 484664
rect 580226 484608 584960 484664
rect 580165 484606 584960 484608
rect 580165 484603 580231 484606
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect 3049 475690 3115 475693
rect -960 475688 3115 475690
rect -960 475632 3054 475688
rect 3110 475632 3115 475688
rect -960 475630 3115 475632
rect -960 475540 480 475630
rect 3049 475627 3115 475630
rect 579981 471474 580047 471477
rect 583520 471474 584960 471564
rect 579981 471472 584960 471474
rect 579981 471416 579986 471472
rect 580042 471416 584960 471472
rect 579981 471414 584960 471416
rect 579981 471411 580047 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 3509 462634 3575 462637
rect -960 462632 3575 462634
rect -960 462576 3514 462632
rect 3570 462576 3575 462632
rect -960 462574 3575 462576
rect -960 462484 480 462574
rect 3509 462571 3575 462574
rect 580165 458146 580231 458149
rect 583520 458146 584960 458236
rect 580165 458144 584960 458146
rect 580165 458088 580170 458144
rect 580226 458088 584960 458144
rect 580165 458086 584960 458088
rect 580165 458083 580231 458086
rect 583520 457996 584960 458086
rect -960 449578 480 449668
rect 3141 449578 3207 449581
rect -960 449576 3207 449578
rect -960 449520 3146 449576
rect 3202 449520 3207 449576
rect -960 449518 3207 449520
rect -960 449428 480 449518
rect 3141 449515 3207 449518
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 580165 431626 580231 431629
rect 583520 431626 584960 431716
rect 580165 431624 584960 431626
rect 580165 431568 580170 431624
rect 580226 431568 584960 431624
rect 580165 431566 584960 431568
rect 580165 431563 580231 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect 3509 423602 3575 423605
rect -960 423600 3575 423602
rect -960 423544 3514 423600
rect 3570 423544 3575 423600
rect -960 423542 3575 423544
rect -960 423452 480 423542
rect 3509 423539 3575 423542
rect 580165 418298 580231 418301
rect 583520 418298 584960 418388
rect 580165 418296 584960 418298
rect 580165 418240 580170 418296
rect 580226 418240 584960 418296
rect 580165 418238 584960 418240
rect 580165 418235 580231 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 2865 410546 2931 410549
rect -960 410544 2931 410546
rect -960 410488 2870 410544
rect 2926 410488 2931 410544
rect -960 410486 2931 410488
rect -960 410396 480 410486
rect 2865 410483 2931 410486
rect 580165 404970 580231 404973
rect 583520 404970 584960 405060
rect 580165 404968 584960 404970
rect 580165 404912 580170 404968
rect 580226 404912 584960 404968
rect 580165 404910 584960 404912
rect 580165 404907 580231 404910
rect 583520 404820 584960 404910
rect -960 397490 480 397580
rect 3509 397490 3575 397493
rect -960 397488 3575 397490
rect -960 397432 3514 397488
rect 3570 397432 3575 397488
rect -960 397430 3575 397432
rect -960 397340 480 397430
rect 3509 397427 3575 397430
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 580165 378450 580231 378453
rect 583520 378450 584960 378540
rect 580165 378448 584960 378450
rect 580165 378392 580170 378448
rect 580226 378392 584960 378448
rect 580165 378390 584960 378392
rect 580165 378387 580231 378390
rect 583520 378300 584960 378390
rect -960 371378 480 371468
rect 3509 371378 3575 371381
rect -960 371376 3575 371378
rect -960 371320 3514 371376
rect 3570 371320 3575 371376
rect -960 371318 3575 371320
rect -960 371228 480 371318
rect 3509 371315 3575 371318
rect 580257 365122 580323 365125
rect 583520 365122 584960 365212
rect 580257 365120 584960 365122
rect 580257 365064 580262 365120
rect 580318 365064 584960 365120
rect 580257 365062 584960 365064
rect 580257 365059 580323 365062
rect 583520 364972 584960 365062
rect -960 358458 480 358548
rect 3141 358458 3207 358461
rect -960 358456 3207 358458
rect -960 358400 3146 358456
rect 3202 358400 3207 358456
rect -960 358398 3207 358400
rect -960 358308 480 358398
rect 3141 358395 3207 358398
rect 580165 351930 580231 351933
rect 583520 351930 584960 352020
rect 580165 351928 584960 351930
rect 580165 351872 580170 351928
rect 580226 351872 584960 351928
rect 580165 351870 584960 351872
rect 580165 351867 580231 351870
rect 583520 351780 584960 351870
rect -960 345402 480 345492
rect 3325 345402 3391 345405
rect -960 345400 3391 345402
rect -960 345344 3330 345400
rect 3386 345344 3391 345400
rect -960 345342 3391 345344
rect -960 345252 480 345342
rect 3325 345339 3391 345342
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 580165 325274 580231 325277
rect 583520 325274 584960 325364
rect 580165 325272 584960 325274
rect 580165 325216 580170 325272
rect 580226 325216 584960 325272
rect 580165 325214 584960 325216
rect 580165 325211 580231 325214
rect 583520 325124 584960 325214
rect -960 319290 480 319380
rect 3325 319290 3391 319293
rect -960 319288 3391 319290
rect -960 319232 3330 319288
rect 3386 319232 3391 319288
rect -960 319230 3391 319232
rect -960 319140 480 319230
rect 3325 319227 3391 319230
rect 579981 312082 580047 312085
rect 583520 312082 584960 312172
rect 579981 312080 584960 312082
rect 579981 312024 579986 312080
rect 580042 312024 584960 312080
rect 579981 312022 584960 312024
rect 579981 312019 580047 312022
rect 583520 311932 584960 312022
rect -960 306234 480 306324
rect 3509 306234 3575 306237
rect -960 306232 3575 306234
rect -960 306176 3514 306232
rect 3570 306176 3575 306232
rect -960 306174 3575 306176
rect -960 306084 480 306174
rect 3509 306171 3575 306174
rect 580165 298754 580231 298757
rect 583520 298754 584960 298844
rect 580165 298752 584960 298754
rect 580165 298696 580170 298752
rect 580226 298696 584960 298752
rect 580165 298694 584960 298696
rect 580165 298691 580231 298694
rect 583520 298604 584960 298694
rect -960 293178 480 293268
rect 3509 293178 3575 293181
rect -960 293176 3575 293178
rect -960 293120 3514 293176
rect 3570 293120 3575 293176
rect -960 293118 3575 293120
rect -960 293028 480 293118
rect 3509 293115 3575 293118
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 265617 276722 265683 276725
rect 190410 276720 265683 276722
rect 190410 276664 265622 276720
rect 265678 276664 265683 276720
rect 190410 276662 265683 276664
rect 154573 276042 154639 276045
rect 189022 276042 189028 276044
rect 154573 276040 189028 276042
rect 154573 275984 154578 276040
rect 154634 275984 189028 276040
rect 154573 275982 189028 275984
rect 154573 275979 154639 275982
rect 189022 275980 189028 275982
rect 189092 276042 189098 276044
rect 190410 276042 190470 276662
rect 265617 276659 265683 276662
rect 189092 275982 190470 276042
rect 189092 275980 189098 275982
rect 580165 272234 580231 272237
rect 583520 272234 584960 272324
rect 580165 272232 584960 272234
rect 580165 272176 580170 272232
rect 580226 272176 584960 272232
rect 580165 272174 584960 272176
rect 580165 272171 580231 272174
rect 583520 272084 584960 272174
rect 186998 271084 187004 271148
rect 187068 271146 187074 271148
rect 428457 271146 428523 271149
rect 187068 271144 428523 271146
rect 187068 271088 428462 271144
rect 428518 271088 428523 271144
rect 187068 271086 428523 271088
rect 187068 271084 187074 271086
rect 428457 271083 428523 271086
rect 151905 270602 151971 270605
rect 186998 270602 187004 270604
rect 151905 270600 187004 270602
rect 151905 270544 151910 270600
rect 151966 270544 187004 270600
rect 151905 270542 187004 270544
rect 151905 270539 151971 270542
rect 186998 270540 187004 270542
rect 187068 270540 187074 270604
rect -960 267202 480 267292
rect 3049 267202 3115 267205
rect -960 267200 3115 267202
rect -960 267144 3054 267200
rect 3110 267144 3115 267200
rect -960 267142 3115 267144
rect -960 267052 480 267142
rect 3049 267139 3115 267142
rect 167637 265298 167703 265301
rect 193254 265298 193260 265300
rect 167637 265296 193260 265298
rect 167637 265240 167642 265296
rect 167698 265240 193260 265296
rect 167637 265238 193260 265240
rect 167637 265235 167703 265238
rect 193254 265236 193260 265238
rect 193324 265236 193330 265300
rect 166257 265162 166323 265165
rect 194542 265162 194548 265164
rect 166257 265160 194548 265162
rect 166257 265104 166262 265160
rect 166318 265104 194548 265160
rect 166257 265102 194548 265104
rect 166257 265099 166323 265102
rect 194542 265100 194548 265102
rect 194612 265100 194618 265164
rect 113030 264964 113036 265028
rect 113100 265026 113106 265028
rect 140129 265026 140195 265029
rect 113100 265024 140195 265026
rect 113100 264968 140134 265024
rect 140190 264968 140195 265024
rect 113100 264966 140195 264968
rect 113100 264964 113106 264966
rect 140129 264963 140195 264966
rect 163405 265026 163471 265029
rect 194726 265026 194732 265028
rect 163405 265024 194732 265026
rect 163405 264968 163410 265024
rect 163466 264968 194732 265024
rect 163405 264966 194732 264968
rect 163405 264963 163471 264966
rect 194726 264964 194732 264966
rect 194796 264964 194802 265028
rect 121126 263740 121132 263804
rect 121196 263802 121202 263804
rect 146937 263802 147003 263805
rect 121196 263800 147003 263802
rect 121196 263744 146942 263800
rect 146998 263744 147003 263800
rect 121196 263742 147003 263744
rect 121196 263740 121202 263742
rect 146937 263739 147003 263742
rect 118550 263604 118556 263668
rect 118620 263666 118626 263668
rect 151077 263666 151143 263669
rect 118620 263664 151143 263666
rect 118620 263608 151082 263664
rect 151138 263608 151143 263664
rect 118620 263606 151143 263608
rect 118620 263604 118626 263606
rect 151077 263603 151143 263606
rect 166073 263258 166139 263261
rect 166349 263258 166415 263261
rect 166073 263256 166415 263258
rect 166073 263200 166078 263256
rect 166134 263200 166354 263256
rect 166410 263200 166415 263256
rect 166073 263198 166415 263200
rect 166073 263195 166139 263198
rect 166349 263195 166415 263198
rect 167545 263122 167611 263125
rect 167729 263122 167795 263125
rect 191966 263122 191972 263124
rect 167545 263120 191972 263122
rect 167545 263064 167550 263120
rect 167606 263064 167734 263120
rect 167790 263064 191972 263120
rect 167545 263062 191972 263064
rect 167545 263059 167611 263062
rect 167729 263059 167795 263062
rect 191966 263060 191972 263062
rect 192036 263060 192042 263124
rect 153009 262986 153075 262989
rect 186589 262986 186655 262989
rect 412633 262986 412699 262989
rect 153009 262984 412699 262986
rect 153009 262928 153014 262984
rect 153070 262928 186594 262984
rect 186650 262928 412638 262984
rect 412694 262928 412699 262984
rect 153009 262926 412699 262928
rect 153009 262923 153075 262926
rect 186589 262923 186655 262926
rect 412633 262923 412699 262926
rect 115790 262788 115796 262852
rect 115860 262850 115866 262852
rect 148317 262850 148383 262853
rect 115860 262848 148383 262850
rect 115860 262792 148322 262848
rect 148378 262792 148383 262848
rect 115860 262790 148383 262792
rect 115860 262788 115866 262790
rect 148317 262787 148383 262790
rect 150433 262850 150499 262853
rect 151353 262850 151419 262853
rect 477493 262850 477559 262853
rect 150433 262848 477559 262850
rect 150433 262792 150438 262848
rect 150494 262792 151358 262848
rect 151414 262792 477498 262848
rect 477554 262792 477559 262848
rect 150433 262790 477559 262792
rect 150433 262787 150499 262790
rect 151353 262787 151419 262790
rect 477493 262787 477559 262790
rect 112846 262652 112852 262716
rect 112916 262714 112922 262716
rect 127893 262714 127959 262717
rect 112916 262712 127959 262714
rect 112916 262656 127898 262712
rect 127954 262656 127959 262712
rect 112916 262654 127959 262656
rect 112916 262652 112922 262654
rect 127893 262651 127959 262654
rect 166073 262714 166139 262717
rect 193438 262714 193444 262716
rect 166073 262712 193444 262714
rect 166073 262656 166078 262712
rect 166134 262656 193444 262712
rect 166073 262654 193444 262656
rect 166073 262651 166139 262654
rect 193438 262652 193444 262654
rect 193508 262652 193514 262716
rect 111558 262516 111564 262580
rect 111628 262578 111634 262580
rect 133321 262578 133387 262581
rect 133689 262578 133755 262581
rect 111628 262576 133755 262578
rect 111628 262520 133326 262576
rect 133382 262520 133694 262576
rect 133750 262520 133755 262576
rect 111628 262518 133755 262520
rect 111628 262516 111634 262518
rect 133321 262515 133387 262518
rect 133689 262515 133755 262518
rect 163681 262578 163747 262581
rect 191782 262578 191788 262580
rect 163681 262576 191788 262578
rect 163681 262520 163686 262576
rect 163742 262520 191788 262576
rect 163681 262518 191788 262520
rect 163681 262515 163747 262518
rect 191782 262516 191788 262518
rect 191852 262516 191858 262580
rect 114134 262380 114140 262444
rect 114204 262442 114210 262444
rect 141417 262442 141483 262445
rect 114204 262440 141483 262442
rect 114204 262384 141422 262440
rect 141478 262384 141483 262440
rect 114204 262382 141483 262384
rect 114204 262380 114210 262382
rect 141417 262379 141483 262382
rect 162117 262442 162183 262445
rect 190494 262442 190500 262444
rect 162117 262440 190500 262442
rect 162117 262384 162122 262440
rect 162178 262384 190500 262440
rect 162117 262382 190500 262384
rect 162117 262379 162183 262382
rect 190494 262380 190500 262382
rect 190564 262380 190570 262444
rect 111374 262244 111380 262308
rect 111444 262306 111450 262308
rect 126237 262306 126303 262309
rect 111444 262304 126303 262306
rect 111444 262248 126242 262304
rect 126298 262248 126303 262304
rect 111444 262246 126303 262248
rect 111444 262244 111450 262246
rect 126237 262243 126303 262246
rect 187969 262306 188035 262309
rect 188102 262306 188108 262308
rect 187969 262304 188108 262306
rect 187969 262248 187974 262304
rect 188030 262248 188108 262304
rect 187969 262246 188108 262248
rect 187969 262243 188035 262246
rect 188102 262244 188108 262246
rect 188172 262244 188178 262308
rect 111190 260884 111196 260948
rect 111260 260946 111266 260948
rect 138289 260946 138355 260949
rect 111260 260944 138355 260946
rect 111260 260888 138294 260944
rect 138350 260888 138355 260944
rect 111260 260886 138355 260888
rect 111260 260884 111266 260886
rect 138289 260883 138355 260886
rect 138013 260810 138079 260813
rect 138933 260810 138999 260813
rect 138013 260808 138999 260810
rect 138013 260752 138018 260808
rect 138074 260752 138938 260808
rect 138994 260752 138999 260808
rect 138013 260750 138999 260752
rect 138013 260747 138079 260750
rect 138933 260747 138999 260750
rect 143809 260810 143875 260813
rect 144453 260810 144519 260813
rect 143809 260808 144519 260810
rect 143809 260752 143814 260808
rect 143870 260752 144458 260808
rect 144514 260752 144519 260808
rect 143809 260750 144519 260752
rect 143809 260747 143875 260750
rect 144453 260747 144519 260750
rect 120942 260476 120948 260540
rect 121012 260538 121018 260540
rect 149237 260538 149303 260541
rect 121012 260536 149303 260538
rect 121012 260480 149242 260536
rect 149298 260480 149303 260536
rect 121012 260478 149303 260480
rect 121012 260476 121018 260478
rect 149237 260475 149303 260478
rect 113582 260340 113588 260404
rect 113652 260402 113658 260404
rect 138013 260402 138079 260405
rect 113652 260400 138079 260402
rect 113652 260344 138018 260400
rect 138074 260344 138079 260400
rect 113652 260342 138079 260344
rect 113652 260340 113658 260342
rect 138013 260339 138079 260342
rect 118366 260204 118372 260268
rect 118436 260266 118442 260268
rect 143717 260266 143783 260269
rect 144913 260266 144979 260269
rect 145879 260266 145945 260269
rect 118436 260264 143783 260266
rect 118436 260208 143722 260264
rect 143778 260208 143783 260264
rect 118436 260206 143783 260208
rect 118436 260204 118442 260206
rect 143717 260203 143783 260206
rect 144686 260264 145945 260266
rect 144686 260208 144918 260264
rect 144974 260208 145884 260264
rect 145940 260208 145945 260264
rect 144686 260206 145945 260208
rect 115606 260068 115612 260132
rect 115676 260130 115682 260132
rect 142245 260130 142311 260133
rect 143119 260130 143185 260133
rect 115676 260128 143185 260130
rect 115676 260072 142250 260128
rect 142306 260072 143124 260128
rect 143180 260072 143185 260128
rect 115676 260070 143185 260072
rect 115676 260068 115682 260070
rect 142245 260067 142311 260070
rect 143119 260067 143185 260070
rect 116894 259932 116900 259996
rect 116964 259994 116970 259996
rect 144545 259994 144611 259997
rect 116964 259992 144611 259994
rect 116964 259936 144550 259992
rect 144606 259936 144611 259992
rect 116964 259934 144611 259936
rect 116964 259932 116970 259934
rect 144545 259931 144611 259934
rect 117078 259796 117084 259860
rect 117148 259858 117154 259860
rect 144686 259858 144746 260206
rect 144913 260203 144979 260206
rect 145879 260203 145945 260206
rect 160093 260266 160159 260269
rect 160783 260266 160849 260269
rect 160093 260264 160849 260266
rect 160093 260208 160098 260264
rect 160154 260208 160788 260264
rect 160844 260208 160849 260264
rect 160093 260206 160849 260208
rect 160093 260203 160159 260206
rect 160783 260203 160849 260206
rect 163497 260266 163563 260269
rect 171041 260266 171107 260269
rect 163497 260264 171107 260266
rect 163497 260208 163502 260264
rect 163558 260208 171046 260264
rect 171102 260208 171107 260264
rect 163497 260206 171107 260208
rect 163497 260203 163563 260206
rect 171041 260203 171107 260206
rect 180885 260266 180951 260269
rect 189349 260266 189415 260269
rect 180885 260264 189415 260266
rect 180885 260208 180890 260264
rect 180946 260208 189354 260264
rect 189410 260208 189415 260264
rect 180885 260206 189415 260208
rect 180885 260203 180951 260206
rect 189349 260203 189415 260206
rect 187969 260130 188035 260133
rect 166766 260128 188035 260130
rect 166766 260072 187974 260128
rect 188030 260072 188035 260128
rect 166766 260070 188035 260072
rect 164233 259994 164299 259997
rect 165061 259994 165127 259997
rect 166766 259994 166826 260070
rect 187969 260067 188035 260070
rect 164233 259992 166826 259994
rect 164233 259936 164238 259992
rect 164294 259936 165066 259992
rect 165122 259936 166826 259992
rect 164233 259934 166826 259936
rect 171041 259994 171107 259997
rect 186865 259994 186931 259997
rect 171041 259992 186931 259994
rect 171041 259936 171046 259992
rect 171102 259936 186870 259992
rect 186926 259936 186931 259992
rect 171041 259934 186931 259936
rect 164233 259931 164299 259934
rect 165061 259931 165127 259934
rect 171041 259931 171107 259934
rect 186865 259931 186931 259934
rect 117148 259798 144746 259858
rect 162117 259858 162183 259861
rect 188153 259858 188219 259861
rect 162117 259856 188219 259858
rect 162117 259800 162122 259856
rect 162178 259800 188158 259856
rect 188214 259800 188219 259856
rect 162117 259798 188219 259800
rect 117148 259796 117154 259798
rect 162117 259795 162183 259798
rect 188153 259795 188219 259798
rect 113950 259660 113956 259724
rect 114020 259722 114026 259724
rect 125685 259722 125751 259725
rect 114020 259720 125751 259722
rect 114020 259664 125690 259720
rect 125746 259664 125751 259720
rect 114020 259662 125751 259664
rect 114020 259660 114026 259662
rect 125685 259659 125751 259662
rect 160921 259722 160987 259725
rect 180885 259722 180951 259725
rect 188429 259722 188495 259725
rect 160921 259720 180951 259722
rect 160921 259664 160926 259720
rect 160982 259664 180890 259720
rect 180946 259664 180951 259720
rect 160921 259662 180951 259664
rect 160921 259659 160987 259662
rect 180885 259659 180951 259662
rect 184614 259720 188495 259722
rect 184614 259664 188434 259720
rect 188490 259664 188495 259720
rect 184614 259662 188495 259664
rect 118233 259588 118299 259589
rect 118182 259586 118188 259588
rect 118142 259526 118188 259586
rect 118252 259584 118299 259588
rect 118294 259528 118299 259584
rect 118182 259524 118188 259526
rect 118252 259524 118299 259528
rect 118233 259523 118299 259524
rect 130837 259586 130903 259589
rect 184614 259586 184674 259662
rect 188429 259659 188495 259662
rect 185393 259588 185459 259589
rect 185342 259586 185348 259588
rect 130837 259584 184674 259586
rect 130837 259528 130842 259584
rect 130898 259528 184674 259584
rect 130837 259526 184674 259528
rect 185302 259526 185348 259586
rect 185412 259584 185459 259588
rect 185454 259528 185459 259584
rect 130837 259523 130903 259526
rect 185342 259524 185348 259526
rect 185412 259524 185459 259528
rect 185393 259523 185459 259524
rect 186037 259588 186103 259589
rect 186037 259584 186084 259588
rect 186148 259586 186154 259588
rect 186037 259528 186042 259584
rect 186037 259524 186084 259528
rect 186148 259526 186194 259586
rect 186148 259524 186154 259526
rect 186037 259523 186103 259524
rect 580165 258906 580231 258909
rect 583520 258906 584960 258996
rect 580165 258904 584960 258906
rect 580165 258848 580170 258904
rect 580226 258848 584960 258904
rect 580165 258846 584960 258848
rect 580165 258843 580231 258846
rect 583520 258756 584960 258846
rect -960 254146 480 254236
rect 3509 254146 3575 254149
rect -960 254144 3575 254146
rect -960 254088 3514 254144
rect 3570 254088 3575 254144
rect -960 254086 3575 254088
rect -960 253996 480 254086
rect 3509 254083 3575 254086
rect 580165 245578 580231 245581
rect 583520 245578 584960 245668
rect 580165 245576 584960 245578
rect 580165 245520 580170 245576
rect 580226 245520 584960 245576
rect 580165 245518 584960 245520
rect 580165 245515 580231 245518
rect 583520 245428 584960 245518
rect -960 241090 480 241180
rect 3509 241090 3575 241093
rect -960 241088 3575 241090
rect -960 241032 3514 241088
rect 3570 241032 3575 241088
rect -960 241030 3575 241032
rect -960 240940 480 241030
rect 3509 241027 3575 241030
rect 580441 232386 580507 232389
rect 583520 232386 584960 232476
rect 580441 232384 584960 232386
rect 580441 232328 580446 232384
rect 580502 232328 584960 232384
rect 580441 232326 584960 232328
rect 580441 232323 580507 232326
rect 583520 232236 584960 232326
rect -960 227884 480 228124
rect 580349 219058 580415 219061
rect 583520 219058 584960 219148
rect 580349 219056 584960 219058
rect 580349 219000 580354 219056
rect 580410 219000 584960 219056
rect 580349 218998 584960 219000
rect 580349 218995 580415 218998
rect 583520 218908 584960 218998
rect -960 214978 480 215068
rect 2773 214978 2839 214981
rect -960 214976 2839 214978
rect -960 214920 2778 214976
rect 2834 214920 2839 214976
rect -960 214918 2839 214920
rect -960 214828 480 214918
rect 2773 214915 2839 214918
rect 186446 210292 186452 210356
rect 186516 210354 186522 210356
rect 199285 210354 199351 210357
rect 186516 210352 199351 210354
rect 186516 210296 199290 210352
rect 199346 210296 199351 210352
rect 186516 210294 199351 210296
rect 186516 210292 186522 210294
rect 199285 210291 199351 210294
rect 579797 205730 579863 205733
rect 583520 205730 584960 205820
rect 579797 205728 584960 205730
rect 579797 205672 579802 205728
rect 579858 205672 584960 205728
rect 579797 205670 584960 205672
rect 579797 205667 579863 205670
rect 583520 205580 584960 205670
rect 186078 202812 186084 202876
rect 186148 202874 186154 202876
rect 187233 202874 187299 202877
rect 186148 202872 187299 202874
rect 186148 202816 187238 202872
rect 187294 202816 187299 202872
rect 186148 202814 187299 202816
rect 186148 202812 186154 202814
rect 187233 202811 187299 202814
rect -960 201922 480 202012
rect 3417 201922 3483 201925
rect -960 201920 3483 201922
rect -960 201864 3422 201920
rect 3478 201864 3483 201920
rect -960 201862 3483 201864
rect -960 201772 480 201862
rect 3417 201859 3483 201862
rect 185342 201724 185348 201788
rect 185412 201786 185418 201788
rect 188337 201786 188403 201789
rect 185412 201784 188403 201786
rect 185412 201728 188342 201784
rect 188398 201728 188403 201784
rect 185412 201726 188403 201728
rect 185412 201724 185418 201726
rect 188337 201723 188403 201726
rect 109953 200698 110019 200701
rect 109953 200696 129750 200698
rect 109953 200640 109958 200696
rect 110014 200640 129750 200696
rect 109953 200638 129750 200640
rect 109953 200635 110019 200638
rect 129690 200426 129750 200638
rect 157190 200636 157196 200700
rect 157260 200698 157266 200700
rect 179822 200698 179828 200700
rect 157260 200638 179828 200698
rect 157260 200636 157266 200638
rect 179822 200636 179828 200638
rect 179892 200636 179898 200700
rect 166206 200500 166212 200564
rect 166276 200562 166282 200564
rect 182950 200562 182956 200564
rect 166276 200502 182956 200562
rect 166276 200500 166282 200502
rect 182950 200500 182956 200502
rect 183020 200500 183026 200564
rect 129690 200366 138076 200426
rect 107193 200290 107259 200293
rect 137870 200290 137876 200292
rect 107193 200288 137876 200290
rect 107193 200232 107198 200288
rect 107254 200232 137876 200288
rect 107193 200230 137876 200232
rect 107193 200227 107259 200230
rect 137870 200228 137876 200230
rect 137940 200228 137946 200292
rect 138016 200290 138076 200366
rect 166574 200364 166580 200428
rect 166644 200426 166650 200428
rect 200297 200426 200363 200429
rect 166644 200424 200363 200426
rect 166644 200368 200302 200424
rect 200358 200368 200363 200424
rect 166644 200366 200363 200368
rect 166644 200364 166650 200366
rect 200297 200363 200363 200366
rect 198917 200290 198983 200293
rect 138016 200230 142354 200290
rect 105629 200154 105695 200157
rect 136398 200154 136404 200156
rect 105629 200152 136404 200154
rect 105629 200096 105634 200152
rect 105690 200096 136404 200152
rect 105629 200094 136404 200096
rect 105629 200091 105695 200094
rect 136398 200092 136404 200094
rect 136468 200092 136474 200156
rect 137502 200092 137508 200156
rect 137572 200154 137578 200156
rect 137572 200094 137938 200154
rect 137572 200092 137578 200094
rect 137878 199919 137938 200094
rect 139526 200092 139532 200156
rect 139596 200092 139602 200156
rect 140814 200092 140820 200156
rect 140884 200154 140890 200156
rect 140884 200094 141802 200154
rect 140884 200092 140890 200094
rect 139534 199919 139594 200092
rect 141742 199919 141802 200094
rect 142294 199919 142354 200230
rect 164742 200288 198983 200290
rect 164742 200232 198922 200288
rect 198978 200232 198983 200288
rect 164742 200230 198983 200232
rect 145414 200092 145420 200156
rect 145484 200154 145490 200156
rect 163446 200154 163452 200156
rect 145484 200094 147874 200154
rect 145484 200092 145490 200094
rect 147814 199919 147874 200094
rect 155634 200094 163452 200154
rect 155634 199919 155694 200094
rect 163446 200092 163452 200094
rect 163516 200092 163522 200156
rect 164742 199919 164802 200230
rect 198917 200227 198983 200230
rect 169150 200092 169156 200156
rect 169220 200154 169226 200156
rect 204253 200154 204319 200157
rect 169220 200094 169586 200154
rect 169220 200092 169226 200094
rect 169526 199919 169586 200094
rect 172470 200152 204319 200154
rect 172470 200096 204258 200152
rect 204314 200096 204319 200152
rect 172470 200094 204319 200096
rect 132723 199914 132789 199919
rect 103237 199882 103303 199885
rect 131665 199882 131731 199885
rect 132723 199884 132728 199914
rect 132784 199884 132789 199914
rect 132907 199914 132973 199919
rect 103237 199880 131731 199882
rect 103237 199824 103242 199880
rect 103298 199824 131670 199880
rect 131726 199824 131731 199880
rect 103237 199822 131731 199824
rect 103237 199819 103303 199822
rect 131665 199819 131731 199822
rect 132718 199820 132724 199884
rect 132788 199882 132794 199884
rect 132788 199822 132846 199882
rect 132907 199858 132912 199914
rect 132968 199882 132973 199914
rect 133459 199914 133525 199919
rect 133459 199884 133464 199914
rect 133520 199884 133525 199914
rect 133919 199916 133985 199919
rect 133919 199914 134258 199916
rect 133086 199882 133092 199884
rect 132968 199858 133092 199882
rect 132907 199853 133092 199858
rect 132910 199822 133092 199853
rect 132788 199820 132794 199822
rect 133086 199820 133092 199822
rect 133156 199820 133162 199884
rect 133454 199820 133460 199884
rect 133524 199882 133530 199884
rect 133524 199822 133582 199882
rect 133919 199858 133924 199914
rect 133980 199884 134258 199914
rect 134747 199914 134813 199919
rect 134379 199884 134445 199885
rect 134747 199884 134752 199914
rect 134808 199884 134813 199914
rect 135115 199914 135181 199919
rect 135115 199884 135120 199914
rect 135176 199884 135181 199914
rect 135299 199914 135365 199919
rect 133980 199858 134196 199884
rect 133919 199856 134196 199858
rect 133919 199853 133985 199856
rect 133524 199820 133530 199822
rect 134190 199820 134196 199856
rect 134260 199820 134266 199884
rect 134374 199820 134380 199884
rect 134444 199882 134450 199884
rect 134444 199822 134536 199882
rect 134444 199820 134450 199822
rect 134742 199820 134748 199884
rect 134812 199882 134818 199884
rect 134812 199822 134870 199882
rect 134812 199820 134818 199822
rect 135110 199820 135116 199884
rect 135180 199882 135186 199884
rect 135180 199822 135238 199882
rect 135299 199858 135304 199914
rect 135360 199882 135365 199914
rect 135851 199914 135917 199919
rect 135851 199884 135856 199914
rect 135912 199884 135917 199914
rect 136587 199914 136653 199919
rect 135478 199882 135484 199884
rect 135360 199858 135484 199882
rect 135299 199853 135484 199858
rect 135302 199822 135484 199853
rect 135180 199820 135186 199822
rect 135478 199820 135484 199822
rect 135548 199820 135554 199884
rect 135846 199820 135852 199884
rect 135916 199882 135922 199884
rect 135916 199822 135974 199882
rect 136587 199858 136592 199914
rect 136648 199882 136653 199914
rect 137139 199914 137205 199919
rect 137139 199884 137144 199914
rect 137200 199884 137205 199914
rect 137323 199914 137389 199919
rect 136950 199882 136956 199884
rect 136648 199858 136956 199882
rect 136587 199853 136956 199858
rect 136590 199822 136956 199853
rect 135916 199820 135922 199822
rect 136950 199820 136956 199822
rect 137020 199820 137026 199884
rect 137134 199820 137140 199884
rect 137204 199882 137210 199884
rect 137204 199822 137262 199882
rect 137323 199858 137328 199914
rect 137384 199882 137389 199914
rect 137875 199914 137941 199919
rect 137686 199882 137692 199884
rect 137384 199858 137692 199882
rect 137323 199853 137692 199858
rect 137326 199822 137692 199853
rect 137204 199820 137210 199822
rect 137686 199820 137692 199822
rect 137756 199820 137762 199884
rect 137875 199858 137880 199914
rect 137936 199858 137941 199914
rect 138059 199914 138125 199919
rect 138059 199884 138064 199914
rect 138120 199884 138125 199914
rect 138427 199914 138493 199919
rect 137875 199853 137941 199858
rect 138054 199820 138060 199884
rect 138124 199882 138130 199884
rect 138124 199822 138182 199882
rect 138427 199858 138432 199914
rect 138488 199882 138493 199914
rect 139163 199914 139229 199919
rect 138606 199882 138612 199884
rect 138488 199858 138612 199882
rect 138427 199853 138612 199858
rect 138430 199822 138612 199853
rect 138124 199820 138130 199822
rect 138606 199820 138612 199822
rect 138676 199820 138682 199884
rect 138790 199820 138796 199884
rect 138860 199882 138866 199884
rect 139163 199882 139168 199914
rect 138860 199858 139168 199882
rect 139224 199858 139229 199914
rect 139347 199914 139413 199919
rect 139347 199884 139352 199914
rect 139408 199884 139413 199914
rect 139531 199914 139597 199919
rect 138860 199853 139229 199858
rect 138860 199822 139226 199853
rect 138860 199820 138866 199822
rect 139342 199820 139348 199884
rect 139412 199882 139418 199884
rect 139412 199822 139470 199882
rect 139531 199858 139536 199914
rect 139592 199858 139597 199914
rect 139715 199914 139781 199919
rect 140175 199916 140241 199919
rect 139715 199884 139720 199914
rect 139776 199884 139781 199914
rect 140132 199914 140241 199916
rect 140132 199884 140180 199914
rect 139531 199853 139597 199858
rect 139412 199820 139418 199822
rect 139710 199820 139716 199884
rect 139780 199882 139786 199884
rect 139780 199822 139838 199882
rect 139780 199820 139786 199822
rect 140078 199820 140084 199884
rect 140148 199858 140180 199884
rect 140236 199858 140241 199914
rect 140451 199914 140517 199919
rect 140451 199884 140456 199914
rect 140512 199884 140517 199914
rect 140727 199914 140793 199919
rect 141279 199916 141345 199919
rect 140148 199853 140241 199858
rect 140148 199822 140192 199853
rect 140148 199820 140154 199822
rect 140446 199820 140452 199884
rect 140516 199882 140522 199884
rect 140516 199822 140574 199882
rect 140727 199858 140732 199914
rect 140788 199882 140793 199914
rect 141236 199914 141345 199916
rect 141236 199884 141284 199914
rect 140998 199882 141004 199884
rect 140788 199858 141004 199882
rect 140727 199853 141004 199858
rect 140730 199822 141004 199853
rect 140516 199820 140522 199822
rect 140998 199820 141004 199822
rect 141068 199820 141074 199884
rect 141182 199820 141188 199884
rect 141252 199858 141284 199884
rect 141340 199858 141345 199914
rect 141252 199853 141345 199858
rect 141739 199914 141805 199919
rect 141739 199858 141744 199914
rect 141800 199858 141805 199914
rect 141739 199853 141805 199858
rect 142291 199914 142357 199919
rect 142291 199858 142296 199914
rect 142352 199858 142357 199914
rect 142475 199914 142541 199919
rect 142475 199884 142480 199914
rect 142536 199884 142541 199914
rect 142659 199914 142725 199919
rect 142291 199853 142357 199858
rect 141252 199822 141296 199853
rect 141252 199820 141258 199822
rect 142470 199820 142476 199884
rect 142540 199882 142546 199884
rect 142540 199822 142598 199882
rect 142659 199858 142664 199914
rect 142720 199858 142725 199914
rect 143027 199914 143093 199919
rect 143027 199884 143032 199914
rect 143088 199884 143093 199914
rect 144499 199914 144565 199919
rect 142659 199853 142725 199858
rect 142540 199820 142546 199822
rect 134379 199819 134445 199820
rect 123477 199746 123543 199749
rect 142662 199748 142722 199853
rect 143022 199820 143028 199884
rect 143092 199882 143098 199884
rect 144499 199882 144504 199914
rect 143092 199822 143150 199882
rect 143214 199858 144504 199882
rect 144560 199858 144565 199914
rect 144683 199914 144749 199919
rect 145695 199916 145761 199919
rect 144683 199884 144688 199914
rect 144744 199884 144749 199914
rect 145652 199914 145761 199916
rect 143214 199853 144565 199858
rect 143214 199822 144562 199853
rect 143092 199820 143098 199822
rect 123477 199744 140790 199746
rect 123477 199688 123482 199744
rect 123538 199688 140790 199744
rect 123477 199686 140790 199688
rect 123477 199683 123543 199686
rect 131297 199610 131363 199613
rect 136449 199612 136515 199613
rect 133086 199610 133092 199612
rect 131297 199608 133092 199610
rect 131297 199552 131302 199608
rect 131358 199552 133092 199608
rect 131297 199550 133092 199552
rect 131297 199547 131363 199550
rect 133086 199548 133092 199550
rect 133156 199548 133162 199612
rect 136398 199610 136404 199612
rect 136358 199550 136404 199610
rect 136468 199608 136515 199612
rect 136510 199552 136515 199608
rect 136398 199548 136404 199550
rect 136468 199548 136515 199552
rect 137870 199548 137876 199612
rect 137940 199610 137946 199612
rect 138013 199610 138079 199613
rect 137940 199608 138079 199610
rect 137940 199552 138018 199608
rect 138074 199552 138079 199608
rect 137940 199550 138079 199552
rect 140730 199610 140790 199686
rect 142654 199684 142660 199748
rect 142724 199684 142730 199748
rect 143073 199746 143139 199749
rect 143214 199746 143274 199822
rect 144678 199820 144684 199884
rect 144748 199882 144754 199884
rect 144748 199822 144806 199882
rect 144748 199820 144754 199822
rect 145046 199820 145052 199884
rect 145116 199882 145122 199884
rect 145652 199882 145700 199914
rect 145116 199858 145700 199882
rect 145756 199858 145761 199914
rect 145116 199853 145761 199858
rect 146339 199914 146405 199919
rect 146339 199858 146344 199914
rect 146400 199882 146405 199914
rect 146707 199914 146773 199919
rect 146707 199884 146712 199914
rect 146768 199884 146773 199914
rect 146891 199914 146957 199919
rect 146518 199882 146524 199884
rect 146400 199858 146524 199882
rect 146339 199853 146524 199858
rect 145116 199822 145712 199853
rect 146342 199822 146524 199853
rect 145116 199820 145122 199822
rect 146518 199820 146524 199822
rect 146588 199820 146594 199884
rect 146702 199820 146708 199884
rect 146772 199882 146778 199884
rect 146772 199822 146830 199882
rect 146891 199858 146896 199914
rect 146952 199858 146957 199914
rect 147075 199914 147141 199919
rect 147075 199884 147080 199914
rect 147136 199884 147141 199914
rect 147811 199914 147877 199919
rect 146891 199853 146957 199858
rect 146772 199820 146778 199822
rect 146894 199748 146954 199853
rect 147070 199820 147076 199884
rect 147140 199882 147146 199884
rect 147140 199822 147198 199882
rect 147811 199858 147816 199914
rect 147872 199858 147877 199914
rect 148179 199914 148245 199919
rect 149007 199916 149073 199919
rect 148179 199884 148184 199914
rect 148240 199884 148245 199914
rect 148964 199914 149073 199916
rect 147811 199853 147877 199858
rect 147140 199820 147146 199822
rect 148174 199820 148180 199884
rect 148244 199882 148250 199884
rect 148244 199822 148302 199882
rect 148964 199858 149012 199914
rect 149068 199858 149073 199914
rect 149283 199914 149349 199919
rect 150295 199916 150361 199919
rect 149283 199884 149288 199914
rect 149344 199884 149349 199914
rect 150252 199914 150361 199916
rect 148964 199853 149073 199858
rect 148244 199820 148250 199822
rect 148964 199749 149024 199853
rect 149278 199820 149284 199884
rect 149348 199882 149354 199884
rect 149348 199822 149406 199882
rect 149348 199820 149354 199822
rect 149646 199820 149652 199884
rect 149716 199882 149722 199884
rect 150252 199882 150300 199914
rect 149716 199858 150300 199882
rect 150356 199858 150361 199914
rect 150939 199914 151005 199919
rect 150939 199884 150944 199914
rect 151000 199884 151005 199914
rect 151123 199914 151189 199919
rect 153055 199916 153121 199919
rect 153791 199916 153857 199919
rect 149716 199853 150361 199858
rect 149716 199822 150312 199853
rect 149716 199820 149722 199822
rect 150934 199820 150940 199884
rect 151004 199882 151010 199884
rect 151004 199822 151062 199882
rect 151123 199858 151128 199914
rect 151184 199858 151189 199914
rect 153012 199914 153121 199916
rect 151123 199853 151189 199858
rect 151004 199820 151010 199822
rect 143073 199744 143274 199746
rect 143073 199688 143078 199744
rect 143134 199688 143274 199744
rect 143073 199686 143274 199688
rect 143073 199683 143139 199686
rect 146886 199684 146892 199748
rect 146956 199684 146962 199748
rect 148961 199744 149027 199749
rect 151126 199748 151186 199853
rect 151494 199822 152474 199882
rect 148961 199688 148966 199744
rect 149022 199688 149027 199744
rect 148961 199683 149027 199688
rect 151118 199684 151124 199748
rect 151188 199684 151194 199748
rect 151494 199610 151554 199822
rect 152414 199746 152474 199822
rect 152590 199820 152596 199884
rect 152660 199882 152666 199884
rect 153012 199882 153060 199914
rect 152660 199858 153060 199882
rect 153116 199858 153121 199914
rect 153748 199914 153857 199916
rect 152660 199853 153121 199858
rect 152660 199822 153072 199853
rect 152660 199820 152666 199822
rect 153326 199820 153332 199884
rect 153396 199882 153402 199884
rect 153748 199882 153796 199914
rect 153396 199858 153796 199882
rect 153852 199858 153857 199914
rect 154435 199914 154501 199919
rect 153396 199853 153857 199858
rect 153396 199822 153808 199853
rect 153396 199820 153402 199822
rect 154062 199820 154068 199884
rect 154132 199882 154138 199884
rect 154435 199882 154440 199914
rect 154132 199858 154440 199882
rect 154496 199858 154501 199914
rect 154987 199914 155053 199919
rect 154132 199853 154501 199858
rect 154132 199822 154498 199853
rect 154132 199820 154138 199822
rect 154614 199820 154620 199884
rect 154684 199882 154690 199884
rect 154987 199882 154992 199914
rect 154684 199858 154992 199882
rect 155048 199858 155053 199914
rect 154684 199853 155053 199858
rect 155631 199914 155697 199919
rect 155999 199916 156065 199919
rect 155631 199858 155636 199914
rect 155692 199858 155697 199914
rect 155956 199914 156065 199916
rect 155956 199884 156004 199914
rect 155631 199853 155697 199858
rect 154684 199822 155050 199853
rect 154684 199820 154690 199822
rect 155902 199820 155908 199884
rect 155972 199858 156004 199884
rect 156060 199858 156065 199914
rect 156459 199914 156525 199919
rect 156459 199882 156464 199914
rect 155972 199853 156065 199858
rect 156278 199858 156464 199882
rect 156520 199858 156525 199914
rect 157195 199914 157261 199919
rect 158023 199916 158089 199919
rect 156278 199853 156525 199858
rect 155972 199822 156016 199853
rect 156278 199822 156522 199853
rect 155972 199820 155978 199822
rect 155953 199746 156019 199749
rect 152414 199744 156019 199746
rect 152414 199688 155958 199744
rect 156014 199688 156019 199744
rect 152414 199686 156019 199688
rect 155953 199683 156019 199686
rect 140730 199550 151554 199610
rect 156278 199610 156338 199822
rect 156638 199820 156644 199884
rect 156708 199882 156714 199884
rect 157195 199882 157200 199914
rect 156708 199858 157200 199882
rect 157256 199858 157261 199914
rect 157980 199914 158089 199916
rect 156708 199853 157261 199858
rect 156708 199822 157258 199853
rect 156708 199820 156714 199822
rect 157742 199820 157748 199884
rect 157812 199882 157818 199884
rect 157980 199882 158028 199914
rect 157812 199858 158028 199882
rect 158084 199858 158089 199914
rect 158299 199914 158365 199919
rect 158299 199882 158304 199914
rect 157812 199853 158089 199858
rect 158164 199858 158304 199882
rect 158360 199858 158365 199914
rect 158164 199853 158365 199858
rect 158575 199916 158641 199919
rect 159679 199916 159745 199919
rect 158575 199914 158776 199916
rect 158575 199858 158580 199914
rect 158636 199858 158776 199914
rect 159636 199914 159745 199916
rect 158575 199856 158776 199858
rect 158575 199853 158641 199856
rect 157812 199822 158040 199853
rect 158164 199822 158362 199853
rect 157812 199820 157818 199822
rect 156454 199684 156460 199748
rect 156524 199746 156530 199748
rect 156689 199746 156755 199749
rect 157149 199748 157215 199749
rect 157149 199746 157196 199748
rect 156524 199744 156755 199746
rect 156524 199688 156694 199744
rect 156750 199688 156755 199744
rect 156524 199686 156755 199688
rect 157104 199744 157196 199746
rect 157104 199688 157154 199744
rect 157104 199686 157196 199688
rect 156524 199684 156530 199686
rect 156689 199683 156755 199686
rect 157149 199684 157196 199686
rect 157260 199684 157266 199748
rect 157926 199684 157932 199748
rect 157996 199746 158002 199748
rect 158164 199746 158224 199822
rect 157996 199686 158224 199746
rect 157996 199684 158002 199686
rect 158294 199684 158300 199748
rect 158364 199746 158370 199748
rect 158716 199746 158776 199856
rect 158846 199820 158852 199884
rect 158916 199882 158922 199884
rect 159636 199882 159684 199914
rect 158916 199858 159684 199882
rect 159740 199858 159745 199914
rect 160139 199914 160205 199919
rect 160139 199884 160144 199914
rect 160200 199884 160205 199914
rect 160875 199914 160941 199919
rect 161335 199916 161401 199919
rect 158916 199853 159745 199858
rect 158916 199822 159696 199853
rect 158916 199820 158922 199822
rect 160134 199820 160140 199884
rect 160204 199882 160210 199884
rect 160204 199822 160262 199882
rect 160875 199858 160880 199914
rect 160936 199858 160941 199914
rect 161292 199914 161401 199916
rect 160875 199853 160941 199858
rect 160204 199820 160210 199822
rect 158364 199686 158776 199746
rect 160878 199746 160938 199853
rect 161054 199820 161060 199884
rect 161124 199882 161130 199884
rect 161292 199882 161340 199914
rect 161124 199858 161340 199882
rect 161396 199858 161401 199914
rect 161611 199914 161677 199919
rect 161611 199884 161616 199914
rect 161672 199884 161677 199914
rect 162071 199916 162137 199919
rect 162623 199916 162689 199919
rect 162071 199914 162180 199916
rect 161124 199853 161401 199858
rect 161124 199822 161352 199853
rect 161124 199820 161130 199822
rect 161606 199820 161612 199884
rect 161676 199882 161682 199884
rect 161676 199822 161734 199882
rect 162071 199858 162076 199914
rect 162132 199858 162180 199914
rect 162580 199914 162689 199916
rect 162071 199853 162180 199858
rect 161676 199820 161682 199822
rect 162120 199749 162180 199853
rect 162342 199820 162348 199884
rect 162412 199882 162418 199884
rect 162580 199882 162628 199914
rect 162412 199858 162628 199882
rect 162684 199858 162689 199914
rect 163267 199914 163333 199919
rect 162991 199882 163057 199885
rect 163267 199884 163272 199914
rect 163328 199884 163333 199914
rect 163727 199916 163793 199919
rect 163727 199914 164066 199916
rect 162412 199853 162689 199858
rect 162948 199880 163057 199882
rect 162412 199822 162640 199853
rect 162948 199824 162996 199880
rect 163052 199824 163057 199880
rect 162412 199820 162418 199822
rect 162948 199819 163057 199824
rect 163262 199820 163268 199884
rect 163332 199882 163338 199884
rect 163332 199822 163390 199882
rect 163451 199880 163517 199885
rect 163451 199824 163456 199880
rect 163512 199824 163517 199880
rect 163727 199858 163732 199914
rect 163788 199858 164066 199914
rect 163727 199856 164066 199858
rect 163727 199853 163793 199856
rect 163332 199820 163338 199822
rect 163451 199819 163517 199824
rect 161565 199746 161631 199749
rect 160878 199744 161631 199746
rect 160878 199688 161570 199744
rect 161626 199688 161631 199744
rect 160878 199686 161631 199688
rect 158364 199684 158370 199686
rect 157149 199683 157215 199684
rect 161565 199683 161631 199686
rect 162117 199744 162183 199749
rect 162948 199748 163008 199819
rect 162117 199688 162122 199744
rect 162178 199688 162183 199744
rect 162117 199683 162183 199688
rect 162894 199684 162900 199748
rect 162964 199686 163008 199748
rect 162964 199684 162970 199686
rect 163078 199684 163084 199748
rect 163148 199746 163154 199748
rect 163454 199746 163514 199819
rect 163148 199686 163514 199746
rect 163773 199746 163839 199749
rect 164006 199746 164066 199856
rect 164739 199914 164805 199919
rect 165199 199916 165265 199919
rect 164739 199858 164744 199914
rect 164800 199858 164805 199914
rect 164926 199914 165265 199916
rect 164926 199884 165204 199914
rect 164739 199853 164805 199858
rect 164918 199820 164924 199884
rect 164988 199858 165204 199884
rect 165260 199858 165265 199914
rect 168051 199914 168117 199919
rect 166947 199884 167013 199885
rect 167867 199884 167933 199885
rect 168051 199884 168056 199914
rect 168112 199884 168117 199914
rect 168235 199914 168301 199919
rect 166942 199882 166948 199884
rect 164988 199856 165265 199858
rect 164988 199820 164994 199856
rect 165199 199853 165265 199856
rect 166856 199822 166948 199882
rect 166942 199820 166948 199822
rect 167012 199820 167018 199884
rect 167862 199882 167868 199884
rect 167776 199822 167868 199882
rect 167862 199820 167868 199822
rect 167932 199820 167938 199884
rect 168046 199820 168052 199884
rect 168116 199882 168122 199884
rect 168116 199822 168174 199882
rect 168235 199858 168240 199914
rect 168296 199858 168301 199914
rect 168603 199914 168669 199919
rect 168603 199884 168608 199914
rect 168664 199884 168669 199914
rect 168879 199916 168945 199919
rect 168879 199914 169172 199916
rect 168235 199853 168301 199858
rect 168116 199820 168122 199822
rect 166947 199819 167013 199820
rect 167867 199819 167933 199820
rect 163773 199744 164066 199746
rect 163773 199688 163778 199744
rect 163834 199688 164066 199744
rect 163773 199686 164066 199688
rect 164693 199746 164759 199749
rect 165470 199746 165476 199748
rect 164693 199744 165476 199746
rect 164693 199688 164698 199744
rect 164754 199688 165476 199744
rect 164693 199686 165476 199688
rect 163148 199684 163154 199686
rect 163773 199683 163839 199686
rect 164693 199683 164759 199686
rect 165470 199684 165476 199686
rect 165540 199684 165546 199748
rect 166257 199746 166323 199749
rect 166809 199748 166875 199749
rect 167545 199748 167611 199749
rect 166574 199746 166580 199748
rect 166257 199744 166580 199746
rect 166257 199688 166262 199744
rect 166318 199688 166580 199744
rect 166257 199686 166580 199688
rect 166257 199683 166323 199686
rect 166574 199684 166580 199686
rect 166644 199684 166650 199748
rect 166758 199746 166764 199748
rect 166718 199686 166764 199746
rect 166828 199744 166875 199748
rect 166870 199688 166875 199744
rect 166758 199684 166764 199686
rect 166828 199684 166875 199688
rect 167494 199684 167500 199748
rect 167564 199746 167611 199748
rect 168097 199746 168163 199749
rect 168238 199746 168298 199853
rect 168598 199820 168604 199884
rect 168668 199882 168674 199884
rect 168668 199822 168726 199882
rect 168879 199858 168884 199914
rect 168940 199882 169172 199914
rect 169523 199914 169589 199919
rect 169334 199882 169340 199884
rect 168940 199858 169340 199882
rect 168879 199856 169340 199858
rect 168879 199853 168945 199856
rect 169112 199822 169340 199856
rect 168668 199820 168674 199822
rect 169334 199820 169340 199822
rect 169404 199820 169410 199884
rect 169523 199858 169528 199914
rect 169584 199858 169589 199914
rect 169523 199853 169589 199858
rect 169707 199914 169773 199919
rect 169707 199858 169712 199914
rect 169768 199858 169773 199914
rect 169707 199853 169773 199858
rect 170535 199914 170601 199919
rect 170535 199858 170540 199914
rect 170596 199858 170601 199914
rect 170995 199914 171061 199919
rect 170995 199884 171000 199914
rect 171056 199884 171061 199914
rect 171179 199914 171245 199919
rect 170535 199853 170601 199858
rect 169710 199749 169770 199853
rect 170538 199749 170598 199853
rect 170990 199820 170996 199884
rect 171060 199882 171066 199884
rect 171060 199822 171118 199882
rect 171179 199858 171184 199914
rect 171240 199858 171245 199914
rect 171179 199853 171245 199858
rect 171547 199882 171613 199885
rect 171726 199882 171732 199884
rect 171547 199880 171732 199882
rect 171060 199820 171066 199822
rect 171182 199749 171242 199853
rect 171547 199824 171552 199880
rect 171608 199824 171732 199880
rect 171547 199822 171732 199824
rect 171547 199819 171613 199822
rect 171726 199820 171732 199822
rect 171796 199820 171802 199884
rect 167564 199744 167656 199746
rect 167606 199688 167656 199744
rect 167564 199686 167656 199688
rect 168097 199744 168298 199746
rect 168097 199688 168102 199744
rect 168158 199688 168298 199744
rect 168097 199686 168298 199688
rect 168741 199746 168807 199749
rect 168966 199746 168972 199748
rect 168741 199744 168972 199746
rect 168741 199688 168746 199744
rect 168802 199688 168972 199744
rect 168741 199686 168972 199688
rect 167564 199684 167611 199686
rect 166809 199683 166875 199684
rect 167545 199683 167611 199684
rect 168097 199683 168163 199686
rect 168741 199683 168807 199686
rect 168966 199684 168972 199686
rect 169036 199684 169042 199748
rect 169710 199744 169819 199749
rect 169710 199688 169758 199744
rect 169814 199688 169819 199744
rect 169710 199686 169819 199688
rect 169753 199683 169819 199686
rect 170029 199748 170095 199749
rect 170029 199744 170076 199748
rect 170140 199746 170146 199748
rect 170029 199688 170034 199744
rect 170029 199684 170076 199688
rect 170140 199686 170186 199746
rect 170489 199744 170598 199749
rect 170489 199688 170494 199744
rect 170550 199688 170598 199744
rect 170489 199686 170598 199688
rect 170673 199746 170739 199749
rect 170857 199746 170923 199749
rect 170673 199744 170923 199746
rect 170673 199688 170678 199744
rect 170734 199688 170862 199744
rect 170918 199688 170923 199744
rect 170673 199686 170923 199688
rect 170140 199684 170146 199686
rect 170029 199683 170095 199684
rect 170489 199683 170555 199686
rect 170673 199683 170739 199686
rect 170857 199683 170923 199686
rect 171133 199744 171242 199749
rect 171133 199688 171138 199744
rect 171194 199688 171242 199744
rect 171133 199686 171242 199688
rect 171501 199746 171567 199749
rect 172470 199746 172530 200094
rect 204253 200091 204319 200094
rect 174307 199914 174373 199919
rect 172830 199820 172836 199884
rect 172900 199882 172906 199884
rect 173203 199882 173269 199885
rect 172900 199880 173269 199882
rect 172900 199824 173208 199880
rect 173264 199824 173269 199880
rect 172900 199822 173269 199824
rect 172900 199820 172906 199822
rect 173203 199819 173269 199822
rect 173387 199880 173453 199885
rect 173387 199824 173392 199880
rect 173448 199824 173453 199880
rect 174307 199858 174312 199914
rect 174368 199882 174373 199914
rect 175411 199914 175477 199919
rect 174486 199882 174492 199884
rect 174368 199858 174492 199882
rect 174307 199853 174492 199858
rect 173387 199819 173453 199824
rect 174310 199822 174492 199853
rect 174486 199820 174492 199822
rect 174556 199820 174562 199884
rect 174859 199882 174925 199885
rect 175411 199884 175416 199914
rect 175472 199884 175477 199914
rect 176515 199914 176581 199919
rect 175038 199882 175044 199884
rect 174859 199880 175044 199882
rect 174859 199824 174864 199880
rect 174920 199824 175044 199880
rect 174859 199822 175044 199824
rect 174859 199819 174925 199822
rect 175038 199820 175044 199822
rect 175108 199820 175114 199884
rect 175406 199820 175412 199884
rect 175476 199882 175482 199884
rect 175963 199882 176029 199885
rect 175476 199822 175534 199882
rect 175782 199880 176029 199882
rect 175782 199824 175968 199880
rect 176024 199824 176029 199880
rect 175782 199822 176029 199824
rect 175476 199820 175482 199822
rect 171501 199744 172530 199746
rect 171501 199688 171506 199744
rect 171562 199688 172530 199744
rect 171501 199686 172530 199688
rect 171133 199683 171199 199686
rect 171501 199683 171567 199686
rect 172646 199684 172652 199748
rect 172716 199746 172722 199748
rect 173249 199746 173315 199749
rect 173390 199748 173450 199819
rect 172716 199744 173315 199746
rect 172716 199688 173254 199744
rect 173310 199688 173315 199744
rect 172716 199686 173315 199688
rect 172716 199684 172722 199686
rect 173249 199683 173315 199686
rect 173382 199684 173388 199748
rect 173452 199684 173458 199748
rect 174118 199684 174124 199748
rect 174188 199746 174194 199748
rect 175181 199746 175247 199749
rect 174188 199744 175247 199746
rect 174188 199688 175186 199744
rect 175242 199688 175247 199744
rect 174188 199686 175247 199688
rect 174188 199684 174194 199686
rect 175181 199683 175247 199686
rect 175457 199746 175523 199749
rect 175782 199748 175842 199822
rect 175963 199819 176029 199822
rect 176331 199880 176397 199885
rect 176515 199884 176520 199914
rect 176576 199884 176581 199914
rect 176883 199914 176949 199919
rect 176331 199824 176336 199880
rect 176392 199824 176397 199880
rect 176331 199819 176397 199824
rect 176510 199820 176516 199884
rect 176580 199882 176586 199884
rect 176580 199822 176638 199882
rect 176883 199858 176888 199914
rect 176944 199882 176949 199914
rect 200982 199882 200988 199884
rect 176944 199858 200988 199882
rect 176883 199853 200988 199858
rect 176886 199822 200988 199853
rect 176580 199820 176586 199822
rect 200982 199820 200988 199822
rect 201052 199820 201058 199884
rect 175590 199746 175596 199748
rect 175457 199744 175596 199746
rect 175457 199688 175462 199744
rect 175518 199688 175596 199744
rect 175457 199686 175596 199688
rect 175457 199683 175523 199686
rect 175590 199684 175596 199686
rect 175660 199684 175666 199748
rect 175774 199684 175780 199748
rect 175844 199684 175850 199748
rect 176334 199746 176394 199819
rect 189206 199746 189212 199748
rect 176334 199686 189212 199746
rect 189206 199684 189212 199686
rect 189276 199684 189282 199748
rect 160369 199610 160435 199613
rect 156278 199608 160435 199610
rect 156278 199552 160374 199608
rect 160430 199552 160435 199608
rect 156278 199550 160435 199552
rect 137940 199548 137946 199550
rect 136449 199547 136515 199548
rect 138013 199547 138079 199550
rect 160369 199547 160435 199550
rect 162393 199610 162459 199613
rect 180742 199610 180748 199612
rect 162393 199608 180748 199610
rect 162393 199552 162398 199608
rect 162454 199552 180748 199608
rect 162393 199550 180748 199552
rect 162393 199547 162459 199550
rect 180742 199548 180748 199550
rect 180812 199548 180818 199612
rect 114369 199474 114435 199477
rect 148961 199474 149027 199477
rect 114369 199472 149027 199474
rect 114369 199416 114374 199472
rect 114430 199416 148966 199472
rect 149022 199416 149027 199472
rect 114369 199414 149027 199416
rect 114369 199411 114435 199414
rect 148961 199411 149027 199414
rect 151169 199474 151235 199477
rect 182582 199474 182588 199476
rect 151169 199472 182588 199474
rect 151169 199416 151174 199472
rect 151230 199416 182588 199472
rect 151169 199414 182588 199416
rect 151169 199411 151235 199414
rect 182582 199412 182588 199414
rect 182652 199412 182658 199476
rect 133965 199338 134031 199341
rect 134190 199338 134196 199340
rect 133965 199336 134196 199338
rect 133965 199280 133970 199336
rect 134026 199280 134196 199336
rect 133965 199278 134196 199280
rect 133965 199275 134031 199278
rect 134190 199276 134196 199278
rect 134260 199276 134266 199340
rect 135253 199338 135319 199341
rect 135478 199338 135484 199340
rect 135253 199336 135484 199338
rect 135253 199280 135258 199336
rect 135314 199280 135484 199336
rect 135253 199278 135484 199280
rect 135253 199275 135319 199278
rect 135478 199276 135484 199278
rect 135548 199276 135554 199340
rect 140405 199338 140471 199341
rect 146886 199338 146892 199340
rect 140405 199336 146892 199338
rect 140405 199280 140410 199336
rect 140466 199280 146892 199336
rect 140405 199278 146892 199280
rect 140405 199275 140471 199278
rect 146886 199276 146892 199278
rect 146956 199276 146962 199340
rect 151721 199338 151787 199341
rect 183502 199338 183508 199340
rect 151721 199336 183508 199338
rect 151721 199280 151726 199336
rect 151782 199280 183508 199336
rect 151721 199278 183508 199280
rect 151721 199275 151787 199278
rect 183502 199276 183508 199278
rect 183572 199276 183578 199340
rect 135478 199140 135484 199204
rect 135548 199202 135554 199204
rect 136541 199202 136607 199205
rect 135548 199200 136607 199202
rect 135548 199144 136546 199200
rect 136602 199144 136607 199200
rect 135548 199142 136607 199144
rect 135548 199140 135554 199142
rect 136541 199139 136607 199142
rect 138933 199202 138999 199205
rect 140078 199202 140084 199204
rect 138933 199200 140084 199202
rect 138933 199144 138938 199200
rect 138994 199144 140084 199200
rect 138933 199142 140084 199144
rect 138933 199139 138999 199142
rect 140078 199140 140084 199142
rect 140148 199140 140154 199204
rect 142613 199202 142679 199205
rect 145046 199202 145052 199204
rect 142613 199200 145052 199202
rect 142613 199144 142618 199200
rect 142674 199144 145052 199200
rect 142613 199142 145052 199144
rect 142613 199139 142679 199142
rect 145046 199140 145052 199142
rect 145116 199140 145122 199204
rect 150934 199140 150940 199204
rect 151004 199202 151010 199204
rect 151004 199142 171150 199202
rect 151004 199140 151010 199142
rect 120717 199066 120783 199069
rect 152917 199066 152983 199069
rect 120717 199064 152983 199066
rect 120717 199008 120722 199064
rect 120778 199008 152922 199064
rect 152978 199008 152983 199064
rect 120717 199006 152983 199008
rect 120717 199003 120783 199006
rect 152917 199003 152983 199006
rect 165429 199066 165495 199069
rect 166206 199066 166212 199068
rect 165429 199064 166212 199066
rect 165429 199008 165434 199064
rect 165490 199008 166212 199064
rect 165429 199006 166212 199008
rect 165429 199003 165495 199006
rect 166206 199004 166212 199006
rect 166276 199004 166282 199068
rect 171090 199066 171150 199142
rect 178166 199066 178172 199068
rect 171090 199006 178172 199066
rect 178166 199004 178172 199006
rect 178236 199004 178242 199068
rect 118601 198930 118667 198933
rect 152365 198930 152431 198933
rect 118601 198928 152431 198930
rect 118601 198872 118606 198928
rect 118662 198872 152370 198928
rect 152426 198872 152431 198928
rect 118601 198870 152431 198872
rect 118601 198867 118667 198870
rect 152365 198867 152431 198870
rect 163446 198868 163452 198932
rect 163516 198930 163522 198932
rect 180425 198930 180491 198933
rect 163516 198928 180491 198930
rect 163516 198872 180430 198928
rect 180486 198872 180491 198928
rect 163516 198870 180491 198872
rect 163516 198868 163522 198870
rect 180425 198867 180491 198870
rect 146109 198794 146175 198797
rect 118650 198792 146175 198794
rect 118650 198736 146114 198792
rect 146170 198736 146175 198792
rect 118650 198734 146175 198736
rect 111701 198658 111767 198661
rect 118650 198658 118710 198734
rect 146109 198731 146175 198734
rect 170489 198794 170555 198797
rect 173433 198794 173499 198797
rect 170489 198792 173499 198794
rect 170489 198736 170494 198792
rect 170550 198736 173438 198792
rect 173494 198736 173499 198792
rect 170489 198734 173499 198736
rect 170489 198731 170555 198734
rect 173433 198731 173499 198734
rect 174813 198794 174879 198797
rect 201718 198794 201724 198796
rect 174813 198792 201724 198794
rect 174813 198736 174818 198792
rect 174874 198736 201724 198792
rect 174813 198734 201724 198736
rect 174813 198731 174879 198734
rect 201718 198732 201724 198734
rect 201788 198732 201794 198796
rect 111701 198656 118710 198658
rect 111701 198600 111706 198656
rect 111762 198600 118710 198656
rect 111701 198598 118710 198600
rect 111701 198595 111767 198598
rect 131021 198522 131087 198525
rect 140446 198522 140452 198524
rect 131021 198520 140452 198522
rect 131021 198464 131026 198520
rect 131082 198464 140452 198520
rect 131021 198462 140452 198464
rect 131021 198459 131087 198462
rect 140446 198460 140452 198462
rect 140516 198460 140522 198524
rect 142337 198522 142403 198525
rect 148174 198522 148180 198524
rect 142337 198520 148180 198522
rect 142337 198464 142342 198520
rect 142398 198464 148180 198520
rect 142337 198462 148180 198464
rect 142337 198459 142403 198462
rect 148174 198460 148180 198462
rect 148244 198460 148250 198524
rect 133873 198388 133939 198389
rect 133822 198386 133828 198388
rect 133782 198326 133828 198386
rect 133892 198384 133939 198388
rect 133934 198328 133939 198384
rect 133822 198324 133828 198326
rect 133892 198324 133939 198328
rect 134190 198324 134196 198388
rect 134260 198386 134266 198388
rect 134333 198386 134399 198389
rect 134260 198384 134399 198386
rect 134260 198328 134338 198384
rect 134394 198328 134399 198384
rect 134260 198326 134399 198328
rect 134260 198324 134266 198326
rect 133873 198323 133939 198324
rect 134333 198323 134399 198326
rect 134977 198386 135043 198389
rect 135110 198386 135116 198388
rect 134977 198384 135116 198386
rect 134977 198328 134982 198384
rect 135038 198328 135116 198384
rect 134977 198326 135116 198328
rect 134977 198323 135043 198326
rect 135110 198324 135116 198326
rect 135180 198324 135186 198388
rect 136081 198386 136147 198389
rect 136214 198386 136220 198388
rect 136081 198384 136220 198386
rect 136081 198328 136086 198384
rect 136142 198328 136220 198384
rect 136081 198326 136220 198328
rect 136081 198323 136147 198326
rect 136214 198324 136220 198326
rect 136284 198324 136290 198388
rect 138933 198386 138999 198389
rect 141182 198386 141188 198388
rect 138933 198384 141188 198386
rect 138933 198328 138938 198384
rect 138994 198328 141188 198384
rect 138933 198326 141188 198328
rect 138933 198323 138999 198326
rect 141182 198324 141188 198326
rect 141252 198324 141258 198388
rect 162761 198386 162827 198389
rect 162894 198386 162900 198388
rect 162761 198384 162900 198386
rect 162761 198328 162766 198384
rect 162822 198328 162900 198384
rect 162761 198326 162900 198328
rect 162761 198323 162827 198326
rect 162894 198324 162900 198326
rect 162964 198324 162970 198388
rect 120349 198250 120415 198253
rect 162945 198252 163011 198253
rect 142654 198250 142660 198252
rect 120349 198248 142660 198250
rect 120349 198192 120354 198248
rect 120410 198192 142660 198248
rect 120349 198190 142660 198192
rect 120349 198187 120415 198190
rect 142654 198188 142660 198190
rect 142724 198188 142730 198252
rect 162894 198250 162900 198252
rect 162854 198190 162900 198250
rect 162964 198248 163011 198252
rect 163006 198192 163011 198248
rect 162894 198188 162900 198190
rect 162964 198188 163011 198192
rect 162945 198187 163011 198188
rect 167637 198252 167703 198253
rect 167637 198248 167684 198252
rect 167748 198250 167754 198252
rect 170213 198250 170279 198253
rect 196382 198250 196388 198252
rect 167637 198192 167642 198248
rect 167637 198188 167684 198192
rect 167748 198190 167794 198250
rect 170213 198248 196388 198250
rect 170213 198192 170218 198248
rect 170274 198192 196388 198248
rect 170213 198190 196388 198192
rect 167748 198188 167754 198190
rect 167637 198187 167703 198188
rect 170213 198187 170279 198190
rect 196382 198188 196388 198190
rect 196452 198188 196458 198252
rect 108757 198114 108823 198117
rect 139853 198114 139919 198117
rect 108757 198112 139919 198114
rect 108757 198056 108762 198112
rect 108818 198056 139858 198112
rect 139914 198056 139919 198112
rect 108757 198054 139919 198056
rect 108757 198051 108823 198054
rect 139853 198051 139919 198054
rect 140313 198114 140379 198117
rect 140446 198114 140452 198116
rect 140313 198112 140452 198114
rect 140313 198056 140318 198112
rect 140374 198056 140452 198112
rect 140313 198054 140452 198056
rect 140313 198051 140379 198054
rect 140446 198052 140452 198054
rect 140516 198052 140522 198116
rect 141785 198114 141851 198117
rect 142429 198116 142495 198117
rect 142286 198114 142292 198116
rect 141785 198112 142292 198114
rect 141785 198056 141790 198112
rect 141846 198056 142292 198112
rect 141785 198054 142292 198056
rect 141785 198051 141851 198054
rect 142286 198052 142292 198054
rect 142356 198052 142362 198116
rect 142429 198112 142476 198116
rect 142540 198114 142546 198116
rect 162945 198114 163011 198117
rect 163313 198116 163379 198117
rect 163078 198114 163084 198116
rect 142429 198056 142434 198112
rect 142429 198052 142476 198056
rect 142540 198054 142586 198114
rect 162945 198112 163084 198114
rect 162945 198056 162950 198112
rect 163006 198056 163084 198112
rect 162945 198054 163084 198056
rect 142540 198052 142546 198054
rect 142429 198051 142495 198052
rect 162945 198051 163011 198054
rect 163078 198052 163084 198054
rect 163148 198052 163154 198116
rect 163262 198052 163268 198116
rect 163332 198114 163379 198116
rect 164601 198114 164667 198117
rect 166993 198116 167059 198117
rect 167913 198116 167979 198117
rect 168097 198116 168163 198117
rect 164918 198114 164924 198116
rect 163332 198112 163424 198114
rect 163374 198056 163424 198112
rect 163332 198054 163424 198056
rect 164601 198112 164924 198114
rect 164601 198056 164606 198112
rect 164662 198056 164924 198112
rect 164601 198054 164924 198056
rect 163332 198052 163379 198054
rect 163313 198051 163379 198052
rect 164601 198051 164667 198054
rect 164918 198052 164924 198054
rect 164988 198052 164994 198116
rect 166942 198052 166948 198116
rect 167012 198114 167059 198116
rect 167862 198114 167868 198116
rect 167012 198112 167104 198114
rect 167054 198056 167104 198112
rect 167012 198054 167104 198056
rect 167822 198054 167868 198114
rect 167932 198112 167979 198116
rect 167974 198056 167979 198112
rect 167012 198052 167059 198054
rect 167862 198052 167868 198054
rect 167932 198052 167979 198056
rect 168046 198052 168052 198116
rect 168116 198114 168163 198116
rect 170765 198114 170831 198117
rect 198774 198114 198780 198116
rect 168116 198112 168208 198114
rect 168158 198056 168208 198112
rect 168116 198054 168208 198056
rect 170765 198112 198780 198114
rect 170765 198056 170770 198112
rect 170826 198056 198780 198112
rect 170765 198054 198780 198056
rect 168116 198052 168163 198054
rect 166993 198051 167059 198052
rect 167913 198051 167979 198052
rect 168097 198051 168163 198052
rect 170765 198051 170831 198054
rect 198774 198052 198780 198054
rect 198844 198052 198850 198116
rect 132769 197980 132835 197981
rect 133505 197980 133571 197981
rect 132718 197916 132724 197980
rect 132788 197978 132835 197980
rect 132788 197976 132880 197978
rect 132830 197920 132880 197976
rect 132788 197918 132880 197920
rect 132788 197916 132835 197918
rect 133454 197916 133460 197980
rect 133524 197978 133571 197980
rect 134333 197978 134399 197981
rect 135846 197978 135852 197980
rect 133524 197976 133616 197978
rect 133566 197920 133616 197976
rect 133524 197918 133616 197920
rect 134333 197976 135852 197978
rect 134333 197920 134338 197976
rect 134394 197920 135852 197976
rect 134333 197918 135852 197920
rect 133524 197916 133571 197918
rect 132769 197915 132835 197916
rect 133505 197915 133571 197916
rect 134333 197915 134399 197918
rect 135846 197916 135852 197918
rect 135916 197916 135922 197980
rect 136265 197978 136331 197981
rect 137134 197978 137140 197980
rect 136265 197976 137140 197978
rect 136265 197920 136270 197976
rect 136326 197920 137140 197976
rect 136265 197918 137140 197920
rect 136265 197915 136331 197918
rect 137134 197916 137140 197918
rect 137204 197916 137210 197980
rect 149605 197978 149671 197981
rect 176745 197978 176811 197981
rect 149605 197976 176811 197978
rect 149605 197920 149610 197976
rect 149666 197920 176750 197976
rect 176806 197920 176811 197976
rect 149605 197918 176811 197920
rect 149605 197915 149671 197918
rect 176745 197915 176811 197918
rect 132309 197844 132375 197845
rect 134517 197844 134583 197845
rect 134793 197844 134859 197845
rect 132309 197840 132356 197844
rect 132420 197842 132426 197844
rect 132309 197784 132314 197840
rect 132309 197780 132356 197784
rect 132420 197782 132466 197842
rect 134517 197840 134564 197844
rect 134628 197842 134634 197844
rect 134517 197784 134522 197840
rect 132420 197780 132426 197782
rect 134517 197780 134564 197784
rect 134628 197782 134674 197842
rect 134628 197780 134634 197782
rect 134742 197780 134748 197844
rect 134812 197842 134859 197844
rect 134812 197840 134904 197842
rect 134854 197784 134904 197840
rect 134812 197782 134904 197784
rect 134812 197780 134859 197782
rect 135110 197780 135116 197844
rect 135180 197842 135186 197844
rect 135345 197842 135411 197845
rect 135180 197840 135411 197842
rect 135180 197784 135350 197840
rect 135406 197784 135411 197840
rect 135180 197782 135411 197784
rect 135180 197780 135186 197782
rect 132309 197779 132375 197780
rect 134517 197779 134583 197780
rect 134793 197779 134859 197780
rect 135345 197779 135411 197782
rect 135846 197780 135852 197844
rect 135916 197842 135922 197844
rect 135989 197842 136055 197845
rect 135916 197840 136055 197842
rect 135916 197784 135994 197840
rect 136050 197784 136055 197840
rect 135916 197782 136055 197784
rect 135916 197780 135922 197782
rect 135989 197779 136055 197782
rect 167494 197780 167500 197844
rect 167564 197842 167570 197844
rect 167729 197842 167795 197845
rect 167564 197840 167795 197842
rect 167564 197784 167734 197840
rect 167790 197784 167795 197840
rect 167564 197782 167795 197784
rect 167564 197780 167570 197782
rect 167729 197779 167795 197782
rect 134149 197706 134215 197709
rect 134374 197706 134380 197708
rect 134149 197704 134380 197706
rect 134149 197648 134154 197704
rect 134210 197648 134380 197704
rect 134149 197646 134380 197648
rect 134149 197643 134215 197646
rect 134374 197644 134380 197646
rect 134444 197644 134450 197708
rect 134241 197570 134307 197573
rect 134374 197570 134380 197572
rect 134241 197568 134380 197570
rect 134241 197512 134246 197568
rect 134302 197512 134380 197568
rect 134241 197510 134380 197512
rect 134241 197507 134307 197510
rect 134374 197508 134380 197510
rect 134444 197508 134450 197572
rect 176745 197570 176811 197573
rect 179454 197570 179460 197572
rect 176745 197568 179460 197570
rect 176745 197512 176750 197568
rect 176806 197512 179460 197568
rect 176745 197510 179460 197512
rect 176745 197507 176811 197510
rect 179454 197508 179460 197510
rect 179524 197508 179530 197572
rect 121310 197236 121316 197300
rect 121380 197298 121386 197300
rect 154297 197298 154363 197301
rect 121380 197296 154363 197298
rect 121380 197240 154302 197296
rect 154358 197240 154363 197296
rect 121380 197238 154363 197240
rect 121380 197236 121386 197238
rect 154297 197235 154363 197238
rect 138657 196890 138723 196893
rect 139342 196890 139348 196892
rect 138657 196888 139348 196890
rect 138657 196832 138662 196888
rect 138718 196832 139348 196888
rect 138657 196830 139348 196832
rect 138657 196827 138723 196830
rect 139342 196828 139348 196830
rect 139412 196828 139418 196892
rect 154573 196890 154639 196893
rect 183686 196890 183692 196892
rect 154573 196888 183692 196890
rect 154573 196832 154578 196888
rect 154634 196832 183692 196888
rect 154573 196830 183692 196832
rect 154573 196827 154639 196830
rect 183686 196828 183692 196830
rect 183756 196828 183762 196892
rect 119981 196754 120047 196757
rect 153101 196754 153167 196757
rect 119981 196752 153167 196754
rect 119981 196696 119986 196752
rect 120042 196696 153106 196752
rect 153162 196696 153167 196752
rect 119981 196694 153167 196696
rect 119981 196691 120047 196694
rect 153101 196691 153167 196694
rect 154021 196754 154087 196757
rect 187734 196754 187740 196756
rect 154021 196752 187740 196754
rect 154021 196696 154026 196752
rect 154082 196696 187740 196752
rect 154021 196694 187740 196696
rect 154021 196691 154087 196694
rect 187734 196692 187740 196694
rect 187804 196692 187810 196756
rect 153745 196618 153811 196621
rect 187918 196618 187924 196620
rect 153745 196616 187924 196618
rect 153745 196560 153750 196616
rect 153806 196560 187924 196616
rect 153745 196558 187924 196560
rect 153745 196555 153811 196558
rect 187918 196556 187924 196558
rect 187988 196556 187994 196620
rect 168598 196420 168604 196484
rect 168668 196482 168674 196484
rect 169937 196482 170003 196485
rect 168668 196480 170003 196482
rect 168668 196424 169942 196480
rect 169998 196424 170003 196480
rect 168668 196422 170003 196424
rect 168668 196420 168674 196422
rect 169937 196419 170003 196422
rect 169334 195876 169340 195940
rect 169404 195938 169410 195940
rect 169937 195938 170003 195941
rect 169404 195936 170003 195938
rect 169404 195880 169942 195936
rect 169998 195880 170003 195936
rect 169404 195878 170003 195880
rect 169404 195876 169410 195878
rect 169937 195875 170003 195878
rect 139853 195802 139919 195805
rect 144678 195802 144684 195804
rect 139853 195800 144684 195802
rect 139853 195744 139858 195800
rect 139914 195744 144684 195800
rect 139853 195742 144684 195744
rect 139853 195739 139919 195742
rect 144678 195740 144684 195742
rect 144748 195740 144754 195804
rect 152181 195666 152247 195669
rect 187182 195666 187188 195668
rect 152181 195664 187188 195666
rect 152181 195608 152186 195664
rect 152242 195608 187188 195664
rect 152181 195606 187188 195608
rect 152181 195603 152247 195606
rect 187182 195604 187188 195606
rect 187252 195604 187258 195668
rect 138657 195394 138723 195397
rect 140998 195394 141004 195396
rect 138657 195392 141004 195394
rect 138657 195336 138662 195392
rect 138718 195336 141004 195392
rect 138657 195334 141004 195336
rect 138657 195331 138723 195334
rect 140998 195332 141004 195334
rect 141068 195332 141074 195396
rect 104801 195122 104867 195125
rect 135110 195122 135116 195124
rect 104801 195120 135116 195122
rect 104801 195064 104806 195120
rect 104862 195064 135116 195120
rect 104801 195062 135116 195064
rect 104801 195059 104867 195062
rect 135110 195060 135116 195062
rect 135180 195060 135186 195124
rect 120165 194850 120231 194853
rect 138790 194850 138796 194852
rect 120165 194848 138796 194850
rect 120165 194792 120170 194848
rect 120226 194792 138796 194848
rect 120165 194790 138796 194792
rect 120165 194787 120231 194790
rect 138790 194788 138796 194790
rect 138860 194788 138866 194852
rect 130326 194244 130332 194308
rect 130396 194306 130402 194308
rect 149421 194306 149487 194309
rect 130396 194304 149487 194306
rect 130396 194248 149426 194304
rect 149482 194248 149487 194304
rect 130396 194246 149487 194248
rect 130396 194244 130402 194246
rect 149421 194243 149487 194246
rect 155033 194034 155099 194037
rect 184974 194034 184980 194036
rect 155033 194032 184980 194034
rect 155033 193976 155038 194032
rect 155094 193976 184980 194032
rect 155033 193974 184980 193976
rect 155033 193971 155099 193974
rect 184974 193972 184980 193974
rect 185044 193972 185050 194036
rect 115565 193898 115631 193901
rect 149697 193898 149763 193901
rect 115565 193896 149763 193898
rect 115565 193840 115570 193896
rect 115626 193840 149702 193896
rect 149758 193840 149763 193896
rect 115565 193838 149763 193840
rect 115565 193835 115631 193838
rect 149697 193835 149763 193838
rect 169385 193898 169451 193901
rect 203006 193898 203012 193900
rect 169385 193896 203012 193898
rect 169385 193840 169390 193896
rect 169446 193840 203012 193896
rect 169385 193838 203012 193840
rect 169385 193835 169451 193838
rect 203006 193836 203012 193838
rect 203076 193836 203082 193900
rect 127566 193700 127572 193764
rect 127636 193762 127642 193764
rect 149237 193762 149303 193765
rect 127636 193760 149303 193762
rect 127636 193704 149242 193760
rect 149298 193704 149303 193760
rect 127636 193702 149303 193704
rect 127636 193700 127642 193702
rect 149237 193699 149303 193702
rect 161657 193354 161723 193357
rect 178350 193354 178356 193356
rect 161657 193352 178356 193354
rect 161657 193296 161662 193352
rect 161718 193296 178356 193352
rect 161657 193294 178356 193296
rect 161657 193291 161723 193294
rect 178350 193292 178356 193294
rect 178420 193292 178426 193356
rect 157517 193082 157583 193085
rect 179638 193082 179644 193084
rect 157517 193080 179644 193082
rect 157517 193024 157522 193080
rect 157578 193024 179644 193080
rect 157517 193022 179644 193024
rect 157517 193019 157583 193022
rect 179638 193020 179644 193022
rect 179708 193020 179714 193084
rect 124990 192884 124996 192948
rect 125060 192946 125066 192948
rect 145649 192946 145715 192949
rect 125060 192944 145715 192946
rect 125060 192888 145654 192944
rect 145710 192888 145715 192944
rect 125060 192886 145715 192888
rect 125060 192884 125066 192886
rect 145649 192883 145715 192886
rect 156413 192946 156479 192949
rect 180926 192946 180932 192948
rect 156413 192944 180932 192946
rect 156413 192888 156418 192944
rect 156474 192888 180932 192944
rect 156413 192886 180932 192888
rect 156413 192883 156479 192886
rect 180926 192884 180932 192886
rect 180996 192884 181002 192948
rect 104249 192810 104315 192813
rect 135437 192810 135503 192813
rect 104249 192808 135503 192810
rect 104249 192752 104254 192808
rect 104310 192752 135442 192808
rect 135498 192752 135503 192808
rect 104249 192750 135503 192752
rect 104249 192747 104315 192750
rect 135437 192747 135503 192750
rect 165245 192810 165311 192813
rect 196198 192810 196204 192812
rect 165245 192808 196204 192810
rect 165245 192752 165250 192808
rect 165306 192752 196204 192808
rect 165245 192750 196204 192752
rect 165245 192747 165311 192750
rect 196198 192748 196204 192750
rect 196268 192748 196274 192812
rect 149462 192612 149468 192676
rect 149532 192674 149538 192676
rect 159081 192674 159147 192677
rect 149532 192672 159147 192674
rect 149532 192616 159086 192672
rect 159142 192616 159147 192672
rect 149532 192614 159147 192616
rect 149532 192612 149538 192614
rect 159081 192611 159147 192614
rect 175406 192612 175412 192676
rect 175476 192674 175482 192676
rect 208669 192674 208735 192677
rect 175476 192672 208735 192674
rect 175476 192616 208674 192672
rect 208730 192616 208735 192672
rect 175476 192614 208735 192616
rect 175476 192612 175482 192614
rect 208669 192611 208735 192614
rect 106733 192538 106799 192541
rect 141601 192538 141667 192541
rect 106733 192536 141667 192538
rect 106733 192480 106738 192536
rect 106794 192480 141606 192536
rect 141662 192480 141667 192536
rect 106733 192478 141667 192480
rect 106733 192475 106799 192478
rect 141601 192475 141667 192478
rect 162853 192538 162919 192541
rect 196014 192538 196020 192540
rect 162853 192536 196020 192538
rect 162853 192480 162858 192536
rect 162914 192480 196020 192536
rect 162853 192478 196020 192480
rect 162853 192475 162919 192478
rect 196014 192476 196020 192478
rect 196084 192476 196090 192540
rect 580165 192538 580231 192541
rect 583520 192538 584960 192628
rect 580165 192536 584960 192538
rect 580165 192480 580170 192536
rect 580226 192480 584960 192536
rect 580165 192478 584960 192480
rect 580165 192475 580231 192478
rect 138013 192404 138079 192405
rect 138013 192400 138060 192404
rect 138124 192402 138130 192404
rect 138013 192344 138018 192400
rect 138013 192340 138060 192344
rect 138124 192342 138170 192402
rect 583520 192388 584960 192478
rect 138124 192340 138130 192342
rect 138013 192339 138079 192340
rect 122966 192204 122972 192268
rect 123036 192266 123042 192268
rect 143349 192266 143415 192269
rect 123036 192264 143415 192266
rect 123036 192208 143354 192264
rect 143410 192208 143415 192264
rect 123036 192206 143415 192208
rect 123036 192204 123042 192206
rect 143349 192203 143415 192206
rect 127750 192068 127756 192132
rect 127820 192130 127826 192132
rect 143441 192130 143507 192133
rect 127820 192128 143507 192130
rect 127820 192072 143446 192128
rect 143502 192072 143507 192128
rect 127820 192070 143507 192072
rect 127820 192068 127826 192070
rect 143441 192067 143507 192070
rect 124806 191796 124812 191860
rect 124876 191858 124882 191860
rect 143533 191858 143599 191861
rect 124876 191856 143599 191858
rect 124876 191800 143538 191856
rect 143594 191800 143599 191856
rect 124876 191798 143599 191800
rect 124876 191796 124882 191798
rect 143533 191795 143599 191798
rect 126830 191388 126836 191452
rect 126900 191450 126906 191452
rect 146661 191450 146727 191453
rect 126900 191448 146727 191450
rect 126900 191392 146666 191448
rect 146722 191392 146727 191448
rect 126900 191390 146727 191392
rect 126900 191388 126906 191390
rect 146661 191387 146727 191390
rect 122230 191252 122236 191316
rect 122300 191314 122306 191316
rect 147673 191314 147739 191317
rect 122300 191312 147739 191314
rect 122300 191256 147678 191312
rect 147734 191256 147739 191312
rect 122300 191254 147739 191256
rect 122300 191252 122306 191254
rect 147673 191251 147739 191254
rect 124070 191116 124076 191180
rect 124140 191178 124146 191180
rect 143625 191178 143691 191181
rect 149329 191180 149395 191181
rect 124140 191176 143691 191178
rect 124140 191120 143630 191176
rect 143686 191120 143691 191176
rect 124140 191118 143691 191120
rect 124140 191116 124146 191118
rect 143625 191115 143691 191118
rect 149278 191116 149284 191180
rect 149348 191178 149395 191180
rect 149348 191176 149440 191178
rect 149390 191120 149440 191176
rect 149348 191118 149440 191120
rect 149348 191116 149395 191118
rect 149329 191115 149395 191116
rect 112897 191042 112963 191045
rect 144729 191042 144795 191045
rect 112897 191040 144795 191042
rect 112897 190984 112902 191040
rect 112958 190984 144734 191040
rect 144790 190984 144795 191040
rect 112897 190982 144795 190984
rect 112897 190979 112963 190982
rect 144729 190979 144795 190982
rect 131982 190844 131988 190908
rect 132052 190906 132058 190908
rect 148041 190906 148107 190909
rect 132052 190904 148107 190906
rect 132052 190848 148046 190904
rect 148102 190848 148107 190904
rect 132052 190846 148107 190848
rect 132052 190844 132058 190846
rect 148041 190843 148107 190846
rect 130878 190708 130884 190772
rect 130948 190770 130954 190772
rect 144453 190770 144519 190773
rect 130948 190768 144519 190770
rect 130948 190712 144458 190768
rect 144514 190712 144519 190768
rect 130948 190710 144519 190712
rect 130948 190708 130954 190710
rect 144453 190707 144519 190710
rect 130694 190572 130700 190636
rect 130764 190634 130770 190636
rect 143809 190634 143875 190637
rect 130764 190632 143875 190634
rect 130764 190576 143814 190632
rect 143870 190576 143875 190632
rect 130764 190574 143875 190576
rect 130764 190572 130770 190574
rect 143809 190571 143875 190574
rect 130510 190436 130516 190500
rect 130580 190498 130586 190500
rect 144085 190498 144151 190501
rect 130580 190496 144151 190498
rect 130580 190440 144090 190496
rect 144146 190440 144151 190496
rect 130580 190438 144151 190440
rect 130580 190436 130586 190438
rect 144085 190435 144151 190438
rect 165797 190498 165863 190501
rect 178534 190498 178540 190500
rect 165797 190496 178540 190498
rect 165797 190440 165802 190496
rect 165858 190440 178540 190496
rect 165797 190438 178540 190440
rect 165797 190435 165863 190438
rect 178534 190436 178540 190438
rect 178604 190436 178610 190500
rect 125174 190300 125180 190364
rect 125244 190362 125250 190364
rect 145741 190362 145807 190365
rect 125244 190360 145807 190362
rect 125244 190304 145746 190360
rect 145802 190304 145807 190360
rect 125244 190302 145807 190304
rect 125244 190300 125250 190302
rect 145741 190299 145807 190302
rect 138473 190090 138539 190093
rect 144310 190090 144316 190092
rect 138473 190088 144316 190090
rect 138473 190032 138478 190088
rect 138534 190032 144316 190088
rect 138473 190030 144316 190032
rect 138473 190027 138539 190030
rect 144310 190028 144316 190030
rect 144380 190028 144386 190092
rect 122598 189892 122604 189956
rect 122668 189954 122674 189956
rect 147121 189954 147187 189957
rect 122668 189952 147187 189954
rect 122668 189896 147126 189952
rect 147182 189896 147187 189952
rect 122668 189894 147187 189896
rect 122668 189892 122674 189894
rect 147121 189891 147187 189894
rect 138933 189818 138999 189821
rect 139710 189818 139716 189820
rect 138933 189816 139716 189818
rect 138933 189760 138938 189816
rect 138994 189760 139716 189816
rect 138933 189758 139716 189760
rect 138933 189755 138999 189758
rect 139710 189756 139716 189758
rect 139780 189756 139786 189820
rect 113766 189620 113772 189684
rect 113836 189682 113842 189684
rect 140497 189682 140563 189685
rect 113836 189680 140563 189682
rect 113836 189624 140502 189680
rect 140558 189624 140563 189680
rect 113836 189622 140563 189624
rect 113836 189620 113842 189622
rect 140497 189619 140563 189622
rect -960 188866 480 188956
rect 3417 188866 3483 188869
rect -960 188864 3483 188866
rect -960 188808 3422 188864
rect 3478 188808 3483 188864
rect -960 188806 3483 188808
rect -960 188716 480 188806
rect 3417 188803 3483 188806
rect 126646 187308 126652 187372
rect 126716 187370 126722 187372
rect 146702 187370 146708 187372
rect 126716 187310 146708 187370
rect 126716 187308 126722 187310
rect 146702 187308 146708 187310
rect 146772 187308 146778 187372
rect 127382 187172 127388 187236
rect 127452 187234 127458 187236
rect 148133 187234 148199 187237
rect 127452 187232 148199 187234
rect 127452 187176 148138 187232
rect 148194 187176 148199 187232
rect 127452 187174 148199 187176
rect 127452 187172 127458 187174
rect 148133 187171 148199 187174
rect 163221 186962 163287 186965
rect 163630 186962 163636 186964
rect 163221 186960 163636 186962
rect 163221 186904 163226 186960
rect 163282 186904 163636 186960
rect 163221 186902 163636 186904
rect 163221 186899 163287 186902
rect 163630 186900 163636 186902
rect 163700 186900 163706 186964
rect 108297 186826 108363 186829
rect 137001 186826 137067 186829
rect 108297 186824 137067 186826
rect 108297 186768 108302 186824
rect 108358 186768 137006 186824
rect 137062 186768 137067 186824
rect 108297 186766 137067 186768
rect 108297 186763 108363 186766
rect 137001 186763 137067 186766
rect 162894 186764 162900 186828
rect 162964 186826 162970 186828
rect 163221 186826 163287 186829
rect 162964 186824 163287 186826
rect 162964 186768 163226 186824
rect 163282 186768 163287 186824
rect 162964 186766 163287 186768
rect 162964 186764 162970 186766
rect 163221 186763 163287 186766
rect 122414 186628 122420 186692
rect 122484 186690 122490 186692
rect 136633 186690 136699 186693
rect 122484 186688 136699 186690
rect 122484 186632 136638 186688
rect 136694 186632 136699 186688
rect 122484 186630 136699 186632
rect 122484 186628 122490 186630
rect 136633 186627 136699 186630
rect 148542 186628 148548 186692
rect 148612 186690 148618 186692
rect 161606 186690 161612 186692
rect 148612 186630 161612 186690
rect 148612 186628 148618 186630
rect 161606 186628 161612 186630
rect 161676 186628 161682 186692
rect 104433 186554 104499 186557
rect 137185 186556 137251 186557
rect 136214 186554 136220 186556
rect 104433 186552 136220 186554
rect 104433 186496 104438 186552
rect 104494 186496 136220 186552
rect 104433 186494 136220 186496
rect 104433 186491 104499 186494
rect 136214 186492 136220 186494
rect 136284 186492 136290 186556
rect 137134 186554 137140 186556
rect 137094 186494 137140 186554
rect 137204 186552 137251 186556
rect 137246 186496 137251 186552
rect 137134 186492 137140 186494
rect 137204 186492 137251 186496
rect 161422 186492 161428 186556
rect 161492 186554 161498 186556
rect 169845 186554 169911 186557
rect 161492 186552 169911 186554
rect 161492 186496 169850 186552
rect 169906 186496 169911 186552
rect 161492 186494 169911 186496
rect 161492 186492 161498 186494
rect 137185 186491 137251 186492
rect 169845 186491 169911 186494
rect 176653 186554 176719 186557
rect 201902 186554 201908 186556
rect 176653 186552 201908 186554
rect 176653 186496 176658 186552
rect 176714 186496 201908 186552
rect 176653 186494 201908 186496
rect 176653 186491 176719 186494
rect 201902 186492 201908 186494
rect 201972 186492 201978 186556
rect 150893 186418 150959 186421
rect 151302 186418 151308 186420
rect 150893 186416 151308 186418
rect 150893 186360 150898 186416
rect 150954 186360 151308 186416
rect 150893 186358 151308 186360
rect 150893 186355 150959 186358
rect 151302 186356 151308 186358
rect 151372 186356 151378 186420
rect 151854 186356 151860 186420
rect 151924 186418 151930 186420
rect 152733 186418 152799 186421
rect 151924 186416 152799 186418
rect 151924 186360 152738 186416
rect 152794 186360 152799 186416
rect 151924 186358 152799 186360
rect 151924 186356 151930 186358
rect 152733 186355 152799 186358
rect 153510 186356 153516 186420
rect 153580 186418 153586 186420
rect 153837 186418 153903 186421
rect 153580 186416 153903 186418
rect 153580 186360 153842 186416
rect 153898 186360 153903 186416
rect 153580 186358 153903 186360
rect 153580 186356 153586 186358
rect 153837 186355 153903 186358
rect 162158 186356 162164 186420
rect 162228 186418 162234 186420
rect 162669 186418 162735 186421
rect 162228 186416 162735 186418
rect 162228 186360 162674 186416
rect 162730 186360 162735 186416
rect 162228 186358 162735 186360
rect 162228 186356 162234 186358
rect 162669 186355 162735 186358
rect 163313 186418 163379 186421
rect 163998 186418 164004 186420
rect 163313 186416 164004 186418
rect 163313 186360 163318 186416
rect 163374 186360 164004 186416
rect 163313 186358 164004 186360
rect 163313 186355 163379 186358
rect 163998 186356 164004 186358
rect 164068 186356 164074 186420
rect 164601 186418 164667 186421
rect 164918 186418 164924 186420
rect 164601 186416 164924 186418
rect 164601 186360 164606 186416
rect 164662 186360 164924 186416
rect 164601 186358 164924 186360
rect 164601 186355 164667 186358
rect 164918 186356 164924 186358
rect 164988 186356 164994 186420
rect 169886 186356 169892 186420
rect 169956 186418 169962 186420
rect 170990 186418 170996 186420
rect 169956 186358 170996 186418
rect 169956 186356 169962 186358
rect 170990 186356 170996 186358
rect 171060 186356 171066 186420
rect 135713 186282 135779 186285
rect 139209 186284 139275 186285
rect 136030 186282 136036 186284
rect 135713 186280 136036 186282
rect 135713 186224 135718 186280
rect 135774 186224 136036 186280
rect 135713 186222 136036 186224
rect 135713 186219 135779 186222
rect 136030 186220 136036 186222
rect 136100 186220 136106 186284
rect 139158 186220 139164 186284
rect 139228 186282 139275 186284
rect 139228 186280 139320 186282
rect 139270 186224 139320 186280
rect 139228 186222 139320 186224
rect 139228 186220 139275 186222
rect 139526 186220 139532 186284
rect 139596 186282 139602 186284
rect 139853 186282 139919 186285
rect 139596 186280 139919 186282
rect 139596 186224 139858 186280
rect 139914 186224 139919 186280
rect 139596 186222 139919 186224
rect 139596 186220 139602 186222
rect 139209 186219 139275 186220
rect 139853 186219 139919 186222
rect 140129 186282 140195 186285
rect 140262 186282 140268 186284
rect 140129 186280 140268 186282
rect 140129 186224 140134 186280
rect 140190 186224 140268 186280
rect 140129 186222 140268 186224
rect 140129 186219 140195 186222
rect 140262 186220 140268 186222
rect 140332 186220 140338 186284
rect 146886 186220 146892 186284
rect 146956 186282 146962 186284
rect 147489 186282 147555 186285
rect 146956 186280 147555 186282
rect 146956 186224 147494 186280
rect 147550 186224 147555 186280
rect 146956 186222 147555 186224
rect 146956 186220 146962 186222
rect 147489 186219 147555 186222
rect 148174 186220 148180 186284
rect 148244 186282 148250 186284
rect 148869 186282 148935 186285
rect 153285 186284 153351 186285
rect 153285 186282 153332 186284
rect 148244 186280 148935 186282
rect 148244 186224 148874 186280
rect 148930 186224 148935 186280
rect 148244 186222 148935 186224
rect 153240 186280 153332 186282
rect 153240 186224 153290 186280
rect 153240 186222 153332 186224
rect 148244 186220 148250 186222
rect 148869 186219 148935 186222
rect 153285 186220 153332 186222
rect 153396 186220 153402 186284
rect 153653 186282 153719 186285
rect 154062 186282 154068 186284
rect 153653 186280 154068 186282
rect 153653 186224 153658 186280
rect 153714 186224 154068 186280
rect 153653 186222 154068 186224
rect 153285 186219 153351 186220
rect 153653 186219 153719 186222
rect 154062 186220 154068 186222
rect 154132 186220 154138 186284
rect 155902 186220 155908 186284
rect 155972 186282 155978 186284
rect 156045 186282 156111 186285
rect 155972 186280 156111 186282
rect 155972 186224 156050 186280
rect 156106 186224 156111 186280
rect 155972 186222 156111 186224
rect 155972 186220 155978 186222
rect 156045 186219 156111 186222
rect 158110 186220 158116 186284
rect 158180 186282 158186 186284
rect 158253 186282 158319 186285
rect 158180 186280 158319 186282
rect 158180 186224 158258 186280
rect 158314 186224 158319 186280
rect 158180 186222 158319 186224
rect 158180 186220 158186 186222
rect 158253 186219 158319 186222
rect 160134 186220 160140 186284
rect 160204 186282 160210 186284
rect 160461 186282 160527 186285
rect 160204 186280 160527 186282
rect 160204 186224 160466 186280
rect 160522 186224 160527 186280
rect 160204 186222 160527 186224
rect 160204 186220 160210 186222
rect 160461 186219 160527 186222
rect 162485 186284 162551 186285
rect 162485 186280 162532 186284
rect 162596 186282 162602 186284
rect 162485 186224 162490 186280
rect 162485 186220 162532 186224
rect 162596 186222 162642 186282
rect 162596 186220 162602 186222
rect 163262 186220 163268 186284
rect 163332 186282 163338 186284
rect 164049 186282 164115 186285
rect 163332 186280 164115 186282
rect 163332 186224 164054 186280
rect 164110 186224 164115 186280
rect 163332 186222 164115 186224
rect 163332 186220 163338 186222
rect 162485 186219 162551 186220
rect 164049 186219 164115 186222
rect 164734 186220 164740 186284
rect 164804 186282 164810 186284
rect 164877 186282 164943 186285
rect 164804 186280 164943 186282
rect 164804 186224 164882 186280
rect 164938 186224 164943 186280
rect 164804 186222 164943 186224
rect 164804 186220 164810 186222
rect 164877 186219 164943 186222
rect 170581 186282 170647 186285
rect 170990 186282 170996 186284
rect 170581 186280 170996 186282
rect 170581 186224 170586 186280
rect 170642 186224 170996 186280
rect 170581 186222 170996 186224
rect 170581 186219 170647 186222
rect 170990 186220 170996 186222
rect 171060 186220 171066 186284
rect 174302 186220 174308 186284
rect 174372 186282 174378 186284
rect 174537 186282 174603 186285
rect 174372 186280 174603 186282
rect 174372 186224 174542 186280
rect 174598 186224 174603 186280
rect 174372 186222 174603 186224
rect 174372 186220 174378 186222
rect 174537 186219 174603 186222
rect 176285 186282 176351 186285
rect 176510 186282 176516 186284
rect 176285 186280 176516 186282
rect 176285 186224 176290 186280
rect 176346 186224 176516 186280
rect 176285 186222 176516 186224
rect 176285 186219 176351 186222
rect 176510 186220 176516 186222
rect 176580 186220 176586 186284
rect 176878 186220 176884 186284
rect 176948 186282 176954 186284
rect 177849 186282 177915 186285
rect 176948 186280 177915 186282
rect 176948 186224 177854 186280
rect 177910 186224 177915 186280
rect 176948 186222 177915 186224
rect 176948 186220 176954 186222
rect 177849 186219 177915 186222
rect 132861 186146 132927 186149
rect 133086 186146 133092 186148
rect 132861 186144 133092 186146
rect 132861 186088 132866 186144
rect 132922 186088 133092 186144
rect 132861 186086 133092 186088
rect 132861 186083 132927 186086
rect 133086 186084 133092 186086
rect 133156 186084 133162 186148
rect 134333 186146 134399 186149
rect 134558 186146 134564 186148
rect 134333 186144 134564 186146
rect 134333 186088 134338 186144
rect 134394 186088 134564 186144
rect 134333 186086 134564 186088
rect 134333 186083 134399 186086
rect 134558 186084 134564 186086
rect 134628 186084 134634 186148
rect 149278 186084 149284 186148
rect 149348 186146 149354 186148
rect 160185 186146 160251 186149
rect 149348 186144 160251 186146
rect 149348 186088 160190 186144
rect 160246 186088 160251 186144
rect 149348 186086 160251 186088
rect 149348 186084 149354 186086
rect 160185 186083 160251 186086
rect 162894 186084 162900 186148
rect 162964 186146 162970 186148
rect 163497 186146 163563 186149
rect 162964 186144 163563 186146
rect 162964 186088 163502 186144
rect 163558 186088 163563 186144
rect 162964 186086 163563 186088
rect 162964 186084 162970 186086
rect 163497 186083 163563 186086
rect 172881 186146 172947 186149
rect 173382 186146 173388 186148
rect 172881 186144 173388 186146
rect 172881 186088 172886 186144
rect 172942 186088 173388 186144
rect 172881 186086 173388 186088
rect 172881 186083 172947 186086
rect 173382 186084 173388 186086
rect 173452 186084 173458 186148
rect 125358 185948 125364 186012
rect 125428 186010 125434 186012
rect 145373 186010 145439 186013
rect 125428 186008 145439 186010
rect 125428 185952 145378 186008
rect 145434 185952 145439 186008
rect 125428 185950 145439 185952
rect 125428 185948 125434 185950
rect 145373 185947 145439 185950
rect 173198 185948 173204 186012
rect 173268 186010 173274 186012
rect 173709 186010 173775 186013
rect 173268 186008 173775 186010
rect 173268 185952 173714 186008
rect 173770 185952 173775 186008
rect 173268 185950 173775 185952
rect 173268 185948 173274 185950
rect 173709 185947 173775 185950
rect 107469 185874 107535 185877
rect 136950 185874 136956 185876
rect 107469 185872 136956 185874
rect 107469 185816 107474 185872
rect 107530 185816 136956 185872
rect 107469 185814 136956 185816
rect 107469 185811 107535 185814
rect 136950 185812 136956 185814
rect 137020 185812 137026 185876
rect 142654 185812 142660 185876
rect 142724 185874 142730 185876
rect 158161 185874 158227 185877
rect 169201 185876 169267 185877
rect 142724 185872 158227 185874
rect 142724 185816 158166 185872
rect 158222 185816 158227 185872
rect 142724 185814 158227 185816
rect 142724 185812 142730 185814
rect 158161 185811 158227 185814
rect 169150 185812 169156 185876
rect 169220 185874 169267 185876
rect 175641 185874 175707 185877
rect 175958 185874 175964 185876
rect 169220 185872 169312 185874
rect 169262 185816 169312 185872
rect 169220 185814 169312 185816
rect 175641 185872 175964 185874
rect 175641 185816 175646 185872
rect 175702 185816 175964 185872
rect 175641 185814 175964 185816
rect 169220 185812 169267 185814
rect 169201 185811 169267 185812
rect 175641 185811 175707 185814
rect 175958 185812 175964 185814
rect 176028 185812 176034 185876
rect 119838 185676 119844 185740
rect 119908 185738 119914 185740
rect 132125 185738 132191 185741
rect 119908 185736 132191 185738
rect 119908 185680 132130 185736
rect 132186 185680 132191 185736
rect 119908 185678 132191 185680
rect 119908 185676 119914 185678
rect 132125 185675 132191 185678
rect 132769 185738 132835 185741
rect 133454 185738 133460 185740
rect 132769 185736 133460 185738
rect 132769 185680 132774 185736
rect 132830 185680 133460 185736
rect 132769 185678 133460 185680
rect 132769 185675 132835 185678
rect 133454 185676 133460 185678
rect 133524 185676 133530 185740
rect 133873 185738 133939 185741
rect 134926 185738 134932 185740
rect 133873 185736 134932 185738
rect 133873 185680 133878 185736
rect 133934 185680 134932 185736
rect 133873 185678 134932 185680
rect 133873 185675 133939 185678
rect 134926 185676 134932 185678
rect 134996 185676 135002 185740
rect 139117 185738 139183 185741
rect 165981 185740 166047 185741
rect 147070 185738 147076 185740
rect 139117 185736 147076 185738
rect 139117 185680 139122 185736
rect 139178 185680 147076 185736
rect 139117 185678 147076 185680
rect 139117 185675 139183 185678
rect 147070 185676 147076 185678
rect 147140 185676 147146 185740
rect 165981 185736 166028 185740
rect 166092 185738 166098 185740
rect 165981 185680 165986 185736
rect 165981 185676 166028 185680
rect 166092 185678 166138 185738
rect 166092 185676 166098 185678
rect 166206 185676 166212 185740
rect 166276 185738 166282 185740
rect 166901 185738 166967 185741
rect 166276 185736 166967 185738
rect 166276 185680 166906 185736
rect 166962 185680 166967 185736
rect 166276 185678 166967 185680
rect 166276 185676 166282 185678
rect 165981 185675 166047 185676
rect 166901 185675 166967 185678
rect 167310 185676 167316 185740
rect 167380 185738 167386 185740
rect 167729 185738 167795 185741
rect 167380 185736 167795 185738
rect 167380 185680 167734 185736
rect 167790 185680 167795 185736
rect 167380 185678 167795 185680
rect 167380 185676 167386 185678
rect 167729 185675 167795 185678
rect 169150 185676 169156 185740
rect 169220 185738 169226 185740
rect 169293 185738 169359 185741
rect 169220 185736 169359 185738
rect 169220 185680 169298 185736
rect 169354 185680 169359 185736
rect 169220 185678 169359 185680
rect 169220 185676 169226 185678
rect 169293 185675 169359 185678
rect 172237 185740 172303 185741
rect 172237 185736 172284 185740
rect 172348 185738 172354 185740
rect 175733 185738 175799 185741
rect 200614 185738 200620 185740
rect 172237 185680 172242 185736
rect 172237 185676 172284 185680
rect 172348 185678 172394 185738
rect 175733 185736 200620 185738
rect 175733 185680 175738 185736
rect 175794 185680 200620 185736
rect 175733 185678 200620 185680
rect 172348 185676 172354 185678
rect 172237 185675 172303 185676
rect 175733 185675 175799 185678
rect 200614 185676 200620 185678
rect 200684 185676 200690 185740
rect 131614 185540 131620 185604
rect 131684 185602 131690 185604
rect 132401 185602 132467 185605
rect 131684 185600 132467 185602
rect 131684 185544 132406 185600
rect 132462 185544 132467 185600
rect 131684 185542 132467 185544
rect 131684 185540 131690 185542
rect 132401 185539 132467 185542
rect 132902 185540 132908 185604
rect 132972 185602 132978 185604
rect 133689 185602 133755 185605
rect 132972 185600 133755 185602
rect 132972 185544 133694 185600
rect 133750 185544 133755 185600
rect 132972 185542 133755 185544
rect 132972 185540 132978 185542
rect 133689 185539 133755 185542
rect 134241 185602 134307 185605
rect 134374 185602 134380 185604
rect 134241 185600 134380 185602
rect 134241 185544 134246 185600
rect 134302 185544 134380 185600
rect 134241 185542 134380 185544
rect 134241 185539 134307 185542
rect 134374 185540 134380 185542
rect 134444 185540 134450 185604
rect 134558 185540 134564 185604
rect 134628 185602 134634 185604
rect 134977 185602 135043 185605
rect 134628 185600 135043 185602
rect 134628 185544 134982 185600
rect 135038 185544 135043 185600
rect 134628 185542 135043 185544
rect 134628 185540 134634 185542
rect 134977 185539 135043 185542
rect 137093 185602 137159 185605
rect 140589 185604 140655 185605
rect 137686 185602 137692 185604
rect 137093 185600 137692 185602
rect 137093 185544 137098 185600
rect 137154 185544 137692 185600
rect 137093 185542 137692 185544
rect 137093 185539 137159 185542
rect 137686 185540 137692 185542
rect 137756 185540 137762 185604
rect 140589 185600 140636 185604
rect 140700 185602 140706 185604
rect 140589 185544 140594 185600
rect 140589 185540 140636 185544
rect 140700 185542 140746 185602
rect 140700 185540 140706 185542
rect 140998 185540 141004 185604
rect 141068 185602 141074 185604
rect 141969 185602 142035 185605
rect 142981 185604 143047 185605
rect 149881 185604 149947 185605
rect 142981 185602 143028 185604
rect 141068 185600 142035 185602
rect 141068 185544 141974 185600
rect 142030 185544 142035 185600
rect 141068 185542 142035 185544
rect 142936 185600 143028 185602
rect 142936 185544 142986 185600
rect 142936 185542 143028 185544
rect 141068 185540 141074 185542
rect 140589 185539 140655 185540
rect 141969 185539 142035 185542
rect 142981 185540 143028 185542
rect 143092 185540 143098 185604
rect 149830 185602 149836 185604
rect 149790 185542 149836 185602
rect 149900 185600 149947 185604
rect 149942 185544 149947 185600
rect 149830 185540 149836 185542
rect 149900 185540 149947 185544
rect 142981 185539 143047 185540
rect 149881 185539 149947 185540
rect 151445 185604 151511 185605
rect 152273 185604 152339 185605
rect 151445 185600 151492 185604
rect 151556 185602 151562 185604
rect 152222 185602 152228 185604
rect 151445 185544 151450 185600
rect 151445 185540 151492 185544
rect 151556 185542 151602 185602
rect 152182 185542 152228 185602
rect 152292 185600 152339 185604
rect 152334 185544 152339 185600
rect 151556 185540 151562 185542
rect 152222 185540 152228 185542
rect 152292 185540 152339 185544
rect 151445 185539 151511 185540
rect 152273 185539 152339 185540
rect 152549 185604 152615 185605
rect 152549 185600 152596 185604
rect 152660 185602 152666 185604
rect 152549 185544 152554 185600
rect 152549 185540 152596 185544
rect 152660 185542 152706 185602
rect 152660 185540 152666 185542
rect 153694 185540 153700 185604
rect 153764 185602 153770 185604
rect 154205 185602 154271 185605
rect 153764 185600 154271 185602
rect 153764 185544 154210 185600
rect 154266 185544 154271 185600
rect 153764 185542 154271 185544
rect 153764 185540 153770 185542
rect 152549 185539 152615 185540
rect 154205 185539 154271 185542
rect 155401 185602 155467 185605
rect 155534 185602 155540 185604
rect 155401 185600 155540 185602
rect 155401 185544 155406 185600
rect 155462 185544 155540 185600
rect 155401 185542 155540 185544
rect 155401 185539 155467 185542
rect 155534 185540 155540 185542
rect 155604 185540 155610 185604
rect 156822 185540 156828 185604
rect 156892 185602 156898 185604
rect 156965 185602 157031 185605
rect 156892 185600 157031 185602
rect 156892 185544 156970 185600
rect 157026 185544 157031 185600
rect 156892 185542 157031 185544
rect 156892 185540 156898 185542
rect 156965 185539 157031 185542
rect 157190 185540 157196 185604
rect 157260 185602 157266 185604
rect 158713 185602 158779 185605
rect 157260 185600 158779 185602
rect 157260 185544 158718 185600
rect 158774 185544 158779 185600
rect 157260 185542 158779 185544
rect 157260 185540 157266 185542
rect 158713 185539 158779 185542
rect 160686 185540 160692 185604
rect 160756 185602 160762 185604
rect 161013 185602 161079 185605
rect 160756 185600 161079 185602
rect 160756 185544 161018 185600
rect 161074 185544 161079 185600
rect 160756 185542 161079 185544
rect 160756 185540 160762 185542
rect 161013 185539 161079 185542
rect 165838 185540 165844 185604
rect 165908 185602 165914 185604
rect 166625 185602 166691 185605
rect 167545 185604 167611 185605
rect 167494 185602 167500 185604
rect 165908 185600 166691 185602
rect 165908 185544 166630 185600
rect 166686 185544 166691 185600
rect 165908 185542 166691 185544
rect 167454 185542 167500 185602
rect 167564 185600 167611 185604
rect 167606 185544 167611 185600
rect 165908 185540 165914 185542
rect 166625 185539 166691 185542
rect 167494 185540 167500 185542
rect 167564 185540 167611 185544
rect 167545 185539 167611 185540
rect 168005 185604 168071 185605
rect 168005 185600 168052 185604
rect 168116 185602 168122 185604
rect 168005 185544 168010 185600
rect 168005 185540 168052 185544
rect 168116 185542 168162 185602
rect 168116 185540 168122 185542
rect 168598 185540 168604 185604
rect 168668 185602 168674 185604
rect 169569 185602 169635 185605
rect 168668 185600 169635 185602
rect 168668 185544 169574 185600
rect 169630 185544 169635 185600
rect 168668 185542 169635 185544
rect 168668 185540 168674 185542
rect 168005 185539 168071 185540
rect 169569 185539 169635 185542
rect 171542 185540 171548 185604
rect 171612 185602 171618 185604
rect 171869 185602 171935 185605
rect 171612 185600 171935 185602
rect 171612 185544 171874 185600
rect 171930 185544 171935 185600
rect 171612 185542 171935 185544
rect 171612 185540 171618 185542
rect 171869 185539 171935 185542
rect 172053 185604 172119 185605
rect 172053 185600 172100 185604
rect 172164 185602 172170 185604
rect 172053 185544 172058 185600
rect 172053 185540 172100 185544
rect 172164 185542 172210 185602
rect 172164 185540 172170 185542
rect 173014 185540 173020 185604
rect 173084 185602 173090 185604
rect 173157 185602 173223 185605
rect 173084 185600 173223 185602
rect 173084 185544 173162 185600
rect 173218 185544 173223 185600
rect 173084 185542 173223 185544
rect 173084 185540 173090 185542
rect 172053 185539 172119 185540
rect 173157 185539 173223 185542
rect 173341 185602 173407 185605
rect 197854 185602 197860 185604
rect 173341 185600 197860 185602
rect 173341 185544 173346 185600
rect 173402 185544 197860 185600
rect 173341 185542 197860 185544
rect 173341 185539 173407 185542
rect 197854 185540 197860 185542
rect 197924 185540 197930 185604
rect 134742 185404 134748 185468
rect 134812 185466 134818 185468
rect 135069 185466 135135 185469
rect 134812 185464 135135 185466
rect 134812 185408 135074 185464
rect 135130 185408 135135 185464
rect 134812 185406 135135 185408
rect 134812 185404 134818 185406
rect 135069 185403 135135 185406
rect 141049 185466 141115 185469
rect 142102 185466 142108 185468
rect 141049 185464 142108 185466
rect 141049 185408 141054 185464
rect 141110 185408 142108 185464
rect 141049 185406 142108 185408
rect 141049 185403 141115 185406
rect 142102 185404 142108 185406
rect 142172 185404 142178 185468
rect 145230 185404 145236 185468
rect 145300 185466 145306 185468
rect 165705 185466 165771 185469
rect 145300 185464 165771 185466
rect 145300 185408 165710 185464
rect 165766 185408 165771 185464
rect 145300 185406 165771 185408
rect 145300 185404 145306 185406
rect 165705 185403 165771 185406
rect 176009 185466 176075 185469
rect 200798 185466 200804 185468
rect 176009 185464 200804 185466
rect 176009 185408 176014 185464
rect 176070 185408 200804 185464
rect 176009 185406 200804 185408
rect 176009 185403 176075 185406
rect 200798 185404 200804 185406
rect 200868 185404 200874 185468
rect 132861 185330 132927 185333
rect 133822 185330 133828 185332
rect 132861 185328 133828 185330
rect 132861 185272 132866 185328
rect 132922 185272 133828 185328
rect 132861 185270 133828 185272
rect 132861 185267 132927 185270
rect 133822 185268 133828 185270
rect 133892 185268 133898 185332
rect 140957 185330 141023 185333
rect 143758 185330 143764 185332
rect 140957 185328 143764 185330
rect 140957 185272 140962 185328
rect 141018 185272 143764 185328
rect 140957 185270 143764 185272
rect 140957 185267 141023 185270
rect 143758 185268 143764 185270
rect 143828 185268 143834 185332
rect 165705 185330 165771 185333
rect 166758 185330 166764 185332
rect 165705 185328 166764 185330
rect 165705 185272 165710 185328
rect 165766 185272 166764 185328
rect 165705 185270 166764 185272
rect 165705 185267 165771 185270
rect 166758 185268 166764 185270
rect 166828 185268 166834 185332
rect 173065 185330 173131 185333
rect 197670 185330 197676 185332
rect 173065 185328 197676 185330
rect 173065 185272 173070 185328
rect 173126 185272 197676 185328
rect 173065 185270 197676 185272
rect 173065 185267 173131 185270
rect 197670 185268 197676 185270
rect 197740 185268 197746 185332
rect 133229 185196 133295 185197
rect 133229 185192 133276 185196
rect 133340 185194 133346 185196
rect 172145 185194 172211 185197
rect 197302 185194 197308 185196
rect 133229 185136 133234 185192
rect 133229 185132 133276 185136
rect 133340 185134 133386 185194
rect 172145 185192 197308 185194
rect 172145 185136 172150 185192
rect 172206 185136 197308 185192
rect 172145 185134 197308 185136
rect 133340 185132 133346 185134
rect 133229 185131 133295 185132
rect 172145 185131 172211 185134
rect 197302 185132 197308 185134
rect 197372 185132 197378 185196
rect 170673 184922 170739 184925
rect 170806 184922 170812 184924
rect 170673 184920 170812 184922
rect 170673 184864 170678 184920
rect 170734 184864 170812 184920
rect 170673 184862 170812 184864
rect 170673 184859 170739 184862
rect 170806 184860 170812 184862
rect 170876 184860 170882 184924
rect 148726 183364 148732 183428
rect 148796 183426 148802 183428
rect 164417 183426 164483 183429
rect 148796 183424 164483 183426
rect 148796 183368 164422 183424
rect 164478 183368 164483 183424
rect 148796 183366 164483 183368
rect 148796 183364 148802 183366
rect 164417 183363 164483 183366
rect 135897 183154 135963 183157
rect 136214 183154 136220 183156
rect 135897 183152 136220 183154
rect 135897 183096 135902 183152
rect 135958 183096 136220 183152
rect 135897 183094 136220 183096
rect 135897 183091 135963 183094
rect 136214 183092 136220 183094
rect 136284 183092 136290 183156
rect 147070 181868 147076 181932
rect 147140 181930 147146 181932
rect 147305 181930 147371 181933
rect 147140 181928 147371 181930
rect 147140 181872 147310 181928
rect 147366 181872 147371 181928
rect 147140 181870 147371 181872
rect 147140 181868 147146 181870
rect 147305 181867 147371 181870
rect 147438 181732 147444 181796
rect 147508 181794 147514 181796
rect 160829 181794 160895 181797
rect 147508 181792 160895 181794
rect 147508 181736 160834 181792
rect 160890 181736 160895 181792
rect 147508 181734 160895 181736
rect 147508 181732 147514 181734
rect 160829 181731 160895 181734
rect 175590 180780 175596 180844
rect 175660 180842 175666 180844
rect 191189 180842 191255 180845
rect 175660 180840 191255 180842
rect 175660 180784 191194 180840
rect 191250 180784 191255 180840
rect 175660 180782 191255 180784
rect 175660 180780 175666 180782
rect 191189 180779 191255 180782
rect 166349 180298 166415 180301
rect 166574 180298 166580 180300
rect 166349 180296 166580 180298
rect 166349 180240 166354 180296
rect 166410 180240 166580 180296
rect 166349 180238 166580 180240
rect 166349 180235 166415 180238
rect 166574 180236 166580 180238
rect 166644 180236 166650 180300
rect 168782 179964 168788 180028
rect 168852 180026 168858 180028
rect 169109 180026 169175 180029
rect 168852 180024 169175 180026
rect 168852 179968 169114 180024
rect 169170 179968 169175 180024
rect 168852 179966 169175 179968
rect 168852 179964 168858 179966
rect 169109 179963 169175 179966
rect 159030 179420 159036 179484
rect 159100 179482 159106 179484
rect 159173 179482 159239 179485
rect 159100 179480 159239 179482
rect 159100 179424 159178 179480
rect 159234 179424 159239 179480
rect 159100 179422 159239 179424
rect 159100 179420 159106 179422
rect 159173 179419 159239 179422
rect 139761 179346 139827 179349
rect 140078 179346 140084 179348
rect 139761 179344 140084 179346
rect 139761 179288 139766 179344
rect 139822 179288 140084 179344
rect 139761 179286 140084 179288
rect 139761 179283 139827 179286
rect 140078 179284 140084 179286
rect 140148 179284 140154 179348
rect 146518 179284 146524 179348
rect 146588 179346 146594 179348
rect 146753 179346 146819 179349
rect 146588 179344 146819 179346
rect 146588 179288 146758 179344
rect 146814 179288 146819 179344
rect 146588 179286 146819 179288
rect 146588 179284 146594 179286
rect 146753 179283 146819 179286
rect 580165 179210 580231 179213
rect 583520 179210 584960 179300
rect 580165 179208 584960 179210
rect 580165 179152 580170 179208
rect 580226 179152 584960 179208
rect 580165 179150 584960 179152
rect 580165 179147 580231 179150
rect 145598 179012 145604 179076
rect 145668 179074 145674 179076
rect 162761 179074 162827 179077
rect 145668 179072 162827 179074
rect 145668 179016 162766 179072
rect 162822 179016 162827 179072
rect 583520 179060 584960 179150
rect 145668 179014 162827 179016
rect 145668 179012 145674 179014
rect 162761 179011 162827 179014
rect 148910 178468 148916 178532
rect 148980 178530 148986 178532
rect 160553 178530 160619 178533
rect 148980 178528 160619 178530
rect 148980 178472 160558 178528
rect 160614 178472 160619 178528
rect 148980 178470 160619 178472
rect 148980 178468 148986 178470
rect 160553 178467 160619 178470
rect 165286 178468 165292 178532
rect 165356 178530 165362 178532
rect 165521 178530 165587 178533
rect 165356 178528 165587 178530
rect 165356 178472 165526 178528
rect 165582 178472 165587 178528
rect 165356 178470 165587 178472
rect 165356 178468 165362 178470
rect 165521 178467 165587 178470
rect 160737 177986 160803 177989
rect 161054 177986 161060 177988
rect 160737 177984 161060 177986
rect 160737 177928 160742 177984
rect 160798 177928 161060 177984
rect 160737 177926 161060 177928
rect 160737 177923 160803 177926
rect 161054 177924 161060 177926
rect 161124 177924 161130 177988
rect 138381 177172 138447 177173
rect 138381 177168 138428 177172
rect 138492 177170 138498 177172
rect 138381 177112 138386 177168
rect 138381 177108 138428 177112
rect 138492 177110 138538 177170
rect 138492 177108 138498 177110
rect 138381 177107 138447 177108
rect 177062 176564 177068 176628
rect 177132 176626 177138 176628
rect 177297 176626 177363 176629
rect 177132 176624 177363 176626
rect 177132 176568 177302 176624
rect 177358 176568 177363 176624
rect 177132 176566 177363 176568
rect 177132 176564 177138 176566
rect 177297 176563 177363 176566
rect -960 175796 480 176036
rect 139025 174996 139091 174997
rect 138974 174994 138980 174996
rect 138934 174934 138980 174994
rect 139044 174992 139091 174996
rect 139086 174936 139091 174992
rect 138974 174932 138980 174934
rect 139044 174932 139091 174936
rect 139025 174931 139091 174932
rect 187233 174586 187299 174589
rect 197486 174586 197492 174588
rect 187233 174584 197492 174586
rect 187233 174528 187238 174584
rect 187294 174528 197492 174584
rect 187233 174526 197492 174528
rect 187233 174523 187299 174526
rect 197486 174524 197492 174526
rect 197556 174524 197562 174588
rect 201493 173500 201559 173501
rect 201493 173496 201540 173500
rect 201604 173498 201610 173500
rect 201493 173440 201498 173496
rect 201493 173436 201540 173440
rect 201604 173438 201650 173498
rect 201604 173436 201610 173438
rect 201493 173435 201559 173436
rect 161289 171186 161355 171189
rect 161422 171186 161428 171188
rect 161289 171184 161428 171186
rect 161289 171128 161294 171184
rect 161350 171128 161428 171184
rect 161289 171126 161428 171128
rect 161289 171123 161355 171126
rect 161422 171124 161428 171126
rect 161492 171124 161498 171188
rect 142061 171052 142127 171053
rect 142061 171050 142108 171052
rect 142016 171048 142108 171050
rect 142172 171050 142178 171052
rect 161289 171050 161355 171053
rect 161422 171050 161428 171052
rect 142016 170992 142066 171048
rect 142016 170990 142108 170992
rect 142061 170988 142108 170990
rect 142172 170990 142254 171050
rect 161289 171048 161428 171050
rect 161289 170992 161294 171048
rect 161350 170992 161428 171048
rect 161289 170990 161428 170992
rect 142172 170988 142178 170990
rect 142061 170987 142127 170988
rect 161289 170987 161355 170990
rect 161422 170988 161428 170990
rect 161492 170988 161498 171052
rect 580165 165882 580231 165885
rect 583520 165882 584960 165972
rect 580165 165880 584960 165882
rect 580165 165824 580170 165880
rect 580226 165824 584960 165880
rect 580165 165822 584960 165824
rect 580165 165819 580231 165822
rect 583520 165732 584960 165822
rect -960 162890 480 162980
rect 3417 162890 3483 162893
rect -960 162888 3483 162890
rect -960 162832 3422 162888
rect 3478 162832 3483 162888
rect -960 162830 3483 162832
rect -960 162740 480 162830
rect 3417 162827 3483 162830
rect 142102 161604 142108 161668
rect 142172 161604 142178 161668
rect 142110 161533 142170 161604
rect 142061 161530 142170 161533
rect 142016 161528 142170 161530
rect 142016 161472 142066 161528
rect 142122 161472 142170 161528
rect 142016 161470 142170 161472
rect 161289 161530 161355 161533
rect 161422 161530 161428 161532
rect 161289 161528 161428 161530
rect 161289 161472 161294 161528
rect 161350 161472 161428 161528
rect 161289 161470 161428 161472
rect 142061 161467 142127 161470
rect 161289 161467 161355 161470
rect 161422 161468 161428 161470
rect 161492 161468 161498 161532
rect 142061 161396 142127 161397
rect 142061 161394 142108 161396
rect 142016 161392 142108 161394
rect 142172 161394 142178 161396
rect 161289 161394 161355 161397
rect 161422 161394 161428 161396
rect 142016 161336 142066 161392
rect 142016 161334 142108 161336
rect 142061 161332 142108 161334
rect 142172 161334 142254 161394
rect 161289 161392 161428 161394
rect 161289 161336 161294 161392
rect 161350 161336 161428 161392
rect 161289 161334 161428 161336
rect 142172 161332 142178 161334
rect 142061 161331 142127 161332
rect 161289 161331 161355 161334
rect 161422 161332 161428 161334
rect 161492 161332 161498 161396
rect 157517 152690 157583 152693
rect 185342 152690 185348 152692
rect 157517 152688 185348 152690
rect 157517 152632 157522 152688
rect 157578 152632 185348 152688
rect 157517 152630 185348 152632
rect 157517 152627 157583 152630
rect 185342 152628 185348 152630
rect 185412 152628 185418 152692
rect 580257 152690 580323 152693
rect 583520 152690 584960 152780
rect 580257 152688 584960 152690
rect 580257 152632 580262 152688
rect 580318 152632 584960 152688
rect 580257 152630 584960 152632
rect 580257 152627 580323 152630
rect 156137 152554 156203 152557
rect 185158 152554 185164 152556
rect 156137 152552 185164 152554
rect 156137 152496 156142 152552
rect 156198 152496 185164 152552
rect 156137 152494 185164 152496
rect 156137 152491 156203 152494
rect 185158 152492 185164 152494
rect 185228 152492 185234 152556
rect 583520 152540 584960 152630
rect 145230 152356 145236 152420
rect 145300 152418 145306 152420
rect 200481 152418 200547 152421
rect 145300 152416 200547 152418
rect 145300 152360 200486 152416
rect 200542 152360 200547 152416
rect 145300 152358 200547 152360
rect 145300 152356 145306 152358
rect 200481 152355 200547 152358
rect 142102 151948 142108 152012
rect 142172 151948 142178 152012
rect 142110 151877 142170 151948
rect 142061 151874 142170 151877
rect 142016 151872 142170 151874
rect 142016 151816 142066 151872
rect 142122 151816 142170 151872
rect 142016 151814 142170 151816
rect 161289 151874 161355 151877
rect 161422 151874 161428 151876
rect 161289 151872 161428 151874
rect 161289 151816 161294 151872
rect 161350 151816 161428 151872
rect 161289 151814 161428 151816
rect 142061 151811 142127 151814
rect 161289 151811 161355 151814
rect 161422 151812 161428 151814
rect 161492 151812 161498 151876
rect 142061 151740 142127 151741
rect 142061 151738 142108 151740
rect 142016 151736 142108 151738
rect 142172 151738 142178 151740
rect 161289 151738 161355 151741
rect 161422 151738 161428 151740
rect 142016 151680 142066 151736
rect 142016 151678 142108 151680
rect 142061 151676 142108 151678
rect 142172 151678 142254 151738
rect 161289 151736 161428 151738
rect 161289 151680 161294 151736
rect 161350 151680 161428 151736
rect 161289 151678 161428 151680
rect 142172 151676 142178 151678
rect 142061 151675 142127 151676
rect 161289 151675 161355 151678
rect 161422 151676 161428 151678
rect 161492 151676 161498 151740
rect 156045 150378 156111 150381
rect 181110 150378 181116 150380
rect 156045 150376 181116 150378
rect 156045 150320 156050 150376
rect 156106 150320 181116 150376
rect 156045 150318 181116 150320
rect 156045 150315 156111 150318
rect 181110 150316 181116 150318
rect 181180 150316 181186 150380
rect 156229 150242 156295 150245
rect 183870 150242 183876 150244
rect 156229 150240 183876 150242
rect 156229 150184 156234 150240
rect 156290 150184 183876 150240
rect 156229 150182 183876 150184
rect 156229 150179 156295 150182
rect 183870 150180 183876 150182
rect 183940 150180 183946 150244
rect 174169 150106 174235 150109
rect 203006 150106 203012 150108
rect 174169 150104 203012 150106
rect 174169 150048 174174 150104
rect 174230 150048 203012 150104
rect 174169 150046 203012 150048
rect 174169 150043 174235 150046
rect 203006 150044 203012 150046
rect 203076 150044 203082 150108
rect 174353 149970 174419 149973
rect 203190 149970 203196 149972
rect 174353 149968 203196 149970
rect -960 149834 480 149924
rect 174353 149912 174358 149968
rect 174414 149912 203196 149968
rect 174353 149910 203196 149912
rect 174353 149907 174419 149910
rect 203190 149908 203196 149910
rect 203260 149908 203266 149972
rect 3417 149834 3483 149837
rect -960 149832 3483 149834
rect -960 149776 3422 149832
rect 3478 149776 3483 149832
rect -960 149774 3483 149776
rect -960 149684 480 149774
rect 3417 149771 3483 149774
rect 153377 149834 153443 149837
rect 182766 149834 182772 149836
rect 153377 149832 182772 149834
rect 153377 149776 153382 149832
rect 153438 149776 182772 149832
rect 153377 149774 182772 149776
rect 153377 149771 153443 149774
rect 182766 149772 182772 149774
rect 182836 149772 182842 149836
rect 154849 149698 154915 149701
rect 187366 149698 187372 149700
rect 154849 149696 187372 149698
rect 154849 149640 154854 149696
rect 154910 149640 187372 149696
rect 154849 149638 187372 149640
rect 154849 149635 154915 149638
rect 187366 149636 187372 149638
rect 187436 149636 187442 149700
rect 186957 149156 187023 149157
rect 186957 149154 187004 149156
rect 186912 149152 187004 149154
rect 186912 149096 186962 149152
rect 186912 149094 187004 149096
rect 186957 149092 187004 149094
rect 187068 149092 187074 149156
rect 186957 149091 187023 149092
rect 123661 148474 123727 148477
rect 143758 148474 143764 148476
rect 123661 148472 143764 148474
rect 123661 148416 123666 148472
rect 123722 148416 143764 148472
rect 123661 148414 143764 148416
rect 123661 148411 123727 148414
rect 143758 148412 143764 148414
rect 143828 148412 143834 148476
rect 165705 148474 165771 148477
rect 191598 148474 191604 148476
rect 165705 148472 191604 148474
rect 165705 148416 165710 148472
rect 165766 148416 191604 148472
rect 165705 148414 191604 148416
rect 165705 148411 165771 148414
rect 191598 148412 191604 148414
rect 191668 148412 191674 148476
rect 100477 148338 100543 148341
rect 132585 148338 132651 148341
rect 100477 148336 132651 148338
rect 100477 148280 100482 148336
rect 100538 148280 132590 148336
rect 132646 148280 132651 148336
rect 100477 148278 132651 148280
rect 100477 148275 100543 148278
rect 132585 148275 132651 148278
rect 163129 148338 163195 148341
rect 188286 148338 188292 148340
rect 163129 148336 188292 148338
rect 163129 148280 163134 148336
rect 163190 148280 188292 148336
rect 163129 148278 188292 148280
rect 163129 148275 163195 148278
rect 188286 148276 188292 148278
rect 188356 148276 188362 148340
rect 196566 147732 196572 147796
rect 196636 147794 196642 147796
rect 196801 147794 196867 147797
rect 196636 147792 196867 147794
rect 196636 147736 196806 147792
rect 196862 147736 196867 147792
rect 196636 147734 196867 147736
rect 196636 147732 196642 147734
rect 196801 147731 196867 147734
rect 198733 147794 198799 147797
rect 199326 147794 199332 147796
rect 198733 147792 199332 147794
rect 198733 147736 198738 147792
rect 198794 147736 199332 147792
rect 198733 147734 199332 147736
rect 198733 147731 198799 147734
rect 199326 147732 199332 147734
rect 199396 147732 199402 147796
rect 137001 147658 137067 147661
rect 142470 147658 142476 147660
rect 137001 147656 142476 147658
rect 137001 147600 137006 147656
rect 137062 147600 142476 147656
rect 137001 147598 142476 147600
rect 137001 147595 137067 147598
rect 142470 147596 142476 147598
rect 142540 147596 142546 147660
rect 180333 147658 180399 147661
rect 193622 147658 193628 147660
rect 180333 147656 193628 147658
rect 180333 147600 180338 147656
rect 180394 147600 193628 147656
rect 180333 147598 193628 147600
rect 180333 147595 180399 147598
rect 193622 147596 193628 147598
rect 193692 147596 193698 147660
rect 169845 147522 169911 147525
rect 189390 147522 189396 147524
rect 169845 147520 189396 147522
rect 169845 147464 169850 147520
rect 169906 147464 189396 147520
rect 169845 147462 189396 147464
rect 169845 147459 169911 147462
rect 189390 147460 189396 147462
rect 189460 147460 189466 147524
rect 171133 147386 171199 147389
rect 192150 147386 192156 147388
rect 171133 147384 192156 147386
rect 171133 147328 171138 147384
rect 171194 147328 192156 147384
rect 171133 147326 192156 147328
rect 171133 147323 171199 147326
rect 192150 147324 192156 147326
rect 192220 147324 192226 147388
rect 173985 147250 174051 147253
rect 198958 147250 198964 147252
rect 173985 147248 198964 147250
rect 173985 147192 173990 147248
rect 174046 147192 198964 147248
rect 173985 147190 198964 147192
rect 173985 147187 174051 147190
rect 198958 147188 198964 147190
rect 199028 147188 199034 147252
rect 157241 147114 157307 147117
rect 183134 147114 183140 147116
rect 157241 147112 183140 147114
rect 157241 147056 157246 147112
rect 157302 147056 183140 147112
rect 157241 147054 183140 147056
rect 157241 147051 157307 147054
rect 183134 147052 183140 147054
rect 183204 147052 183210 147116
rect 116209 146978 116275 146981
rect 142286 146978 142292 146980
rect 116209 146976 142292 146978
rect 116209 146920 116214 146976
rect 116270 146920 142292 146976
rect 116209 146918 142292 146920
rect 116209 146915 116275 146918
rect 142286 146916 142292 146918
rect 142356 146916 142362 146980
rect 151997 146978 152063 146981
rect 181294 146978 181300 146980
rect 151997 146976 181300 146978
rect 151997 146920 152002 146976
rect 152058 146920 181300 146976
rect 151997 146918 181300 146920
rect 151997 146915 152063 146918
rect 181294 146916 181300 146918
rect 181364 146916 181370 146980
rect 173893 146162 173959 146165
rect 191281 146162 191347 146165
rect 173893 146160 191347 146162
rect 173893 146104 173898 146160
rect 173954 146104 191286 146160
rect 191342 146104 191347 146160
rect 173893 146102 191347 146104
rect 173893 146099 173959 146102
rect 191281 146099 191347 146102
rect 164233 146026 164299 146029
rect 195145 146026 195211 146029
rect 164233 146024 195211 146026
rect 164233 145968 164238 146024
rect 164294 145968 195150 146024
rect 195206 145968 195211 146024
rect 164233 145966 195211 145968
rect 164233 145963 164299 145966
rect 195145 145963 195211 145966
rect 112846 145828 112852 145892
rect 112916 145890 112922 145892
rect 126973 145890 127039 145893
rect 112916 145888 127039 145890
rect 112916 145832 126978 145888
rect 127034 145832 127039 145888
rect 112916 145830 127039 145832
rect 112916 145828 112922 145830
rect 126973 145827 127039 145830
rect 162945 145890 163011 145893
rect 194726 145890 194732 145892
rect 162945 145888 194732 145890
rect 162945 145832 162950 145888
rect 163006 145832 194732 145888
rect 162945 145830 194732 145832
rect 162945 145827 163011 145830
rect 194726 145828 194732 145830
rect 194796 145828 194802 145892
rect 111190 145692 111196 145756
rect 111260 145754 111266 145756
rect 131849 145754 131915 145757
rect 111260 145752 131915 145754
rect 111260 145696 131854 145752
rect 131910 145696 131915 145752
rect 111260 145694 131915 145696
rect 111260 145692 111266 145694
rect 131849 145691 131915 145694
rect 158805 145754 158871 145757
rect 191465 145754 191531 145757
rect 158805 145752 191531 145754
rect 158805 145696 158810 145752
rect 158866 145696 191470 145752
rect 191526 145696 191531 145752
rect 158805 145694 191531 145696
rect 158805 145691 158871 145694
rect 191465 145691 191531 145694
rect 120574 145556 120580 145620
rect 120644 145618 120650 145620
rect 153285 145618 153351 145621
rect 120644 145616 153351 145618
rect 120644 145560 153290 145616
rect 153346 145560 153351 145616
rect 120644 145558 153351 145560
rect 120644 145556 120650 145558
rect 153285 145555 153351 145558
rect 160921 145618 160987 145621
rect 193213 145618 193279 145621
rect 160921 145616 193279 145618
rect 160921 145560 160926 145616
rect 160982 145560 193218 145616
rect 193274 145560 193279 145616
rect 160921 145558 193279 145560
rect 160921 145555 160987 145558
rect 193213 145555 193279 145558
rect 119654 144876 119660 144940
rect 119724 144938 119730 144940
rect 182449 144938 182515 144941
rect 183461 144938 183527 144941
rect 119724 144936 183527 144938
rect 119724 144880 182454 144936
rect 182510 144880 183466 144936
rect 183522 144880 183527 144936
rect 119724 144878 183527 144880
rect 119724 144876 119730 144878
rect 182449 144875 182515 144878
rect 183461 144875 183527 144878
rect 115606 144740 115612 144804
rect 115676 144802 115682 144804
rect 142797 144802 142863 144805
rect 115676 144800 142863 144802
rect 115676 144744 142802 144800
rect 142858 144744 142863 144800
rect 115676 144742 142863 144744
rect 115676 144740 115682 144742
rect 142797 144739 142863 144742
rect 182950 144740 182956 144804
rect 183020 144802 183026 144804
rect 191557 144802 191623 144805
rect 183020 144800 191623 144802
rect 183020 144744 191562 144800
rect 191618 144744 191623 144800
rect 183020 144742 191623 144744
rect 183020 144740 183026 144742
rect 191557 144739 191623 144742
rect 116894 144604 116900 144668
rect 116964 144666 116970 144668
rect 144453 144666 144519 144669
rect 116964 144664 144519 144666
rect 116964 144608 144458 144664
rect 144514 144608 144519 144664
rect 116964 144606 144519 144608
rect 116964 144604 116970 144606
rect 144453 144603 144519 144606
rect 167729 144666 167795 144669
rect 191966 144666 191972 144668
rect 167729 144664 191972 144666
rect 167729 144608 167734 144664
rect 167790 144608 191972 144664
rect 167729 144606 191972 144608
rect 167729 144603 167795 144606
rect 191966 144604 191972 144606
rect 192036 144604 192042 144668
rect 114134 144468 114140 144532
rect 114204 144530 114210 144532
rect 141141 144530 141207 144533
rect 114204 144528 141207 144530
rect 114204 144472 141146 144528
rect 141202 144472 141207 144528
rect 114204 144470 141207 144472
rect 114204 144468 114210 144470
rect 141141 144467 141207 144470
rect 164141 144530 164207 144533
rect 191782 144530 191788 144532
rect 164141 144528 191788 144530
rect 164141 144472 164146 144528
rect 164202 144472 191788 144528
rect 164141 144470 191788 144472
rect 164141 144467 164207 144470
rect 191782 144468 191788 144470
rect 191852 144468 191858 144532
rect 117078 144332 117084 144396
rect 117148 144394 117154 144396
rect 145557 144394 145623 144397
rect 117148 144392 145623 144394
rect 117148 144336 145562 144392
rect 145618 144336 145623 144392
rect 117148 144334 145623 144336
rect 117148 144332 117154 144334
rect 145557 144331 145623 144334
rect 166625 144394 166691 144397
rect 194542 144394 194548 144396
rect 166625 144392 194548 144394
rect 166625 144336 166630 144392
rect 166686 144336 194548 144392
rect 166625 144334 194548 144336
rect 166625 144331 166691 144334
rect 194542 144332 194548 144334
rect 194612 144332 194618 144396
rect 118182 144196 118188 144260
rect 118252 144258 118258 144260
rect 147213 144258 147279 144261
rect 118252 144256 147279 144258
rect 118252 144200 147218 144256
rect 147274 144200 147279 144256
rect 118252 144198 147279 144200
rect 118252 144196 118258 144198
rect 147213 144195 147279 144198
rect 162761 144258 162827 144261
rect 190494 144258 190500 144260
rect 162761 144256 190500 144258
rect 162761 144200 162766 144256
rect 162822 144200 190500 144256
rect 162761 144198 190500 144200
rect 162761 144195 162827 144198
rect 190494 144196 190500 144198
rect 190564 144196 190570 144260
rect 115790 144060 115796 144124
rect 115860 144122 115866 144124
rect 147765 144122 147831 144125
rect 115860 144120 147831 144122
rect 115860 144064 147770 144120
rect 147826 144064 147831 144120
rect 115860 144062 147831 144064
rect 115860 144060 115866 144062
rect 147765 144059 147831 144062
rect 157701 144122 157767 144125
rect 188102 144122 188108 144124
rect 157701 144120 188108 144122
rect 157701 144064 157706 144120
rect 157762 144064 188108 144120
rect 157701 144062 188108 144064
rect 157701 144059 157767 144062
rect 188102 144060 188108 144062
rect 188172 144060 188178 144124
rect 113582 143924 113588 143988
rect 113652 143986 113658 143988
rect 138933 143986 138999 143989
rect 113652 143984 138999 143986
rect 113652 143928 138938 143984
rect 138994 143928 138999 143984
rect 113652 143926 138999 143928
rect 113652 143924 113658 143926
rect 138933 143923 138999 143926
rect 185577 143578 185643 143581
rect 190494 143578 190500 143580
rect 185577 143576 190500 143578
rect 185577 143520 185582 143576
rect 185638 143520 190500 143576
rect 185577 143518 190500 143520
rect 185577 143515 185643 143518
rect 190494 143516 190500 143518
rect 190564 143516 190570 143580
rect 111374 143380 111380 143444
rect 111444 143442 111450 143444
rect 125593 143442 125659 143445
rect 111444 143440 125659 143442
rect 111444 143384 125598 143440
rect 125654 143384 125659 143440
rect 111444 143382 125659 143384
rect 111444 143380 111450 143382
rect 125593 143379 125659 143382
rect 163865 143442 163931 143445
rect 186865 143442 186931 143445
rect 163865 143440 186931 143442
rect 163865 143384 163870 143440
rect 163926 143384 186870 143440
rect 186926 143384 186931 143440
rect 163865 143382 186931 143384
rect 163865 143379 163931 143382
rect 186865 143379 186931 143382
rect 111558 143244 111564 143308
rect 111628 143306 111634 143308
rect 132861 143306 132927 143309
rect 111628 143304 132927 143306
rect 111628 143248 132866 143304
rect 132922 143248 132927 143304
rect 111628 143246 132927 143248
rect 111628 143244 111634 143246
rect 132861 143243 132927 143246
rect 162209 143306 162275 143309
rect 188153 143306 188219 143309
rect 162209 143304 188219 143306
rect 162209 143248 162214 143304
rect 162270 143248 188158 143304
rect 188214 143248 188219 143304
rect 162209 143246 188219 143248
rect 162209 143243 162275 143246
rect 188153 143243 188219 143246
rect 121126 143108 121132 143172
rect 121196 143170 121202 143172
rect 146661 143170 146727 143173
rect 121196 143168 146727 143170
rect 121196 143112 146666 143168
rect 146722 143112 146727 143168
rect 121196 143110 146727 143112
rect 121196 143108 121202 143110
rect 146661 143107 146727 143110
rect 157241 143170 157307 143173
rect 187693 143170 187759 143173
rect 157241 143168 187759 143170
rect 157241 143112 157246 143168
rect 157302 143112 187698 143168
rect 187754 143112 187759 143168
rect 157241 143110 187759 143112
rect 157241 143107 157307 143110
rect 187693 143107 187759 143110
rect 119153 143034 119219 143037
rect 145097 143034 145163 143037
rect 119153 143032 145163 143034
rect 119153 142976 119158 143032
rect 119214 142976 145102 143032
rect 145158 142976 145163 143032
rect 119153 142974 145163 142976
rect 119153 142971 119219 142974
rect 145097 142971 145163 142974
rect 155401 143034 155467 143037
rect 187785 143034 187851 143037
rect 155401 143032 187851 143034
rect 155401 142976 155406 143032
rect 155462 142976 187790 143032
rect 187846 142976 187851 143032
rect 155401 142974 187851 142976
rect 155401 142971 155467 142974
rect 187785 142971 187851 142974
rect 120901 142898 120967 142901
rect 149973 142898 150039 142901
rect 120901 142896 150039 142898
rect 120901 142840 120906 142896
rect 120962 142840 149978 142896
rect 150034 142840 150039 142896
rect 120901 142838 150039 142840
rect 120901 142835 120967 142838
rect 149973 142835 150039 142838
rect 153837 142898 153903 142901
rect 186497 142898 186563 142901
rect 153837 142896 186563 142898
rect 153837 142840 153842 142896
rect 153898 142840 186502 142896
rect 186558 142840 186563 142896
rect 153837 142838 186563 142840
rect 153837 142835 153903 142838
rect 186497 142835 186563 142838
rect 119337 142762 119403 142765
rect 148317 142762 148383 142765
rect 119337 142760 148383 142762
rect 119337 142704 119342 142760
rect 119398 142704 148322 142760
rect 148378 142704 148383 142760
rect 119337 142702 148383 142704
rect 119337 142699 119403 142702
rect 148317 142699 148383 142702
rect 152273 142762 152339 142765
rect 186957 142762 187023 142765
rect 152273 142760 187023 142762
rect 152273 142704 152278 142760
rect 152334 142704 186962 142760
rect 187018 142704 187023 142760
rect 152273 142702 187023 142704
rect 152273 142699 152339 142702
rect 186957 142699 187023 142702
rect 113950 142564 113956 142628
rect 114020 142626 114026 142628
rect 125685 142626 125751 142629
rect 114020 142624 125751 142626
rect 114020 142568 125690 142624
rect 125746 142568 125751 142624
rect 114020 142566 125751 142568
rect 114020 142564 114026 142566
rect 125685 142563 125751 142566
rect 142061 142354 142127 142357
rect 142286 142354 142292 142356
rect 142016 142352 142292 142354
rect 142016 142296 142066 142352
rect 142122 142296 142292 142352
rect 142016 142294 142292 142296
rect 142061 142291 142127 142294
rect 142286 142292 142292 142294
rect 142356 142292 142362 142356
rect 161289 142354 161355 142357
rect 161606 142354 161612 142356
rect 161289 142352 161612 142354
rect 161289 142296 161294 142352
rect 161350 142296 161612 142352
rect 161289 142294 161612 142296
rect 161289 142291 161355 142294
rect 161606 142292 161612 142294
rect 161676 142292 161682 142356
rect 126973 142218 127039 142221
rect 128169 142218 128235 142221
rect 189022 142218 189028 142220
rect 126973 142216 189028 142218
rect 126973 142160 126978 142216
rect 127034 142160 128174 142216
rect 128230 142160 189028 142216
rect 126973 142158 189028 142160
rect 126973 142155 127039 142158
rect 128169 142155 128235 142158
rect 189022 142156 189028 142158
rect 189092 142156 189098 142220
rect 157333 142082 157399 142085
rect 188838 142082 188844 142084
rect 157333 142080 188844 142082
rect 157333 142024 157338 142080
rect 157394 142024 188844 142080
rect 157333 142022 188844 142024
rect 157333 142019 157399 142022
rect 188838 142020 188844 142022
rect 188908 142020 188914 142084
rect 130653 141946 130719 141949
rect 142654 141946 142660 141948
rect 130653 141944 142660 141946
rect 130653 141888 130658 141944
rect 130714 141888 142660 141944
rect 130653 141886 142660 141888
rect 130653 141883 130719 141886
rect 142654 141884 142660 141886
rect 142724 141884 142730 141948
rect 118366 141748 118372 141812
rect 118436 141810 118442 141812
rect 143901 141810 143967 141813
rect 118436 141808 143967 141810
rect 118436 141752 143906 141808
rect 143962 141752 143967 141808
rect 118436 141750 143967 141752
rect 118436 141748 118442 141750
rect 143901 141747 143967 141750
rect 117078 141612 117084 141676
rect 117148 141674 117154 141676
rect 130653 141674 130719 141677
rect 141417 141676 141483 141677
rect 141366 141674 141372 141676
rect 117148 141672 130719 141674
rect 117148 141616 130658 141672
rect 130714 141616 130719 141672
rect 117148 141614 130719 141616
rect 141326 141614 141372 141674
rect 141436 141672 141483 141676
rect 141478 141616 141483 141672
rect 117148 141612 117154 141614
rect 130653 141611 130719 141614
rect 141366 141612 141372 141614
rect 141436 141612 141483 141616
rect 141417 141611 141483 141612
rect 176745 141674 176811 141677
rect 177614 141674 177620 141676
rect 176745 141672 177620 141674
rect 176745 141616 176750 141672
rect 176806 141616 177620 141672
rect 176745 141614 177620 141616
rect 176745 141611 176811 141614
rect 177614 141612 177620 141614
rect 177684 141612 177690 141676
rect 120942 141476 120948 141540
rect 121012 141538 121018 141540
rect 149053 141538 149119 141541
rect 121012 141536 149119 141538
rect 121012 141480 149058 141536
rect 149114 141480 149119 141536
rect 121012 141478 149119 141480
rect 121012 141476 121018 141478
rect 149053 141475 149119 141478
rect 166073 141538 166139 141541
rect 193438 141538 193444 141540
rect 166073 141536 193444 141538
rect 166073 141480 166078 141536
rect 166134 141480 193444 141536
rect 166073 141478 193444 141480
rect 166073 141475 166139 141478
rect 193438 141476 193444 141478
rect 193508 141476 193514 141540
rect 118550 141340 118556 141404
rect 118620 141402 118626 141404
rect 150525 141402 150591 141405
rect 118620 141400 150591 141402
rect 118620 141344 150530 141400
rect 150586 141344 150591 141400
rect 118620 141342 150591 141344
rect 118620 141340 118626 141342
rect 150525 141339 150591 141342
rect 152825 141402 152891 141405
rect 186405 141402 186471 141405
rect 152825 141400 186471 141402
rect 152825 141344 152830 141400
rect 152886 141344 186410 141400
rect 186466 141344 186471 141400
rect 152825 141342 186471 141344
rect 152825 141339 152891 141342
rect 186405 141339 186471 141342
rect 141509 141268 141575 141269
rect 141509 141266 141556 141268
rect 141464 141264 141556 141266
rect 141464 141208 141514 141264
rect 141464 141206 141556 141208
rect 141509 141204 141556 141206
rect 141620 141204 141626 141268
rect 176653 141266 176719 141269
rect 177246 141266 177252 141268
rect 176653 141264 177252 141266
rect 176653 141208 176658 141264
rect 176714 141208 177252 141264
rect 176653 141206 177252 141208
rect 141509 141203 141575 141204
rect 176653 141203 176719 141206
rect 177246 141204 177252 141206
rect 177316 141204 177322 141268
rect 189574 141266 189580 141268
rect 180750 141206 189580 141266
rect 124213 141130 124279 141133
rect 180750 141130 180810 141206
rect 189574 141204 189580 141206
rect 189644 141204 189650 141268
rect 192334 141266 192340 141268
rect 190410 141206 192340 141266
rect 124213 141128 180810 141130
rect 124213 141072 124218 141128
rect 124274 141072 180810 141128
rect 124213 141070 180810 141072
rect 184473 141130 184539 141133
rect 188102 141130 188108 141132
rect 184473 141128 188108 141130
rect 184473 141072 184478 141128
rect 184534 141072 188108 141128
rect 184473 141070 188108 141072
rect 124213 141067 124279 141070
rect 184473 141067 184539 141070
rect 188102 141068 188108 141070
rect 188172 141068 188178 141132
rect 125133 140994 125199 140997
rect 190410 140994 190470 141206
rect 192334 141204 192340 141206
rect 192404 141204 192410 141268
rect 125133 140992 190470 140994
rect 125133 140936 125138 140992
rect 125194 140936 190470 140992
rect 125133 140934 190470 140936
rect 125133 140931 125199 140934
rect 116526 140796 116532 140860
rect 116596 140858 116602 140860
rect 184289 140858 184355 140861
rect 116596 140856 184355 140858
rect 116596 140800 184294 140856
rect 184350 140800 184355 140856
rect 116596 140798 184355 140800
rect 116596 140796 116602 140798
rect 184289 140795 184355 140798
rect 186313 140858 186379 140861
rect 186814 140858 186820 140860
rect 186313 140856 186820 140858
rect 186313 140800 186318 140856
rect 186374 140800 186820 140856
rect 186313 140798 186820 140800
rect 186313 140795 186379 140798
rect 186814 140796 186820 140798
rect 186884 140796 186890 140860
rect 190862 140796 190868 140860
rect 190932 140858 190938 140860
rect 191281 140858 191347 140861
rect 190932 140856 191347 140858
rect 190932 140800 191286 140856
rect 191342 140800 191347 140856
rect 190932 140798 191347 140800
rect 190932 140796 190938 140798
rect 191281 140795 191347 140798
rect 120758 140660 120764 140724
rect 120828 140722 120834 140724
rect 123477 140722 123543 140725
rect 120828 140720 123543 140722
rect 120828 140664 123482 140720
rect 123538 140664 123543 140720
rect 120828 140662 123543 140664
rect 120828 140660 120834 140662
rect 123477 140659 123543 140662
rect 178585 140722 178651 140725
rect 193254 140722 193260 140724
rect 178585 140720 193260 140722
rect 178585 140664 178590 140720
rect 178646 140664 193260 140720
rect 178585 140662 193260 140664
rect 178585 140659 178651 140662
rect 193254 140660 193260 140662
rect 193324 140660 193330 140724
rect 193438 140660 193444 140724
rect 193508 140722 193514 140724
rect 193673 140722 193739 140725
rect 193508 140720 193739 140722
rect 193508 140664 193678 140720
rect 193734 140664 193739 140720
rect 193508 140662 193739 140664
rect 193508 140660 193514 140662
rect 193673 140659 193739 140662
rect 117814 140524 117820 140588
rect 117884 140586 117890 140588
rect 184933 140586 184999 140589
rect 193213 140588 193279 140589
rect 193213 140586 193260 140588
rect 117884 140584 184999 140586
rect 117884 140528 184938 140584
rect 184994 140528 184999 140584
rect 117884 140526 184999 140528
rect 193168 140584 193260 140586
rect 193168 140528 193218 140584
rect 193168 140526 193260 140528
rect 117884 140524 117890 140526
rect 184933 140523 184999 140526
rect 193213 140524 193260 140526
rect 193324 140524 193330 140588
rect 193213 140523 193279 140524
rect 108246 140388 108252 140452
rect 108316 140450 108322 140452
rect 185025 140450 185091 140453
rect 185945 140450 186011 140453
rect 108316 140448 186011 140450
rect 108316 140392 185030 140448
rect 185086 140392 185950 140448
rect 186006 140392 186011 140448
rect 108316 140390 186011 140392
rect 108316 140388 108322 140390
rect 185025 140387 185091 140390
rect 185945 140387 186011 140390
rect 117865 140314 117931 140317
rect 127750 140314 127756 140316
rect 117865 140312 127756 140314
rect 117865 140256 117870 140312
rect 117926 140256 127756 140312
rect 117865 140254 127756 140256
rect 117865 140251 117931 140254
rect 127750 140252 127756 140254
rect 127820 140252 127826 140316
rect 154757 140314 154823 140317
rect 174813 140314 174879 140317
rect 180793 140314 180859 140317
rect 181437 140314 181503 140317
rect 154757 140312 174738 140314
rect 154757 140256 154762 140312
rect 154818 140256 174738 140312
rect 154757 140254 174738 140256
rect 154757 140251 154823 140254
rect 150341 140178 150407 140181
rect 153929 140178 153995 140181
rect 173934 140178 173940 140180
rect 150341 140176 151830 140178
rect 150341 140120 150346 140176
rect 150402 140120 151830 140176
rect 150341 140118 151830 140120
rect 150341 140115 150407 140118
rect 113030 139980 113036 140044
rect 113100 140042 113106 140044
rect 139485 140042 139551 140045
rect 113100 140040 139551 140042
rect 113100 139984 139490 140040
rect 139546 139984 139551 140040
rect 113100 139982 139551 139984
rect 151770 140042 151830 140118
rect 153929 140176 173940 140178
rect 153929 140120 153934 140176
rect 153990 140120 173940 140176
rect 153929 140118 173940 140120
rect 153929 140115 153995 140118
rect 173934 140116 173940 140118
rect 174004 140116 174010 140180
rect 174678 140178 174738 140254
rect 174813 140312 181503 140314
rect 174813 140256 174818 140312
rect 174874 140256 180798 140312
rect 180854 140256 181442 140312
rect 181498 140256 181503 140312
rect 174813 140254 181503 140256
rect 174813 140251 174879 140254
rect 180793 140251 180859 140254
rect 181437 140251 181503 140254
rect 185025 140314 185091 140317
rect 186078 140314 186084 140316
rect 185025 140312 186084 140314
rect 185025 140256 185030 140312
rect 185086 140256 186084 140312
rect 185025 140254 186084 140256
rect 185025 140251 185091 140254
rect 186078 140252 186084 140254
rect 186148 140252 186154 140316
rect 178718 140178 178724 140180
rect 174678 140118 178724 140178
rect 178718 140116 178724 140118
rect 178788 140116 178794 140180
rect 182081 140178 182147 140181
rect 576117 140178 576183 140181
rect 182081 140176 576183 140178
rect 182081 140120 182086 140176
rect 182142 140120 576122 140176
rect 576178 140120 576183 140176
rect 182081 140118 576183 140120
rect 182081 140115 182147 140118
rect 576117 140115 576183 140118
rect 179822 140042 179828 140044
rect 151770 139982 179828 140042
rect 113100 139980 113106 139982
rect 139485 139979 139551 139982
rect 179822 139980 179828 139982
rect 179892 139980 179898 140044
rect 183185 140042 183251 140045
rect 184749 140044 184815 140045
rect 183318 140042 183324 140044
rect 183185 140040 183324 140042
rect 183185 139984 183190 140040
rect 183246 139984 183324 140040
rect 183185 139982 183324 139984
rect 183185 139979 183251 139982
rect 183318 139980 183324 139982
rect 183388 139980 183394 140044
rect 184749 140042 184796 140044
rect 184704 140040 184796 140042
rect 184704 139984 184754 140040
rect 184704 139982 184796 139984
rect 184749 139980 184796 139982
rect 184860 139980 184866 140044
rect 184749 139979 184815 139980
rect 119286 139844 119292 139908
rect 119356 139906 119362 139908
rect 182173 139906 182239 139909
rect 119356 139904 182239 139906
rect 119356 139848 182178 139904
rect 182234 139848 182239 139904
rect 119356 139846 182239 139848
rect 119356 139844 119362 139846
rect 182173 139843 182239 139846
rect 185301 139906 185367 139909
rect 186078 139906 186084 139908
rect 185301 139904 186084 139906
rect 185301 139848 185306 139904
rect 185362 139848 186084 139904
rect 185301 139846 186084 139848
rect 185301 139843 185367 139846
rect 186078 139844 186084 139846
rect 186148 139844 186154 139908
rect 173934 139708 173940 139772
rect 174004 139770 174010 139772
rect 180006 139770 180012 139772
rect 174004 139710 180012 139770
rect 174004 139708 174010 139710
rect 180006 139708 180012 139710
rect 180076 139708 180082 139772
rect 180425 139770 180491 139773
rect 286317 139770 286383 139773
rect 180425 139768 286383 139770
rect 180425 139712 180430 139768
rect 180486 139712 286322 139768
rect 286378 139712 286383 139768
rect 180425 139710 286383 139712
rect 180425 139707 180491 139710
rect 286317 139707 286383 139710
rect 179873 139634 179939 139637
rect 327717 139634 327783 139637
rect 179873 139632 327783 139634
rect 179873 139576 179878 139632
rect 179934 139576 327722 139632
rect 327778 139576 327783 139632
rect 179873 139574 327783 139576
rect 179873 139571 179939 139574
rect 327717 139571 327783 139574
rect 31017 139498 31083 139501
rect 174813 139498 174879 139501
rect 31017 139496 174879 139498
rect 31017 139440 31022 139496
rect 31078 139440 174818 139496
rect 174874 139440 174879 139496
rect 31017 139438 174879 139440
rect 31017 139435 31083 139438
rect 174813 139435 174879 139438
rect 180190 139436 180196 139500
rect 180260 139498 180266 139500
rect 180260 139438 180810 139498
rect 180260 139436 180266 139438
rect 121913 139362 121979 139365
rect 118650 139360 121979 139362
rect 118650 139304 121918 139360
rect 121974 139304 121979 139360
rect 118650 139302 121979 139304
rect 115013 139226 115079 139229
rect 118650 139226 118710 139302
rect 121913 139299 121979 139302
rect 122046 139300 122052 139364
rect 122116 139362 122122 139364
rect 122741 139362 122807 139365
rect 122116 139360 122807 139362
rect 122116 139304 122746 139360
rect 122802 139304 122807 139360
rect 122116 139302 122807 139304
rect 122116 139300 122122 139302
rect 122741 139299 122807 139302
rect 122925 139362 122991 139365
rect 124121 139362 124187 139365
rect 122925 139360 124187 139362
rect 122925 139304 122930 139360
rect 122986 139304 124126 139360
rect 124182 139304 124187 139360
rect 122925 139302 124187 139304
rect 122925 139299 122991 139302
rect 124121 139299 124187 139302
rect 126462 139300 126468 139364
rect 126532 139362 126538 139364
rect 126881 139362 126947 139365
rect 129641 139364 129707 139365
rect 129590 139362 129596 139364
rect 126532 139360 126947 139362
rect 126532 139304 126886 139360
rect 126942 139304 126947 139360
rect 126532 139302 126947 139304
rect 129550 139302 129596 139362
rect 129660 139360 129707 139364
rect 131665 139362 131731 139365
rect 132217 139362 132283 139365
rect 138289 139362 138355 139365
rect 129702 139304 129707 139360
rect 126532 139300 126538 139302
rect 126881 139299 126947 139302
rect 129590 139300 129596 139302
rect 129660 139300 129707 139304
rect 129641 139299 129707 139300
rect 131622 139360 131731 139362
rect 131622 139304 131670 139360
rect 131726 139304 131731 139360
rect 131622 139299 131731 139304
rect 131806 139360 132283 139362
rect 131806 139304 132222 139360
rect 132278 139304 132283 139360
rect 131806 139302 132283 139304
rect 115013 139224 118710 139226
rect 115013 139168 115018 139224
rect 115074 139168 118710 139224
rect 115013 139166 118710 139168
rect 115013 139163 115079 139166
rect 120022 139164 120028 139228
rect 120092 139226 120098 139228
rect 122189 139226 122255 139229
rect 120092 139224 122255 139226
rect 120092 139168 122194 139224
rect 122250 139168 122255 139224
rect 120092 139166 122255 139168
rect 120092 139164 120098 139166
rect 122189 139163 122255 139166
rect 120942 139028 120948 139092
rect 121012 139090 121018 139092
rect 131622 139090 131682 139299
rect 121012 139030 131682 139090
rect 121012 139028 121018 139030
rect 115105 138954 115171 138957
rect 131806 138954 131866 139302
rect 132217 139299 132283 139302
rect 137970 139360 138355 139362
rect 137970 139304 138294 139360
rect 138350 139304 138355 139360
rect 137970 139302 138355 139304
rect 115105 138952 131866 138954
rect 115105 138896 115110 138952
rect 115166 138896 131866 138952
rect 115105 138894 131866 138896
rect 115105 138891 115171 138894
rect 116761 138818 116827 138821
rect 137970 138818 138030 139302
rect 138289 139299 138355 139302
rect 150934 139300 150940 139364
rect 151004 139362 151010 139364
rect 151077 139362 151143 139365
rect 152365 139362 152431 139365
rect 151004 139360 151143 139362
rect 151004 139304 151082 139360
rect 151138 139304 151143 139360
rect 151004 139302 151143 139304
rect 151004 139300 151010 139302
rect 151077 139299 151143 139302
rect 151770 139360 152431 139362
rect 151770 139304 152370 139360
rect 152426 139304 152431 139360
rect 151770 139302 152431 139304
rect 116761 138816 138030 138818
rect 116761 138760 116766 138816
rect 116822 138760 138030 138816
rect 116761 138758 138030 138760
rect 116761 138755 116827 138758
rect 118550 138620 118556 138684
rect 118620 138682 118626 138684
rect 151770 138682 151830 139302
rect 152365 139299 152431 139302
rect 154798 139300 154804 139364
rect 154868 139362 154874 139364
rect 155125 139362 155191 139365
rect 154868 139360 155191 139362
rect 154868 139304 155130 139360
rect 155186 139304 155191 139360
rect 154868 139302 155191 139304
rect 154868 139300 154874 139302
rect 155125 139299 155191 139302
rect 155350 139300 155356 139364
rect 155420 139362 155426 139364
rect 155677 139362 155743 139365
rect 155420 139360 155743 139362
rect 155420 139304 155682 139360
rect 155738 139304 155743 139360
rect 155420 139302 155743 139304
rect 155420 139300 155426 139302
rect 155677 139299 155743 139302
rect 159214 139300 159220 139364
rect 159284 139362 159290 139364
rect 159541 139362 159607 139365
rect 160001 139364 160067 139365
rect 159950 139362 159956 139364
rect 159284 139360 159607 139362
rect 159284 139304 159546 139360
rect 159602 139304 159607 139360
rect 159284 139302 159607 139304
rect 159910 139302 159956 139362
rect 160020 139360 160067 139364
rect 160062 139304 160067 139360
rect 159284 139300 159290 139302
rect 159541 139299 159607 139302
rect 159950 139300 159956 139302
rect 160020 139300 160067 139304
rect 160001 139299 160067 139300
rect 163957 139362 164023 139365
rect 179689 139362 179755 139365
rect 180517 139362 180583 139365
rect 180750 139362 180810 139438
rect 195094 139436 195100 139500
rect 195164 139498 195170 139500
rect 195605 139498 195671 139501
rect 195164 139496 195671 139498
rect 195164 139440 195610 139496
rect 195666 139440 195671 139496
rect 195164 139438 195671 139440
rect 195164 139436 195170 139438
rect 195605 139435 195671 139438
rect 189257 139362 189323 139365
rect 194041 139362 194107 139365
rect 163957 139360 171150 139362
rect 163957 139304 163962 139360
rect 164018 139304 171150 139360
rect 163957 139302 171150 139304
rect 163957 139299 164023 139302
rect 118620 138622 151830 138682
rect 171090 138682 171150 139302
rect 179689 139360 179890 139362
rect 179689 139304 179694 139360
rect 179750 139304 179890 139360
rect 179689 139302 179890 139304
rect 179689 139299 179755 139302
rect 179830 138954 179890 139302
rect 180517 139360 180626 139362
rect 180517 139304 180522 139360
rect 180578 139304 180626 139360
rect 180517 139299 180626 139304
rect 180750 139360 189323 139362
rect 180750 139304 189262 139360
rect 189318 139304 189323 139360
rect 180750 139302 189323 139304
rect 189257 139299 189323 139302
rect 190410 139360 194107 139362
rect 190410 139304 194046 139360
rect 194102 139304 194107 139360
rect 190410 139302 194107 139304
rect 180566 139090 180626 139299
rect 186405 139226 186471 139229
rect 190410 139226 190470 139302
rect 194041 139299 194107 139302
rect 580349 139362 580415 139365
rect 583520 139362 584960 139452
rect 580349 139360 584960 139362
rect 580349 139304 580354 139360
rect 580410 139304 584960 139360
rect 580349 139302 584960 139304
rect 580349 139299 580415 139302
rect 186405 139224 190470 139226
rect 186405 139168 186410 139224
rect 186466 139168 190470 139224
rect 583520 139212 584960 139302
rect 186405 139166 190470 139168
rect 186405 139163 186471 139166
rect 189441 139090 189507 139093
rect 180566 139088 189507 139090
rect 180566 139032 189446 139088
rect 189502 139032 189507 139088
rect 180566 139030 189507 139032
rect 189441 139027 189507 139030
rect 179830 138894 180810 138954
rect 180750 138818 180810 138894
rect 183318 138892 183324 138956
rect 183388 138954 183394 138956
rect 193673 138954 193739 138957
rect 183388 138952 193739 138954
rect 183388 138896 193678 138952
rect 193734 138896 193739 138952
rect 183388 138894 193739 138896
rect 183388 138892 183394 138894
rect 193673 138891 193739 138894
rect 190913 138818 190979 138821
rect 180750 138816 190979 138818
rect 180750 138760 190918 138816
rect 190974 138760 190979 138816
rect 180750 138758 190979 138760
rect 190913 138755 190979 138758
rect 196525 138682 196591 138685
rect 171090 138680 196591 138682
rect 171090 138624 196530 138680
rect 196586 138624 196591 138680
rect 171090 138622 196591 138624
rect 118620 138620 118626 138622
rect 196525 138619 196591 138622
rect 119245 138546 119311 138549
rect 122373 138546 122439 138549
rect 119245 138544 122439 138546
rect 119245 138488 119250 138544
rect 119306 138488 122378 138544
rect 122434 138488 122439 138544
rect 119245 138486 122439 138488
rect 119245 138483 119311 138486
rect 122373 138483 122439 138486
rect 184790 138484 184796 138548
rect 184860 138546 184866 138548
rect 191097 138546 191163 138549
rect 184860 138544 191163 138546
rect 184860 138488 191102 138544
rect 191158 138488 191163 138544
rect 184860 138486 191163 138488
rect 184860 138484 184866 138486
rect 191097 138483 191163 138486
rect 187049 138140 187115 138141
rect 186998 138138 187004 138140
rect 186958 138078 187004 138138
rect 187068 138136 187115 138140
rect 187110 138080 187115 138136
rect 186998 138076 187004 138078
rect 187068 138076 187115 138080
rect 187049 138075 187115 138076
rect 122741 138004 122807 138005
rect 122741 138000 122788 138004
rect 122852 138002 122858 138004
rect 122741 137944 122746 138000
rect 122741 137940 122788 137944
rect 122852 137942 122898 138002
rect 122852 137940 122858 137942
rect 122741 137939 122807 137940
rect 186078 137396 186084 137460
rect 186148 137458 186154 137460
rect 197721 137458 197787 137461
rect 186148 137456 197787 137458
rect 186148 137400 197726 137456
rect 197782 137400 197787 137456
rect 186148 137398 197787 137400
rect 186148 137396 186154 137398
rect 197721 137395 197787 137398
rect 189022 137260 189028 137324
rect 189092 137322 189098 137324
rect 580349 137322 580415 137325
rect 189092 137320 580415 137322
rect 189092 137264 580354 137320
rect 580410 137264 580415 137320
rect 189092 137262 580415 137264
rect 189092 137260 189098 137262
rect 580349 137259 580415 137262
rect -960 136778 480 136868
rect 3509 136778 3575 136781
rect -960 136776 3575 136778
rect -960 136720 3514 136776
rect 3570 136720 3575 136776
rect -960 136718 3575 136720
rect -960 136628 480 136718
rect 3509 136715 3575 136718
rect 119654 130324 119660 130388
rect 119724 130386 119730 130388
rect 120022 130386 120028 130388
rect 119724 130326 120028 130386
rect 119724 130324 119730 130326
rect 120022 130324 120028 130326
rect 120092 130324 120098 130388
rect 122741 128484 122807 128485
rect 122741 128482 122788 128484
rect 122696 128480 122788 128482
rect 122696 128424 122746 128480
rect 122696 128422 122788 128424
rect 122741 128420 122788 128422
rect 122852 128420 122858 128484
rect 122741 128419 122807 128420
rect 580533 126034 580599 126037
rect 583520 126034 584960 126124
rect 580533 126032 584960 126034
rect 580533 125976 580538 126032
rect 580594 125976 584960 126032
rect 580533 125974 584960 125976
rect 580533 125971 580599 125974
rect 583520 125884 584960 125974
rect -960 123572 480 123812
rect 122741 122908 122807 122909
rect 122741 122906 122788 122908
rect 122696 122904 122788 122906
rect 122852 122906 122858 122908
rect 122696 122848 122746 122904
rect 122696 122846 122788 122848
rect 122741 122844 122788 122846
rect 122852 122846 122934 122906
rect 122852 122844 122858 122846
rect 122741 122843 122807 122844
rect 122741 122772 122807 122773
rect 122741 122770 122788 122772
rect 122696 122768 122788 122770
rect 122852 122770 122858 122772
rect 122696 122712 122746 122768
rect 122696 122710 122788 122712
rect 122741 122708 122788 122710
rect 122852 122710 122934 122770
rect 122852 122708 122858 122710
rect 122741 122707 122807 122708
rect 191046 114412 191052 114476
rect 191116 114474 191122 114476
rect 191189 114474 191255 114477
rect 191116 114472 191255 114474
rect 191116 114416 191194 114472
rect 191250 114416 191255 114472
rect 191116 114414 191255 114416
rect 191116 114412 191122 114414
rect 191189 114411 191255 114414
rect 122782 113324 122788 113388
rect 122852 113324 122858 113388
rect 122790 113253 122850 113324
rect 122741 113250 122850 113253
rect 122696 113248 122850 113250
rect 122696 113192 122746 113248
rect 122802 113192 122850 113248
rect 122696 113190 122850 113192
rect 122741 113187 122807 113190
rect 122741 113114 122807 113117
rect 122696 113112 122850 113114
rect 122696 113056 122746 113112
rect 122802 113056 122850 113112
rect 122696 113054 122850 113056
rect 122741 113051 122850 113054
rect 122790 112980 122850 113051
rect 122782 112916 122788 112980
rect 122852 112916 122858 112980
rect 580441 112842 580507 112845
rect 583520 112842 584960 112932
rect 580441 112840 584960 112842
rect 580441 112784 580446 112840
rect 580502 112784 584960 112840
rect 580441 112782 584960 112784
rect 580441 112779 580507 112782
rect 583520 112692 584960 112782
rect -960 110666 480 110756
rect 3141 110666 3207 110669
rect -960 110664 3207 110666
rect -960 110608 3146 110664
rect 3202 110608 3207 110664
rect -960 110606 3207 110608
rect -960 110516 480 110606
rect 3141 110603 3207 110606
rect 122741 103596 122807 103597
rect 122741 103594 122788 103596
rect 122696 103592 122788 103594
rect 122852 103594 122858 103596
rect 122696 103536 122746 103592
rect 122696 103534 122788 103536
rect 122741 103532 122788 103534
rect 122852 103534 122934 103594
rect 122852 103532 122858 103534
rect 122741 103531 122807 103532
rect 122741 103458 122807 103461
rect 122696 103456 122850 103458
rect 122696 103400 122746 103456
rect 122802 103400 122850 103456
rect 122696 103398 122850 103400
rect 122741 103395 122850 103398
rect 122790 103324 122850 103395
rect 122782 103260 122788 103324
rect 122852 103260 122858 103324
rect 580349 99514 580415 99517
rect 583520 99514 584960 99604
rect 580349 99512 584960 99514
rect 580349 99456 580354 99512
rect 580410 99456 584960 99512
rect 580349 99454 584960 99456
rect 580349 99451 580415 99454
rect 583520 99364 584960 99454
rect -960 97610 480 97700
rect -960 97550 674 97610
rect -960 97474 480 97550
rect 614 97474 674 97550
rect -960 97460 674 97474
rect 246 97414 674 97460
rect 246 96930 306 97414
rect 246 96870 6930 96930
rect 6870 96658 6930 96870
rect 119470 96658 119476 96660
rect 6870 96598 119476 96658
rect 119470 96596 119476 96598
rect 119540 96596 119546 96660
rect 122741 93940 122807 93941
rect 122741 93938 122788 93940
rect 122696 93936 122788 93938
rect 122852 93938 122858 93940
rect 122696 93880 122746 93936
rect 122696 93878 122788 93880
rect 122741 93876 122788 93878
rect 122852 93878 122934 93938
rect 122852 93876 122858 93878
rect 122741 93875 122807 93876
rect 122741 93802 122807 93805
rect 122696 93800 122850 93802
rect 122696 93744 122746 93800
rect 122802 93744 122850 93800
rect 122696 93742 122850 93744
rect 122741 93739 122850 93742
rect 122790 93668 122850 93739
rect 122782 93604 122788 93668
rect 122852 93604 122858 93668
rect 122741 89724 122807 89725
rect 122741 89722 122788 89724
rect 122696 89720 122788 89722
rect 122696 89664 122746 89720
rect 122696 89662 122788 89664
rect 122741 89660 122788 89662
rect 122852 89660 122858 89724
rect 122741 89659 122807 89660
rect 580165 86186 580231 86189
rect 583520 86186 584960 86276
rect 580165 86184 584960 86186
rect 580165 86128 580170 86184
rect 580226 86128 584960 86184
rect 580165 86126 584960 86128
rect 580165 86123 580231 86126
rect 583520 86036 584960 86126
rect -960 84690 480 84780
rect -960 84630 6930 84690
rect -960 84540 480 84630
rect 6870 84282 6930 84630
rect 119286 84282 119292 84284
rect 6870 84222 119292 84282
rect 119286 84220 119292 84222
rect 119356 84220 119362 84284
rect 119654 83404 119660 83468
rect 119724 83466 119730 83468
rect 120022 83466 120028 83468
rect 119724 83406 120028 83466
rect 119724 83404 119730 83406
rect 120022 83404 120028 83406
rect 120092 83404 120098 83468
rect 127566 81908 127572 81972
rect 127636 81970 127642 81972
rect 145782 81970 145788 81972
rect 127636 81910 145788 81970
rect 127636 81908 127642 81910
rect 145782 81908 145788 81910
rect 145852 81908 145858 81972
rect 160686 81908 160692 81972
rect 160756 81970 160762 81972
rect 161238 81970 161244 81972
rect 160756 81910 161244 81970
rect 160756 81908 160762 81910
rect 161238 81908 161244 81910
rect 161308 81908 161314 81972
rect 185342 81908 185348 81972
rect 185412 81970 185418 81972
rect 191189 81970 191255 81973
rect 185412 81968 191255 81970
rect 185412 81912 191194 81968
rect 191250 81912 191255 81968
rect 185412 81910 191255 81912
rect 185412 81908 185418 81910
rect 191189 81907 191255 81910
rect 122230 81364 122236 81428
rect 122300 81426 122306 81428
rect 122465 81426 122531 81429
rect 122300 81424 122531 81426
rect 122300 81368 122470 81424
rect 122526 81368 122531 81424
rect 122300 81366 122531 81368
rect 122300 81364 122306 81366
rect 122465 81363 122531 81366
rect 140814 81364 140820 81428
rect 140884 81426 140890 81428
rect 141734 81426 141740 81428
rect 140884 81366 141740 81426
rect 140884 81364 140890 81366
rect 141734 81364 141740 81366
rect 141804 81364 141810 81428
rect 130694 81228 130700 81292
rect 130764 81290 130770 81292
rect 143022 81290 143028 81292
rect 130764 81230 143028 81290
rect 130764 81228 130770 81230
rect 143022 81228 143028 81230
rect 143092 81228 143098 81292
rect 172462 81228 172468 81292
rect 172532 81290 172538 81292
rect 195329 81290 195395 81293
rect 172532 81288 195395 81290
rect 172532 81232 195334 81288
rect 195390 81232 195395 81288
rect 172532 81230 195395 81232
rect 172532 81228 172538 81230
rect 195329 81227 195395 81230
rect 130510 81092 130516 81156
rect 130580 81154 130586 81156
rect 143390 81154 143396 81156
rect 130580 81094 143396 81154
rect 130580 81092 130586 81094
rect 143390 81092 143396 81094
rect 143460 81092 143466 81156
rect 171910 81092 171916 81156
rect 171980 81154 171986 81156
rect 196985 81154 197051 81157
rect 171980 81152 197051 81154
rect 171980 81096 196990 81152
rect 197046 81096 197051 81152
rect 171980 81094 197051 81096
rect 171980 81092 171986 81094
rect 196985 81091 197051 81094
rect 122966 80956 122972 81020
rect 123036 81018 123042 81020
rect 143206 81018 143212 81020
rect 123036 80958 143212 81018
rect 123036 80956 123042 80958
rect 143206 80956 143212 80958
rect 143276 80956 143282 81020
rect 145414 80956 145420 81020
rect 145484 81018 145490 81020
rect 147622 81018 147628 81020
rect 145484 80958 147628 81018
rect 145484 80956 145490 80958
rect 147622 80956 147628 80958
rect 147692 80956 147698 81020
rect 155902 80956 155908 81020
rect 155972 81018 155978 81020
rect 186497 81018 186563 81021
rect 155972 81016 186563 81018
rect 155972 80960 186502 81016
rect 186558 80960 186563 81016
rect 155972 80958 186563 80960
rect 155972 80956 155978 80958
rect 186497 80955 186563 80958
rect 187141 81020 187207 81021
rect 187141 81016 187188 81020
rect 187252 81018 187258 81020
rect 187417 81018 187483 81021
rect 198089 81018 198155 81021
rect 187141 80960 187146 81016
rect 187141 80956 187188 80960
rect 187252 80958 187298 81018
rect 187417 81016 198155 81018
rect 187417 80960 187422 81016
rect 187478 80960 198094 81016
rect 198150 80960 198155 81016
rect 187417 80958 198155 80960
rect 187252 80956 187258 80958
rect 187141 80955 187207 80956
rect 187417 80955 187483 80958
rect 198089 80955 198155 80958
rect 126646 80820 126652 80884
rect 126716 80882 126722 80884
rect 146518 80882 146524 80884
rect 126716 80822 146524 80882
rect 126716 80820 126722 80822
rect 146518 80820 146524 80822
rect 146588 80820 146594 80884
rect 148358 80820 148364 80884
rect 148428 80882 148434 80884
rect 161422 80882 161428 80884
rect 148428 80822 161428 80882
rect 148428 80820 148434 80822
rect 161422 80820 161428 80822
rect 161492 80820 161498 80884
rect 180006 80882 180012 80884
rect 162672 80822 180012 80882
rect 146702 80746 146708 80748
rect 128310 80686 146708 80746
rect 122414 80548 122420 80612
rect 122484 80610 122490 80612
rect 128310 80610 128370 80686
rect 146702 80684 146708 80686
rect 146772 80684 146778 80748
rect 154430 80684 154436 80748
rect 154500 80746 154506 80748
rect 162672 80746 162732 80822
rect 180006 80820 180012 80822
rect 180076 80820 180082 80884
rect 154500 80686 162732 80746
rect 154500 80684 154506 80686
rect 177246 80684 177252 80748
rect 177316 80746 177322 80748
rect 177757 80746 177823 80749
rect 178401 80748 178467 80749
rect 178350 80746 178356 80748
rect 177316 80744 177823 80746
rect 177316 80688 177762 80744
rect 177818 80688 177823 80744
rect 177316 80686 177823 80688
rect 178310 80686 178356 80746
rect 178420 80744 178467 80748
rect 200941 80746 201007 80749
rect 178462 80688 178467 80744
rect 177316 80684 177322 80686
rect 177757 80683 177823 80686
rect 178350 80684 178356 80686
rect 178420 80684 178467 80688
rect 178401 80683 178467 80684
rect 179370 80744 201007 80746
rect 179370 80688 200946 80744
rect 201002 80688 201007 80744
rect 179370 80686 201007 80688
rect 122484 80550 128370 80610
rect 132033 80610 132099 80613
rect 133086 80610 133092 80612
rect 132033 80608 133092 80610
rect 132033 80552 132038 80608
rect 132094 80552 133092 80608
rect 132033 80550 133092 80552
rect 122484 80548 122490 80550
rect 132033 80547 132099 80550
rect 133086 80548 133092 80550
rect 133156 80548 133162 80612
rect 147438 80548 147444 80612
rect 147508 80610 147514 80612
rect 147508 80550 158132 80610
rect 147508 80548 147514 80550
rect 131941 80474 132007 80477
rect 133454 80474 133460 80476
rect 131941 80472 133460 80474
rect 131941 80416 131946 80472
rect 132002 80416 133460 80472
rect 131941 80414 133460 80416
rect 131941 80411 132007 80414
rect 133454 80412 133460 80414
rect 133524 80412 133530 80476
rect 138606 80412 138612 80476
rect 138676 80474 138682 80476
rect 147254 80474 147260 80476
rect 138676 80414 147260 80474
rect 138676 80412 138682 80414
rect 147254 80412 147260 80414
rect 147324 80412 147330 80476
rect 149462 80412 149468 80476
rect 149532 80474 149538 80476
rect 158072 80474 158132 80550
rect 159214 80548 159220 80612
rect 159284 80610 159290 80612
rect 177849 80610 177915 80613
rect 159284 80608 177915 80610
rect 159284 80552 177854 80608
rect 177910 80552 177915 80608
rect 159284 80550 177915 80552
rect 159284 80548 159290 80550
rect 177849 80547 177915 80550
rect 161790 80474 161796 80476
rect 149532 80414 150450 80474
rect 158072 80414 161796 80474
rect 149532 80412 149538 80414
rect 122833 80340 122899 80341
rect 122782 80338 122788 80340
rect 122742 80278 122788 80338
rect 122852 80336 122899 80340
rect 122894 80280 122899 80336
rect 122782 80276 122788 80278
rect 122852 80276 122899 80280
rect 122833 80275 122899 80276
rect 131757 80338 131823 80341
rect 140814 80338 140820 80340
rect 131757 80336 140820 80338
rect 131757 80280 131762 80336
rect 131818 80280 140820 80336
rect 131757 80278 140820 80280
rect 131757 80275 131823 80278
rect 140814 80276 140820 80278
rect 140884 80338 140890 80340
rect 141918 80338 141924 80340
rect 140884 80278 141924 80338
rect 140884 80276 140890 80278
rect 141918 80276 141924 80278
rect 141988 80276 141994 80340
rect 117773 80202 117839 80205
rect 138606 80202 138612 80204
rect 117773 80200 138612 80202
rect 117773 80144 117778 80200
rect 117834 80144 138612 80200
rect 117773 80142 138612 80144
rect 117773 80139 117839 80142
rect 138606 80140 138612 80142
rect 138676 80140 138682 80204
rect 150390 80202 150450 80414
rect 161790 80412 161796 80414
rect 161860 80412 161866 80476
rect 178534 80474 178540 80476
rect 173022 80414 178540 80474
rect 150934 80276 150940 80340
rect 151004 80338 151010 80340
rect 151670 80338 151676 80340
rect 151004 80278 151676 80338
rect 151004 80276 151010 80278
rect 151670 80276 151676 80278
rect 151740 80276 151746 80340
rect 158846 80276 158852 80340
rect 158916 80338 158922 80340
rect 173022 80338 173082 80414
rect 178534 80412 178540 80414
rect 178604 80412 178610 80476
rect 158916 80278 159788 80338
rect 158916 80276 158922 80278
rect 150390 80142 159190 80202
rect 134926 80066 134932 80068
rect 133922 80006 134932 80066
rect 132539 79962 132605 79967
rect 131614 79868 131620 79932
rect 131684 79930 131690 79932
rect 132309 79930 132375 79933
rect 131684 79928 132375 79930
rect 131684 79872 132314 79928
rect 132370 79872 132375 79928
rect 132539 79906 132544 79962
rect 132600 79906 132605 79962
rect 132539 79901 132605 79906
rect 133091 79962 133157 79967
rect 133091 79906 133096 79962
rect 133152 79906 133157 79962
rect 133922 79933 133982 80006
rect 134926 80004 134932 80006
rect 134996 80004 135002 80068
rect 135110 80004 135116 80068
rect 135180 80066 135186 80068
rect 137870 80066 137876 80068
rect 135180 80006 136512 80066
rect 135180 80004 135186 80006
rect 136452 79967 136512 80006
rect 137326 80006 137876 80066
rect 136452 79962 136561 79967
rect 133091 79901 133157 79906
rect 131684 79870 132375 79872
rect 131684 79868 131690 79870
rect 132309 79867 132375 79870
rect 126462 79732 126468 79796
rect 126532 79794 126538 79796
rect 130653 79794 130719 79797
rect 126532 79792 130719 79794
rect 126532 79736 130658 79792
rect 130714 79736 130719 79792
rect 126532 79734 130719 79736
rect 126532 79732 126538 79734
rect 130653 79731 130719 79734
rect 130929 79794 130995 79797
rect 132542 79794 132602 79901
rect 133094 79831 133154 79901
rect 133454 79868 133460 79932
rect 133524 79930 133530 79932
rect 133919 79930 133985 79933
rect 133524 79928 133985 79930
rect 133524 79872 133924 79928
rect 133980 79872 133985 79928
rect 133524 79870 133985 79872
rect 133524 79868 133530 79870
rect 133919 79867 133985 79870
rect 134190 79868 134196 79932
rect 134260 79930 134266 79932
rect 134471 79930 134537 79933
rect 134260 79928 134537 79930
rect 134260 79872 134476 79928
rect 134532 79872 134537 79928
rect 134260 79870 134537 79872
rect 134260 79868 134266 79870
rect 134471 79867 134537 79870
rect 134742 79868 134748 79932
rect 134812 79930 134818 79932
rect 134812 79899 134856 79930
rect 134812 79894 134905 79899
rect 134812 79868 134844 79894
rect 134796 79838 134844 79868
rect 134900 79838 134905 79894
rect 135478 79868 135484 79932
rect 135548 79930 135554 79932
rect 135759 79930 135825 79933
rect 136452 79932 136500 79962
rect 135548 79928 135825 79930
rect 135548 79872 135764 79928
rect 135820 79872 135825 79928
rect 135548 79870 135825 79872
rect 135548 79868 135554 79870
rect 135759 79867 135825 79870
rect 136398 79868 136404 79932
rect 136468 79906 136500 79932
rect 136556 79906 136561 79962
rect 136955 79932 137021 79933
rect 136950 79930 136956 79932
rect 136468 79901 136561 79906
rect 136468 79870 136512 79901
rect 136864 79870 136956 79930
rect 136468 79868 136474 79870
rect 136950 79868 136956 79870
rect 137020 79868 137026 79932
rect 136955 79867 137021 79868
rect 134796 79836 134905 79838
rect 134839 79833 134905 79836
rect 137326 79831 137386 80006
rect 137870 80004 137876 80006
rect 137940 80004 137946 80068
rect 138790 80066 138796 80068
rect 138430 80006 138796 80066
rect 138243 79962 138309 79967
rect 137502 79868 137508 79932
rect 137572 79930 137578 79932
rect 137875 79930 137941 79933
rect 137572 79928 137941 79930
rect 137572 79872 137880 79928
rect 137936 79872 137941 79928
rect 137572 79870 137941 79872
rect 137572 79868 137578 79870
rect 137875 79867 137941 79870
rect 138054 79868 138060 79932
rect 138124 79930 138130 79932
rect 138243 79930 138248 79962
rect 138124 79906 138248 79930
rect 138304 79906 138309 79962
rect 138430 79933 138490 80006
rect 138790 80004 138796 80006
rect 138860 80004 138866 80068
rect 140262 80066 140268 80068
rect 140086 80006 140268 80066
rect 140086 79933 140146 80006
rect 140262 80004 140268 80006
rect 140332 80004 140338 80068
rect 140446 80066 140452 80068
rect 140408 80004 140452 80066
rect 140516 80004 140522 80068
rect 151854 80004 151860 80068
rect 151924 80066 151930 80068
rect 154062 80066 154068 80068
rect 151924 80006 152474 80066
rect 151924 80004 151930 80006
rect 140408 79933 140468 80004
rect 142567 79964 142633 79967
rect 142524 79962 142633 79964
rect 138124 79901 138309 79906
rect 138427 79928 138493 79933
rect 138979 79932 139045 79933
rect 139531 79932 139597 79933
rect 138974 79930 138980 79932
rect 138124 79870 138306 79901
rect 138427 79872 138432 79928
rect 138488 79872 138493 79928
rect 138124 79868 138130 79870
rect 138427 79867 138493 79872
rect 138888 79870 138980 79930
rect 138974 79868 138980 79870
rect 139044 79868 139050 79932
rect 139526 79930 139532 79932
rect 139440 79870 139532 79930
rect 139526 79868 139532 79870
rect 139596 79868 139602 79932
rect 139715 79930 139781 79933
rect 139894 79930 139900 79932
rect 139715 79928 139900 79930
rect 139715 79872 139720 79928
rect 139776 79872 139900 79928
rect 139715 79870 139900 79872
rect 138979 79867 139045 79868
rect 139531 79867 139597 79868
rect 139715 79867 139781 79870
rect 139894 79868 139900 79870
rect 139964 79868 139970 79932
rect 140083 79928 140149 79933
rect 140083 79872 140088 79928
rect 140144 79872 140149 79928
rect 140083 79867 140149 79872
rect 140359 79928 140468 79933
rect 140635 79932 140701 79933
rect 140359 79872 140364 79928
rect 140420 79872 140468 79928
rect 140359 79867 140468 79872
rect 140630 79868 140636 79932
rect 140700 79930 140706 79932
rect 141187 79930 141253 79933
rect 141739 79932 141805 79933
rect 141550 79930 141556 79932
rect 140700 79870 140792 79930
rect 141187 79928 141556 79930
rect 141187 79872 141192 79928
rect 141248 79872 141556 79928
rect 141187 79870 141556 79872
rect 140700 79868 140706 79870
rect 140635 79867 140701 79868
rect 141187 79867 141253 79870
rect 141550 79868 141556 79870
rect 141620 79868 141626 79932
rect 141734 79868 141740 79932
rect 141804 79930 141810 79932
rect 141804 79870 141896 79930
rect 142524 79906 142572 79962
rect 142628 79930 142633 79962
rect 142843 79962 142909 79967
rect 142628 79906 142722 79930
rect 142524 79870 142722 79906
rect 142843 79906 142848 79962
rect 142904 79906 142909 79962
rect 142843 79901 142909 79906
rect 143027 79962 143093 79967
rect 143027 79906 143032 79962
rect 143088 79906 143093 79962
rect 143395 79962 143461 79967
rect 145879 79964 145945 79967
rect 143027 79901 143093 79906
rect 141804 79868 141810 79870
rect 141739 79867 141805 79868
rect 130929 79792 132602 79794
rect 130929 79736 130934 79792
rect 130990 79736 132602 79792
rect 133091 79826 133157 79831
rect 133091 79770 133096 79826
rect 133152 79770 133157 79826
rect 137323 79826 137389 79831
rect 133551 79794 133617 79797
rect 134333 79796 134399 79797
rect 133091 79765 133157 79770
rect 133508 79792 133617 79794
rect 130929 79734 132602 79736
rect 133508 79736 133556 79792
rect 133612 79736 133617 79792
rect 130929 79731 130995 79734
rect 133508 79731 133617 79736
rect 133822 79732 133828 79796
rect 133892 79794 133898 79796
rect 134333 79794 134380 79796
rect 133892 79792 134380 79794
rect 133892 79736 134338 79792
rect 133892 79734 134380 79736
rect 133892 79732 133898 79734
rect 134333 79732 134380 79734
rect 134444 79732 134450 79796
rect 135662 79732 135668 79796
rect 135732 79794 135738 79796
rect 135897 79794 135963 79797
rect 137323 79794 137328 79826
rect 135732 79792 135963 79794
rect 135732 79736 135902 79792
rect 135958 79736 135963 79792
rect 135732 79734 135963 79736
rect 135732 79732 135738 79734
rect 134333 79731 134399 79732
rect 135897 79731 135963 79734
rect 136820 79770 137328 79794
rect 137384 79770 137389 79826
rect 136820 79765 137389 79770
rect 137878 79797 137938 79867
rect 140408 79797 140468 79867
rect 142662 79797 142722 79870
rect 142846 79797 142906 79901
rect 143030 79797 143090 79901
rect 143206 79868 143212 79932
rect 143276 79930 143282 79932
rect 143395 79930 143400 79962
rect 143276 79906 143400 79930
rect 143456 79906 143461 79962
rect 145836 79962 145945 79964
rect 143947 79932 144013 79933
rect 143942 79930 143948 79932
rect 143276 79901 143461 79906
rect 143276 79870 143458 79901
rect 143856 79870 143948 79930
rect 143276 79868 143282 79870
rect 143942 79868 143948 79870
rect 144012 79868 144018 79932
rect 145414 79868 145420 79932
rect 145484 79930 145490 79932
rect 145836 79930 145884 79962
rect 145484 79906 145884 79930
rect 145940 79906 145945 79962
rect 147627 79962 147693 79967
rect 145484 79901 145945 79906
rect 145484 79870 145896 79901
rect 145484 79868 145490 79870
rect 146518 79868 146524 79932
rect 146588 79930 146594 79932
rect 146707 79930 146773 79933
rect 146588 79928 146773 79930
rect 146588 79872 146712 79928
rect 146768 79872 146773 79928
rect 146588 79870 146773 79872
rect 146588 79868 146594 79870
rect 143947 79867 144013 79868
rect 146707 79867 146773 79870
rect 146886 79868 146892 79932
rect 146956 79930 146962 79932
rect 147438 79930 147444 79932
rect 146956 79870 147444 79930
rect 146956 79868 146962 79870
rect 147438 79868 147444 79870
rect 147508 79868 147514 79932
rect 147627 79906 147632 79962
rect 147688 79930 147693 79962
rect 149283 79962 149349 79967
rect 147806 79930 147812 79932
rect 147688 79906 147812 79930
rect 147627 79901 147812 79906
rect 147630 79870 147812 79901
rect 147806 79868 147812 79870
rect 147876 79868 147882 79932
rect 148547 79928 148613 79933
rect 148547 79872 148552 79928
rect 148608 79872 148613 79928
rect 148547 79867 148613 79872
rect 148731 79930 148797 79933
rect 149094 79930 149100 79932
rect 148731 79928 149100 79930
rect 148731 79872 148736 79928
rect 148792 79872 149100 79928
rect 148731 79870 149100 79872
rect 148731 79867 148797 79870
rect 149094 79868 149100 79870
rect 149164 79868 149170 79932
rect 149283 79906 149288 79962
rect 149344 79906 149349 79962
rect 150019 79962 150085 79967
rect 149283 79901 149349 79906
rect 148550 79797 148610 79867
rect 137878 79792 137987 79797
rect 136820 79734 137386 79765
rect 137878 79736 137926 79792
rect 137982 79736 137987 79792
rect 137878 79734 137987 79736
rect 120758 79596 120764 79660
rect 120828 79658 120834 79660
rect 124121 79658 124187 79661
rect 120828 79656 124187 79658
rect 120828 79600 124126 79656
rect 124182 79600 124187 79656
rect 120828 79598 124187 79600
rect 120828 79596 120834 79598
rect 124121 79595 124187 79598
rect 132902 79596 132908 79660
rect 132972 79658 132978 79660
rect 133508 79658 133568 79731
rect 136820 79661 136880 79734
rect 137921 79731 137987 79734
rect 138059 79794 138125 79797
rect 138841 79796 138907 79797
rect 138422 79794 138428 79796
rect 138059 79792 138428 79794
rect 138059 79736 138064 79792
rect 138120 79736 138428 79792
rect 138059 79734 138428 79736
rect 138059 79731 138125 79734
rect 138422 79732 138428 79734
rect 138492 79732 138498 79796
rect 138790 79732 138796 79796
rect 138860 79794 138907 79796
rect 139071 79794 139137 79797
rect 139301 79794 139367 79797
rect 138860 79792 138952 79794
rect 138902 79736 138952 79792
rect 138860 79734 138952 79736
rect 139071 79792 139367 79794
rect 139071 79736 139076 79792
rect 139132 79736 139306 79792
rect 139362 79736 139367 79792
rect 139071 79734 139367 79736
rect 138860 79732 138907 79734
rect 138841 79731 138907 79732
rect 139071 79731 139137 79734
rect 139301 79731 139367 79734
rect 139807 79794 139873 79797
rect 140078 79794 140084 79796
rect 139807 79792 140084 79794
rect 139807 79736 139812 79792
rect 139868 79736 140084 79792
rect 139807 79734 140084 79736
rect 139807 79731 139873 79734
rect 140078 79732 140084 79734
rect 140148 79732 140154 79796
rect 140405 79792 140471 79797
rect 140405 79736 140410 79792
rect 140466 79736 140471 79792
rect 140405 79731 140471 79736
rect 140681 79794 140747 79797
rect 140814 79794 140820 79796
rect 140681 79792 140820 79794
rect 140681 79736 140686 79792
rect 140742 79736 140820 79792
rect 140681 79734 140820 79736
rect 140681 79731 140747 79734
rect 140814 79732 140820 79734
rect 140884 79732 140890 79796
rect 142662 79792 142771 79797
rect 142662 79736 142710 79792
rect 142766 79736 142771 79792
rect 142662 79734 142771 79736
rect 142846 79792 142955 79797
rect 142846 79736 142894 79792
rect 142950 79736 142955 79792
rect 142846 79734 142955 79736
rect 143030 79792 143139 79797
rect 143030 79736 143078 79792
rect 143134 79736 143139 79792
rect 143030 79734 143139 79736
rect 142705 79731 142771 79734
rect 142889 79731 142955 79734
rect 143073 79731 143139 79734
rect 144126 79732 144132 79796
rect 144196 79794 144202 79796
rect 144821 79794 144887 79797
rect 145833 79796 145899 79797
rect 144196 79792 144887 79794
rect 144196 79736 144826 79792
rect 144882 79736 144887 79792
rect 144196 79734 144887 79736
rect 144196 79732 144202 79734
rect 144821 79731 144887 79734
rect 145782 79732 145788 79796
rect 145852 79794 145899 79796
rect 145852 79792 145944 79794
rect 145894 79736 145944 79792
rect 145852 79734 145944 79736
rect 145852 79732 145899 79734
rect 146702 79732 146708 79796
rect 146772 79794 146778 79796
rect 146891 79794 146957 79797
rect 146772 79792 146957 79794
rect 146772 79736 146896 79792
rect 146952 79736 146957 79792
rect 146772 79734 146957 79736
rect 146772 79732 146778 79734
rect 145833 79731 145899 79732
rect 146891 79731 146957 79734
rect 147254 79732 147260 79796
rect 147324 79794 147330 79796
rect 147443 79794 147509 79797
rect 147995 79796 148061 79797
rect 147324 79792 147509 79794
rect 147324 79736 147448 79792
rect 147504 79736 147509 79792
rect 147324 79734 147509 79736
rect 147324 79732 147330 79734
rect 147443 79731 147509 79734
rect 147990 79732 147996 79796
rect 148060 79794 148066 79796
rect 148060 79734 148152 79794
rect 148501 79792 148610 79797
rect 148501 79736 148506 79792
rect 148562 79736 148610 79792
rect 148501 79734 148610 79736
rect 149286 79797 149346 79901
rect 149830 79868 149836 79932
rect 149900 79930 149906 79932
rect 150019 79930 150024 79962
rect 149900 79906 150024 79930
rect 150080 79906 150085 79962
rect 150847 79964 150913 79967
rect 151123 79964 151189 79967
rect 151399 79964 151465 79967
rect 150847 79962 150956 79964
rect 150295 79930 150361 79933
rect 149900 79901 150085 79906
rect 150252 79928 150361 79930
rect 149900 79870 150082 79901
rect 150252 79872 150300 79928
rect 150356 79872 150361 79928
rect 150847 79906 150852 79962
rect 150908 79906 150956 79962
rect 151123 79962 151246 79964
rect 151123 79932 151128 79962
rect 151184 79932 151246 79962
rect 150847 79901 150956 79906
rect 149900 79868 149906 79870
rect 150252 79867 150361 79872
rect 149286 79792 149395 79797
rect 149286 79736 149334 79792
rect 149390 79736 149395 79792
rect 149286 79734 149395 79736
rect 148060 79732 148066 79734
rect 147995 79731 148061 79732
rect 148501 79731 148567 79734
rect 149329 79731 149395 79734
rect 149646 79732 149652 79796
rect 149716 79794 149722 79796
rect 150252 79794 150312 79867
rect 149716 79734 150312 79794
rect 150896 79794 150956 79901
rect 151118 79868 151124 79932
rect 151188 79904 151246 79932
rect 151399 79962 151508 79964
rect 151399 79906 151404 79962
rect 151460 79932 151508 79962
rect 151675 79932 151741 79933
rect 152227 79932 152293 79933
rect 151460 79906 151492 79932
rect 151188 79868 151194 79904
rect 151399 79901 151492 79906
rect 151448 79870 151492 79901
rect 151486 79868 151492 79870
rect 151556 79868 151562 79932
rect 151670 79868 151676 79932
rect 151740 79930 151746 79932
rect 152222 79930 152228 79932
rect 151740 79870 151832 79930
rect 152136 79870 152228 79930
rect 151740 79868 151746 79870
rect 152222 79868 152228 79870
rect 152292 79868 152298 79932
rect 152414 79930 152474 80006
rect 153656 80006 154068 80066
rect 153656 79933 153716 80006
rect 154062 80004 154068 80006
rect 154132 80004 154138 80068
rect 157190 80004 157196 80068
rect 157260 80066 157266 80068
rect 157260 80006 158914 80066
rect 157260 80004 157266 80006
rect 154343 79964 154409 79967
rect 154343 79962 154452 79964
rect 152779 79930 152845 79933
rect 152963 79930 153029 79933
rect 152414 79928 152845 79930
rect 152414 79872 152784 79928
rect 152840 79872 152845 79928
rect 152414 79870 152845 79872
rect 151675 79867 151741 79868
rect 152227 79867 152293 79868
rect 152779 79867 152845 79870
rect 152920 79928 153029 79930
rect 152920 79872 152968 79928
rect 153024 79872 153029 79928
rect 152920 79867 153029 79872
rect 153607 79928 153716 79933
rect 153607 79872 153612 79928
rect 153668 79872 153716 79928
rect 153607 79867 153716 79872
rect 153883 79930 153949 79933
rect 154062 79930 154068 79932
rect 153883 79928 154068 79930
rect 153883 79872 153888 79928
rect 153944 79872 154068 79928
rect 153883 79870 154068 79872
rect 153883 79867 153949 79870
rect 154062 79868 154068 79870
rect 154132 79868 154138 79932
rect 154343 79906 154348 79962
rect 154404 79932 154452 79962
rect 155355 79962 155421 79967
rect 155631 79964 155697 79967
rect 154404 79906 154436 79932
rect 154343 79901 154436 79906
rect 154392 79870 154436 79901
rect 154430 79868 154436 79870
rect 154500 79868 154506 79932
rect 154614 79868 154620 79932
rect 154684 79930 154690 79932
rect 154987 79930 155053 79933
rect 154684 79928 155053 79930
rect 154684 79872 154992 79928
rect 155048 79872 155053 79928
rect 154684 79870 155053 79872
rect 154684 79868 154690 79870
rect 151302 79794 151308 79796
rect 150896 79734 151308 79794
rect 149716 79732 149722 79734
rect 151302 79732 151308 79734
rect 151372 79732 151378 79796
rect 151537 79794 151603 79797
rect 152043 79796 152109 79797
rect 151670 79794 151676 79796
rect 151537 79792 151676 79794
rect 151537 79736 151542 79792
rect 151598 79736 151676 79792
rect 151537 79734 151676 79736
rect 151537 79731 151603 79734
rect 151670 79732 151676 79734
rect 151740 79732 151746 79796
rect 152038 79794 152044 79796
rect 151952 79734 152044 79794
rect 152038 79732 152044 79734
rect 152108 79732 152114 79796
rect 152590 79732 152596 79796
rect 152660 79794 152666 79796
rect 152920 79794 152980 79867
rect 152660 79734 152980 79794
rect 153656 79794 153716 79867
rect 154113 79794 154179 79797
rect 153656 79792 154179 79794
rect 153656 79736 154118 79792
rect 154174 79736 154179 79792
rect 153656 79734 154179 79736
rect 152660 79732 152666 79734
rect 152043 79731 152109 79732
rect 154113 79731 154179 79734
rect 133638 79658 133644 79660
rect 132972 79598 133644 79658
rect 132972 79596 132978 79598
rect 133638 79596 133644 79598
rect 133708 79596 133714 79660
rect 134609 79658 134675 79661
rect 134793 79658 134859 79661
rect 134609 79656 134859 79658
rect 134609 79600 134614 79656
rect 134670 79600 134798 79656
rect 134854 79600 134859 79656
rect 134609 79598 134859 79600
rect 134609 79595 134675 79598
rect 134793 79595 134859 79598
rect 135621 79658 135687 79661
rect 135846 79658 135852 79660
rect 135621 79656 135852 79658
rect 135621 79600 135626 79656
rect 135682 79600 135852 79656
rect 135621 79598 135852 79600
rect 135621 79595 135687 79598
rect 135846 79596 135852 79598
rect 135916 79596 135922 79660
rect 136030 79596 136036 79660
rect 136100 79658 136106 79660
rect 136633 79658 136699 79661
rect 136100 79656 136699 79658
rect 136100 79600 136638 79656
rect 136694 79600 136699 79656
rect 136100 79598 136699 79600
rect 136100 79596 136106 79598
rect 136633 79595 136699 79598
rect 136817 79656 136883 79661
rect 137093 79660 137159 79661
rect 137093 79658 137140 79660
rect 136817 79600 136822 79656
rect 136878 79600 136883 79656
rect 136817 79595 136883 79600
rect 137048 79656 137140 79658
rect 137048 79600 137098 79656
rect 137048 79598 137140 79600
rect 137093 79596 137140 79598
rect 137204 79596 137210 79660
rect 137277 79658 137343 79661
rect 137686 79658 137692 79660
rect 137277 79656 137692 79658
rect 137277 79600 137282 79656
rect 137338 79600 137692 79656
rect 137277 79598 137692 79600
rect 137093 79595 137159 79596
rect 137277 79595 137343 79598
rect 137686 79596 137692 79598
rect 137756 79596 137762 79660
rect 152089 79658 152155 79661
rect 137970 79656 152155 79658
rect 137970 79600 152094 79656
rect 152150 79600 152155 79656
rect 137970 79598 152155 79600
rect 120717 79522 120783 79525
rect 137970 79522 138030 79598
rect 152089 79595 152155 79598
rect 152406 79596 152412 79660
rect 152476 79658 152482 79660
rect 153009 79658 153075 79661
rect 152476 79656 153075 79658
rect 152476 79600 153014 79656
rect 153070 79600 153075 79656
rect 152476 79598 153075 79600
rect 152476 79596 152482 79598
rect 153009 79595 153075 79598
rect 153510 79596 153516 79660
rect 153580 79658 153586 79660
rect 154062 79658 154068 79660
rect 153580 79598 154068 79658
rect 153580 79596 153586 79598
rect 154062 79596 154068 79598
rect 154132 79596 154138 79660
rect 154297 79658 154363 79661
rect 154438 79658 154498 79868
rect 154987 79867 155053 79870
rect 155166 79868 155172 79932
rect 155236 79930 155242 79932
rect 155355 79930 155360 79962
rect 155236 79906 155360 79930
rect 155416 79906 155421 79962
rect 155588 79962 155697 79964
rect 155588 79932 155636 79962
rect 155236 79901 155421 79906
rect 155236 79870 155418 79901
rect 155236 79868 155242 79870
rect 155534 79868 155540 79932
rect 155604 79906 155636 79932
rect 155692 79906 155697 79962
rect 158854 79933 158914 80006
rect 159130 79933 159190 80142
rect 159728 79967 159788 80278
rect 165846 80278 173082 80338
rect 165846 80202 165906 80278
rect 173198 80276 173204 80340
rect 173268 80338 173274 80340
rect 179370 80338 179430 80686
rect 200941 80683 201007 80686
rect 190862 80610 190868 80612
rect 190410 80550 190868 80610
rect 183737 80340 183803 80341
rect 183686 80338 183692 80340
rect 173268 80278 179430 80338
rect 183646 80278 183692 80338
rect 183756 80336 183803 80340
rect 190410 80338 190470 80550
rect 190862 80548 190868 80550
rect 190932 80548 190938 80612
rect 183798 80280 183803 80336
rect 173268 80276 173274 80278
rect 183686 80276 183692 80278
rect 183756 80276 183803 80280
rect 183737 80275 183803 80276
rect 189030 80278 190470 80338
rect 166942 80202 166948 80204
rect 165754 80142 165906 80202
rect 165984 80142 166948 80202
rect 162158 80004 162164 80068
rect 162228 80004 162234 80068
rect 163262 80004 163268 80068
rect 163332 80066 163338 80068
rect 163332 80006 163836 80066
rect 163332 80004 163338 80006
rect 159679 79962 159788 79967
rect 155907 79932 155973 79933
rect 155902 79930 155908 79932
rect 155604 79901 155697 79906
rect 155604 79870 155648 79901
rect 155816 79870 155908 79930
rect 155604 79868 155610 79870
rect 155902 79868 155908 79870
rect 155972 79868 155978 79932
rect 156454 79868 156460 79932
rect 156524 79930 156530 79932
rect 156643 79930 156709 79933
rect 156524 79928 156709 79930
rect 156524 79872 156648 79928
rect 156704 79872 156709 79928
rect 156524 79870 156709 79872
rect 156524 79868 156530 79870
rect 155907 79867 155973 79868
rect 156600 79867 156709 79870
rect 157011 79930 157077 79933
rect 157190 79930 157196 79932
rect 157011 79928 157196 79930
rect 157011 79872 157016 79928
rect 157072 79872 157196 79928
rect 157011 79870 157196 79872
rect 157011 79867 157077 79870
rect 157190 79868 157196 79870
rect 157260 79868 157266 79932
rect 157471 79930 157537 79933
rect 157471 79928 157672 79930
rect 157471 79872 157476 79928
rect 157532 79872 157672 79928
rect 157471 79870 157672 79872
rect 157471 79867 157537 79870
rect 155401 79660 155467 79661
rect 155350 79658 155356 79660
rect 154297 79656 154498 79658
rect 154297 79600 154302 79656
rect 154358 79600 154498 79656
rect 154297 79598 154498 79600
rect 155310 79598 155356 79658
rect 155420 79656 155467 79660
rect 155462 79600 155467 79656
rect 154297 79595 154363 79598
rect 155350 79596 155356 79598
rect 155420 79596 155467 79600
rect 155401 79595 155467 79596
rect 155769 79658 155835 79661
rect 155910 79658 155970 79867
rect 156600 79661 156660 79867
rect 157006 79732 157012 79796
rect 157076 79794 157082 79796
rect 157333 79794 157399 79797
rect 157076 79792 157399 79794
rect 157076 79736 157338 79792
rect 157394 79736 157399 79792
rect 157076 79734 157399 79736
rect 157076 79732 157082 79734
rect 157333 79731 157399 79734
rect 157612 79661 157672 79870
rect 158294 79868 158300 79932
rect 158364 79930 158370 79932
rect 158575 79930 158641 79933
rect 158364 79928 158641 79930
rect 158364 79872 158580 79928
rect 158636 79872 158641 79928
rect 158364 79870 158641 79872
rect 158364 79868 158370 79870
rect 158575 79867 158641 79870
rect 158851 79928 158917 79933
rect 158851 79872 158856 79928
rect 158912 79872 158917 79928
rect 158851 79867 158917 79872
rect 159127 79930 159193 79933
rect 159127 79928 159374 79930
rect 159127 79872 159132 79928
rect 159188 79872 159374 79928
rect 159679 79906 159684 79962
rect 159740 79906 159788 79962
rect 159679 79901 159788 79906
rect 159863 79964 159929 79967
rect 161335 79964 161401 79967
rect 159863 79962 160064 79964
rect 159863 79906 159868 79962
rect 159924 79930 160064 79962
rect 161292 79962 161401 79964
rect 160134 79930 160140 79932
rect 159924 79906 160140 79930
rect 159863 79904 160140 79906
rect 159863 79901 159929 79904
rect 159127 79870 159374 79872
rect 159127 79867 159193 79870
rect 158854 79797 158914 79867
rect 157747 79794 157813 79797
rect 158110 79794 158116 79796
rect 157747 79792 158116 79794
rect 157747 79736 157752 79792
rect 157808 79736 158116 79792
rect 157747 79734 158116 79736
rect 157747 79731 157813 79734
rect 158110 79732 158116 79734
rect 158180 79732 158186 79796
rect 158391 79794 158457 79797
rect 158391 79792 158500 79794
rect 158391 79736 158396 79792
rect 158452 79736 158500 79792
rect 158391 79731 158500 79736
rect 158805 79792 158914 79797
rect 158805 79736 158810 79792
rect 158866 79736 158914 79792
rect 158805 79734 158914 79736
rect 158805 79731 158871 79734
rect 159030 79732 159036 79796
rect 159100 79794 159106 79796
rect 159173 79794 159239 79797
rect 159100 79792 159239 79794
rect 159100 79736 159178 79792
rect 159234 79736 159239 79792
rect 159100 79734 159239 79736
rect 159100 79732 159106 79734
rect 159173 79731 159239 79734
rect 155769 79656 155970 79658
rect 155769 79600 155774 79656
rect 155830 79600 155970 79656
rect 155769 79598 155970 79600
rect 156597 79656 156663 79661
rect 156597 79600 156602 79656
rect 156658 79600 156663 79656
rect 155769 79595 155835 79598
rect 156597 79595 156663 79600
rect 156822 79596 156828 79660
rect 156892 79658 156898 79660
rect 156965 79658 157031 79661
rect 156892 79656 157031 79658
rect 156892 79600 156970 79656
rect 157026 79600 157031 79656
rect 156892 79598 157031 79600
rect 156892 79596 156898 79598
rect 156965 79595 157031 79598
rect 157609 79656 157675 79661
rect 157609 79600 157614 79656
rect 157670 79600 157675 79656
rect 157609 79595 157675 79600
rect 158440 79660 158500 79731
rect 158440 79598 158484 79660
rect 158478 79596 158484 79598
rect 158548 79596 158554 79660
rect 158621 79658 158687 79661
rect 159314 79658 159374 79870
rect 159728 79794 159788 79901
rect 160004 79870 160140 79904
rect 160134 79868 160140 79870
rect 160204 79868 160210 79932
rect 160323 79928 160389 79933
rect 161292 79932 161340 79962
rect 160323 79872 160328 79928
rect 160384 79872 160389 79928
rect 160323 79867 160389 79872
rect 160870 79868 160876 79932
rect 160940 79930 160946 79932
rect 161238 79930 161244 79932
rect 160940 79870 161244 79930
rect 160940 79868 160946 79870
rect 161238 79868 161244 79870
rect 161308 79906 161340 79932
rect 161396 79906 161401 79962
rect 161979 79962 162045 79967
rect 161308 79901 161401 79906
rect 161611 79928 161677 79933
rect 161979 79932 161984 79962
rect 162040 79932 162045 79962
rect 161308 79870 161352 79901
rect 161611 79872 161616 79928
rect 161672 79872 161677 79928
rect 161308 79868 161314 79870
rect 161611 79867 161677 79872
rect 161974 79868 161980 79932
rect 162044 79930 162050 79932
rect 162166 79930 162226 80004
rect 162899 79962 162965 79967
rect 162715 79930 162781 79933
rect 162044 79870 162102 79930
rect 162166 79928 162781 79930
rect 162166 79872 162720 79928
rect 162776 79872 162781 79928
rect 162899 79906 162904 79962
rect 162960 79906 162965 79962
rect 162899 79901 162965 79906
rect 163267 79928 163333 79933
rect 162166 79870 162781 79872
rect 162044 79868 162050 79870
rect 162715 79867 162781 79870
rect 159909 79794 159975 79797
rect 159728 79792 159975 79794
rect 159728 79736 159914 79792
rect 159970 79736 159975 79792
rect 159728 79734 159975 79736
rect 159909 79731 159975 79734
rect 160139 79792 160205 79797
rect 160139 79736 160144 79792
rect 160200 79736 160205 79792
rect 160139 79731 160205 79736
rect 160142 79661 160202 79731
rect 159817 79660 159883 79661
rect 159766 79658 159772 79660
rect 158621 79656 159374 79658
rect 158621 79600 158626 79656
rect 158682 79600 159374 79656
rect 158621 79598 159374 79600
rect 159726 79598 159772 79658
rect 159836 79656 159883 79660
rect 159878 79600 159883 79656
rect 158621 79595 158687 79598
rect 159766 79596 159772 79598
rect 159836 79596 159883 79600
rect 159817 79595 159883 79596
rect 160093 79656 160202 79661
rect 160093 79600 160098 79656
rect 160154 79600 160202 79656
rect 160093 79598 160202 79600
rect 160093 79595 160159 79598
rect 120717 79520 138030 79522
rect 120717 79464 120722 79520
rect 120778 79464 138030 79520
rect 120717 79462 138030 79464
rect 120717 79459 120783 79462
rect 138238 79460 138244 79524
rect 138308 79522 138314 79524
rect 146937 79522 147003 79525
rect 147121 79524 147187 79525
rect 138308 79520 147003 79522
rect 138308 79464 146942 79520
rect 146998 79464 147003 79520
rect 138308 79462 147003 79464
rect 138308 79460 138314 79462
rect 146937 79459 147003 79462
rect 147070 79460 147076 79524
rect 147140 79522 147187 79524
rect 147397 79524 147463 79525
rect 147673 79524 147739 79525
rect 147397 79522 147444 79524
rect 147140 79520 147232 79522
rect 147182 79464 147232 79520
rect 147140 79462 147232 79464
rect 147352 79520 147444 79522
rect 147352 79464 147402 79520
rect 147352 79462 147444 79464
rect 147140 79460 147187 79462
rect 147121 79459 147187 79460
rect 147397 79460 147444 79462
rect 147508 79460 147514 79524
rect 147622 79460 147628 79524
rect 147692 79522 147739 79524
rect 148133 79524 148199 79525
rect 148133 79522 148180 79524
rect 147692 79520 147784 79522
rect 147734 79464 147784 79520
rect 147692 79462 147784 79464
rect 148088 79520 148180 79522
rect 148244 79522 148250 79524
rect 148542 79522 148548 79524
rect 148088 79464 148138 79520
rect 148088 79462 148180 79464
rect 147692 79460 147739 79462
rect 147397 79459 147463 79460
rect 147673 79459 147739 79460
rect 148133 79460 148180 79462
rect 148244 79462 148548 79522
rect 148244 79460 148250 79462
rect 148542 79460 148548 79462
rect 148612 79460 148618 79524
rect 149278 79460 149284 79524
rect 149348 79522 149354 79524
rect 153653 79522 153719 79525
rect 149348 79520 153719 79522
rect 149348 79464 153658 79520
rect 153714 79464 153719 79520
rect 149348 79462 153719 79464
rect 149348 79460 149354 79462
rect 148133 79459 148199 79460
rect 153653 79459 153719 79462
rect 153878 79460 153884 79524
rect 153948 79522 153954 79524
rect 154389 79522 154455 79525
rect 154573 79522 154639 79525
rect 153948 79520 154639 79522
rect 153948 79464 154394 79520
rect 154450 79464 154578 79520
rect 154634 79464 154639 79520
rect 153948 79462 154639 79464
rect 153948 79460 153954 79462
rect 154389 79459 154455 79462
rect 154573 79459 154639 79462
rect 155125 79522 155191 79525
rect 159214 79522 159220 79524
rect 155125 79520 159220 79522
rect 155125 79464 155130 79520
rect 155186 79464 159220 79520
rect 155125 79462 159220 79464
rect 155125 79459 155191 79462
rect 159214 79460 159220 79462
rect 159284 79460 159290 79524
rect 160326 79522 160386 79867
rect 160599 79828 160665 79831
rect 160556 79826 160665 79828
rect 160556 79770 160604 79826
rect 160660 79794 160665 79826
rect 160870 79794 160876 79796
rect 160660 79770 160876 79794
rect 160556 79734 160876 79770
rect 160870 79732 160876 79734
rect 160940 79732 160946 79796
rect 161422 79732 161428 79796
rect 161492 79794 161498 79796
rect 161614 79794 161674 79867
rect 162347 79794 162413 79797
rect 161492 79734 161674 79794
rect 161492 79732 161498 79734
rect 160502 79596 160508 79660
rect 160572 79658 160578 79660
rect 161197 79658 161263 79661
rect 160572 79656 161263 79658
rect 160572 79600 161202 79656
rect 161258 79600 161263 79656
rect 160572 79598 161263 79600
rect 160572 79596 160578 79598
rect 161197 79595 161263 79598
rect 160461 79522 160527 79525
rect 160326 79520 160527 79522
rect 160326 79464 160466 79520
rect 160522 79464 160527 79520
rect 160326 79462 160527 79464
rect 160461 79459 160527 79462
rect 160737 79522 160803 79525
rect 161054 79522 161060 79524
rect 160737 79520 161060 79522
rect 160737 79464 160742 79520
rect 160798 79464 161060 79520
rect 160737 79462 161060 79464
rect 160737 79459 160803 79462
rect 161054 79460 161060 79462
rect 161124 79460 161130 79524
rect 161614 79522 161674 79734
rect 162212 79792 162413 79794
rect 162212 79736 162352 79792
rect 162408 79736 162413 79792
rect 162212 79734 162413 79736
rect 162212 79661 162272 79734
rect 162347 79731 162413 79734
rect 162902 79661 162962 79901
rect 163267 79872 163272 79928
rect 163328 79872 163333 79928
rect 163267 79867 163333 79872
rect 163446 79868 163452 79932
rect 163516 79930 163522 79932
rect 163635 79930 163701 79933
rect 163516 79928 163701 79930
rect 163516 79872 163640 79928
rect 163696 79872 163701 79928
rect 163516 79870 163701 79872
rect 163776 79930 163836 80006
rect 165754 79967 165814 80142
rect 165984 79967 166044 80142
rect 166942 80140 166948 80142
rect 167012 80140 167018 80204
rect 169150 80202 169156 80204
rect 168606 80142 169156 80202
rect 168606 79967 168666 80142
rect 169150 80140 169156 80142
rect 169220 80140 169226 80204
rect 169886 80140 169892 80204
rect 169956 80202 169962 80204
rect 189030 80202 189090 80278
rect 169956 80142 171058 80202
rect 169956 80140 169962 80142
rect 170806 80066 170812 80068
rect 170446 80006 170812 80066
rect 165751 79962 165817 79967
rect 164095 79930 164161 79933
rect 163776 79928 164161 79930
rect 163776 79872 164100 79928
rect 164156 79872 164161 79928
rect 163776 79870 164161 79872
rect 163516 79868 163522 79870
rect 163635 79867 163701 79870
rect 164095 79867 164161 79870
rect 164371 79930 164437 79933
rect 164550 79930 164556 79932
rect 164371 79928 164556 79930
rect 164371 79872 164376 79928
rect 164432 79872 164556 79928
rect 164371 79870 164556 79872
rect 164371 79867 164437 79870
rect 164550 79868 164556 79870
rect 164620 79868 164626 79932
rect 164734 79868 164740 79932
rect 164804 79930 164810 79932
rect 164923 79930 164989 79933
rect 164804 79928 164989 79930
rect 164804 79872 164928 79928
rect 164984 79872 164989 79928
rect 164804 79870 164989 79872
rect 164804 79868 164810 79870
rect 164923 79867 164989 79870
rect 165286 79868 165292 79932
rect 165356 79930 165362 79932
rect 165475 79930 165541 79933
rect 165356 79928 165541 79930
rect 165356 79872 165480 79928
rect 165536 79872 165541 79928
rect 165751 79906 165756 79962
rect 165812 79906 165817 79962
rect 165751 79901 165817 79906
rect 165935 79962 166044 79967
rect 165935 79906 165940 79962
rect 165996 79906 166044 79962
rect 168235 79964 168301 79967
rect 168235 79962 168358 79964
rect 165935 79904 166044 79906
rect 165935 79901 166001 79904
rect 165356 79870 165541 79872
rect 165356 79868 165362 79870
rect 165475 79867 165541 79870
rect 166206 79868 166212 79932
rect 166276 79930 166282 79932
rect 166855 79930 166921 79933
rect 166276 79928 166921 79930
rect 166276 79872 166860 79928
rect 166916 79872 166921 79928
rect 166276 79870 166921 79872
rect 166276 79868 166282 79870
rect 166855 79867 166921 79870
rect 167407 79930 167473 79933
rect 168235 79932 168240 79962
rect 168296 79932 168358 79962
rect 168603 79962 168669 79967
rect 167678 79930 167684 79932
rect 167407 79928 167684 79930
rect 167407 79872 167412 79928
rect 167468 79872 167684 79928
rect 167407 79870 167684 79872
rect 167407 79867 167473 79870
rect 167678 79868 167684 79870
rect 167748 79868 167754 79932
rect 168230 79868 168236 79932
rect 168300 79904 168358 79932
rect 168419 79928 168485 79933
rect 168300 79868 168306 79904
rect 168419 79872 168424 79928
rect 168480 79872 168485 79928
rect 168603 79906 168608 79962
rect 168664 79906 168669 79962
rect 169707 79962 169773 79967
rect 168603 79901 168669 79906
rect 168419 79867 168485 79872
rect 168782 79868 168788 79932
rect 168852 79930 168858 79932
rect 169063 79930 169129 79933
rect 169707 79932 169712 79962
rect 169768 79932 169773 79962
rect 170446 79933 170506 80006
rect 170806 80004 170812 80006
rect 170876 80004 170882 80068
rect 170998 79967 171058 80142
rect 173942 80142 189090 80202
rect 173750 80066 173756 80068
rect 172746 80006 173756 80066
rect 170995 79962 171061 79967
rect 168852 79928 169129 79930
rect 168852 79872 169068 79928
rect 169124 79872 169129 79928
rect 168852 79870 169129 79872
rect 168852 79868 168858 79870
rect 169063 79867 169129 79870
rect 169702 79868 169708 79932
rect 169772 79930 169778 79932
rect 169772 79870 169830 79930
rect 170443 79928 170509 79933
rect 170443 79872 170448 79928
rect 170504 79872 170509 79928
rect 169772 79868 169778 79870
rect 170443 79867 170509 79872
rect 170719 79928 170785 79933
rect 170719 79872 170724 79928
rect 170780 79872 170785 79928
rect 170995 79906 171000 79962
rect 171056 79906 171061 79962
rect 171363 79962 171429 79967
rect 172007 79964 172073 79967
rect 171363 79932 171368 79962
rect 171424 79932 171429 79962
rect 171964 79962 172073 79964
rect 170995 79901 171061 79906
rect 170719 79867 170785 79872
rect 171358 79868 171364 79932
rect 171428 79930 171434 79932
rect 171547 79930 171613 79933
rect 171964 79932 172012 79962
rect 171726 79930 171732 79932
rect 171428 79870 171486 79930
rect 171547 79928 171732 79930
rect 171547 79872 171552 79928
rect 171608 79872 171732 79928
rect 171547 79870 171732 79872
rect 171428 79868 171434 79870
rect 171547 79867 171613 79870
rect 171726 79868 171732 79870
rect 171796 79868 171802 79932
rect 171910 79868 171916 79932
rect 171980 79906 172012 79932
rect 172068 79906 172073 79962
rect 171980 79901 172073 79906
rect 172283 79962 172349 79967
rect 172283 79906 172288 79962
rect 172344 79930 172349 79962
rect 172746 79933 172806 80006
rect 173750 80004 173756 80006
rect 173820 80004 173826 80068
rect 173942 79933 174002 80142
rect 197670 80004 197676 80068
rect 197740 80066 197746 80068
rect 197997 80066 198063 80069
rect 197740 80064 198063 80066
rect 197740 80008 198002 80064
rect 198058 80008 198063 80064
rect 197740 80006 198063 80008
rect 197740 80004 197746 80006
rect 197997 80003 198063 80006
rect 176699 79962 176765 79967
rect 172462 79930 172468 79932
rect 172344 79906 172468 79930
rect 172283 79901 172468 79906
rect 171980 79870 172024 79901
rect 172286 79870 172468 79901
rect 171980 79868 171986 79870
rect 172462 79868 172468 79870
rect 172532 79868 172538 79932
rect 172743 79928 172809 79933
rect 172743 79872 172748 79928
rect 172804 79872 172809 79928
rect 172743 79867 172809 79872
rect 173939 79928 174005 79933
rect 173939 79872 173944 79928
rect 174000 79872 174005 79928
rect 173939 79867 174005 79872
rect 174123 79928 174189 79933
rect 174123 79872 174128 79928
rect 174184 79872 174189 79928
rect 174123 79867 174189 79872
rect 174302 79868 174308 79932
rect 174372 79930 174378 79932
rect 174583 79930 174649 79933
rect 174372 79928 174649 79930
rect 174372 79872 174588 79928
rect 174644 79872 174649 79928
rect 174372 79870 174649 79872
rect 174372 79868 174378 79870
rect 174583 79867 174649 79870
rect 174859 79930 174925 79933
rect 175038 79930 175044 79932
rect 174859 79928 175044 79930
rect 174859 79872 174864 79928
rect 174920 79872 175044 79928
rect 174859 79870 175044 79872
rect 174859 79867 174925 79870
rect 175038 79868 175044 79870
rect 175108 79868 175114 79932
rect 175227 79928 175293 79933
rect 175411 79932 175477 79933
rect 175227 79872 175232 79928
rect 175288 79872 175293 79928
rect 175227 79867 175293 79872
rect 175406 79868 175412 79932
rect 175476 79930 175482 79932
rect 175476 79870 175568 79930
rect 175476 79868 175482 79870
rect 175774 79868 175780 79932
rect 175844 79930 175850 79932
rect 175963 79930 176029 79933
rect 175844 79928 176029 79930
rect 175844 79872 175968 79928
rect 176024 79872 176029 79928
rect 175844 79870 176029 79872
rect 175844 79868 175850 79870
rect 175411 79867 175477 79868
rect 175963 79867 176029 79870
rect 176142 79868 176148 79932
rect 176212 79930 176218 79932
rect 176515 79930 176581 79933
rect 176212 79928 176581 79930
rect 176212 79872 176520 79928
rect 176576 79872 176581 79928
rect 176699 79906 176704 79962
rect 176760 79906 176765 79962
rect 177343 79962 177409 79967
rect 176699 79901 176765 79906
rect 176212 79870 176581 79872
rect 176212 79868 176218 79870
rect 176515 79867 176581 79870
rect 163270 79794 163330 79867
rect 165478 79797 165538 79867
rect 163998 79794 164004 79796
rect 163270 79734 164004 79794
rect 163998 79732 164004 79734
rect 164068 79732 164074 79796
rect 165429 79792 165538 79797
rect 166027 79796 166093 79797
rect 166022 79794 166028 79796
rect 165429 79736 165434 79792
rect 165490 79736 165538 79792
rect 165429 79734 165538 79736
rect 165936 79734 166028 79794
rect 165429 79731 165495 79734
rect 166022 79732 166028 79734
rect 166092 79732 166098 79796
rect 166390 79732 166396 79796
rect 166460 79794 166466 79796
rect 166579 79794 166645 79797
rect 166460 79792 166645 79794
rect 166460 79736 166584 79792
rect 166640 79736 166645 79792
rect 166460 79734 166645 79736
rect 166460 79732 166466 79734
rect 166027 79731 166093 79732
rect 166579 79731 166645 79734
rect 167494 79732 167500 79796
rect 167564 79794 167570 79796
rect 168097 79794 168163 79797
rect 167564 79792 168163 79794
rect 167564 79736 168102 79792
rect 168158 79736 168163 79792
rect 167564 79734 168163 79736
rect 168422 79794 168482 79867
rect 169334 79794 169340 79796
rect 168422 79734 169340 79794
rect 167564 79732 167570 79734
rect 168097 79731 168163 79734
rect 169334 79732 169340 79734
rect 169404 79732 169410 79796
rect 170075 79794 170141 79797
rect 170722 79794 170782 79867
rect 174126 79797 174186 79867
rect 174862 79797 174922 79867
rect 170990 79794 170996 79796
rect 170075 79792 170644 79794
rect 170075 79736 170080 79792
rect 170136 79736 170644 79792
rect 170075 79734 170644 79736
rect 170722 79734 170996 79794
rect 170075 79731 170141 79734
rect 161841 79660 161907 79661
rect 161790 79596 161796 79660
rect 161860 79658 161907 79660
rect 161860 79656 161952 79658
rect 161902 79600 161952 79656
rect 161860 79598 161952 79600
rect 162209 79656 162275 79661
rect 162209 79600 162214 79656
rect 162270 79600 162275 79656
rect 161860 79596 161907 79598
rect 161841 79595 161907 79596
rect 162209 79595 162275 79600
rect 162342 79596 162348 79660
rect 162412 79658 162418 79660
rect 162577 79658 162643 79661
rect 162412 79656 162643 79658
rect 162412 79600 162582 79656
rect 162638 79600 162643 79656
rect 162412 79598 162643 79600
rect 162902 79656 163011 79661
rect 162902 79600 162950 79656
rect 163006 79600 163011 79656
rect 162902 79598 163011 79600
rect 162412 79596 162418 79598
rect 162577 79595 162643 79598
rect 162945 79595 163011 79598
rect 163630 79596 163636 79660
rect 163700 79658 163706 79660
rect 163773 79658 163839 79661
rect 163700 79656 163839 79658
rect 163700 79600 163778 79656
rect 163834 79600 163839 79656
rect 163700 79598 163839 79600
rect 163700 79596 163706 79598
rect 163773 79595 163839 79598
rect 164918 79596 164924 79660
rect 164988 79658 164994 79660
rect 165061 79658 165127 79661
rect 164988 79656 165127 79658
rect 164988 79600 165066 79656
rect 165122 79600 165127 79656
rect 164988 79598 165127 79600
rect 164988 79596 164994 79598
rect 165061 79595 165127 79598
rect 166809 79658 166875 79661
rect 166993 79658 167059 79661
rect 166809 79656 167059 79658
rect 166809 79600 166814 79656
rect 166870 79600 166998 79656
rect 167054 79600 167059 79656
rect 166809 79598 167059 79600
rect 166809 79595 166875 79598
rect 166993 79595 167059 79598
rect 167678 79596 167684 79660
rect 167748 79658 167754 79660
rect 167913 79658 167979 79661
rect 167748 79656 167979 79658
rect 167748 79600 167918 79656
rect 167974 79600 167979 79656
rect 167748 79598 167979 79600
rect 167748 79596 167754 79598
rect 167913 79595 167979 79598
rect 168966 79596 168972 79660
rect 169036 79658 169042 79660
rect 169293 79658 169359 79661
rect 169036 79656 169359 79658
rect 169036 79600 169298 79656
rect 169354 79600 169359 79656
rect 169036 79598 169359 79600
rect 169036 79596 169042 79598
rect 169293 79595 169359 79598
rect 169477 79660 169543 79661
rect 169477 79656 169524 79660
rect 169588 79658 169594 79660
rect 169477 79600 169482 79656
rect 169477 79596 169524 79600
rect 169588 79598 169634 79658
rect 169588 79596 169594 79598
rect 170070 79596 170076 79660
rect 170140 79658 170146 79660
rect 170213 79658 170279 79661
rect 170140 79656 170279 79658
rect 170140 79600 170218 79656
rect 170274 79600 170279 79656
rect 170140 79598 170279 79600
rect 170584 79660 170644 79734
rect 170952 79732 170996 79734
rect 171060 79732 171066 79796
rect 171542 79732 171548 79796
rect 171612 79794 171618 79796
rect 171777 79794 171843 79797
rect 171612 79792 171843 79794
rect 171612 79736 171782 79792
rect 171838 79736 171843 79792
rect 171612 79734 171843 79736
rect 171612 79732 171618 79734
rect 170952 79661 171012 79732
rect 171777 79731 171843 79734
rect 172053 79796 172119 79797
rect 172053 79792 172100 79796
rect 172164 79794 172170 79796
rect 172053 79736 172058 79792
rect 172053 79732 172100 79736
rect 172164 79734 172210 79794
rect 172164 79732 172170 79734
rect 172830 79732 172836 79796
rect 172900 79794 172906 79796
rect 173203 79794 173269 79797
rect 172900 79792 173269 79794
rect 172900 79736 173208 79792
rect 173264 79736 173269 79792
rect 172900 79734 173269 79736
rect 172900 79732 172906 79734
rect 172053 79731 172119 79732
rect 173203 79731 173269 79734
rect 174077 79792 174186 79797
rect 174077 79736 174082 79792
rect 174138 79736 174186 79792
rect 174077 79734 174186 79736
rect 174353 79794 174419 79797
rect 174491 79794 174557 79797
rect 174353 79792 174557 79794
rect 174353 79736 174358 79792
rect 174414 79736 174496 79792
rect 174552 79736 174557 79792
rect 174353 79734 174557 79736
rect 174862 79792 174971 79797
rect 174862 79736 174910 79792
rect 174966 79736 174971 79792
rect 174862 79734 174971 79736
rect 174077 79731 174143 79734
rect 174353 79731 174419 79734
rect 174491 79731 174557 79734
rect 174905 79731 174971 79734
rect 175038 79732 175044 79796
rect 175108 79794 175114 79796
rect 175230 79794 175290 79867
rect 175917 79796 175983 79797
rect 176147 79796 176213 79797
rect 175912 79794 175918 79796
rect 175108 79734 175290 79794
rect 175826 79734 175918 79794
rect 175108 79732 175114 79734
rect 175912 79732 175918 79734
rect 175982 79732 175988 79796
rect 176142 79794 176148 79796
rect 176056 79734 176148 79794
rect 176142 79732 176148 79734
rect 176212 79732 176218 79796
rect 176285 79794 176351 79797
rect 176510 79794 176516 79796
rect 176285 79792 176516 79794
rect 176285 79736 176290 79792
rect 176346 79736 176516 79792
rect 176285 79734 176516 79736
rect 175917 79731 175983 79732
rect 176147 79731 176213 79732
rect 176285 79731 176351 79734
rect 176510 79732 176516 79734
rect 176580 79732 176586 79796
rect 170584 79598 170628 79660
rect 170140 79596 170146 79598
rect 169477 79595 169543 79596
rect 170213 79595 170279 79598
rect 170622 79596 170628 79598
rect 170692 79596 170698 79660
rect 170949 79656 171015 79661
rect 176101 79658 176167 79661
rect 170949 79600 170954 79656
rect 171010 79600 171015 79656
rect 170949 79595 171015 79600
rect 171550 79656 176167 79658
rect 171550 79600 176106 79656
rect 176162 79600 176167 79656
rect 171550 79598 176167 79600
rect 176702 79658 176762 79901
rect 176878 79868 176884 79932
rect 176948 79930 176954 79932
rect 177343 79930 177348 79962
rect 176948 79906 177348 79930
rect 177404 79906 177409 79962
rect 177573 79932 177639 79933
rect 177573 79930 177620 79932
rect 176948 79901 177409 79906
rect 177528 79928 177620 79930
rect 176948 79870 177406 79901
rect 177528 79872 177578 79928
rect 177528 79870 177620 79872
rect 176948 79868 176954 79870
rect 177573 79868 177620 79870
rect 177684 79868 177690 79932
rect 177849 79930 177915 79933
rect 180885 79930 180951 79933
rect 177849 79928 180951 79930
rect 177849 79872 177854 79928
rect 177910 79872 180890 79928
rect 180946 79872 180951 79928
rect 177849 79870 180951 79872
rect 177573 79867 177639 79868
rect 177849 79867 177915 79870
rect 180885 79867 180951 79870
rect 197629 79930 197695 79933
rect 197854 79930 197860 79932
rect 197629 79928 197860 79930
rect 197629 79872 197634 79928
rect 197690 79872 197860 79928
rect 197629 79870 197860 79872
rect 197629 79867 197695 79870
rect 197854 79868 197860 79870
rect 197924 79868 197930 79932
rect 177062 79732 177068 79796
rect 177132 79794 177138 79796
rect 177481 79794 177547 79797
rect 177132 79792 177547 79794
rect 177132 79736 177486 79792
rect 177542 79736 177547 79792
rect 177132 79734 177547 79736
rect 177132 79732 177138 79734
rect 177481 79731 177547 79734
rect 177062 79658 177068 79660
rect 176702 79598 177068 79658
rect 161933 79522 161999 79525
rect 161614 79520 161999 79522
rect 161614 79464 161938 79520
rect 161994 79464 161999 79520
rect 161614 79462 161999 79464
rect 161933 79459 161999 79462
rect 162393 79522 162459 79525
rect 162526 79522 162532 79524
rect 162393 79520 162532 79522
rect 162393 79464 162398 79520
rect 162454 79464 162532 79520
rect 162393 79462 162532 79464
rect 162393 79459 162459 79462
rect 162526 79460 162532 79462
rect 162596 79522 162602 79524
rect 162669 79522 162735 79525
rect 162596 79520 162735 79522
rect 162596 79464 162674 79520
rect 162730 79464 162735 79520
rect 162596 79462 162735 79464
rect 162596 79460 162602 79462
rect 162669 79459 162735 79462
rect 162894 79460 162900 79524
rect 162964 79522 162970 79524
rect 163589 79522 163655 79525
rect 171550 79522 171610 79598
rect 176101 79595 176167 79598
rect 177062 79596 177068 79598
rect 177132 79596 177138 79660
rect 177297 79658 177363 79661
rect 177852 79658 177912 79867
rect 178217 79796 178283 79797
rect 178166 79794 178172 79796
rect 178126 79734 178172 79794
rect 178236 79792 178283 79796
rect 178278 79736 178283 79792
rect 178166 79732 178172 79734
rect 178236 79732 178283 79736
rect 178217 79731 178283 79732
rect 177297 79656 177912 79658
rect 177297 79600 177302 79656
rect 177358 79600 177912 79656
rect 177297 79598 177912 79600
rect 177297 79595 177363 79598
rect 178534 79596 178540 79660
rect 178604 79658 178610 79660
rect 180057 79658 180123 79661
rect 178604 79656 180123 79658
rect 178604 79600 180062 79656
rect 180118 79600 180123 79656
rect 178604 79598 180123 79600
rect 178604 79596 178610 79598
rect 180057 79595 180123 79598
rect 382273 79522 382339 79525
rect 162964 79520 171610 79522
rect 162964 79464 163594 79520
rect 163650 79464 171610 79520
rect 162964 79462 171610 79464
rect 171688 79520 382339 79522
rect 171688 79464 382278 79520
rect 382334 79464 382339 79520
rect 171688 79462 382339 79464
rect 162964 79460 162970 79462
rect 163589 79459 163655 79462
rect 132350 79324 132356 79388
rect 132420 79386 132426 79388
rect 150709 79386 150775 79389
rect 152825 79388 152891 79389
rect 152774 79386 152780 79388
rect 132420 79384 150775 79386
rect 132420 79328 150714 79384
rect 150770 79328 150775 79384
rect 132420 79326 150775 79328
rect 152734 79326 152780 79386
rect 152844 79384 152891 79388
rect 152886 79328 152891 79384
rect 132420 79324 132426 79326
rect 150709 79323 150775 79326
rect 152774 79324 152780 79326
rect 152844 79324 152891 79328
rect 153694 79324 153700 79388
rect 153764 79386 153770 79388
rect 153837 79386 153903 79389
rect 153764 79384 153903 79386
rect 153764 79328 153842 79384
rect 153898 79328 153903 79384
rect 153764 79326 153903 79328
rect 153764 79324 153770 79326
rect 152825 79323 152891 79324
rect 153837 79323 153903 79326
rect 154798 79324 154804 79388
rect 154868 79386 154874 79388
rect 155401 79386 155467 79389
rect 154868 79384 155467 79386
rect 154868 79328 155406 79384
rect 155462 79328 155467 79384
rect 154868 79326 155467 79328
rect 154868 79324 154874 79326
rect 155401 79323 155467 79326
rect 155677 79388 155743 79389
rect 155677 79384 155724 79388
rect 155788 79386 155794 79388
rect 157057 79386 157123 79389
rect 157742 79386 157748 79388
rect 155677 79328 155682 79384
rect 155677 79324 155724 79328
rect 155788 79326 155834 79386
rect 157057 79384 157748 79386
rect 157057 79328 157062 79384
rect 157118 79328 157748 79384
rect 157057 79326 157748 79328
rect 155788 79324 155794 79326
rect 155677 79323 155743 79324
rect 157057 79323 157123 79326
rect 157742 79324 157748 79326
rect 157812 79324 157818 79388
rect 157926 79324 157932 79388
rect 157996 79386 158002 79388
rect 158253 79386 158319 79389
rect 157996 79384 158319 79386
rect 157996 79328 158258 79384
rect 158314 79328 158319 79384
rect 157996 79326 158319 79328
rect 157996 79324 158002 79326
rect 158253 79323 158319 79326
rect 161606 79324 161612 79388
rect 161676 79386 161682 79388
rect 162117 79386 162183 79389
rect 171688 79386 171748 79462
rect 382273 79459 382339 79462
rect 161676 79384 171748 79386
rect 161676 79328 162122 79384
rect 162178 79328 171748 79384
rect 161676 79326 171748 79328
rect 171961 79386 172027 79389
rect 172329 79388 172395 79389
rect 171961 79384 172208 79386
rect 171961 79328 171966 79384
rect 172022 79328 172208 79384
rect 171961 79326 172208 79328
rect 161676 79324 161682 79326
rect 162117 79323 162183 79326
rect 171961 79323 172027 79326
rect 125358 79188 125364 79252
rect 125428 79250 125434 79252
rect 145281 79250 145347 79253
rect 125428 79248 145347 79250
rect 125428 79192 145286 79248
rect 145342 79192 145347 79248
rect 125428 79190 145347 79192
rect 125428 79188 125434 79190
rect 145281 79187 145347 79190
rect 148910 79188 148916 79252
rect 148980 79250 148986 79252
rect 148980 79190 151922 79250
rect 148980 79188 148986 79190
rect 129590 79052 129596 79116
rect 129660 79114 129666 79116
rect 150157 79114 150223 79117
rect 129660 79112 150223 79114
rect 129660 79056 150162 79112
rect 150218 79056 150223 79112
rect 129660 79054 150223 79056
rect 129660 79052 129666 79054
rect 150157 79051 150223 79054
rect 150801 79114 150867 79117
rect 151353 79116 151419 79117
rect 151118 79114 151124 79116
rect 150801 79112 151124 79114
rect 150801 79056 150806 79112
rect 150862 79056 151124 79112
rect 150801 79054 151124 79056
rect 150801 79051 150867 79054
rect 151118 79052 151124 79054
rect 151188 79052 151194 79116
rect 151302 79052 151308 79116
rect 151372 79114 151419 79116
rect 151862 79114 151922 79190
rect 152038 79188 152044 79252
rect 152108 79250 152114 79252
rect 164233 79250 164299 79253
rect 152108 79248 164299 79250
rect 152108 79192 164238 79248
rect 164294 79192 164299 79248
rect 152108 79190 164299 79192
rect 152108 79188 152114 79190
rect 164233 79187 164299 79190
rect 164734 79188 164740 79252
rect 164804 79250 164810 79252
rect 165153 79250 165219 79253
rect 164804 79248 165219 79250
rect 164804 79192 165158 79248
rect 165214 79192 165219 79248
rect 164804 79190 165219 79192
rect 164804 79188 164810 79190
rect 165153 79187 165219 79190
rect 165286 79188 165292 79252
rect 165356 79250 165362 79252
rect 165521 79250 165587 79253
rect 165356 79248 165587 79250
rect 165356 79192 165526 79248
rect 165582 79192 165587 79248
rect 165356 79190 165587 79192
rect 165356 79188 165362 79190
rect 165521 79187 165587 79190
rect 165797 79250 165863 79253
rect 167269 79252 167335 79253
rect 168189 79252 168255 79253
rect 166574 79250 166580 79252
rect 165797 79248 166580 79250
rect 165797 79192 165802 79248
rect 165858 79192 166580 79248
rect 165797 79190 166580 79192
rect 165797 79187 165863 79190
rect 166574 79188 166580 79190
rect 166644 79188 166650 79252
rect 167269 79250 167316 79252
rect 167224 79248 167316 79250
rect 167380 79250 167386 79252
rect 168046 79250 168052 79252
rect 167224 79192 167274 79248
rect 167224 79190 167316 79192
rect 167269 79188 167316 79190
rect 167380 79190 168052 79250
rect 167380 79188 167386 79190
rect 168046 79188 168052 79190
rect 168116 79188 168122 79252
rect 168189 79248 168236 79252
rect 168300 79250 168306 79252
rect 168189 79192 168194 79248
rect 168189 79188 168236 79192
rect 168300 79190 168346 79250
rect 168300 79188 168306 79190
rect 168598 79188 168604 79252
rect 168668 79250 168674 79252
rect 169661 79250 169727 79253
rect 168668 79248 169727 79250
rect 168668 79192 169666 79248
rect 169722 79192 169727 79248
rect 168668 79190 169727 79192
rect 168668 79188 168674 79190
rect 167269 79187 167335 79188
rect 168189 79187 168255 79188
rect 169661 79187 169727 79190
rect 171726 79188 171732 79252
rect 171796 79250 171802 79252
rect 171961 79250 172027 79253
rect 171796 79248 172027 79250
rect 171796 79192 171966 79248
rect 172022 79192 172027 79248
rect 171796 79190 172027 79192
rect 172148 79250 172208 79326
rect 172278 79324 172284 79388
rect 172348 79386 172395 79388
rect 172973 79388 173039 79389
rect 174445 79388 174511 79389
rect 172973 79386 173020 79388
rect 172348 79384 172440 79386
rect 172390 79328 172440 79384
rect 172348 79326 172440 79328
rect 172928 79384 173020 79386
rect 172928 79328 172978 79384
rect 172928 79326 173020 79328
rect 172348 79324 172395 79326
rect 172329 79323 172395 79324
rect 172973 79324 173020 79326
rect 173084 79324 173090 79388
rect 174445 79386 174492 79388
rect 174400 79384 174492 79386
rect 174400 79328 174450 79384
rect 174400 79326 174492 79328
rect 174445 79324 174492 79326
rect 174556 79324 174562 79388
rect 175733 79386 175799 79389
rect 176142 79386 176148 79388
rect 175733 79384 176148 79386
rect 175733 79328 175738 79384
rect 175794 79328 176148 79384
rect 175733 79326 176148 79328
rect 172973 79323 173039 79324
rect 174445 79323 174511 79324
rect 175733 79323 175799 79326
rect 176142 79324 176148 79326
rect 176212 79324 176218 79388
rect 176653 79386 176719 79389
rect 177246 79386 177252 79388
rect 176653 79384 177252 79386
rect 176653 79328 176658 79384
rect 176714 79328 177252 79384
rect 176653 79326 177252 79328
rect 176653 79323 176719 79326
rect 177246 79324 177252 79326
rect 177316 79324 177322 79388
rect 180885 79386 180951 79389
rect 191046 79386 191052 79388
rect 180885 79384 191052 79386
rect 180885 79328 180890 79384
rect 180946 79328 191052 79384
rect 180885 79326 191052 79328
rect 180885 79323 180951 79326
rect 191046 79324 191052 79326
rect 191116 79324 191122 79388
rect 172278 79250 172284 79252
rect 172148 79190 172284 79250
rect 171796 79188 171802 79190
rect 171961 79187 172027 79190
rect 172278 79188 172284 79190
rect 172348 79188 172354 79252
rect 173249 79250 173315 79253
rect 175641 79250 175707 79253
rect 173249 79248 175707 79250
rect 173249 79192 173254 79248
rect 173310 79192 175646 79248
rect 175702 79192 175707 79248
rect 173249 79190 175707 79192
rect 173249 79187 173315 79190
rect 175641 79187 175707 79190
rect 175917 79250 175983 79253
rect 178677 79250 178743 79253
rect 189206 79250 189212 79252
rect 175917 79248 189212 79250
rect 175917 79192 175922 79248
rect 175978 79192 178682 79248
rect 178738 79192 189212 79248
rect 175917 79190 189212 79192
rect 175917 79187 175983 79190
rect 178677 79187 178743 79190
rect 189206 79188 189212 79190
rect 189276 79188 189282 79252
rect 160369 79114 160435 79117
rect 151372 79112 151464 79114
rect 151414 79056 151464 79112
rect 151372 79054 151464 79056
rect 151862 79112 160435 79114
rect 151862 79056 160374 79112
rect 160430 79056 160435 79112
rect 151862 79054 160435 79056
rect 151372 79052 151419 79054
rect 151353 79051 151419 79052
rect 160369 79051 160435 79054
rect 165613 79114 165679 79117
rect 166574 79114 166580 79116
rect 165613 79112 166580 79114
rect 165613 79056 165618 79112
rect 165674 79056 166580 79112
rect 165613 79054 166580 79056
rect 165613 79051 165679 79054
rect 166574 79052 166580 79054
rect 166644 79052 166650 79116
rect 168373 79114 168439 79117
rect 190494 79114 190500 79116
rect 168373 79112 190500 79114
rect 168373 79056 168378 79112
rect 168434 79056 190500 79112
rect 168373 79054 190500 79056
rect 168373 79051 168439 79054
rect 190494 79052 190500 79054
rect 190564 79052 190570 79116
rect 139209 78980 139275 78981
rect 122598 78916 122604 78980
rect 122668 78978 122674 78980
rect 138054 78978 138060 78980
rect 122668 78918 138060 78978
rect 122668 78916 122674 78918
rect 138054 78916 138060 78918
rect 138124 78916 138130 78980
rect 139158 78916 139164 78980
rect 139228 78978 139275 78980
rect 139577 78978 139643 78981
rect 140630 78978 140636 78980
rect 139228 78976 139320 78978
rect 139270 78920 139320 78976
rect 139228 78918 139320 78920
rect 139577 78976 140636 78978
rect 139577 78920 139582 78976
rect 139638 78920 140636 78976
rect 139577 78918 140636 78920
rect 139228 78916 139275 78918
rect 139209 78915 139275 78916
rect 139577 78915 139643 78918
rect 140630 78916 140636 78918
rect 140700 78916 140706 78980
rect 141141 78978 141207 78981
rect 142429 78980 142495 78981
rect 141366 78978 141372 78980
rect 141141 78976 141372 78978
rect 141141 78920 141146 78976
rect 141202 78920 141372 78976
rect 141141 78918 141372 78920
rect 141141 78915 141207 78918
rect 141366 78916 141372 78918
rect 141436 78916 141442 78980
rect 142429 78978 142476 78980
rect 142384 78976 142476 78978
rect 142384 78920 142434 78976
rect 142384 78918 142476 78920
rect 142429 78916 142476 78918
rect 142540 78916 142546 78980
rect 143390 78916 143396 78980
rect 143460 78978 143466 78980
rect 144085 78978 144151 78981
rect 143460 78976 144151 78978
rect 143460 78920 144090 78976
rect 144146 78920 144151 78976
rect 143460 78918 144151 78920
rect 143460 78916 143466 78918
rect 142429 78915 142495 78916
rect 144085 78915 144151 78918
rect 149830 78916 149836 78980
rect 149900 78978 149906 78980
rect 150341 78978 150407 78981
rect 149900 78976 150407 78978
rect 149900 78920 150346 78976
rect 150402 78920 150407 78976
rect 149900 78918 150407 78920
rect 149900 78916 149906 78918
rect 150341 78915 150407 78918
rect 154614 78916 154620 78980
rect 154684 78978 154690 78980
rect 155769 78978 155835 78981
rect 154684 78976 155835 78978
rect 154684 78920 155774 78976
rect 155830 78920 155835 78976
rect 154684 78918 155835 78920
rect 154684 78916 154690 78918
rect 155769 78915 155835 78918
rect 157517 78978 157583 78981
rect 158294 78978 158300 78980
rect 157517 78976 158300 78978
rect 157517 78920 157522 78976
rect 157578 78920 158300 78976
rect 157517 78918 158300 78920
rect 157517 78915 157583 78918
rect 158294 78916 158300 78918
rect 158364 78916 158370 78980
rect 159950 78916 159956 78980
rect 160020 78978 160026 78980
rect 171409 78978 171475 78981
rect 160020 78976 171475 78978
rect 160020 78920 171414 78976
rect 171470 78920 171475 78976
rect 160020 78918 171475 78920
rect 160020 78916 160026 78918
rect 171409 78915 171475 78918
rect 172789 78978 172855 78981
rect 173198 78978 173204 78980
rect 172789 78976 173204 78978
rect 172789 78920 172794 78976
rect 172850 78920 173204 78976
rect 172789 78918 173204 78920
rect 172789 78915 172855 78918
rect 173198 78916 173204 78918
rect 173268 78916 173274 78980
rect 173433 78978 173499 78981
rect 173566 78978 173572 78980
rect 173433 78976 173572 78978
rect 173433 78920 173438 78976
rect 173494 78920 173572 78976
rect 173433 78918 173572 78920
rect 173433 78915 173499 78918
rect 173566 78916 173572 78918
rect 173636 78916 173642 78980
rect 174261 78978 174327 78981
rect 203190 78978 203196 78980
rect 174261 78976 203196 78978
rect 174261 78920 174266 78976
rect 174322 78920 203196 78976
rect 174261 78918 203196 78920
rect 174261 78915 174327 78918
rect 203190 78916 203196 78918
rect 203260 78916 203266 78980
rect 122046 78780 122052 78844
rect 122116 78842 122122 78844
rect 149237 78842 149303 78845
rect 122116 78840 149303 78842
rect 122116 78784 149242 78840
rect 149298 78784 149303 78840
rect 122116 78782 149303 78784
rect 122116 78780 122122 78782
rect 149237 78779 149303 78782
rect 158110 78780 158116 78844
rect 158180 78842 158186 78844
rect 158713 78842 158779 78845
rect 158180 78840 158779 78842
rect 158180 78784 158718 78840
rect 158774 78784 158779 78840
rect 158180 78782 158779 78784
rect 158180 78780 158186 78782
rect 158713 78779 158779 78782
rect 160686 78780 160692 78844
rect 160756 78842 160762 78844
rect 169845 78842 169911 78845
rect 160756 78840 169911 78842
rect 160756 78784 169850 78840
rect 169906 78784 169911 78840
rect 160756 78782 169911 78784
rect 160756 78780 160762 78782
rect 169845 78779 169911 78782
rect 171225 78842 171291 78845
rect 171910 78842 171916 78844
rect 171225 78840 171916 78842
rect 171225 78784 171230 78840
rect 171286 78784 171916 78840
rect 171225 78782 171916 78784
rect 171225 78779 171291 78782
rect 171910 78780 171916 78782
rect 171980 78780 171986 78844
rect 172646 78780 172652 78844
rect 172716 78842 172722 78844
rect 173617 78842 173683 78845
rect 172716 78840 173683 78842
rect 172716 78784 173622 78840
rect 173678 78784 173683 78840
rect 172716 78782 173683 78784
rect 172716 78780 172722 78782
rect 173617 78779 173683 78782
rect 174486 78780 174492 78844
rect 174556 78842 174562 78844
rect 174813 78842 174879 78845
rect 175273 78842 175339 78845
rect 174556 78840 174879 78842
rect 174556 78784 174818 78840
rect 174874 78784 174879 78840
rect 174556 78782 174879 78784
rect 174556 78780 174562 78782
rect 174813 78779 174879 78782
rect 175046 78840 175339 78842
rect 175046 78784 175278 78840
rect 175334 78784 175339 78840
rect 175046 78782 175339 78784
rect 130878 78644 130884 78708
rect 130948 78706 130954 78708
rect 143533 78706 143599 78709
rect 144361 78706 144427 78709
rect 130948 78704 144427 78706
rect 130948 78648 143538 78704
rect 143594 78648 144366 78704
rect 144422 78648 144427 78704
rect 130948 78646 144427 78648
rect 130948 78644 130954 78646
rect 143533 78643 143599 78646
rect 144361 78643 144427 78646
rect 151261 78708 151327 78709
rect 151261 78704 151308 78708
rect 151372 78706 151378 78708
rect 156137 78706 156203 78709
rect 156454 78706 156460 78708
rect 151261 78648 151266 78704
rect 151261 78644 151308 78648
rect 151372 78646 151418 78706
rect 156137 78704 156460 78706
rect 156137 78648 156142 78704
rect 156198 78648 156460 78704
rect 156137 78646 156460 78648
rect 151372 78644 151378 78646
rect 151261 78643 151327 78644
rect 156137 78643 156203 78646
rect 156454 78644 156460 78646
rect 156524 78644 156530 78708
rect 163446 78644 163452 78708
rect 163516 78706 163522 78708
rect 163865 78706 163931 78709
rect 163516 78704 163931 78706
rect 163516 78648 163870 78704
rect 163926 78648 163931 78704
rect 163516 78646 163931 78648
rect 163516 78644 163522 78646
rect 163865 78643 163931 78646
rect 165613 78706 165679 78709
rect 165838 78706 165844 78708
rect 165613 78704 165844 78706
rect 165613 78648 165618 78704
rect 165674 78648 165844 78704
rect 165613 78646 165844 78648
rect 165613 78643 165679 78646
rect 165838 78644 165844 78646
rect 165908 78706 165914 78708
rect 166390 78706 166396 78708
rect 165908 78646 166396 78706
rect 165908 78644 165914 78646
rect 166390 78644 166396 78646
rect 166460 78644 166466 78708
rect 174670 78644 174676 78708
rect 174740 78706 174746 78708
rect 175046 78706 175106 78782
rect 175273 78779 175339 78782
rect 175733 78842 175799 78845
rect 177941 78842 178007 78845
rect 206369 78842 206435 78845
rect 175733 78840 206435 78842
rect 175733 78784 175738 78840
rect 175794 78784 177946 78840
rect 178002 78784 206374 78840
rect 206430 78784 206435 78840
rect 175733 78782 206435 78784
rect 175733 78779 175799 78782
rect 177941 78779 178007 78782
rect 206369 78779 206435 78782
rect 174740 78646 175106 78706
rect 175273 78706 175339 78709
rect 175774 78706 175780 78708
rect 175273 78704 175780 78706
rect 175273 78648 175278 78704
rect 175334 78648 175780 78704
rect 175273 78646 175780 78648
rect 174740 78644 174746 78646
rect 175273 78643 175339 78646
rect 175774 78644 175780 78646
rect 175844 78644 175850 78708
rect 175958 78644 175964 78708
rect 176028 78706 176034 78708
rect 176377 78706 176443 78709
rect 187417 78706 187483 78709
rect 176028 78704 176443 78706
rect 176028 78648 176382 78704
rect 176438 78648 176443 78704
rect 176028 78646 176443 78648
rect 176028 78644 176034 78646
rect 176377 78643 176443 78646
rect 179370 78704 187483 78706
rect 179370 78648 187422 78704
rect 187478 78648 187483 78704
rect 179370 78646 187483 78648
rect 130377 78572 130443 78573
rect 130326 78570 130332 78572
rect 130286 78510 130332 78570
rect 130396 78568 130443 78572
rect 130438 78512 130443 78568
rect 130326 78508 130332 78510
rect 130396 78508 130443 78512
rect 130377 78507 130443 78508
rect 131941 78570 132007 78573
rect 133454 78570 133460 78572
rect 131941 78568 133460 78570
rect 131941 78512 131946 78568
rect 132002 78512 133460 78568
rect 131941 78510 133460 78512
rect 131941 78507 132007 78510
rect 133454 78508 133460 78510
rect 133524 78508 133530 78572
rect 134558 78508 134564 78572
rect 134628 78570 134634 78572
rect 134793 78570 134859 78573
rect 134628 78568 134859 78570
rect 134628 78512 134798 78568
rect 134854 78512 134859 78568
rect 134628 78510 134859 78512
rect 134628 78508 134634 78510
rect 134793 78507 134859 78510
rect 136173 78572 136239 78573
rect 136173 78568 136220 78572
rect 136284 78570 136290 78572
rect 136173 78512 136178 78568
rect 136173 78508 136220 78512
rect 136284 78510 136330 78570
rect 136284 78508 136290 78510
rect 136582 78508 136588 78572
rect 136652 78570 136658 78572
rect 136725 78570 136791 78573
rect 136909 78572 136975 78573
rect 136909 78570 136956 78572
rect 136652 78568 136791 78570
rect 136652 78512 136730 78568
rect 136786 78512 136791 78568
rect 136652 78510 136791 78512
rect 136864 78568 136956 78570
rect 136864 78512 136914 78568
rect 136864 78510 136956 78512
rect 136652 78508 136658 78510
rect 136173 78507 136239 78508
rect 136725 78507 136791 78510
rect 136909 78508 136956 78510
rect 137020 78508 137026 78572
rect 137185 78570 137251 78573
rect 137553 78570 137619 78573
rect 137185 78568 137619 78570
rect 137185 78512 137190 78568
rect 137246 78512 137558 78568
rect 137614 78512 137619 78568
rect 137185 78510 137619 78512
rect 136909 78507 136975 78508
rect 137185 78507 137251 78510
rect 137553 78507 137619 78510
rect 138013 78572 138079 78573
rect 138013 78568 138060 78572
rect 138124 78570 138130 78572
rect 138013 78512 138018 78568
rect 138013 78508 138060 78512
rect 138124 78510 138170 78570
rect 138124 78508 138130 78510
rect 140998 78508 141004 78572
rect 141068 78570 141074 78572
rect 141233 78570 141299 78573
rect 141068 78568 141299 78570
rect 141068 78512 141238 78568
rect 141294 78512 141299 78568
rect 141068 78510 141299 78512
rect 141068 78508 141074 78510
rect 138013 78507 138079 78508
rect 141233 78507 141299 78510
rect 143022 78508 143028 78572
rect 143092 78570 143098 78572
rect 143809 78570 143875 78573
rect 143092 78568 143875 78570
rect 143092 78512 143814 78568
rect 143870 78512 143875 78568
rect 143092 78510 143875 78512
rect 143092 78508 143098 78510
rect 143809 78507 143875 78510
rect 151486 78508 151492 78572
rect 151556 78570 151562 78572
rect 151721 78570 151787 78573
rect 151556 78568 151787 78570
rect 151556 78512 151726 78568
rect 151782 78512 151787 78568
rect 151556 78510 151787 78512
rect 151556 78508 151562 78510
rect 151721 78507 151787 78510
rect 156638 78508 156644 78572
rect 156708 78570 156714 78572
rect 157241 78570 157307 78573
rect 156708 78568 157307 78570
rect 156708 78512 157246 78568
rect 157302 78512 157307 78568
rect 156708 78510 157307 78512
rect 156708 78508 156714 78510
rect 157241 78507 157307 78510
rect 157701 78570 157767 78573
rect 161105 78572 161171 78573
rect 162761 78572 162827 78573
rect 158294 78570 158300 78572
rect 157701 78568 158300 78570
rect 157701 78512 157706 78568
rect 157762 78512 158300 78568
rect 157701 78510 158300 78512
rect 157701 78507 157767 78510
rect 158294 78508 158300 78510
rect 158364 78508 158370 78572
rect 161054 78570 161060 78572
rect 161014 78510 161060 78570
rect 161124 78568 161171 78572
rect 162710 78570 162716 78572
rect 161166 78512 161171 78568
rect 161054 78508 161060 78510
rect 161124 78508 161171 78512
rect 162670 78510 162716 78570
rect 162780 78568 162827 78572
rect 162822 78512 162827 78568
rect 162710 78508 162716 78510
rect 162780 78508 162827 78512
rect 161105 78507 161171 78508
rect 162761 78507 162827 78508
rect 171685 78570 171751 78573
rect 179370 78570 179430 78646
rect 187417 78643 187483 78646
rect 171685 78568 179430 78570
rect 171685 78512 171690 78568
rect 171746 78512 179430 78568
rect 171685 78510 179430 78512
rect 184473 78570 184539 78573
rect 184974 78570 184980 78572
rect 184473 78568 184980 78570
rect 184473 78512 184478 78568
rect 184534 78512 184980 78568
rect 184473 78510 184980 78512
rect 171685 78507 171751 78510
rect 184473 78507 184539 78510
rect 184974 78508 184980 78510
rect 185044 78508 185050 78572
rect 186405 78570 186471 78573
rect 187417 78572 187483 78573
rect 186814 78570 186820 78572
rect 186405 78568 186820 78570
rect 186405 78512 186410 78568
rect 186466 78512 186820 78568
rect 186405 78510 186820 78512
rect 186405 78507 186471 78510
rect 186814 78508 186820 78510
rect 186884 78508 186890 78572
rect 187366 78570 187372 78572
rect 187326 78510 187372 78570
rect 187436 78568 187483 78572
rect 187478 78512 187483 78568
rect 187366 78508 187372 78510
rect 187436 78508 187483 78512
rect 187417 78507 187483 78508
rect 193581 78572 193647 78573
rect 193581 78568 193628 78572
rect 193692 78570 193698 78572
rect 193581 78512 193586 78568
rect 193581 78508 193628 78512
rect 193692 78510 193738 78570
rect 193692 78508 193698 78510
rect 193581 78507 193647 78508
rect 125174 78372 125180 78436
rect 125244 78434 125250 78436
rect 138105 78434 138171 78437
rect 141693 78436 141759 78437
rect 141693 78434 141740 78436
rect 125244 78432 138171 78434
rect 125244 78376 138110 78432
rect 138166 78376 138171 78432
rect 125244 78374 138171 78376
rect 141648 78432 141740 78434
rect 141648 78376 141698 78432
rect 141648 78374 141740 78376
rect 125244 78372 125250 78374
rect 138105 78371 138171 78374
rect 141693 78372 141740 78374
rect 141804 78372 141810 78436
rect 142521 78434 142587 78437
rect 165521 78436 165587 78437
rect 143206 78434 143212 78436
rect 142521 78432 143212 78434
rect 142521 78376 142526 78432
rect 142582 78376 143212 78432
rect 142521 78374 143212 78376
rect 141693 78371 141759 78372
rect 142521 78371 142587 78374
rect 143206 78372 143212 78374
rect 143276 78372 143282 78436
rect 165470 78434 165476 78436
rect 165430 78374 165476 78434
rect 165540 78432 165587 78436
rect 165582 78376 165587 78432
rect 165470 78372 165476 78374
rect 165540 78372 165587 78376
rect 171358 78372 171364 78436
rect 171428 78434 171434 78436
rect 195237 78434 195303 78437
rect 171428 78432 195303 78434
rect 171428 78376 195242 78432
rect 195298 78376 195303 78432
rect 171428 78374 195303 78376
rect 171428 78372 171434 78374
rect 165521 78371 165587 78372
rect 195237 78371 195303 78374
rect 126830 78236 126836 78300
rect 126900 78298 126906 78300
rect 137829 78298 137895 78301
rect 138565 78300 138631 78301
rect 138565 78298 138612 78300
rect 126900 78296 137895 78298
rect 126900 78240 137834 78296
rect 137890 78240 137895 78296
rect 126900 78238 137895 78240
rect 138520 78296 138612 78298
rect 138520 78240 138570 78296
rect 138520 78238 138612 78240
rect 126900 78236 126906 78238
rect 137829 78235 137895 78238
rect 138565 78236 138612 78238
rect 138676 78236 138682 78300
rect 138749 78298 138815 78301
rect 145741 78298 145807 78301
rect 138749 78296 145807 78298
rect 138749 78240 138754 78296
rect 138810 78240 145746 78296
rect 145802 78240 145807 78296
rect 138749 78238 145807 78240
rect 138565 78235 138631 78236
rect 138749 78235 138815 78238
rect 145741 78235 145807 78238
rect 148174 78236 148180 78300
rect 148244 78298 148250 78300
rect 148685 78298 148751 78301
rect 148244 78296 148751 78298
rect 148244 78240 148690 78296
rect 148746 78240 148751 78296
rect 148244 78238 148751 78240
rect 148244 78236 148250 78238
rect 148685 78235 148751 78238
rect 149605 78298 149671 78301
rect 150014 78298 150020 78300
rect 149605 78296 150020 78298
rect 149605 78240 149610 78296
rect 149666 78240 150020 78296
rect 149605 78238 150020 78240
rect 149605 78235 149671 78238
rect 150014 78236 150020 78238
rect 150084 78236 150090 78300
rect 164550 78298 164556 78300
rect 157290 78238 164556 78298
rect 124070 78100 124076 78164
rect 124140 78162 124146 78164
rect 143441 78162 143507 78165
rect 155125 78164 155191 78165
rect 155125 78162 155172 78164
rect 124140 78160 143507 78162
rect 124140 78104 143446 78160
rect 143502 78104 143507 78160
rect 124140 78102 143507 78104
rect 155080 78160 155172 78162
rect 155080 78104 155130 78160
rect 155080 78102 155172 78104
rect 124140 78100 124146 78102
rect 143441 78099 143507 78102
rect 155125 78100 155172 78102
rect 155236 78100 155242 78164
rect 155125 78099 155191 78100
rect 127382 77964 127388 78028
rect 127452 78026 127458 78028
rect 148593 78026 148659 78029
rect 127452 78024 148659 78026
rect 127452 77968 148598 78024
rect 148654 77968 148659 78024
rect 127452 77966 148659 77968
rect 127452 77964 127458 77966
rect 148593 77963 148659 77966
rect 148726 77964 148732 78028
rect 148796 78026 148802 78028
rect 157290 78026 157350 78238
rect 164550 78236 164556 78238
rect 164620 78236 164626 78300
rect 169937 78298 170003 78301
rect 198089 78298 198155 78301
rect 169937 78296 198155 78298
rect 169937 78240 169942 78296
rect 169998 78240 198094 78296
rect 198150 78240 198155 78296
rect 169937 78238 198155 78240
rect 169937 78235 170003 78238
rect 198089 78235 198155 78238
rect 163865 78162 163931 78165
rect 163998 78162 164004 78164
rect 163865 78160 164004 78162
rect 163865 78104 163870 78160
rect 163926 78104 164004 78160
rect 163865 78102 164004 78104
rect 163865 78099 163931 78102
rect 163998 78100 164004 78102
rect 164068 78100 164074 78164
rect 167729 78162 167795 78165
rect 167862 78162 167868 78164
rect 167729 78160 167868 78162
rect 167729 78104 167734 78160
rect 167790 78104 167868 78160
rect 167729 78102 167868 78104
rect 167729 78099 167795 78102
rect 167862 78100 167868 78102
rect 167932 78100 167938 78164
rect 170806 78100 170812 78164
rect 170876 78162 170882 78164
rect 171133 78162 171199 78165
rect 170876 78160 171199 78162
rect 170876 78104 171138 78160
rect 171194 78104 171199 78160
rect 170876 78102 171199 78104
rect 170876 78100 170882 78102
rect 171133 78099 171199 78102
rect 177849 78162 177915 78165
rect 204897 78162 204963 78165
rect 177849 78160 204963 78162
rect 177849 78104 177854 78160
rect 177910 78104 204902 78160
rect 204958 78104 204963 78160
rect 177849 78102 204963 78104
rect 177849 78099 177915 78102
rect 204897 78099 204963 78102
rect 148796 77966 157350 78026
rect 148796 77964 148802 77966
rect 173750 77964 173756 78028
rect 173820 78026 173826 78028
rect 199193 78026 199259 78029
rect 173820 78024 200130 78026
rect 173820 77968 199198 78024
rect 199254 77968 200130 78024
rect 173820 77966 200130 77968
rect 173820 77964 173826 77966
rect 199193 77963 199259 77966
rect 119838 77828 119844 77892
rect 119908 77890 119914 77892
rect 132033 77890 132099 77893
rect 133229 77892 133295 77893
rect 133229 77890 133276 77892
rect 119908 77888 132099 77890
rect 119908 77832 132038 77888
rect 132094 77832 132099 77888
rect 119908 77830 132099 77832
rect 133184 77888 133276 77890
rect 133184 77832 133234 77888
rect 133184 77830 133276 77832
rect 119908 77828 119914 77830
rect 132033 77827 132099 77830
rect 133229 77828 133276 77830
rect 133340 77828 133346 77892
rect 133413 77890 133479 77893
rect 134742 77890 134748 77892
rect 133413 77888 134748 77890
rect 133413 77832 133418 77888
rect 133474 77832 134748 77888
rect 133413 77830 134748 77832
rect 133229 77827 133295 77828
rect 133413 77827 133479 77830
rect 134742 77828 134748 77830
rect 134812 77828 134818 77892
rect 135713 77890 135779 77893
rect 136030 77890 136036 77892
rect 135713 77888 136036 77890
rect 135713 77832 135718 77888
rect 135774 77832 136036 77888
rect 135713 77830 136036 77832
rect 135713 77827 135779 77830
rect 136030 77828 136036 77830
rect 136100 77828 136106 77892
rect 136725 77890 136791 77893
rect 137870 77890 137876 77892
rect 136725 77888 137876 77890
rect 136725 77832 136730 77888
rect 136786 77832 137876 77888
rect 136725 77830 137876 77832
rect 136725 77827 136791 77830
rect 137870 77828 137876 77830
rect 137940 77828 137946 77892
rect 138105 77890 138171 77893
rect 138974 77890 138980 77892
rect 138105 77888 138980 77890
rect 138105 77832 138110 77888
rect 138166 77832 138980 77888
rect 138105 77830 138980 77832
rect 138105 77827 138171 77830
rect 138974 77828 138980 77830
rect 139044 77828 139050 77892
rect 139393 77890 139459 77893
rect 140037 77892 140103 77893
rect 139710 77890 139716 77892
rect 139393 77888 139716 77890
rect 139393 77832 139398 77888
rect 139454 77832 139716 77888
rect 139393 77830 139716 77832
rect 139393 77827 139459 77830
rect 139710 77828 139716 77830
rect 139780 77828 139786 77892
rect 140037 77888 140084 77892
rect 140148 77890 140154 77892
rect 140037 77832 140042 77888
rect 140037 77828 140084 77832
rect 140148 77830 140194 77890
rect 140148 77828 140154 77830
rect 140814 77828 140820 77892
rect 140884 77890 140890 77892
rect 141325 77890 141391 77893
rect 140884 77888 141391 77890
rect 140884 77832 141330 77888
rect 141386 77832 141391 77888
rect 140884 77830 141391 77832
rect 140884 77828 140890 77830
rect 140037 77827 140103 77828
rect 141325 77827 141391 77830
rect 147070 77828 147076 77892
rect 147140 77890 147146 77892
rect 147305 77890 147371 77893
rect 147140 77888 147371 77890
rect 147140 77832 147310 77888
rect 147366 77832 147371 77888
rect 147140 77830 147371 77832
rect 147140 77828 147146 77830
rect 147305 77827 147371 77830
rect 147990 77828 147996 77892
rect 148060 77890 148066 77892
rect 148685 77890 148751 77893
rect 148060 77888 148751 77890
rect 148060 77832 148690 77888
rect 148746 77832 148751 77888
rect 148060 77830 148751 77832
rect 148060 77828 148066 77830
rect 148685 77827 148751 77830
rect 149094 77828 149100 77892
rect 149164 77890 149170 77892
rect 150433 77890 150499 77893
rect 149164 77888 150499 77890
rect 149164 77832 150438 77888
rect 150494 77832 150499 77888
rect 149164 77830 150499 77832
rect 149164 77828 149170 77830
rect 150433 77827 150499 77830
rect 160318 77828 160324 77892
rect 160388 77890 160394 77892
rect 171593 77890 171659 77893
rect 160388 77888 171659 77890
rect 160388 77832 171598 77888
rect 171654 77832 171659 77888
rect 160388 77830 171659 77832
rect 160388 77828 160394 77830
rect 171593 77827 171659 77830
rect 176326 77828 176332 77892
rect 176396 77890 176402 77892
rect 176561 77890 176627 77893
rect 176396 77888 176627 77890
rect 176396 77832 176566 77888
rect 176622 77832 176627 77888
rect 176396 77830 176627 77832
rect 200070 77890 200130 77966
rect 291837 77890 291903 77893
rect 200070 77888 291903 77890
rect 200070 77832 291842 77888
rect 291898 77832 291903 77888
rect 200070 77830 291903 77832
rect 176396 77828 176402 77830
rect 176561 77827 176627 77830
rect 291837 77827 291903 77830
rect 124806 77692 124812 77756
rect 124876 77754 124882 77756
rect 140497 77754 140563 77757
rect 142337 77756 142403 77757
rect 142286 77754 142292 77756
rect 124876 77752 140563 77754
rect 124876 77696 140502 77752
rect 140558 77696 140563 77752
rect 124876 77694 140563 77696
rect 142246 77694 142292 77754
rect 142356 77752 142403 77756
rect 142398 77696 142403 77752
rect 124876 77692 124882 77694
rect 140497 77691 140563 77694
rect 142286 77692 142292 77694
rect 142356 77692 142403 77696
rect 145046 77692 145052 77756
rect 145116 77754 145122 77756
rect 146109 77754 146175 77757
rect 145116 77752 146175 77754
rect 145116 77696 146114 77752
rect 146170 77696 146175 77752
rect 145116 77694 146175 77696
rect 145116 77692 145122 77694
rect 142337 77691 142403 77692
rect 146109 77691 146175 77694
rect 146886 77692 146892 77756
rect 146956 77754 146962 77756
rect 147806 77754 147812 77756
rect 146956 77694 147812 77754
rect 146956 77692 146962 77694
rect 147806 77692 147812 77694
rect 147876 77692 147882 77756
rect 149278 77692 149284 77756
rect 149348 77754 149354 77756
rect 149881 77754 149947 77757
rect 149348 77752 149947 77754
rect 149348 77696 149886 77752
rect 149942 77696 149947 77752
rect 149348 77694 149947 77696
rect 149348 77692 149354 77694
rect 149881 77691 149947 77694
rect 165245 77754 165311 77757
rect 165470 77754 165476 77756
rect 165245 77752 165476 77754
rect 165245 77696 165250 77752
rect 165306 77696 165476 77752
rect 165245 77694 165476 77696
rect 165245 77691 165311 77694
rect 165470 77692 165476 77694
rect 165540 77692 165546 77756
rect 171869 77754 171935 77757
rect 172462 77754 172468 77756
rect 171869 77752 172468 77754
rect 171869 77696 171874 77752
rect 171930 77696 172468 77752
rect 171869 77694 172468 77696
rect 171869 77691 171935 77694
rect 172462 77692 172468 77694
rect 172532 77692 172538 77756
rect 180425 77754 180491 77757
rect 207013 77754 207079 77757
rect 180425 77752 207079 77754
rect 180425 77696 180430 77752
rect 180486 77696 207018 77752
rect 207074 77696 207079 77752
rect 180425 77694 207079 77696
rect 180425 77691 180491 77694
rect 207013 77691 207079 77694
rect 131982 77556 131988 77620
rect 132052 77618 132058 77620
rect 133965 77618 134031 77621
rect 132052 77616 134031 77618
rect 132052 77560 133970 77616
rect 134026 77560 134031 77616
rect 132052 77558 134031 77560
rect 132052 77556 132058 77558
rect 133965 77555 134031 77558
rect 135989 77618 136055 77621
rect 137553 77620 137619 77621
rect 136398 77618 136404 77620
rect 135989 77616 136404 77618
rect 135989 77560 135994 77616
rect 136050 77560 136404 77616
rect 135989 77558 136404 77560
rect 135989 77555 136055 77558
rect 136398 77556 136404 77558
rect 136468 77556 136474 77620
rect 137502 77618 137508 77620
rect 137462 77558 137508 77618
rect 137572 77616 137619 77620
rect 145373 77618 145439 77621
rect 137614 77560 137619 77616
rect 137502 77556 137508 77558
rect 137572 77556 137619 77560
rect 137553 77555 137619 77556
rect 137970 77616 145439 77618
rect 137970 77560 145378 77616
rect 145434 77560 145439 77616
rect 137970 77558 145439 77560
rect 137553 77482 137619 77485
rect 137686 77482 137692 77484
rect 137553 77480 137692 77482
rect 137553 77424 137558 77480
rect 137614 77424 137692 77480
rect 137553 77422 137692 77424
rect 137553 77419 137619 77422
rect 137686 77420 137692 77422
rect 137756 77420 137762 77484
rect 124990 77284 124996 77348
rect 125060 77346 125066 77348
rect 137970 77346 138030 77558
rect 145373 77555 145439 77558
rect 145598 77556 145604 77620
rect 145668 77618 145674 77620
rect 156137 77618 156203 77621
rect 145668 77616 156203 77618
rect 145668 77560 156142 77616
rect 156198 77560 156203 77616
rect 145668 77558 156203 77560
rect 145668 77556 145674 77558
rect 156137 77555 156203 77558
rect 156781 77618 156847 77621
rect 157006 77618 157012 77620
rect 156781 77616 157012 77618
rect 156781 77560 156786 77616
rect 156842 77560 157012 77616
rect 156781 77558 157012 77560
rect 156781 77555 156847 77558
rect 157006 77556 157012 77558
rect 157076 77556 157082 77620
rect 163630 77556 163636 77620
rect 163700 77618 163706 77620
rect 164141 77618 164207 77621
rect 163700 77616 164207 77618
rect 163700 77560 164146 77616
rect 164202 77560 164207 77616
rect 163700 77558 164207 77560
rect 163700 77556 163706 77558
rect 164141 77555 164207 77558
rect 164550 77556 164556 77620
rect 164620 77618 164626 77620
rect 165245 77618 165311 77621
rect 164620 77616 165311 77618
rect 164620 77560 165250 77616
rect 165306 77560 165311 77616
rect 164620 77558 165311 77560
rect 164620 77556 164626 77558
rect 165245 77555 165311 77558
rect 173934 77556 173940 77620
rect 174004 77618 174010 77620
rect 174905 77618 174971 77621
rect 175089 77618 175155 77621
rect 174004 77616 175155 77618
rect 174004 77560 174910 77616
rect 174966 77560 175094 77616
rect 175150 77560 175155 77616
rect 174004 77558 175155 77560
rect 174004 77556 174010 77558
rect 174905 77555 174971 77558
rect 175089 77555 175155 77558
rect 177665 77618 177731 77621
rect 468569 77618 468635 77621
rect 177665 77616 468635 77618
rect 177665 77560 177670 77616
rect 177726 77560 468574 77616
rect 468630 77560 468635 77616
rect 177665 77558 468635 77560
rect 177665 77555 177731 77558
rect 468569 77555 468635 77558
rect 138238 77420 138244 77484
rect 138308 77482 138314 77484
rect 138933 77482 138999 77485
rect 138308 77480 138999 77482
rect 138308 77424 138938 77480
rect 138994 77424 138999 77480
rect 138308 77422 138999 77424
rect 138308 77420 138314 77422
rect 138933 77419 138999 77422
rect 140037 77482 140103 77485
rect 147990 77482 147996 77484
rect 140037 77480 147996 77482
rect 140037 77424 140042 77480
rect 140098 77424 147996 77480
rect 140037 77422 147996 77424
rect 140037 77419 140103 77422
rect 147990 77420 147996 77422
rect 148060 77420 148066 77484
rect 148358 77420 148364 77484
rect 148428 77482 148434 77484
rect 148961 77482 149027 77485
rect 148428 77480 149027 77482
rect 148428 77424 148966 77480
rect 149022 77424 149027 77480
rect 148428 77422 149027 77424
rect 148428 77420 148434 77422
rect 148961 77419 149027 77422
rect 153285 77482 153351 77485
rect 154062 77482 154068 77484
rect 153285 77480 154068 77482
rect 153285 77424 153290 77480
rect 153346 77424 154068 77480
rect 153285 77422 154068 77424
rect 153285 77419 153351 77422
rect 154062 77420 154068 77422
rect 154132 77420 154138 77484
rect 164785 77482 164851 77485
rect 170857 77484 170923 77485
rect 165102 77482 165108 77484
rect 164785 77480 165108 77482
rect 164785 77424 164790 77480
rect 164846 77424 165108 77480
rect 164785 77422 165108 77424
rect 164785 77419 164851 77422
rect 165102 77420 165108 77422
rect 165172 77420 165178 77484
rect 170806 77482 170812 77484
rect 170766 77422 170812 77482
rect 170876 77480 170923 77484
rect 170918 77424 170923 77480
rect 170806 77420 170812 77422
rect 170876 77420 170923 77424
rect 170857 77419 170923 77420
rect 178953 77482 179019 77485
rect 201401 77482 201467 77485
rect 178953 77480 201467 77482
rect 178953 77424 178958 77480
rect 179014 77424 201406 77480
rect 201462 77424 201467 77480
rect 178953 77422 201467 77424
rect 178953 77419 179019 77422
rect 201401 77419 201467 77422
rect 125060 77286 138030 77346
rect 138289 77346 138355 77349
rect 154481 77348 154547 77349
rect 170489 77348 170555 77349
rect 144310 77346 144316 77348
rect 138289 77344 144316 77346
rect 138289 77288 138294 77344
rect 138350 77288 144316 77344
rect 138289 77286 144316 77288
rect 125060 77284 125066 77286
rect 138289 77283 138355 77286
rect 144310 77284 144316 77286
rect 144380 77284 144386 77348
rect 154430 77284 154436 77348
rect 154500 77346 154547 77348
rect 170438 77346 170444 77348
rect 154500 77344 154592 77346
rect 154542 77288 154592 77344
rect 154500 77286 154592 77288
rect 170398 77286 170444 77346
rect 170508 77344 170555 77348
rect 170550 77288 170555 77344
rect 154500 77284 154547 77286
rect 170438 77284 170444 77286
rect 170508 77284 170555 77288
rect 154481 77283 154547 77284
rect 170489 77283 170555 77284
rect 170765 77346 170831 77349
rect 170990 77346 170996 77348
rect 170765 77344 170996 77346
rect 170765 77288 170770 77344
rect 170826 77288 170996 77344
rect 170765 77286 170996 77288
rect 170765 77283 170831 77286
rect 170990 77284 170996 77286
rect 171060 77284 171066 77348
rect 177757 77346 177823 77349
rect 177941 77346 178007 77349
rect 180425 77346 180491 77349
rect 177757 77344 180491 77346
rect 177757 77288 177762 77344
rect 177818 77288 177946 77344
rect 178002 77288 180430 77344
rect 180486 77288 180491 77344
rect 177757 77286 180491 77288
rect 177757 77283 177823 77286
rect 177941 77283 178007 77286
rect 180425 77283 180491 77286
rect 112621 77210 112687 77213
rect 146886 77210 146892 77212
rect 112621 77208 146892 77210
rect 112621 77152 112626 77208
rect 112682 77152 146892 77208
rect 112621 77150 146892 77152
rect 112621 77147 112687 77150
rect 146886 77148 146892 77150
rect 146956 77148 146962 77212
rect 155585 77210 155651 77213
rect 178718 77210 178724 77212
rect 155585 77208 178724 77210
rect 155585 77152 155590 77208
rect 155646 77152 178724 77208
rect 155585 77150 178724 77152
rect 155585 77147 155651 77150
rect 178718 77148 178724 77150
rect 178788 77148 178794 77212
rect 114369 77074 114435 77077
rect 148358 77074 148364 77076
rect 114369 77072 148364 77074
rect 114369 77016 114374 77072
rect 114430 77016 148364 77072
rect 114369 77014 148364 77016
rect 114369 77011 114435 77014
rect 148358 77012 148364 77014
rect 148428 77012 148434 77076
rect 155861 77074 155927 77077
rect 181478 77074 181484 77076
rect 155861 77072 181484 77074
rect 155861 77016 155866 77072
rect 155922 77016 181484 77072
rect 155861 77014 181484 77016
rect 155861 77011 155927 77014
rect 181478 77012 181484 77014
rect 181548 77074 181554 77076
rect 183277 77074 183343 77077
rect 181548 77072 183343 77074
rect 181548 77016 183282 77072
rect 183338 77016 183343 77072
rect 181548 77014 183343 77016
rect 181548 77012 181554 77014
rect 183277 77011 183343 77014
rect 116577 76938 116643 76941
rect 146293 76938 146359 76941
rect 146937 76938 147003 76941
rect 116577 76936 147003 76938
rect 116577 76880 116582 76936
rect 116638 76880 146298 76936
rect 146354 76880 146942 76936
rect 146998 76880 147003 76936
rect 116577 76878 147003 76880
rect 116577 76875 116643 76878
rect 146293 76875 146359 76878
rect 146937 76875 147003 76878
rect 170581 76938 170647 76941
rect 193438 76938 193444 76940
rect 170581 76936 193444 76938
rect 170581 76880 170586 76936
rect 170642 76880 193444 76936
rect 170581 76878 193444 76880
rect 170581 76875 170647 76878
rect 193438 76876 193444 76878
rect 193508 76876 193514 76940
rect 112253 76802 112319 76805
rect 140865 76802 140931 76805
rect 112253 76800 140931 76802
rect 112253 76744 112258 76800
rect 112314 76744 140870 76800
rect 140926 76744 140931 76800
rect 112253 76742 140931 76744
rect 112253 76739 112319 76742
rect 140865 76739 140931 76742
rect 171501 76802 171567 76805
rect 192150 76802 192156 76804
rect 171501 76800 192156 76802
rect 171501 76744 171506 76800
rect 171562 76744 192156 76800
rect 171501 76742 192156 76744
rect 171501 76739 171567 76742
rect 192150 76740 192156 76742
rect 192220 76740 192226 76804
rect 125593 76666 125659 76669
rect 141877 76666 141943 76669
rect 125593 76664 141943 76666
rect 125593 76608 125598 76664
rect 125654 76608 141882 76664
rect 141938 76608 141943 76664
rect 125593 76606 141943 76608
rect 125593 76603 125659 76606
rect 141877 76603 141943 76606
rect 177573 76666 177639 76669
rect 180057 76666 180123 76669
rect 177573 76664 180123 76666
rect 177573 76608 177578 76664
rect 177634 76608 180062 76664
rect 180118 76608 180123 76664
rect 177573 76606 180123 76608
rect 177573 76603 177639 76606
rect 180057 76603 180123 76606
rect 183277 76666 183343 76669
rect 260833 76666 260899 76669
rect 183277 76664 260899 76666
rect 183277 76608 183282 76664
rect 183338 76608 260838 76664
rect 260894 76608 260899 76664
rect 183277 76606 260899 76608
rect 183277 76603 183343 76606
rect 260833 76603 260899 76606
rect 4797 76530 4863 76533
rect 4797 76528 103530 76530
rect 4797 76472 4802 76528
rect 4858 76472 103530 76528
rect 4797 76470 103530 76472
rect 4797 76467 4863 76470
rect 103470 76258 103530 76470
rect 135478 76468 135484 76532
rect 135548 76530 135554 76532
rect 135805 76530 135871 76533
rect 135548 76528 135871 76530
rect 135548 76472 135810 76528
rect 135866 76472 135871 76528
rect 135548 76470 135871 76472
rect 135548 76468 135554 76470
rect 135805 76467 135871 76470
rect 170765 76530 170831 76533
rect 189390 76530 189396 76532
rect 170765 76528 189396 76530
rect 170765 76472 170770 76528
rect 170826 76472 189396 76528
rect 170765 76470 189396 76472
rect 170765 76467 170831 76470
rect 189390 76468 189396 76470
rect 189460 76468 189466 76532
rect 553393 76530 553459 76533
rect 209730 76528 553459 76530
rect 209730 76472 553398 76528
rect 553454 76472 553459 76528
rect 209730 76470 553459 76472
rect 173709 76394 173775 76397
rect 179321 76394 179387 76397
rect 193254 76394 193260 76396
rect 173709 76392 193260 76394
rect 173709 76336 173714 76392
rect 173770 76336 179326 76392
rect 179382 76336 193260 76392
rect 173709 76334 193260 76336
rect 173709 76331 173775 76334
rect 179321 76331 179387 76334
rect 193254 76332 193260 76334
rect 193324 76332 193330 76396
rect 104157 76258 104223 76261
rect 132585 76258 132651 76261
rect 103470 76256 132651 76258
rect 103470 76200 104162 76256
rect 104218 76200 132590 76256
rect 132646 76200 132651 76256
rect 103470 76198 132651 76200
rect 104157 76195 104223 76198
rect 132585 76195 132651 76198
rect 175406 76196 175412 76260
rect 175476 76258 175482 76260
rect 208669 76258 208735 76261
rect 209730 76258 209790 76470
rect 553393 76467 553459 76470
rect 175476 76256 209790 76258
rect 175476 76200 208674 76256
rect 208730 76200 209790 76256
rect 175476 76198 209790 76200
rect 175476 76196 175482 76198
rect 208669 76195 208735 76198
rect 172145 76124 172211 76125
rect 172094 76122 172100 76124
rect 172054 76062 172100 76122
rect 172164 76120 172211 76124
rect 172206 76064 172211 76120
rect 172094 76060 172100 76062
rect 172164 76060 172211 76064
rect 173566 76060 173572 76124
rect 173636 76122 173642 76124
rect 173801 76122 173867 76125
rect 173636 76120 173867 76122
rect 173636 76064 173806 76120
rect 173862 76064 173867 76120
rect 173636 76062 173867 76064
rect 173636 76060 173642 76062
rect 172145 76059 172211 76060
rect 173801 76059 173867 76062
rect 130377 75986 130443 75989
rect 131573 75986 131639 75989
rect 130377 75984 131639 75986
rect 130377 75928 130382 75984
rect 130438 75928 131578 75984
rect 131634 75928 131639 75984
rect 130377 75926 131639 75928
rect 130377 75923 130443 75926
rect 131573 75923 131639 75926
rect 157926 75924 157932 75988
rect 157996 75986 158002 75988
rect 158069 75986 158135 75989
rect 169385 75988 169451 75989
rect 169334 75986 169340 75988
rect 157996 75984 158135 75986
rect 157996 75928 158074 75984
rect 158130 75928 158135 75984
rect 157996 75926 158135 75928
rect 169294 75926 169340 75986
rect 169404 75984 169451 75988
rect 169446 75928 169451 75984
rect 157996 75924 158002 75926
rect 158069 75923 158135 75926
rect 169334 75924 169340 75926
rect 169404 75924 169451 75928
rect 171910 75924 171916 75988
rect 171980 75986 171986 75988
rect 172237 75986 172303 75989
rect 171980 75984 172303 75986
rect 171980 75928 172242 75984
rect 172298 75928 172303 75984
rect 171980 75926 172303 75928
rect 171980 75924 171986 75926
rect 169385 75923 169451 75924
rect 172237 75923 172303 75926
rect 172605 75986 172671 75989
rect 172605 75984 179430 75986
rect 172605 75928 172610 75984
rect 172666 75928 179430 75984
rect 172605 75926 179430 75928
rect 172605 75923 172671 75926
rect 117078 75788 117084 75852
rect 117148 75850 117154 75852
rect 157977 75850 158043 75853
rect 117148 75848 158043 75850
rect 117148 75792 157982 75848
rect 158038 75792 158043 75848
rect 117148 75790 158043 75792
rect 117148 75788 117154 75790
rect 157977 75787 158043 75790
rect 174445 75850 174511 75853
rect 174854 75850 174860 75852
rect 174445 75848 174860 75850
rect 174445 75792 174450 75848
rect 174506 75792 174860 75848
rect 174445 75790 174860 75792
rect 174445 75787 174511 75790
rect 174854 75788 174860 75790
rect 174924 75788 174930 75852
rect 179370 75850 179430 75926
rect 205725 75850 205791 75853
rect 179370 75848 209790 75850
rect 179370 75792 205730 75848
rect 205786 75792 209790 75848
rect 179370 75790 209790 75792
rect 205725 75787 205791 75790
rect 112989 75714 113055 75717
rect 176561 75716 176627 75717
rect 147070 75714 147076 75716
rect 112989 75712 147076 75714
rect 112989 75656 112994 75712
rect 113050 75656 147076 75712
rect 112989 75654 147076 75656
rect 112989 75651 113055 75654
rect 147070 75652 147076 75654
rect 147140 75652 147146 75716
rect 176510 75714 176516 75716
rect 176434 75654 176516 75714
rect 176580 75714 176627 75716
rect 206093 75714 206159 75717
rect 176580 75712 206159 75714
rect 176622 75656 206098 75712
rect 206154 75656 206159 75712
rect 176510 75652 176516 75654
rect 176580 75654 206159 75656
rect 176580 75652 176627 75654
rect 176561 75651 176627 75652
rect 206093 75651 206159 75654
rect 118417 75578 118483 75581
rect 148910 75578 148916 75580
rect 118417 75576 148916 75578
rect 118417 75520 118422 75576
rect 118478 75520 148916 75576
rect 118417 75518 148916 75520
rect 118417 75515 118483 75518
rect 148910 75516 148916 75518
rect 148980 75516 148986 75580
rect 175181 75578 175247 75581
rect 203006 75578 203012 75580
rect 175181 75576 203012 75578
rect 175181 75520 175186 75576
rect 175242 75520 203012 75576
rect 175181 75518 203012 75520
rect 175181 75515 175247 75518
rect 203006 75516 203012 75518
rect 203076 75516 203082 75580
rect 120993 75442 121059 75445
rect 141509 75442 141575 75445
rect 120993 75440 141575 75442
rect 120993 75384 120998 75440
rect 121054 75384 141514 75440
rect 141570 75384 141575 75440
rect 120993 75382 141575 75384
rect 120993 75379 121059 75382
rect 141509 75379 141575 75382
rect 170305 75442 170371 75445
rect 179229 75442 179295 75445
rect 196382 75442 196388 75444
rect 170305 75440 196388 75442
rect 170305 75384 170310 75440
rect 170366 75384 179234 75440
rect 179290 75384 196388 75440
rect 170305 75382 196388 75384
rect 170305 75379 170371 75382
rect 179229 75379 179295 75382
rect 196382 75380 196388 75382
rect 196452 75380 196458 75444
rect 209730 75442 209790 75790
rect 486417 75442 486483 75445
rect 209730 75440 486483 75442
rect 209730 75384 486422 75440
rect 486478 75384 486483 75440
rect 209730 75382 486483 75384
rect 486417 75379 486483 75382
rect 113449 75306 113515 75309
rect 129733 75306 129799 75309
rect 130929 75306 130995 75309
rect 113449 75304 130995 75306
rect 113449 75248 113454 75304
rect 113510 75248 129738 75304
rect 129794 75248 130934 75304
rect 130990 75248 130995 75304
rect 113449 75246 130995 75248
rect 113449 75243 113515 75246
rect 129733 75243 129799 75246
rect 130929 75243 130995 75246
rect 172973 75306 173039 75309
rect 521653 75306 521719 75309
rect 172973 75304 521719 75306
rect 172973 75248 172978 75304
rect 173034 75248 521658 75304
rect 521714 75248 521719 75304
rect 172973 75246 521719 75248
rect 172973 75243 173039 75246
rect 521653 75243 521719 75246
rect 7557 75170 7623 75173
rect 119838 75170 119844 75172
rect 7557 75168 119844 75170
rect 7557 75112 7562 75168
rect 7618 75112 119844 75168
rect 7557 75110 119844 75112
rect 7557 75107 7623 75110
rect 119838 75108 119844 75110
rect 119908 75108 119914 75172
rect 174905 75170 174971 75173
rect 549253 75170 549319 75173
rect 174905 75168 549319 75170
rect 174905 75112 174910 75168
rect 174966 75112 549258 75168
rect 549314 75112 549319 75168
rect 174905 75110 549319 75112
rect 174905 75107 174971 75110
rect 549253 75107 549319 75110
rect 159030 74972 159036 75036
rect 159100 75034 159106 75036
rect 160001 75034 160067 75037
rect 159100 75032 160067 75034
rect 159100 74976 160006 75032
rect 160062 74976 160067 75032
rect 159100 74974 160067 74976
rect 159100 74972 159106 74974
rect 160001 74971 160067 74974
rect 154021 74626 154087 74629
rect 154246 74626 154252 74628
rect 154021 74624 154252 74626
rect 154021 74568 154026 74624
rect 154082 74568 154252 74624
rect 154021 74566 154252 74568
rect 154021 74563 154087 74566
rect 154246 74564 154252 74566
rect 154316 74564 154322 74628
rect 120574 74428 120580 74492
rect 120644 74490 120650 74492
rect 153929 74490 153995 74493
rect 120644 74488 153995 74490
rect 120644 74432 153934 74488
rect 153990 74432 153995 74488
rect 120644 74430 153995 74432
rect 120644 74428 120650 74430
rect 153929 74427 153995 74430
rect 156454 74428 156460 74492
rect 156524 74490 156530 74492
rect 189625 74490 189691 74493
rect 156524 74488 189691 74490
rect 156524 74432 189630 74488
rect 189686 74432 189691 74488
rect 156524 74430 189691 74432
rect 156524 74428 156530 74430
rect 189625 74427 189691 74430
rect 100201 74354 100267 74357
rect 133781 74354 133847 74357
rect 100201 74352 133847 74354
rect 100201 74296 100206 74352
rect 100262 74296 133786 74352
rect 133842 74296 133847 74352
rect 100201 74294 133847 74296
rect 100201 74291 100267 74294
rect 133781 74291 133847 74294
rect 143901 74356 143967 74357
rect 143901 74352 143948 74356
rect 144012 74354 144018 74356
rect 156045 74354 156111 74357
rect 156781 74354 156847 74357
rect 181110 74354 181116 74356
rect 143901 74296 143906 74352
rect 143901 74292 143948 74296
rect 144012 74294 144058 74354
rect 156045 74352 181116 74354
rect 156045 74296 156050 74352
rect 156106 74296 156786 74352
rect 156842 74296 181116 74352
rect 156045 74294 181116 74296
rect 144012 74292 144018 74294
rect 143901 74291 143967 74292
rect 156045 74291 156111 74294
rect 156781 74291 156847 74294
rect 181110 74292 181116 74294
rect 181180 74292 181186 74356
rect 107285 74218 107351 74221
rect 136265 74218 136331 74221
rect 103470 74216 136331 74218
rect 103470 74160 107290 74216
rect 107346 74160 136270 74216
rect 136326 74160 136331 74216
rect 103470 74158 136331 74160
rect 54477 73946 54543 73949
rect 103470 73946 103530 74158
rect 107285 74155 107351 74158
rect 136265 74155 136331 74158
rect 161197 74220 161263 74221
rect 161197 74216 161244 74220
rect 161308 74218 161314 74220
rect 174721 74218 174787 74221
rect 175089 74218 175155 74221
rect 198958 74218 198964 74220
rect 161197 74160 161202 74216
rect 161197 74156 161244 74160
rect 161308 74158 161354 74218
rect 174721 74216 198964 74218
rect 174721 74160 174726 74216
rect 174782 74160 175094 74216
rect 175150 74160 198964 74216
rect 174721 74158 198964 74160
rect 161308 74156 161314 74158
rect 161197 74155 161263 74156
rect 174721 74155 174787 74158
rect 175089 74155 175155 74158
rect 198958 74156 198964 74158
rect 199028 74156 199034 74220
rect 116853 74082 116919 74085
rect 144126 74082 144132 74084
rect 116853 74080 144132 74082
rect 116853 74024 116858 74080
rect 116914 74024 144132 74080
rect 116853 74022 144132 74024
rect 116853 74019 116919 74022
rect 144126 74020 144132 74022
rect 144196 74020 144202 74084
rect 54477 73944 103530 73946
rect 54477 73888 54482 73944
rect 54538 73888 103530 73944
rect 54477 73886 103530 73888
rect 135069 73946 135135 73949
rect 135662 73946 135668 73948
rect 135069 73944 135668 73946
rect 135069 73888 135074 73944
rect 135130 73888 135668 73944
rect 135069 73886 135668 73888
rect 54477 73883 54543 73886
rect 135069 73883 135135 73886
rect 135662 73884 135668 73886
rect 135732 73884 135738 73948
rect 149646 73884 149652 73948
rect 149716 73946 149722 73948
rect 229737 73946 229803 73949
rect 149716 73944 229803 73946
rect 149716 73888 229742 73944
rect 229798 73888 229803 73944
rect 149716 73886 229803 73888
rect 149716 73884 149722 73886
rect 229737 73883 229803 73886
rect 21357 73810 21423 73813
rect 100201 73810 100267 73813
rect 21357 73808 100267 73810
rect 21357 73752 21362 73808
rect 21418 73752 100206 73808
rect 100262 73752 100267 73808
rect 21357 73750 100267 73752
rect 21357 73747 21423 73750
rect 100201 73747 100267 73750
rect 135294 73748 135300 73812
rect 135364 73810 135370 73812
rect 136449 73810 136515 73813
rect 135364 73808 136515 73810
rect 135364 73752 136454 73808
rect 136510 73752 136515 73808
rect 135364 73750 136515 73752
rect 135364 73748 135370 73750
rect 136449 73747 136515 73750
rect 152641 73810 152707 73813
rect 152958 73810 152964 73812
rect 152641 73808 152964 73810
rect 152641 73752 152646 73808
rect 152702 73752 152964 73808
rect 152641 73750 152964 73752
rect 152641 73747 152707 73750
rect 152958 73748 152964 73750
rect 153028 73748 153034 73812
rect 167453 73810 167519 73813
rect 167678 73810 167684 73812
rect 167453 73808 167684 73810
rect 167453 73752 167458 73808
rect 167514 73752 167684 73808
rect 167453 73750 167684 73752
rect 167453 73747 167519 73750
rect 167678 73748 167684 73750
rect 167748 73748 167754 73812
rect 173157 73810 173223 73813
rect 173750 73810 173756 73812
rect 173157 73808 173756 73810
rect 173157 73752 173162 73808
rect 173218 73752 173756 73808
rect 173157 73750 173756 73752
rect 173157 73747 173223 73750
rect 173750 73748 173756 73750
rect 173820 73748 173826 73812
rect 189625 73810 189691 73813
rect 304993 73810 305059 73813
rect 189625 73808 305059 73810
rect 189625 73752 189630 73808
rect 189686 73752 304998 73808
rect 305054 73752 305059 73808
rect 189625 73750 305059 73752
rect 189625 73747 189691 73750
rect 304993 73747 305059 73750
rect 166625 73674 166691 73677
rect 166758 73674 166764 73676
rect 166625 73672 166764 73674
rect 166625 73616 166630 73672
rect 166686 73616 166764 73672
rect 166625 73614 166764 73616
rect 166625 73611 166691 73614
rect 166758 73612 166764 73614
rect 166828 73612 166834 73676
rect 152590 73476 152596 73540
rect 152660 73538 152666 73540
rect 152917 73538 152983 73541
rect 152660 73536 152983 73538
rect 152660 73480 152922 73536
rect 152978 73480 152983 73536
rect 152660 73478 152983 73480
rect 152660 73476 152666 73478
rect 152917 73475 152983 73478
rect 168046 73476 168052 73540
rect 168116 73538 168122 73540
rect 180241 73538 180307 73541
rect 168116 73536 180307 73538
rect 168116 73480 180246 73536
rect 180302 73480 180307 73536
rect 168116 73478 180307 73480
rect 168116 73476 168122 73478
rect 180241 73475 180307 73478
rect 167545 73402 167611 73405
rect 168046 73402 168052 73404
rect 167545 73400 168052 73402
rect 167545 73344 167550 73400
rect 167606 73344 168052 73400
rect 167545 73342 168052 73344
rect 167545 73339 167611 73342
rect 168046 73340 168052 73342
rect 168116 73340 168122 73404
rect 121310 73068 121316 73132
rect 121380 73130 121386 73132
rect 154021 73130 154087 73133
rect 121380 73128 154087 73130
rect 121380 73072 154026 73128
rect 154082 73072 154087 73128
rect 121380 73070 154087 73072
rect 121380 73068 121386 73070
rect 154021 73067 154087 73070
rect 156229 73130 156295 73133
rect 156965 73130 157031 73133
rect 179689 73132 179755 73133
rect 179638 73130 179644 73132
rect 156229 73128 157031 73130
rect 156229 73072 156234 73128
rect 156290 73072 156970 73128
rect 157026 73072 157031 73128
rect 156229 73070 157031 73072
rect 179598 73070 179644 73130
rect 179708 73128 179755 73132
rect 179750 73072 179755 73128
rect 156229 73067 156295 73070
rect 156965 73067 157031 73070
rect 179638 73068 179644 73070
rect 179708 73068 179755 73072
rect 180926 73068 180932 73132
rect 180996 73130 181002 73132
rect 181253 73130 181319 73133
rect 180996 73128 181319 73130
rect 180996 73072 181258 73128
rect 181314 73072 181319 73128
rect 180996 73070 181319 73072
rect 180996 73068 181002 73070
rect 179689 73067 179755 73068
rect 181253 73067 181319 73070
rect 119981 72994 120047 72997
rect 152590 72994 152596 72996
rect 119981 72992 152596 72994
rect 119981 72936 119986 72992
rect 120042 72936 152596 72992
rect 119981 72934 152596 72936
rect 119981 72931 120047 72934
rect 152590 72932 152596 72934
rect 152660 72932 152666 72996
rect 156505 72994 156571 72997
rect 183870 72994 183876 72996
rect 156505 72992 183876 72994
rect 156505 72936 156510 72992
rect 156566 72936 183876 72992
rect 156505 72934 183876 72936
rect 156505 72931 156571 72934
rect 183870 72932 183876 72934
rect 183940 72932 183946 72996
rect 579981 72994 580047 72997
rect 583520 72994 584960 73084
rect 579981 72992 584960 72994
rect 579981 72936 579986 72992
rect 580042 72936 584960 72992
rect 579981 72934 584960 72936
rect 579981 72931 580047 72934
rect 119889 72858 119955 72861
rect 149278 72858 149284 72860
rect 119889 72856 149284 72858
rect 119889 72800 119894 72856
rect 119950 72800 149284 72856
rect 119889 72798 149284 72800
rect 119889 72795 119955 72798
rect 149278 72796 149284 72798
rect 149348 72858 149354 72860
rect 149830 72858 149836 72860
rect 149348 72798 149836 72858
rect 149348 72796 149354 72798
rect 149830 72796 149836 72798
rect 149900 72796 149906 72860
rect 156873 72858 156939 72861
rect 183134 72858 183140 72860
rect 156830 72856 183140 72858
rect 156830 72800 156878 72856
rect 156934 72800 183140 72856
rect 156830 72798 183140 72800
rect 156830 72795 156939 72798
rect 183134 72796 183140 72798
rect 183204 72796 183210 72860
rect 583520 72844 584960 72934
rect 131021 72586 131087 72589
rect 142286 72586 142292 72588
rect 131021 72584 142292 72586
rect 131021 72528 131026 72584
rect 131082 72528 142292 72584
rect 131021 72526 142292 72528
rect 131021 72523 131087 72526
rect 142286 72524 142292 72526
rect 142356 72524 142362 72588
rect 11053 72450 11119 72453
rect 133229 72450 133295 72453
rect 11053 72448 133295 72450
rect 11053 72392 11058 72448
rect 11114 72392 133234 72448
rect 133290 72392 133295 72448
rect 11053 72390 133295 72392
rect 156830 72450 156890 72795
rect 156965 72722 157031 72725
rect 179822 72722 179828 72724
rect 156965 72720 179828 72722
rect 156965 72664 156970 72720
rect 157026 72664 179828 72720
rect 156965 72662 179828 72664
rect 156965 72659 157031 72662
rect 179822 72660 179828 72662
rect 179892 72660 179898 72724
rect 157057 72586 157123 72589
rect 185158 72586 185164 72588
rect 157057 72584 185164 72586
rect 157057 72528 157062 72584
rect 157118 72528 185164 72584
rect 157057 72526 185164 72528
rect 157057 72523 157123 72526
rect 185158 72524 185164 72526
rect 185228 72524 185234 72588
rect 157057 72450 157123 72453
rect 156830 72448 157123 72450
rect 156830 72392 157062 72448
rect 157118 72392 157123 72448
rect 156830 72390 157123 72392
rect 11053 72387 11119 72390
rect 133229 72387 133295 72390
rect 157057 72387 157123 72390
rect 169702 72388 169708 72452
rect 169772 72450 169778 72452
rect 178401 72450 178467 72453
rect 169772 72448 178467 72450
rect 169772 72392 178406 72448
rect 178462 72392 178467 72448
rect 169772 72390 178467 72392
rect 169772 72388 169778 72390
rect 178401 72387 178467 72390
rect 156505 72314 156571 72317
rect 156965 72314 157031 72317
rect 156505 72312 157031 72314
rect 156505 72256 156510 72312
rect 156566 72256 156970 72312
rect 157026 72256 157031 72312
rect 156505 72254 157031 72256
rect 156505 72251 156571 72254
rect 156965 72251 157031 72254
rect 158846 71844 158852 71908
rect 158916 71906 158922 71908
rect 159725 71906 159791 71909
rect 158916 71904 159791 71906
rect 158916 71848 159730 71904
rect 159786 71848 159791 71904
rect 158916 71846 159791 71848
rect 158916 71844 158922 71846
rect 159725 71843 159791 71846
rect 114921 71770 114987 71773
rect 162485 71772 162551 71773
rect 149094 71770 149100 71772
rect 114921 71768 149100 71770
rect -960 71634 480 71724
rect 114921 71712 114926 71768
rect 114982 71712 149100 71768
rect 114921 71710 149100 71712
rect 114921 71707 114987 71710
rect 149094 71708 149100 71710
rect 149164 71708 149170 71772
rect 162485 71768 162532 71772
rect 162596 71770 162602 71772
rect 175457 71770 175523 71773
rect 202413 71770 202479 71773
rect 202781 71770 202847 71773
rect 162485 71712 162490 71768
rect 162485 71708 162532 71712
rect 162596 71710 162642 71770
rect 175457 71768 202847 71770
rect 175457 71712 175462 71768
rect 175518 71712 202418 71768
rect 202474 71712 202786 71768
rect 202842 71712 202847 71768
rect 175457 71710 202847 71712
rect 162596 71708 162602 71710
rect 162485 71707 162551 71708
rect 175457 71707 175523 71710
rect 202413 71707 202479 71710
rect 202781 71707 202847 71710
rect 3509 71634 3575 71637
rect -960 71632 3575 71634
rect -960 71576 3514 71632
rect 3570 71576 3575 71632
rect -960 71574 3575 71576
rect -960 71484 480 71574
rect 3509 71571 3575 71574
rect 120022 71572 120028 71636
rect 120092 71634 120098 71636
rect 153561 71634 153627 71637
rect 120092 71632 153627 71634
rect 120092 71576 153566 71632
rect 153622 71576 153627 71632
rect 120092 71574 153627 71576
rect 120092 71572 120098 71574
rect 153561 71571 153627 71574
rect 118550 71436 118556 71500
rect 118620 71498 118626 71500
rect 152406 71498 152412 71500
rect 118620 71438 152412 71498
rect 118620 71436 118626 71438
rect 152406 71436 152412 71438
rect 152476 71436 152482 71500
rect 111701 71362 111767 71365
rect 145046 71362 145052 71364
rect 111701 71360 145052 71362
rect 111701 71304 111706 71360
rect 111762 71304 145052 71360
rect 111701 71302 145052 71304
rect 111701 71299 111767 71302
rect 145046 71300 145052 71302
rect 145116 71300 145122 71364
rect 166942 71300 166948 71364
rect 167012 71362 167018 71364
rect 172421 71362 172487 71365
rect 167012 71360 172487 71362
rect 167012 71304 172426 71360
rect 172482 71304 172487 71360
rect 167012 71302 172487 71304
rect 167012 71300 167018 71302
rect 172421 71299 172487 71302
rect 112805 71226 112871 71229
rect 145598 71226 145604 71228
rect 112805 71224 145604 71226
rect 112805 71168 112810 71224
rect 112866 71168 145604 71224
rect 112805 71166 145604 71168
rect 112805 71163 112871 71166
rect 145598 71164 145604 71166
rect 145668 71164 145674 71228
rect 148910 71028 148916 71092
rect 148980 71090 148986 71092
rect 200757 71090 200823 71093
rect 148980 71088 200823 71090
rect 148980 71032 200762 71088
rect 200818 71032 200823 71088
rect 148980 71030 200823 71032
rect 148980 71028 148986 71030
rect 200757 71027 200823 71030
rect 202781 71090 202847 71093
rect 543733 71090 543799 71093
rect 202781 71088 543799 71090
rect 202781 71032 202786 71088
rect 202842 71032 543738 71088
rect 543794 71032 543799 71088
rect 202781 71030 543799 71032
rect 202781 71027 202847 71030
rect 543733 71027 543799 71030
rect 144310 70546 144316 70548
rect 122790 70486 144316 70546
rect 113909 70274 113975 70277
rect 122790 70274 122850 70486
rect 144310 70484 144316 70486
rect 144380 70546 144386 70548
rect 144821 70546 144887 70549
rect 144380 70544 144887 70546
rect 144380 70488 144826 70544
rect 144882 70488 144887 70544
rect 144380 70486 144887 70488
rect 144380 70484 144386 70486
rect 144821 70483 144887 70486
rect 195145 70412 195211 70413
rect 195094 70410 195100 70412
rect 195054 70350 195100 70410
rect 195164 70408 195211 70412
rect 195206 70352 195211 70408
rect 195094 70348 195100 70350
rect 195164 70348 195211 70352
rect 195145 70347 195211 70348
rect 113909 70272 122850 70274
rect 113909 70216 113914 70272
rect 113970 70216 122850 70272
rect 113909 70214 122850 70216
rect 166441 70274 166507 70277
rect 166901 70274 166967 70277
rect 191598 70274 191604 70276
rect 166441 70272 191604 70274
rect 166441 70216 166446 70272
rect 166502 70216 166906 70272
rect 166962 70216 191604 70272
rect 166441 70214 191604 70216
rect 113909 70211 113975 70214
rect 166441 70211 166507 70214
rect 166901 70211 166967 70214
rect 191598 70212 191604 70214
rect 191668 70212 191674 70276
rect 166625 70138 166691 70141
rect 166942 70138 166948 70140
rect 166625 70136 166948 70138
rect 166625 70080 166630 70136
rect 166686 70080 166948 70136
rect 166625 70078 166948 70080
rect 166625 70075 166691 70078
rect 166942 70076 166948 70078
rect 167012 70076 167018 70140
rect 176101 70138 176167 70141
rect 176101 70136 200130 70138
rect 176101 70080 176106 70136
rect 176162 70080 200130 70136
rect 176101 70078 200130 70080
rect 176101 70075 176167 70078
rect 200070 69594 200130 70078
rect 200798 69594 200804 69596
rect 200070 69534 200804 69594
rect 200798 69532 200804 69534
rect 200868 69594 200874 69596
rect 561673 69594 561739 69597
rect 200868 69592 561739 69594
rect 200868 69536 561678 69592
rect 561734 69536 561739 69592
rect 200868 69534 561739 69536
rect 200868 69532 200874 69534
rect 561673 69531 561739 69534
rect 169150 68988 169156 69052
rect 169220 69050 169226 69052
rect 183829 69050 183895 69053
rect 169220 69048 183895 69050
rect 169220 68992 183834 69048
rect 183890 68992 183895 69048
rect 169220 68990 183895 68992
rect 169220 68988 169226 68990
rect 183829 68987 183895 68990
rect 120942 68852 120948 68916
rect 121012 68914 121018 68916
rect 154757 68914 154823 68917
rect 121012 68912 154823 68914
rect 121012 68856 154762 68912
rect 154818 68856 154823 68912
rect 121012 68854 154823 68856
rect 121012 68852 121018 68854
rect 154757 68851 154823 68854
rect 171777 68914 171843 68917
rect 199193 68914 199259 68917
rect 171777 68912 199259 68914
rect 171777 68856 171782 68912
rect 171838 68856 199198 68912
rect 199254 68856 199259 68912
rect 171777 68854 199259 68856
rect 171777 68851 171843 68854
rect 199193 68851 199259 68854
rect 200982 68852 200988 68916
rect 201052 68914 201058 68916
rect 201401 68914 201467 68917
rect 201052 68912 201467 68914
rect 201052 68856 201406 68912
rect 201462 68856 201467 68912
rect 201052 68854 201467 68856
rect 201052 68852 201058 68854
rect 201401 68851 201467 68854
rect 111333 68778 111399 68781
rect 144545 68780 144611 68781
rect 188245 68780 188311 68781
rect 144494 68778 144500 68780
rect 111333 68776 144500 68778
rect 144564 68776 144611 68780
rect 111333 68720 111338 68776
rect 111394 68720 144500 68776
rect 144606 68720 144611 68776
rect 111333 68718 144500 68720
rect 111333 68715 111399 68718
rect 144494 68716 144500 68718
rect 144564 68716 144611 68720
rect 150014 68716 150020 68780
rect 150084 68778 150090 68780
rect 179454 68778 179460 68780
rect 150084 68718 179460 68778
rect 150084 68716 150090 68718
rect 179454 68716 179460 68718
rect 179524 68778 179530 68780
rect 179524 68718 180810 68778
rect 179524 68716 179530 68718
rect 144545 68715 144611 68716
rect 115841 68642 115907 68645
rect 148174 68642 148180 68644
rect 115841 68640 148180 68642
rect 115841 68584 115846 68640
rect 115902 68584 148180 68640
rect 115841 68582 148180 68584
rect 115841 68579 115907 68582
rect 148174 68580 148180 68582
rect 148244 68580 148250 68644
rect 112897 68506 112963 68509
rect 143349 68506 143415 68509
rect 144678 68506 144684 68508
rect 112897 68504 144684 68506
rect 112897 68448 112902 68504
rect 112958 68448 143354 68504
rect 143410 68448 144684 68504
rect 112897 68446 144684 68448
rect 112897 68443 112963 68446
rect 143349 68443 143415 68446
rect 144678 68444 144684 68446
rect 144748 68444 144754 68508
rect 110045 68370 110111 68373
rect 115933 68370 115999 68373
rect 140814 68370 140820 68372
rect 110045 68368 140820 68370
rect 110045 68312 110050 68368
rect 110106 68312 115938 68368
rect 115994 68312 140820 68368
rect 110045 68310 140820 68312
rect 110045 68307 110111 68310
rect 115933 68307 115999 68310
rect 140814 68308 140820 68310
rect 140884 68308 140890 68372
rect 180750 68370 180810 68718
rect 188245 68776 188292 68780
rect 188356 68778 188362 68780
rect 188245 68720 188250 68776
rect 188245 68716 188292 68720
rect 188356 68718 188402 68778
rect 188356 68716 188362 68718
rect 188245 68715 188311 68716
rect 220813 68370 220879 68373
rect 180750 68368 220879 68370
rect 180750 68312 220818 68368
rect 220874 68312 220879 68368
rect 180750 68310 220879 68312
rect 220813 68307 220879 68310
rect 8937 68234 9003 68237
rect 131614 68234 131620 68236
rect 8937 68232 131620 68234
rect 8937 68176 8942 68232
rect 8998 68176 131620 68232
rect 8937 68174 131620 68176
rect 8937 68171 9003 68174
rect 131614 68172 131620 68174
rect 131684 68172 131690 68236
rect 147070 68172 147076 68236
rect 147140 68234 147146 68236
rect 189717 68234 189783 68237
rect 147140 68232 189783 68234
rect 147140 68176 189722 68232
rect 189778 68176 189783 68232
rect 147140 68174 189783 68176
rect 147140 68172 147146 68174
rect 189717 68171 189783 68174
rect 199193 68234 199259 68237
rect 504357 68234 504423 68237
rect 199193 68232 504423 68234
rect 199193 68176 199198 68232
rect 199254 68176 504362 68232
rect 504418 68176 504423 68232
rect 199193 68174 504423 68176
rect 199193 68171 199259 68174
rect 504357 68171 504423 68174
rect 160921 67692 160987 67693
rect 160870 67690 160876 67692
rect 160830 67630 160876 67690
rect 160940 67688 160987 67692
rect 160982 67632 160987 67688
rect 160870 67628 160876 67630
rect 160940 67628 160987 67632
rect 160921 67627 160987 67628
rect 107377 67554 107443 67557
rect 138606 67554 138612 67556
rect 103470 67552 138612 67554
rect 103470 67496 107382 67552
rect 107438 67496 138612 67552
rect 103470 67494 138612 67496
rect 80053 67010 80119 67013
rect 103470 67010 103530 67494
rect 107377 67491 107443 67494
rect 138606 67492 138612 67494
rect 138676 67492 138682 67556
rect 161013 67554 161079 67557
rect 161238 67554 161244 67556
rect 161013 67552 161244 67554
rect 161013 67496 161018 67552
rect 161074 67496 161244 67552
rect 161013 67494 161244 67496
rect 161013 67491 161079 67494
rect 161238 67492 161244 67494
rect 161308 67492 161314 67556
rect 165981 67554 166047 67557
rect 200297 67554 200363 67557
rect 201401 67554 201467 67557
rect 165981 67552 201467 67554
rect 165981 67496 165986 67552
rect 166042 67496 200302 67552
rect 200358 67496 201406 67552
rect 201462 67496 201467 67552
rect 165981 67494 201467 67496
rect 165981 67491 166047 67494
rect 200297 67491 200363 67494
rect 201401 67491 201467 67494
rect 151302 67356 151308 67420
rect 151372 67418 151378 67420
rect 182582 67418 182588 67420
rect 151372 67358 182588 67418
rect 151372 67356 151378 67358
rect 182582 67356 182588 67358
rect 182652 67418 182658 67420
rect 242893 67418 242959 67421
rect 182652 67416 242959 67418
rect 182652 67360 242898 67416
rect 242954 67360 242959 67416
rect 182652 67358 242959 67360
rect 182652 67356 182658 67358
rect 242893 67355 242959 67358
rect 148358 67220 148364 67284
rect 148428 67282 148434 67284
rect 213913 67282 213979 67285
rect 148428 67280 213979 67282
rect 148428 67224 213918 67280
rect 213974 67224 213979 67280
rect 148428 67222 213979 67224
rect 148428 67220 148434 67222
rect 213913 67219 213979 67222
rect 165889 67146 165955 67149
rect 197905 67146 197971 67149
rect 423673 67146 423739 67149
rect 165889 67144 423739 67146
rect 165889 67088 165894 67144
rect 165950 67088 197910 67144
rect 197966 67088 423678 67144
rect 423734 67088 423739 67144
rect 165889 67086 423739 67088
rect 165889 67083 165955 67086
rect 197905 67083 197971 67086
rect 423673 67083 423739 67086
rect 80053 67008 103530 67010
rect 80053 66952 80058 67008
rect 80114 66952 103530 67008
rect 80053 66950 103530 66952
rect 112345 67010 112411 67013
rect 133873 67010 133939 67013
rect 137502 67010 137508 67012
rect 112345 67008 137508 67010
rect 112345 66952 112350 67008
rect 112406 66952 133878 67008
rect 133934 66952 137508 67008
rect 112345 66950 137508 66952
rect 80053 66947 80119 66950
rect 112345 66947 112411 66950
rect 133873 66947 133939 66950
rect 137502 66948 137508 66950
rect 137572 66948 137578 67012
rect 201401 67010 201467 67013
rect 430573 67010 430639 67013
rect 201401 67008 430639 67010
rect 201401 66952 201406 67008
rect 201462 66952 430578 67008
rect 430634 66952 430639 67008
rect 201401 66950 430639 66952
rect 201401 66947 201467 66950
rect 430573 66947 430639 66950
rect 24853 66874 24919 66877
rect 133822 66874 133828 66876
rect 24853 66872 133828 66874
rect 24853 66816 24858 66872
rect 24914 66816 133828 66872
rect 24853 66814 133828 66816
rect 24853 66811 24919 66814
rect 133822 66812 133828 66814
rect 133892 66812 133898 66876
rect 146886 66812 146892 66876
rect 146956 66874 146962 66876
rect 193857 66874 193923 66877
rect 200614 66874 200620 66876
rect 146956 66872 193923 66874
rect 146956 66816 193862 66872
rect 193918 66816 193923 66872
rect 146956 66814 193923 66816
rect 146956 66812 146962 66814
rect 193857 66811 193923 66814
rect 200070 66814 200620 66874
rect 176142 66676 176148 66740
rect 176212 66738 176218 66740
rect 200070 66738 200130 66814
rect 200614 66812 200620 66814
rect 200684 66874 200690 66876
rect 557533 66874 557599 66877
rect 200684 66872 557599 66874
rect 200684 66816 557538 66872
rect 557594 66816 557599 66872
rect 200684 66814 557599 66816
rect 200684 66812 200690 66814
rect 557533 66811 557599 66814
rect 176212 66678 200130 66738
rect 176212 66676 176218 66678
rect 108849 66194 108915 66197
rect 139894 66194 139900 66196
rect 103470 66192 139900 66194
rect 103470 66136 108854 66192
rect 108910 66136 139900 66192
rect 103470 66134 139900 66136
rect 93853 65786 93919 65789
rect 103470 65786 103530 66134
rect 108849 66131 108915 66134
rect 139894 66132 139900 66134
rect 139964 66132 139970 66196
rect 181161 66194 181227 66197
rect 188061 66196 188127 66197
rect 187918 66194 187924 66196
rect 181161 66192 187924 66194
rect 181161 66136 181166 66192
rect 181222 66136 187924 66192
rect 181161 66134 187924 66136
rect 181161 66131 181227 66134
rect 187918 66132 187924 66134
rect 187988 66132 187994 66196
rect 188061 66192 188108 66196
rect 188172 66194 188178 66196
rect 188061 66136 188066 66192
rect 188061 66132 188108 66136
rect 188172 66134 188218 66194
rect 188172 66132 188178 66134
rect 188061 66131 188127 66132
rect 139710 66058 139716 66060
rect 93853 65784 103530 65786
rect 93853 65728 93858 65784
rect 93914 65728 103530 65784
rect 93853 65726 103530 65728
rect 113130 65998 139716 66058
rect 93853 65723 93919 65726
rect 93117 65650 93183 65653
rect 111517 65650 111583 65653
rect 113130 65650 113190 65998
rect 139710 65996 139716 65998
rect 139780 65996 139786 66060
rect 161974 65996 161980 66060
rect 162044 66058 162050 66060
rect 196157 66058 196223 66061
rect 196433 66058 196499 66061
rect 162044 66056 196499 66058
rect 162044 66000 196162 66056
rect 196218 66000 196438 66056
rect 196494 66000 196499 66056
rect 162044 65998 196499 66000
rect 162044 65996 162050 65998
rect 196157 65995 196223 65998
rect 196433 65995 196499 65998
rect 93117 65648 113190 65650
rect 93117 65592 93122 65648
rect 93178 65592 111522 65648
rect 111578 65592 113190 65648
rect 93117 65590 113190 65592
rect 93117 65587 93183 65590
rect 111517 65587 111583 65590
rect 187918 65588 187924 65652
rect 187988 65650 187994 65652
rect 274633 65650 274699 65653
rect 187988 65648 274699 65650
rect 187988 65592 274638 65648
rect 274694 65592 274699 65648
rect 187988 65590 274699 65592
rect 187988 65588 187994 65590
rect 274633 65587 274699 65590
rect 7649 65514 7715 65517
rect 133086 65514 133092 65516
rect 7649 65512 133092 65514
rect 7649 65456 7654 65512
rect 7710 65456 133092 65512
rect 7649 65454 133092 65456
rect 7649 65451 7715 65454
rect 133086 65452 133092 65454
rect 133156 65452 133162 65516
rect 196433 65514 196499 65517
rect 380893 65514 380959 65517
rect 196433 65512 380959 65514
rect 196433 65456 196438 65512
rect 196494 65456 380898 65512
rect 380954 65456 380959 65512
rect 196433 65454 380959 65456
rect 196433 65451 196499 65454
rect 380893 65451 380959 65454
rect 188102 65044 188108 65108
rect 188172 65106 188178 65108
rect 188613 65106 188679 65109
rect 197537 65108 197603 65109
rect 188172 65104 188679 65106
rect 188172 65048 188618 65104
rect 188674 65048 188679 65104
rect 188172 65046 188679 65048
rect 188172 65044 188178 65046
rect 188613 65043 188679 65046
rect 197486 65044 197492 65108
rect 197556 65106 197603 65108
rect 197556 65104 197648 65106
rect 197598 65048 197648 65104
rect 197556 65046 197648 65048
rect 197556 65044 197603 65046
rect 197537 65043 197603 65044
rect 102225 64834 102291 64837
rect 103329 64834 103395 64837
rect 135846 64834 135852 64836
rect 102225 64832 135852 64834
rect 102225 64776 102230 64832
rect 102286 64776 103334 64832
rect 103390 64776 135852 64832
rect 102225 64774 135852 64776
rect 102225 64771 102291 64774
rect 103329 64771 103395 64774
rect 135846 64772 135852 64774
rect 135916 64772 135922 64836
rect 152958 64772 152964 64836
rect 153028 64834 153034 64836
rect 208393 64834 208459 64837
rect 153028 64832 208459 64834
rect 153028 64776 208398 64832
rect 208454 64776 208459 64832
rect 153028 64774 208459 64776
rect 153028 64772 153034 64774
rect 208393 64771 208459 64774
rect 174670 64636 174676 64700
rect 174740 64698 174746 64700
rect 201718 64698 201724 64700
rect 174740 64638 201724 64698
rect 174740 64636 174746 64638
rect 201718 64636 201724 64638
rect 201788 64636 201794 64700
rect 171910 64500 171916 64564
rect 171980 64562 171986 64564
rect 197302 64562 197308 64564
rect 171980 64502 197308 64562
rect 171980 64500 171986 64502
rect 197302 64500 197308 64502
rect 197372 64562 197378 64564
rect 197372 64502 200130 64562
rect 197372 64500 197378 64502
rect 200070 64290 200130 64502
rect 208393 64426 208459 64429
rect 259453 64426 259519 64429
rect 208393 64424 259519 64426
rect 208393 64368 208398 64424
rect 208454 64368 259458 64424
rect 259514 64368 259519 64424
rect 208393 64366 259519 64368
rect 208393 64363 208459 64366
rect 259453 64363 259519 64366
rect 511993 64290 512059 64293
rect 200070 64288 512059 64290
rect 200070 64232 511998 64288
rect 512054 64232 512059 64288
rect 200070 64230 512059 64232
rect 511993 64227 512059 64230
rect 46197 64154 46263 64157
rect 102225 64154 102291 64157
rect 46197 64152 102291 64154
rect 46197 64096 46202 64152
rect 46258 64096 102230 64152
rect 102286 64096 102291 64152
rect 46197 64094 102291 64096
rect 46197 64091 46263 64094
rect 102225 64091 102291 64094
rect 201718 64092 201724 64156
rect 201788 64154 201794 64156
rect 547873 64154 547939 64157
rect 201788 64152 547939 64154
rect 201788 64096 547878 64152
rect 547934 64096 547939 64152
rect 201788 64094 547939 64096
rect 201788 64092 201794 64094
rect 547873 64091 547939 64094
rect 108113 63474 108179 63477
rect 139526 63474 139532 63476
rect 108113 63472 139532 63474
rect 108113 63416 108118 63472
rect 108174 63416 139532 63472
rect 108113 63414 139532 63416
rect 108113 63411 108179 63414
rect 139526 63412 139532 63414
rect 139596 63412 139602 63476
rect 157926 63412 157932 63476
rect 157996 63474 158002 63476
rect 192017 63474 192083 63477
rect 193121 63474 193187 63477
rect 157996 63472 193187 63474
rect 157996 63416 192022 63472
rect 192078 63416 193126 63472
rect 193182 63416 193187 63472
rect 157996 63414 193187 63416
rect 157996 63412 158002 63414
rect 192017 63411 192083 63414
rect 193121 63411 193187 63414
rect 110321 63338 110387 63341
rect 138422 63338 138428 63340
rect 110321 63336 138428 63338
rect 110321 63280 110326 63336
rect 110382 63280 138428 63336
rect 110321 63278 138428 63280
rect 110321 63275 110387 63278
rect 138422 63276 138428 63278
rect 138492 63276 138498 63340
rect 155033 63338 155099 63341
rect 189073 63338 189139 63341
rect 292573 63338 292639 63341
rect 155033 63336 292639 63338
rect 155033 63280 155038 63336
rect 155094 63280 189078 63336
rect 189134 63280 292578 63336
rect 292634 63280 292639 63336
rect 155033 63278 292639 63280
rect 155033 63275 155099 63278
rect 189073 63275 189139 63278
rect 292573 63275 292639 63278
rect 193121 63202 193187 63205
rect 331213 63202 331279 63205
rect 193121 63200 331279 63202
rect 193121 63144 193126 63200
rect 193182 63144 331218 63200
rect 331274 63144 331279 63200
rect 193121 63142 331279 63144
rect 193121 63139 193187 63142
rect 331213 63139 331279 63142
rect 165102 63004 165108 63068
rect 165172 63066 165178 63068
rect 198917 63066 198983 63069
rect 414657 63066 414723 63069
rect 165172 63064 414723 63066
rect 165172 63008 198922 63064
rect 198978 63008 414662 63064
rect 414718 63008 414723 63064
rect 165172 63006 414723 63008
rect 165172 63004 165178 63006
rect 198917 63003 198983 63006
rect 414657 63003 414723 63006
rect 92473 62930 92539 62933
rect 108113 62930 108179 62933
rect 92473 62928 108179 62930
rect 92473 62872 92478 62928
rect 92534 62872 108118 62928
rect 108174 62872 108179 62928
rect 92473 62870 108179 62872
rect 92473 62867 92539 62870
rect 108113 62867 108179 62870
rect 172094 62868 172100 62932
rect 172164 62930 172170 62932
rect 196566 62930 196572 62932
rect 172164 62870 196572 62930
rect 172164 62868 172170 62870
rect 196566 62868 196572 62870
rect 196636 62930 196642 62932
rect 514017 62930 514083 62933
rect 196636 62928 514083 62930
rect 196636 62872 514022 62928
rect 514078 62872 514083 62928
rect 196636 62870 514083 62872
rect 196636 62868 196642 62870
rect 514017 62867 514083 62870
rect 75177 62794 75243 62797
rect 110321 62794 110387 62797
rect 75177 62792 110387 62794
rect 75177 62736 75182 62792
rect 75238 62736 110326 62792
rect 110382 62736 110387 62792
rect 75177 62734 110387 62736
rect 75177 62731 75243 62734
rect 110321 62731 110387 62734
rect 176326 62732 176332 62796
rect 176396 62794 176402 62796
rect 201902 62794 201908 62796
rect 176396 62734 201908 62794
rect 176396 62732 176402 62734
rect 201902 62732 201908 62734
rect 201972 62794 201978 62796
rect 567837 62794 567903 62797
rect 201972 62792 567903 62794
rect 201972 62736 567842 62792
rect 567898 62736 567903 62792
rect 201972 62734 567903 62736
rect 201972 62732 201978 62734
rect 567837 62731 567903 62734
rect 151486 62052 151492 62116
rect 151556 62114 151562 62116
rect 183686 62114 183692 62116
rect 151556 62054 183692 62114
rect 151556 62052 151562 62054
rect 183686 62052 183692 62054
rect 183756 62114 183762 62116
rect 249793 62114 249859 62117
rect 183756 62112 249859 62114
rect 183756 62056 249798 62112
rect 249854 62056 249859 62112
rect 183756 62054 249859 62056
rect 183756 62052 183762 62054
rect 249793 62051 249859 62054
rect 154941 61978 155007 61981
rect 187734 61978 187740 61980
rect 154941 61976 187740 61978
rect 154941 61920 154946 61976
rect 155002 61920 187740 61976
rect 154941 61918 187740 61920
rect 154941 61915 155007 61918
rect 187734 61916 187740 61918
rect 187804 61978 187810 61980
rect 277393 61978 277459 61981
rect 187804 61976 277459 61978
rect 187804 61920 277398 61976
rect 277454 61920 277459 61976
rect 187804 61918 277459 61920
rect 187804 61916 187810 61918
rect 277393 61915 277459 61918
rect 156822 61780 156828 61844
rect 156892 61842 156898 61844
rect 191373 61842 191439 61845
rect 320173 61842 320239 61845
rect 156892 61840 320239 61842
rect 156892 61784 191378 61840
rect 191434 61784 320178 61840
rect 320234 61784 320239 61840
rect 156892 61782 320239 61784
rect 156892 61780 156898 61782
rect 191373 61779 191439 61782
rect 320173 61779 320239 61782
rect 163589 61706 163655 61709
rect 196065 61706 196131 61709
rect 382917 61706 382983 61709
rect 163589 61704 382983 61706
rect 163589 61648 163594 61704
rect 163650 61648 196070 61704
rect 196126 61648 382922 61704
rect 382978 61648 382983 61704
rect 163589 61646 382983 61648
rect 163589 61643 163655 61646
rect 196065 61643 196131 61646
rect 382917 61643 382983 61646
rect 183737 61570 183803 61573
rect 193673 61570 193739 61573
rect 437473 61570 437539 61573
rect 183737 61568 437539 61570
rect 183737 61512 183742 61568
rect 183798 61512 193678 61568
rect 193734 61512 437478 61568
rect 437534 61512 437539 61568
rect 183737 61510 437539 61512
rect 183737 61507 183803 61510
rect 193673 61507 193739 61510
rect 437473 61507 437539 61510
rect 168557 61434 168623 61437
rect 202045 61434 202111 61437
rect 459553 61434 459619 61437
rect 168557 61432 459619 61434
rect 168557 61376 168562 61432
rect 168618 61376 202050 61432
rect 202106 61376 459558 61432
rect 459614 61376 459619 61432
rect 168557 61374 459619 61376
rect 168557 61371 168623 61374
rect 202045 61371 202111 61374
rect 459553 61371 459619 61374
rect 151670 61236 151676 61300
rect 151740 61298 151746 61300
rect 180558 61298 180564 61300
rect 151740 61238 180564 61298
rect 151740 61236 151746 61238
rect 180558 61236 180564 61238
rect 180628 61298 180634 61300
rect 245653 61298 245719 61301
rect 180628 61296 245719 61298
rect 180628 61240 245658 61296
rect 245714 61240 245719 61296
rect 180628 61238 245719 61240
rect 180628 61236 180634 61238
rect 245653 61235 245719 61238
rect 103881 60618 103947 60621
rect 104801 60618 104867 60621
rect 138238 60618 138244 60620
rect 103881 60616 138244 60618
rect 103881 60560 103886 60616
rect 103942 60560 104806 60616
rect 104862 60560 138244 60616
rect 103881 60558 138244 60560
rect 103881 60555 103947 60558
rect 104801 60555 104867 60558
rect 138238 60556 138244 60558
rect 138308 60556 138314 60620
rect 155718 60556 155724 60620
rect 155788 60618 155794 60620
rect 189441 60618 189507 60621
rect 189625 60618 189691 60621
rect 155788 60616 189691 60618
rect 155788 60560 189446 60616
rect 189502 60560 189630 60616
rect 189686 60560 189691 60616
rect 155788 60558 189691 60560
rect 155788 60556 155794 60558
rect 189441 60555 189507 60558
rect 189625 60555 189691 60558
rect 158110 60420 158116 60484
rect 158180 60482 158186 60484
rect 190913 60482 190979 60485
rect 191741 60482 191807 60485
rect 158180 60480 191807 60482
rect 158180 60424 190918 60480
rect 190974 60424 191746 60480
rect 191802 60424 191807 60480
rect 158180 60422 191807 60424
rect 158180 60420 158186 60422
rect 190913 60419 190979 60422
rect 191741 60419 191807 60422
rect 173566 60284 173572 60348
rect 173636 60346 173642 60348
rect 198958 60346 198964 60348
rect 173636 60286 198964 60346
rect 173636 60284 173642 60286
rect 198958 60284 198964 60286
rect 199028 60284 199034 60348
rect 189625 60210 189691 60213
rect 299473 60210 299539 60213
rect 189625 60208 299539 60210
rect 189625 60152 189630 60208
rect 189686 60152 299478 60208
rect 299534 60152 299539 60208
rect 189625 60150 299539 60152
rect 189625 60147 189691 60150
rect 299473 60147 299539 60150
rect 191741 60074 191807 60077
rect 338113 60074 338179 60077
rect 191741 60072 338179 60074
rect 191741 60016 191746 60072
rect 191802 60016 338118 60072
rect 338174 60016 338179 60072
rect 191741 60014 338179 60016
rect 191741 60011 191807 60014
rect 338113 60011 338179 60014
rect 84193 59938 84259 59941
rect 103881 59938 103947 59941
rect 84193 59936 103947 59938
rect 84193 59880 84198 59936
rect 84254 59880 103886 59936
rect 103942 59880 103947 59936
rect 84193 59878 103947 59880
rect 84193 59875 84259 59878
rect 103881 59875 103947 59878
rect 147254 59876 147260 59940
rect 147324 59938 147330 59940
rect 193397 59938 193463 59941
rect 147324 59936 193463 59938
rect 147324 59880 193402 59936
rect 193458 59880 193463 59936
rect 147324 59878 193463 59880
rect 147324 59876 147330 59878
rect 193397 59875 193463 59878
rect 198958 59876 198964 59940
rect 199028 59938 199034 59940
rect 525057 59938 525123 59941
rect 199028 59936 525123 59938
rect 199028 59880 525062 59936
rect 525118 59880 525123 59936
rect 199028 59878 525123 59880
rect 199028 59876 199034 59878
rect 525057 59875 525123 59878
rect 580257 59666 580323 59669
rect 583520 59666 584960 59756
rect 580257 59664 584960 59666
rect 580257 59608 580262 59664
rect 580318 59608 584960 59664
rect 580257 59606 584960 59608
rect 580257 59603 580323 59606
rect 583520 59516 584960 59606
rect 107561 59258 107627 59261
rect 140078 59258 140084 59260
rect 107561 59256 140084 59258
rect 107561 59200 107566 59256
rect 107622 59200 140084 59256
rect 107561 59198 140084 59200
rect 107561 59195 107627 59198
rect 140078 59196 140084 59198
rect 140148 59196 140154 59260
rect 160686 59196 160692 59260
rect 160756 59258 160762 59260
rect 194685 59258 194751 59261
rect 195053 59258 195119 59261
rect 160756 59256 195119 59258
rect 160756 59200 194690 59256
rect 194746 59200 195058 59256
rect 195114 59200 195119 59256
rect 160756 59198 195119 59200
rect 160756 59196 160762 59198
rect 194685 59195 194751 59198
rect 195053 59195 195119 59198
rect 158294 59060 158300 59124
rect 158364 59122 158370 59124
rect 192109 59122 192175 59125
rect 193121 59122 193187 59125
rect 158364 59120 193187 59122
rect 158364 59064 192114 59120
rect 192170 59064 193126 59120
rect 193182 59064 193187 59120
rect 158364 59062 193187 59064
rect 158364 59060 158370 59062
rect 192109 59059 192175 59062
rect 193121 59059 193187 59062
rect 174854 58924 174860 58988
rect 174924 58986 174930 58988
rect 201677 58986 201743 58989
rect 202781 58986 202847 58989
rect 174924 58984 202847 58986
rect 174924 58928 201682 58984
rect 201738 58928 202786 58984
rect 202842 58928 202847 58984
rect 174924 58926 202847 58928
rect 174924 58924 174930 58926
rect 201677 58923 201743 58926
rect 202781 58923 202847 58926
rect 193121 58850 193187 58853
rect 327073 58850 327139 58853
rect 193121 58848 327139 58850
rect 193121 58792 193126 58848
rect 193182 58792 327078 58848
rect 327134 58792 327139 58848
rect 193121 58790 327139 58792
rect 193121 58787 193187 58790
rect 327073 58787 327139 58790
rect 195053 58714 195119 58717
rect 362953 58714 363019 58717
rect 195053 58712 363019 58714
rect -960 58578 480 58668
rect 195053 58656 195058 58712
rect 195114 58656 362958 58712
rect 363014 58656 363019 58712
rect 195053 58654 363019 58656
rect 195053 58651 195119 58654
rect 362953 58651 363019 58654
rect 3509 58578 3575 58581
rect -960 58576 3575 58578
rect -960 58520 3514 58576
rect 3570 58520 3575 58576
rect -960 58518 3575 58520
rect -960 58428 480 58518
rect 3509 58515 3575 58518
rect 97993 58578 98059 58581
rect 107561 58578 107627 58581
rect 97993 58576 107627 58578
rect 97993 58520 97998 58576
rect 98054 58520 107566 58576
rect 107622 58520 107627 58576
rect 97993 58518 107627 58520
rect 97993 58515 98059 58518
rect 107561 58515 107627 58518
rect 202781 58578 202847 58581
rect 539685 58578 539751 58581
rect 202781 58576 539751 58578
rect 202781 58520 202786 58576
rect 202842 58520 539690 58576
rect 539746 58520 539751 58576
rect 202781 58518 539751 58520
rect 202781 58515 202847 58518
rect 539685 58515 539751 58518
rect 105813 57898 105879 57901
rect 106181 57898 106247 57901
rect 138054 57898 138060 57900
rect 105813 57896 138060 57898
rect 105813 57840 105818 57896
rect 105874 57840 106186 57896
rect 106242 57840 138060 57896
rect 105813 57838 138060 57840
rect 105813 57835 105879 57838
rect 106181 57835 106247 57838
rect 138054 57836 138060 57838
rect 138124 57836 138130 57900
rect 157006 57836 157012 57900
rect 157076 57898 157082 57900
rect 190545 57898 190611 57901
rect 191741 57898 191807 57901
rect 157076 57896 191807 57898
rect 157076 57840 190550 57896
rect 190606 57840 191746 57896
rect 191802 57840 191807 57896
rect 157076 57838 191807 57840
rect 157076 57836 157082 57838
rect 190545 57835 190611 57838
rect 191741 57835 191807 57838
rect 165286 57700 165292 57764
rect 165356 57762 165362 57764
rect 194777 57762 194843 57765
rect 195053 57762 195119 57765
rect 165356 57760 195119 57762
rect 165356 57704 194782 57760
rect 194838 57704 195058 57760
rect 195114 57704 195119 57760
rect 165356 57702 195119 57704
rect 165356 57700 165362 57702
rect 194777 57699 194843 57702
rect 195053 57699 195119 57702
rect 175038 57564 175044 57628
rect 175108 57626 175114 57628
rect 201534 57626 201540 57628
rect 175108 57566 201540 57626
rect 175108 57564 175114 57566
rect 201534 57564 201540 57566
rect 201604 57626 201610 57628
rect 202822 57626 202828 57628
rect 201604 57566 202828 57626
rect 201604 57564 201610 57566
rect 202822 57564 202828 57566
rect 202892 57564 202898 57628
rect 191741 57490 191807 57493
rect 313273 57490 313339 57493
rect 191741 57488 313339 57490
rect 191741 57432 191746 57488
rect 191802 57432 313278 57488
rect 313334 57432 313339 57488
rect 191741 57430 313339 57432
rect 191741 57427 191807 57430
rect 313273 57427 313339 57430
rect 195053 57354 195119 57357
rect 418797 57354 418863 57357
rect 195053 57352 418863 57354
rect 195053 57296 195058 57352
rect 195114 57296 418802 57352
rect 418858 57296 418863 57352
rect 195053 57294 418863 57296
rect 195053 57291 195119 57294
rect 418797 57291 418863 57294
rect 77293 57218 77359 57221
rect 105813 57218 105879 57221
rect 77293 57216 105879 57218
rect 77293 57160 77298 57216
rect 77354 57160 105818 57216
rect 105874 57160 105879 57216
rect 77293 57158 105879 57160
rect 77293 57155 77359 57158
rect 105813 57155 105879 57158
rect 202822 57156 202828 57220
rect 202892 57218 202898 57220
rect 545757 57218 545823 57221
rect 202892 57216 545823 57218
rect 202892 57160 545762 57216
rect 545818 57160 545823 57216
rect 202892 57158 545823 57160
rect 202892 57156 202898 57158
rect 545757 57155 545823 57158
rect 163262 56476 163268 56540
rect 163332 56538 163338 56540
rect 197445 56538 197511 56541
rect 163332 56536 197511 56538
rect 163332 56480 197450 56536
rect 197506 56480 197511 56536
rect 163332 56478 197511 56480
rect 163332 56476 163338 56478
rect 197445 56475 197511 56478
rect 149830 56340 149836 56404
rect 149900 56402 149906 56404
rect 231853 56402 231919 56405
rect 149900 56400 231919 56402
rect 149900 56344 231858 56400
rect 231914 56344 231919 56400
rect 149900 56342 231919 56344
rect 149900 56340 149906 56342
rect 231853 56339 231919 56342
rect 157190 56204 157196 56268
rect 157260 56266 157266 56268
rect 189257 56266 189323 56269
rect 315297 56266 315363 56269
rect 157260 56264 315363 56266
rect 157260 56208 189262 56264
rect 189318 56208 315302 56264
rect 315358 56208 315363 56264
rect 157260 56206 315363 56208
rect 157260 56204 157266 56206
rect 189257 56203 189323 56206
rect 315297 56203 315363 56206
rect 197445 56130 197511 56133
rect 400949 56130 401015 56133
rect 197445 56128 401015 56130
rect 197445 56072 197450 56128
rect 197506 56072 400954 56128
rect 401010 56072 401015 56128
rect 197445 56070 401015 56072
rect 197445 56067 197511 56070
rect 400949 56067 401015 56070
rect 167678 55932 167684 55996
rect 167748 55994 167754 55996
rect 201769 55994 201835 55997
rect 450537 55994 450603 55997
rect 167748 55992 450603 55994
rect 167748 55936 201774 55992
rect 201830 55936 450542 55992
rect 450598 55936 450603 55992
rect 167748 55934 450603 55936
rect 167748 55932 167754 55934
rect 201769 55931 201835 55934
rect 450537 55931 450603 55934
rect 170438 55796 170444 55860
rect 170508 55858 170514 55860
rect 198825 55858 198891 55861
rect 489913 55858 489979 55861
rect 170508 55856 489979 55858
rect 170508 55800 198830 55856
rect 198886 55800 489918 55856
rect 489974 55800 489979 55856
rect 170508 55798 489979 55800
rect 170508 55796 170514 55798
rect 198825 55795 198891 55798
rect 489913 55795 489979 55798
rect 103973 55178 104039 55181
rect 136582 55178 136588 55180
rect 103973 55176 136588 55178
rect 103973 55120 103978 55176
rect 104034 55120 136588 55176
rect 103973 55118 136588 55120
rect 103973 55115 104039 55118
rect 136582 55116 136588 55118
rect 136652 55116 136658 55180
rect 160870 55116 160876 55180
rect 160940 55178 160946 55180
rect 194593 55178 194659 55181
rect 160940 55176 194659 55178
rect 160940 55120 194598 55176
rect 194654 55120 194659 55176
rect 160940 55118 194659 55120
rect 160940 55116 160946 55118
rect 194593 55115 194659 55118
rect 113817 55044 113883 55045
rect 113766 55042 113772 55044
rect 113726 54982 113772 55042
rect 113836 55040 113883 55044
rect 113878 54984 113883 55040
rect 113766 54980 113772 54982
rect 113836 54980 113883 54984
rect 158478 54980 158484 55044
rect 158548 55042 158554 55044
rect 191833 55042 191899 55045
rect 158548 55040 191899 55042
rect 158548 54984 191838 55040
rect 191894 54984 191899 55040
rect 158548 54982 191899 54984
rect 158548 54980 158554 54982
rect 113817 54979 113883 54980
rect 191833 54979 191899 54982
rect 148174 54844 148180 54908
rect 148244 54906 148250 54908
rect 209865 54906 209931 54909
rect 148244 54904 209931 54906
rect 148244 54848 209870 54904
rect 209926 54848 209931 54904
rect 148244 54846 209931 54848
rect 148244 54844 148250 54846
rect 209865 54843 209931 54846
rect 191833 54770 191899 54773
rect 333973 54770 334039 54773
rect 191833 54768 334039 54770
rect 191833 54712 191838 54768
rect 191894 54712 333978 54768
rect 334034 54712 334039 54768
rect 191833 54710 334039 54712
rect 191833 54707 191899 54710
rect 333973 54707 334039 54710
rect 194593 54634 194659 54637
rect 364977 54634 365043 54637
rect 194593 54632 365043 54634
rect 194593 54576 194598 54632
rect 194654 54576 364982 54632
rect 365038 54576 365043 54632
rect 194593 54574 365043 54576
rect 194593 54571 194659 54574
rect 364977 54571 365043 54574
rect 56593 54498 56659 54501
rect 103973 54498 104039 54501
rect 56593 54496 104039 54498
rect 56593 54440 56598 54496
rect 56654 54440 103978 54496
rect 104034 54440 104039 54496
rect 56593 54438 104039 54440
rect 56593 54435 56659 54438
rect 103973 54435 104039 54438
rect 104893 54498 104959 54501
rect 113817 54498 113883 54501
rect 104893 54496 113883 54498
rect 104893 54440 104898 54496
rect 104954 54440 113822 54496
rect 113878 54440 113883 54496
rect 104893 54438 113883 54440
rect 104893 54435 104959 54438
rect 113817 54435 113883 54438
rect 165470 54436 165476 54500
rect 165540 54498 165546 54500
rect 196198 54498 196204 54500
rect 165540 54438 196204 54498
rect 165540 54436 165546 54438
rect 196198 54436 196204 54438
rect 196268 54498 196274 54500
rect 423765 54498 423831 54501
rect 196268 54496 423831 54498
rect 196268 54440 423770 54496
rect 423826 54440 423831 54496
rect 196268 54438 423831 54440
rect 196268 54436 196274 54438
rect 423765 54435 423831 54438
rect 166574 53756 166580 53820
rect 166644 53818 166650 53820
rect 200205 53818 200271 53821
rect 201401 53818 201467 53821
rect 166644 53816 201467 53818
rect 166644 53760 200210 53816
rect 200266 53760 201406 53816
rect 201462 53760 201467 53816
rect 166644 53758 201467 53760
rect 166644 53756 166650 53758
rect 200205 53755 200271 53758
rect 201401 53755 201467 53758
rect 162526 53620 162532 53684
rect 162596 53682 162602 53684
rect 195973 53682 196039 53685
rect 162596 53680 196039 53682
rect 162596 53624 195978 53680
rect 196034 53624 196039 53680
rect 162596 53622 196039 53624
rect 162596 53620 162602 53622
rect 195973 53619 196039 53622
rect 154246 53484 154252 53548
rect 154316 53546 154322 53548
rect 182766 53546 182772 53548
rect 154316 53486 182772 53546
rect 154316 53484 154322 53486
rect 182766 53484 182772 53486
rect 182836 53546 182842 53548
rect 278773 53546 278839 53549
rect 182836 53544 278839 53546
rect 182836 53488 278778 53544
rect 278834 53488 278839 53544
rect 182836 53486 278839 53488
rect 182836 53484 182842 53486
rect 278773 53483 278839 53486
rect 158846 53348 158852 53412
rect 158916 53410 158922 53412
rect 192845 53410 192911 53413
rect 351913 53410 351979 53413
rect 158916 53408 351979 53410
rect 158916 53352 192850 53408
rect 192906 53352 351918 53408
rect 351974 53352 351979 53408
rect 158916 53350 351979 53352
rect 158916 53348 158922 53350
rect 192845 53347 192911 53350
rect 351913 53347 351979 53350
rect 195973 53274 196039 53277
rect 387793 53274 387859 53277
rect 195973 53272 387859 53274
rect 195973 53216 195978 53272
rect 196034 53216 387798 53272
rect 387854 53216 387859 53272
rect 195973 53214 387859 53216
rect 195973 53211 196039 53214
rect 387793 53211 387859 53214
rect 201401 53138 201467 53141
rect 432597 53138 432663 53141
rect 201401 53136 432663 53138
rect 201401 53080 201406 53136
rect 201462 53080 432602 53136
rect 432658 53080 432663 53136
rect 201401 53078 432663 53080
rect 201401 53075 201467 53078
rect 432597 53075 432663 53078
rect 100753 52458 100819 52461
rect 101765 52458 101831 52461
rect 134190 52458 134196 52460
rect 100753 52456 134196 52458
rect 100753 52400 100758 52456
rect 100814 52400 101770 52456
rect 101826 52400 134196 52456
rect 100753 52398 134196 52400
rect 100753 52395 100819 52398
rect 101765 52395 101831 52398
rect 134190 52396 134196 52398
rect 134260 52396 134266 52460
rect 170622 52396 170628 52460
rect 170692 52458 170698 52460
rect 204621 52458 204687 52461
rect 170692 52456 204687 52458
rect 170692 52400 204626 52456
rect 204682 52400 204687 52456
rect 170692 52398 204687 52400
rect 170692 52396 170698 52398
rect 204621 52395 204687 52398
rect 169334 52260 169340 52324
rect 169404 52322 169410 52324
rect 203006 52322 203012 52324
rect 169404 52262 203012 52322
rect 169404 52260 169410 52262
rect 203006 52260 203012 52262
rect 203076 52322 203082 52324
rect 204110 52322 204116 52324
rect 203076 52262 204116 52322
rect 203076 52260 203082 52262
rect 204110 52260 204116 52262
rect 204180 52260 204186 52324
rect 161238 52124 161244 52188
rect 161308 52186 161314 52188
rect 191557 52186 191623 52189
rect 369853 52186 369919 52189
rect 161308 52184 369919 52186
rect 161308 52128 191562 52184
rect 191618 52128 369858 52184
rect 369914 52128 369919 52184
rect 161308 52126 369919 52128
rect 161308 52124 161314 52126
rect 191557 52123 191623 52126
rect 369853 52123 369919 52126
rect 161054 51988 161060 52052
rect 161124 52050 161130 52052
rect 194225 52050 194291 52053
rect 373993 52050 374059 52053
rect 161124 52048 374059 52050
rect 161124 51992 194230 52048
rect 194286 51992 373998 52048
rect 374054 51992 374059 52048
rect 161124 51990 374059 51992
rect 161124 51988 161130 51990
rect 194225 51987 194291 51990
rect 373993 51987 374059 51990
rect 204110 51852 204116 51916
rect 204180 51914 204186 51916
rect 476113 51914 476179 51917
rect 204180 51912 476179 51914
rect 204180 51856 476118 51912
rect 476174 51856 476179 51912
rect 204180 51854 476179 51856
rect 204180 51852 204186 51854
rect 476113 51851 476179 51854
rect 27705 51778 27771 51781
rect 100753 51778 100819 51781
rect 27705 51776 100819 51778
rect 27705 51720 27710 51776
rect 27766 51720 100758 51776
rect 100814 51720 100819 51776
rect 27705 51718 100819 51720
rect 27705 51715 27771 51718
rect 100753 51715 100819 51718
rect 204621 51778 204687 51781
rect 484393 51778 484459 51781
rect 204621 51776 484459 51778
rect 204621 51720 204626 51776
rect 204682 51720 484398 51776
rect 484454 51720 484459 51776
rect 204621 51718 484459 51720
rect 204621 51715 204687 51718
rect 484393 51715 484459 51718
rect 159030 50900 159036 50964
rect 159100 50962 159106 50964
rect 193305 50962 193371 50965
rect 159100 50960 209790 50962
rect 159100 50904 193310 50960
rect 193366 50904 209790 50960
rect 159100 50902 209790 50904
rect 159100 50900 159106 50902
rect 193305 50899 193371 50902
rect 166758 50764 166764 50828
rect 166828 50826 166834 50828
rect 200113 50826 200179 50829
rect 201401 50826 201467 50829
rect 166828 50824 201467 50826
rect 166828 50768 200118 50824
rect 200174 50768 201406 50824
rect 201462 50768 201467 50824
rect 166828 50766 201467 50768
rect 166828 50764 166834 50766
rect 200113 50763 200179 50766
rect 201401 50763 201467 50766
rect 163446 50628 163452 50692
rect 163516 50690 163522 50692
rect 209730 50690 209790 50902
rect 356053 50690 356119 50693
rect 163516 50630 180810 50690
rect 209730 50688 356119 50690
rect 209730 50632 356058 50688
rect 356114 50632 356119 50688
rect 209730 50630 356119 50632
rect 163516 50628 163522 50630
rect 180750 50554 180810 50630
rect 356053 50627 356119 50630
rect 192201 50554 192267 50557
rect 405733 50554 405799 50557
rect 180750 50552 405799 50554
rect 180750 50496 192206 50552
rect 192262 50496 405738 50552
rect 405794 50496 405799 50552
rect 180750 50494 405799 50496
rect 192201 50491 192267 50494
rect 405733 50491 405799 50494
rect 201401 50418 201467 50421
rect 440233 50418 440299 50421
rect 201401 50416 440299 50418
rect 201401 50360 201406 50416
rect 201462 50360 440238 50416
rect 440294 50360 440299 50416
rect 201401 50358 440299 50360
rect 201401 50355 201467 50358
rect 440233 50355 440299 50358
rect 177062 50220 177068 50284
rect 177132 50282 177138 50284
rect 205817 50282 205883 50285
rect 569953 50282 570019 50285
rect 177132 50280 570019 50282
rect 177132 50224 205822 50280
rect 205878 50224 569958 50280
rect 570014 50224 570019 50280
rect 177132 50222 570019 50224
rect 177132 50220 177138 50222
rect 205817 50219 205883 50222
rect 569953 50219 570019 50222
rect 100753 49602 100819 49605
rect 102041 49602 102107 49605
rect 135662 49602 135668 49604
rect 100753 49600 135668 49602
rect 100753 49544 100758 49600
rect 100814 49544 102046 49600
rect 102102 49544 135668 49600
rect 100753 49542 135668 49544
rect 100753 49539 100819 49542
rect 102041 49539 102107 49542
rect 135662 49540 135668 49542
rect 135732 49540 135738 49604
rect 167862 49540 167868 49604
rect 167932 49602 167938 49604
rect 202505 49602 202571 49605
rect 167932 49600 209790 49602
rect 167932 49544 202510 49600
rect 202566 49544 209790 49600
rect 167932 49542 209790 49544
rect 167932 49540 167938 49542
rect 202505 49539 202571 49542
rect 170806 49404 170812 49468
rect 170876 49466 170882 49468
rect 198774 49466 198780 49468
rect 170876 49406 198780 49466
rect 170876 49404 170882 49406
rect 198774 49404 198780 49406
rect 198844 49404 198850 49468
rect 175958 49268 175964 49332
rect 176028 49330 176034 49332
rect 204437 49330 204503 49333
rect 204713 49330 204779 49333
rect 176028 49328 204779 49330
rect 176028 49272 204442 49328
rect 204498 49272 204718 49328
rect 204774 49272 204779 49328
rect 176028 49270 204779 49272
rect 176028 49268 176034 49270
rect 204437 49267 204503 49270
rect 204713 49267 204779 49270
rect 209730 49194 209790 49542
rect 454677 49194 454743 49197
rect 209730 49192 454743 49194
rect 209730 49136 454682 49192
rect 454738 49136 454743 49192
rect 209730 49134 454743 49136
rect 454677 49131 454743 49134
rect 198774 48996 198780 49060
rect 198844 49058 198850 49060
rect 494053 49058 494119 49061
rect 198844 49056 494119 49058
rect 198844 49000 494058 49056
rect 494114 49000 494119 49056
rect 198844 48998 494119 49000
rect 198844 48996 198850 48998
rect 494053 48995 494119 48998
rect 39297 48922 39363 48925
rect 100753 48922 100819 48925
rect 39297 48920 100819 48922
rect 39297 48864 39302 48920
rect 39358 48864 100758 48920
rect 100814 48864 100819 48920
rect 39297 48862 100819 48864
rect 39297 48859 39363 48862
rect 100753 48859 100819 48862
rect 204713 48922 204779 48925
rect 565813 48922 565879 48925
rect 204713 48920 565879 48922
rect 204713 48864 204718 48920
rect 204774 48864 565818 48920
rect 565874 48864 565879 48920
rect 204713 48862 565879 48864
rect 204713 48859 204779 48862
rect 565813 48859 565879 48862
rect 100753 48242 100819 48245
rect 101949 48242 102015 48245
rect 135478 48242 135484 48244
rect 100753 48240 135484 48242
rect 100753 48184 100758 48240
rect 100814 48184 101954 48240
rect 102010 48184 135484 48240
rect 100753 48182 135484 48184
rect 100753 48179 100819 48182
rect 101949 48179 102015 48182
rect 135478 48180 135484 48182
rect 135548 48180 135554 48244
rect 162710 48180 162716 48244
rect 162780 48242 162786 48244
rect 196014 48242 196020 48244
rect 162780 48182 196020 48242
rect 162780 48180 162786 48182
rect 196014 48180 196020 48182
rect 196084 48180 196090 48244
rect 173750 48044 173756 48108
rect 173820 48106 173826 48108
rect 204529 48106 204595 48109
rect 204805 48106 204871 48109
rect 173820 48104 204871 48106
rect 173820 48048 204534 48104
rect 204590 48048 204810 48104
rect 204866 48048 204871 48104
rect 173820 48046 204871 48048
rect 173820 48044 173826 48046
rect 204529 48043 204595 48046
rect 204805 48043 204871 48046
rect 196014 47636 196020 47700
rect 196084 47698 196090 47700
rect 390553 47698 390619 47701
rect 196084 47696 390619 47698
rect 196084 47640 390558 47696
rect 390614 47640 390619 47696
rect 196084 47638 390619 47640
rect 196084 47636 196090 47638
rect 390553 47635 390619 47638
rect 44173 47562 44239 47565
rect 100753 47562 100819 47565
rect 44173 47560 100819 47562
rect 44173 47504 44178 47560
rect 44234 47504 100758 47560
rect 100814 47504 100819 47560
rect 44173 47502 100819 47504
rect 44173 47499 44239 47502
rect 100753 47499 100819 47502
rect 147438 47500 147444 47564
rect 147508 47562 147514 47564
rect 194593 47562 194659 47565
rect 147508 47560 194659 47562
rect 147508 47504 194598 47560
rect 194654 47504 194659 47560
rect 147508 47502 194659 47504
rect 147508 47500 147514 47502
rect 194593 47499 194659 47502
rect 204805 47562 204871 47565
rect 520917 47562 520983 47565
rect 204805 47560 520983 47562
rect 204805 47504 204810 47560
rect 204866 47504 520922 47560
rect 520978 47504 520983 47560
rect 204805 47502 520983 47504
rect 204805 47499 204871 47502
rect 520917 47499 520983 47502
rect 102225 46882 102291 46885
rect 102685 46882 102751 46885
rect 135294 46882 135300 46884
rect 102225 46880 135300 46882
rect 102225 46824 102230 46880
rect 102286 46824 102690 46880
rect 102746 46824 135300 46880
rect 102225 46822 135300 46824
rect 102225 46819 102291 46822
rect 102685 46819 102751 46822
rect 135294 46820 135300 46822
rect 135364 46820 135370 46884
rect 169518 46820 169524 46884
rect 169588 46882 169594 46884
rect 203241 46882 203307 46885
rect 169588 46880 209790 46882
rect 169588 46824 203246 46880
rect 203302 46824 209790 46880
rect 169588 46822 209790 46824
rect 169588 46820 169594 46822
rect 203241 46819 203307 46822
rect 170990 46684 170996 46748
rect 171060 46746 171066 46748
rect 197077 46746 197143 46749
rect 171060 46744 200130 46746
rect 171060 46688 197082 46744
rect 197138 46688 200130 46744
rect 171060 46686 200130 46688
rect 171060 46684 171066 46686
rect 197077 46683 197143 46686
rect 49693 46202 49759 46205
rect 102225 46202 102291 46205
rect 49693 46200 102291 46202
rect 49693 46144 49698 46200
rect 49754 46144 102230 46200
rect 102286 46144 102291 46200
rect 49693 46142 102291 46144
rect 200070 46202 200130 46686
rect 209730 46338 209790 46822
rect 463693 46338 463759 46341
rect 583520 46338 584960 46428
rect 209730 46336 463759 46338
rect 209730 46280 463698 46336
rect 463754 46280 463759 46336
rect 209730 46278 463759 46280
rect 463693 46275 463759 46278
rect 583342 46278 584960 46338
rect 495433 46202 495499 46205
rect 200070 46200 495499 46202
rect 200070 46144 495438 46200
rect 495494 46144 495499 46200
rect 200070 46142 495499 46144
rect 583342 46202 583402 46278
rect 583520 46202 584960 46278
rect 583342 46188 584960 46202
rect 583342 46142 583586 46188
rect 49693 46139 49759 46142
rect 102225 46139 102291 46142
rect 495433 46139 495499 46142
rect -960 45522 480 45612
rect 192334 45596 192340 45660
rect 192404 45658 192410 45660
rect 583526 45658 583586 46142
rect 192404 45598 583586 45658
rect 192404 45596 192410 45598
rect -960 45462 674 45522
rect -960 45386 480 45462
rect 614 45386 674 45462
rect 163630 45460 163636 45524
rect 163700 45522 163706 45524
rect 197353 45522 197419 45525
rect 163700 45520 197419 45522
rect 163700 45464 197358 45520
rect 197414 45464 197419 45520
rect 163700 45462 197419 45464
rect 163700 45460 163706 45462
rect 197353 45459 197419 45462
rect -960 45372 674 45386
rect 246 45326 674 45372
rect 246 44842 306 45326
rect 148910 45052 148916 45116
rect 148980 45114 148986 45116
rect 212533 45114 212599 45117
rect 148980 45112 212599 45114
rect 148980 45056 212538 45112
rect 212594 45056 212599 45112
rect 148980 45054 212599 45056
rect 148980 45052 148986 45054
rect 212533 45051 212599 45054
rect 152590 44916 152596 44980
rect 152660 44978 152666 44980
rect 267733 44978 267799 44981
rect 152660 44976 267799 44978
rect 152660 44920 267738 44976
rect 267794 44920 267799 44976
rect 152660 44918 267799 44920
rect 152660 44916 152666 44918
rect 267733 44915 267799 44918
rect 197353 44842 197419 44845
rect 408493 44842 408559 44845
rect 246 44782 6930 44842
rect 6870 44298 6930 44782
rect 197353 44840 408559 44842
rect 197353 44784 197358 44840
rect 197414 44784 408498 44840
rect 408554 44784 408559 44840
rect 197353 44782 408559 44784
rect 197353 44779 197419 44782
rect 408493 44779 408559 44782
rect 116526 44298 116532 44300
rect 6870 44238 116532 44298
rect 116526 44236 116532 44238
rect 116596 44236 116602 44300
rect 168046 44100 168052 44164
rect 168116 44162 168122 44164
rect 201769 44162 201835 44165
rect 202781 44162 202847 44165
rect 168116 44160 202847 44162
rect 168116 44104 201774 44160
rect 201830 44104 202786 44160
rect 202842 44104 202847 44160
rect 168116 44102 202847 44104
rect 168116 44100 168122 44102
rect 201769 44099 201835 44102
rect 202781 44099 202847 44102
rect 154430 43964 154436 44028
rect 154500 44026 154506 44028
rect 186998 44026 187004 44028
rect 154500 43966 187004 44026
rect 154500 43964 154506 43966
rect 186998 43964 187004 43966
rect 187068 43964 187074 44028
rect 186998 43556 187004 43620
rect 187068 43618 187074 43620
rect 284385 43618 284451 43621
rect 187068 43616 284451 43618
rect 187068 43560 284390 43616
rect 284446 43560 284451 43616
rect 187068 43558 284451 43560
rect 187068 43556 187074 43558
rect 284385 43555 284451 43558
rect 202781 43482 202847 43485
rect 452653 43482 452719 43485
rect 202781 43480 452719 43482
rect 202781 43424 202786 43480
rect 202842 43424 452658 43480
rect 452714 43424 452719 43480
rect 202781 43422 452719 43424
rect 202781 43419 202847 43422
rect 452653 43419 452719 43422
rect 172278 42740 172284 42804
rect 172348 42802 172354 42804
rect 205633 42802 205699 42805
rect 172348 42800 205699 42802
rect 172348 42744 205638 42800
rect 205694 42744 205699 42800
rect 172348 42742 205699 42744
rect 172348 42740 172354 42742
rect 205633 42739 205699 42742
rect 205633 42122 205699 42125
rect 507853 42122 507919 42125
rect 205633 42120 507919 42122
rect 205633 42064 205638 42120
rect 205694 42064 507858 42120
rect 507914 42064 507919 42120
rect 205633 42062 507919 42064
rect 205633 42059 205699 42062
rect 507853 42059 507919 42062
rect 145598 37844 145604 37908
rect 145668 37906 145674 37908
rect 170397 37906 170463 37909
rect 145668 37904 170463 37906
rect 145668 37848 170402 37904
rect 170458 37848 170463 37904
rect 145668 37846 170463 37848
rect 145668 37844 145674 37846
rect 170397 37843 170463 37846
rect 17217 33826 17283 33829
rect 133638 33826 133644 33828
rect 17217 33824 133644 33826
rect 17217 33768 17222 33824
rect 17278 33768 133644 33824
rect 17217 33766 133644 33768
rect 17217 33763 17283 33766
rect 133638 33764 133644 33766
rect 133708 33764 133714 33828
rect 144678 33764 144684 33828
rect 144748 33826 144754 33828
rect 160369 33826 160435 33829
rect 144748 33824 160435 33826
rect 144748 33768 160374 33824
rect 160430 33768 160435 33824
rect 144748 33766 160435 33768
rect 144748 33764 144754 33766
rect 160369 33763 160435 33766
rect 583520 33146 584960 33236
rect 583342 33086 584960 33146
rect 583342 33010 583402 33086
rect 583520 33010 584960 33086
rect 583342 32996 584960 33010
rect 583342 32950 583586 32996
rect -960 32466 480 32556
rect -960 32406 674 32466
rect -960 32330 480 32406
rect 614 32330 674 32406
rect -960 32316 674 32330
rect 246 32270 674 32316
rect 246 31786 306 32270
rect 117814 31786 117820 31788
rect 246 31726 117820 31786
rect 117814 31724 117820 31726
rect 117884 31724 117890 31788
rect 189574 31724 189580 31788
rect 189644 31786 189650 31788
rect 583526 31786 583586 32950
rect 189644 31726 583586 31786
rect 189644 31724 189650 31726
rect 149646 30908 149652 30972
rect 149716 30970 149722 30972
rect 229093 30970 229159 30973
rect 149716 30968 229159 30970
rect 149716 30912 229098 30968
rect 229154 30912 229159 30968
rect 149716 30910 229159 30912
rect 149716 30908 149722 30910
rect 229093 30907 229159 30910
rect 152406 28188 152412 28252
rect 152476 28250 152482 28252
rect 264973 28250 265039 28253
rect 152476 28248 265039 28250
rect 152476 28192 264978 28248
rect 265034 28192 265039 28248
rect 152476 28190 265039 28192
rect 152476 28188 152482 28190
rect 264973 28187 265039 28190
rect 144494 26828 144500 26892
rect 144564 26890 144570 26892
rect 155953 26890 156019 26893
rect 144564 26888 156019 26890
rect 144564 26832 155958 26888
rect 156014 26832 156019 26888
rect 144564 26830 156019 26832
rect 144564 26828 144570 26830
rect 155953 26827 156019 26830
rect 579981 19818 580047 19821
rect 583520 19818 584960 19908
rect 579981 19816 584960 19818
rect 579981 19760 579986 19816
rect 580042 19760 584960 19816
rect 579981 19758 584960 19760
rect 579981 19755 580047 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 108246 19410 108252 19412
rect -960 19350 108252 19410
rect -960 19260 480 19350
rect 108246 19348 108252 19350
rect 108316 19348 108322 19412
rect 145414 17172 145420 17236
rect 145484 17234 145490 17236
rect 171869 17234 171935 17237
rect 145484 17232 171935 17234
rect 145484 17176 171874 17232
rect 171930 17176 171935 17232
rect 145484 17174 171935 17176
rect 145484 17172 145490 17174
rect 171869 17171 171935 17174
rect 144126 15812 144132 15876
rect 144196 15874 144202 15876
rect 161289 15874 161355 15877
rect 144196 15872 161355 15874
rect 144196 15816 161294 15872
rect 161350 15816 161355 15872
rect 144196 15814 161355 15816
rect 144196 15812 144202 15814
rect 161289 15811 161355 15814
rect 144310 11596 144316 11660
rect 144380 11658 144386 11660
rect 158897 11658 158963 11661
rect 144380 11656 158963 11658
rect 144380 11600 158902 11656
rect 158958 11600 158963 11656
rect 144380 11598 158963 11600
rect 144380 11596 144386 11598
rect 158897 11595 158963 11598
rect 580165 6626 580231 6629
rect 583520 6626 584960 6716
rect 580165 6624 584960 6626
rect -960 6490 480 6580
rect 580165 6568 580170 6624
rect 580226 6568 584960 6624
rect 580165 6566 584960 6568
rect 580165 6563 580231 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect 583520 6476 584960 6566
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
<< via3 >>
rect 189028 275980 189092 276044
rect 187004 271084 187068 271148
rect 187004 270540 187068 270604
rect 193260 265236 193324 265300
rect 194548 265100 194612 265164
rect 113036 264964 113100 265028
rect 194732 264964 194796 265028
rect 121132 263740 121196 263804
rect 118556 263604 118620 263668
rect 191972 263060 192036 263124
rect 115796 262788 115860 262852
rect 112852 262652 112916 262716
rect 193444 262652 193508 262716
rect 111564 262516 111628 262580
rect 191788 262516 191852 262580
rect 114140 262380 114204 262444
rect 190500 262380 190564 262444
rect 111380 262244 111444 262308
rect 188108 262244 188172 262308
rect 111196 260884 111260 260948
rect 120948 260476 121012 260540
rect 113588 260340 113652 260404
rect 118372 260204 118436 260268
rect 115612 260068 115676 260132
rect 116900 259932 116964 259996
rect 117084 259796 117148 259860
rect 113956 259660 114020 259724
rect 118188 259584 118252 259588
rect 118188 259528 118238 259584
rect 118238 259528 118252 259584
rect 118188 259524 118252 259528
rect 185348 259584 185412 259588
rect 185348 259528 185398 259584
rect 185398 259528 185412 259584
rect 185348 259524 185412 259528
rect 186084 259584 186148 259588
rect 186084 259528 186098 259584
rect 186098 259528 186148 259584
rect 186084 259524 186148 259528
rect 186452 210292 186516 210356
rect 186084 202812 186148 202876
rect 185348 201724 185412 201788
rect 157196 200636 157260 200700
rect 179828 200636 179892 200700
rect 166212 200500 166276 200564
rect 182956 200500 183020 200564
rect 137876 200228 137940 200292
rect 166580 200364 166644 200428
rect 136404 200092 136468 200156
rect 137508 200092 137572 200156
rect 139532 200092 139596 200156
rect 140820 200092 140884 200156
rect 145420 200092 145484 200156
rect 163452 200092 163516 200156
rect 169156 200092 169220 200156
rect 132724 199858 132728 199884
rect 132728 199858 132784 199884
rect 132784 199858 132788 199884
rect 132724 199820 132788 199858
rect 133092 199820 133156 199884
rect 133460 199858 133464 199884
rect 133464 199858 133520 199884
rect 133520 199858 133524 199884
rect 133460 199820 133524 199858
rect 134196 199820 134260 199884
rect 134380 199880 134444 199884
rect 134380 199824 134384 199880
rect 134384 199824 134440 199880
rect 134440 199824 134444 199880
rect 134380 199820 134444 199824
rect 134748 199858 134752 199884
rect 134752 199858 134808 199884
rect 134808 199858 134812 199884
rect 134748 199820 134812 199858
rect 135116 199858 135120 199884
rect 135120 199858 135176 199884
rect 135176 199858 135180 199884
rect 135116 199820 135180 199858
rect 135484 199820 135548 199884
rect 135852 199858 135856 199884
rect 135856 199858 135912 199884
rect 135912 199858 135916 199884
rect 135852 199820 135916 199858
rect 136956 199820 137020 199884
rect 137140 199858 137144 199884
rect 137144 199858 137200 199884
rect 137200 199858 137204 199884
rect 137140 199820 137204 199858
rect 137692 199820 137756 199884
rect 138060 199858 138064 199884
rect 138064 199858 138120 199884
rect 138120 199858 138124 199884
rect 138060 199820 138124 199858
rect 138612 199820 138676 199884
rect 138796 199820 138860 199884
rect 139348 199858 139352 199884
rect 139352 199858 139408 199884
rect 139408 199858 139412 199884
rect 139348 199820 139412 199858
rect 139716 199858 139720 199884
rect 139720 199858 139776 199884
rect 139776 199858 139780 199884
rect 139716 199820 139780 199858
rect 140084 199820 140148 199884
rect 140452 199858 140456 199884
rect 140456 199858 140512 199884
rect 140512 199858 140516 199884
rect 140452 199820 140516 199858
rect 141004 199820 141068 199884
rect 141188 199820 141252 199884
rect 142476 199858 142480 199884
rect 142480 199858 142536 199884
rect 142536 199858 142540 199884
rect 142476 199820 142540 199858
rect 143028 199858 143032 199884
rect 143032 199858 143088 199884
rect 143088 199858 143092 199884
rect 143028 199820 143092 199858
rect 133092 199548 133156 199612
rect 136404 199608 136468 199612
rect 136404 199552 136454 199608
rect 136454 199552 136468 199608
rect 136404 199548 136468 199552
rect 137876 199548 137940 199612
rect 142660 199684 142724 199748
rect 144684 199858 144688 199884
rect 144688 199858 144744 199884
rect 144744 199858 144748 199884
rect 144684 199820 144748 199858
rect 145052 199820 145116 199884
rect 146524 199820 146588 199884
rect 146708 199858 146712 199884
rect 146712 199858 146768 199884
rect 146768 199858 146772 199884
rect 146708 199820 146772 199858
rect 147076 199858 147080 199884
rect 147080 199858 147136 199884
rect 147136 199858 147140 199884
rect 147076 199820 147140 199858
rect 148180 199858 148184 199884
rect 148184 199858 148240 199884
rect 148240 199858 148244 199884
rect 148180 199820 148244 199858
rect 149284 199858 149288 199884
rect 149288 199858 149344 199884
rect 149344 199858 149348 199884
rect 149284 199820 149348 199858
rect 149652 199820 149716 199884
rect 150940 199858 150944 199884
rect 150944 199858 151000 199884
rect 151000 199858 151004 199884
rect 150940 199820 151004 199858
rect 146892 199684 146956 199748
rect 151124 199684 151188 199748
rect 152596 199820 152660 199884
rect 153332 199820 153396 199884
rect 154068 199820 154132 199884
rect 154620 199820 154684 199884
rect 155908 199820 155972 199884
rect 156644 199820 156708 199884
rect 157748 199820 157812 199884
rect 156460 199684 156524 199748
rect 157196 199744 157260 199748
rect 157196 199688 157210 199744
rect 157210 199688 157260 199744
rect 157196 199684 157260 199688
rect 157932 199684 157996 199748
rect 158300 199684 158364 199748
rect 158852 199820 158916 199884
rect 160140 199858 160144 199884
rect 160144 199858 160200 199884
rect 160200 199858 160204 199884
rect 160140 199820 160204 199858
rect 161060 199820 161124 199884
rect 161612 199858 161616 199884
rect 161616 199858 161672 199884
rect 161672 199858 161676 199884
rect 161612 199820 161676 199858
rect 162348 199820 162412 199884
rect 163268 199858 163272 199884
rect 163272 199858 163328 199884
rect 163328 199858 163332 199884
rect 163268 199820 163332 199858
rect 162900 199684 162964 199748
rect 163084 199684 163148 199748
rect 164924 199820 164988 199884
rect 166948 199880 167012 199884
rect 166948 199824 166952 199880
rect 166952 199824 167008 199880
rect 167008 199824 167012 199880
rect 166948 199820 167012 199824
rect 167868 199880 167932 199884
rect 167868 199824 167872 199880
rect 167872 199824 167928 199880
rect 167928 199824 167932 199880
rect 167868 199820 167932 199824
rect 168052 199858 168056 199884
rect 168056 199858 168112 199884
rect 168112 199858 168116 199884
rect 168052 199820 168116 199858
rect 165476 199684 165540 199748
rect 166580 199684 166644 199748
rect 166764 199744 166828 199748
rect 166764 199688 166814 199744
rect 166814 199688 166828 199744
rect 166764 199684 166828 199688
rect 167500 199744 167564 199748
rect 168604 199858 168608 199884
rect 168608 199858 168664 199884
rect 168664 199858 168668 199884
rect 168604 199820 168668 199858
rect 169340 199820 169404 199884
rect 170996 199858 171000 199884
rect 171000 199858 171056 199884
rect 171056 199858 171060 199884
rect 170996 199820 171060 199858
rect 171732 199820 171796 199884
rect 167500 199688 167550 199744
rect 167550 199688 167564 199744
rect 167500 199684 167564 199688
rect 168972 199684 169036 199748
rect 170076 199744 170140 199748
rect 170076 199688 170090 199744
rect 170090 199688 170140 199744
rect 170076 199684 170140 199688
rect 172836 199820 172900 199884
rect 174492 199820 174556 199884
rect 175044 199820 175108 199884
rect 175412 199858 175416 199884
rect 175416 199858 175472 199884
rect 175472 199858 175476 199884
rect 175412 199820 175476 199858
rect 172652 199684 172716 199748
rect 173388 199684 173452 199748
rect 174124 199684 174188 199748
rect 176516 199858 176520 199884
rect 176520 199858 176576 199884
rect 176576 199858 176580 199884
rect 176516 199820 176580 199858
rect 200988 199820 201052 199884
rect 175596 199684 175660 199748
rect 175780 199684 175844 199748
rect 189212 199684 189276 199748
rect 180748 199548 180812 199612
rect 182588 199412 182652 199476
rect 134196 199276 134260 199340
rect 135484 199276 135548 199340
rect 146892 199276 146956 199340
rect 183508 199276 183572 199340
rect 135484 199140 135548 199204
rect 140084 199140 140148 199204
rect 145052 199140 145116 199204
rect 150940 199140 151004 199204
rect 166212 199004 166276 199068
rect 178172 199004 178236 199068
rect 163452 198868 163516 198932
rect 201724 198732 201788 198796
rect 140452 198460 140516 198524
rect 148180 198460 148244 198524
rect 133828 198384 133892 198388
rect 133828 198328 133878 198384
rect 133878 198328 133892 198384
rect 133828 198324 133892 198328
rect 134196 198324 134260 198388
rect 135116 198324 135180 198388
rect 136220 198324 136284 198388
rect 141188 198324 141252 198388
rect 162900 198324 162964 198388
rect 142660 198188 142724 198252
rect 162900 198248 162964 198252
rect 162900 198192 162950 198248
rect 162950 198192 162964 198248
rect 162900 198188 162964 198192
rect 167684 198248 167748 198252
rect 167684 198192 167698 198248
rect 167698 198192 167748 198248
rect 167684 198188 167748 198192
rect 196388 198188 196452 198252
rect 140452 198052 140516 198116
rect 142292 198052 142356 198116
rect 142476 198112 142540 198116
rect 142476 198056 142490 198112
rect 142490 198056 142540 198112
rect 142476 198052 142540 198056
rect 163084 198052 163148 198116
rect 163268 198112 163332 198116
rect 163268 198056 163318 198112
rect 163318 198056 163332 198112
rect 163268 198052 163332 198056
rect 164924 198052 164988 198116
rect 166948 198112 167012 198116
rect 166948 198056 166998 198112
rect 166998 198056 167012 198112
rect 166948 198052 167012 198056
rect 167868 198112 167932 198116
rect 167868 198056 167918 198112
rect 167918 198056 167932 198112
rect 167868 198052 167932 198056
rect 168052 198112 168116 198116
rect 168052 198056 168102 198112
rect 168102 198056 168116 198112
rect 168052 198052 168116 198056
rect 198780 198052 198844 198116
rect 132724 197976 132788 197980
rect 132724 197920 132774 197976
rect 132774 197920 132788 197976
rect 132724 197916 132788 197920
rect 133460 197976 133524 197980
rect 133460 197920 133510 197976
rect 133510 197920 133524 197976
rect 133460 197916 133524 197920
rect 135852 197916 135916 197980
rect 137140 197916 137204 197980
rect 132356 197840 132420 197844
rect 132356 197784 132370 197840
rect 132370 197784 132420 197840
rect 132356 197780 132420 197784
rect 134564 197840 134628 197844
rect 134564 197784 134578 197840
rect 134578 197784 134628 197840
rect 134564 197780 134628 197784
rect 134748 197840 134812 197844
rect 134748 197784 134798 197840
rect 134798 197784 134812 197840
rect 134748 197780 134812 197784
rect 135116 197780 135180 197844
rect 135852 197780 135916 197844
rect 167500 197780 167564 197844
rect 134380 197644 134444 197708
rect 134380 197508 134444 197572
rect 179460 197508 179524 197572
rect 121316 197236 121380 197300
rect 139348 196828 139412 196892
rect 183692 196828 183756 196892
rect 187740 196692 187804 196756
rect 187924 196556 187988 196620
rect 168604 196420 168668 196484
rect 169340 195876 169404 195940
rect 144684 195740 144748 195804
rect 187188 195604 187252 195668
rect 141004 195332 141068 195396
rect 135116 195060 135180 195124
rect 138796 194788 138860 194852
rect 130332 194244 130396 194308
rect 184980 193972 185044 194036
rect 203012 193836 203076 193900
rect 127572 193700 127636 193764
rect 178356 193292 178420 193356
rect 179644 193020 179708 193084
rect 124996 192884 125060 192948
rect 180932 192884 180996 192948
rect 196204 192748 196268 192812
rect 149468 192612 149532 192676
rect 175412 192612 175476 192676
rect 196020 192476 196084 192540
rect 138060 192400 138124 192404
rect 138060 192344 138074 192400
rect 138074 192344 138124 192400
rect 138060 192340 138124 192344
rect 122972 192204 123036 192268
rect 127756 192068 127820 192132
rect 124812 191796 124876 191860
rect 126836 191388 126900 191452
rect 122236 191252 122300 191316
rect 124076 191116 124140 191180
rect 149284 191176 149348 191180
rect 149284 191120 149334 191176
rect 149334 191120 149348 191176
rect 149284 191116 149348 191120
rect 131988 190844 132052 190908
rect 130884 190708 130948 190772
rect 130700 190572 130764 190636
rect 130516 190436 130580 190500
rect 178540 190436 178604 190500
rect 125180 190300 125244 190364
rect 144316 190028 144380 190092
rect 122604 189892 122668 189956
rect 139716 189756 139780 189820
rect 113772 189620 113836 189684
rect 126652 187308 126716 187372
rect 146708 187308 146772 187372
rect 127388 187172 127452 187236
rect 163636 186900 163700 186964
rect 162900 186764 162964 186828
rect 122420 186628 122484 186692
rect 148548 186628 148612 186692
rect 161612 186628 161676 186692
rect 136220 186492 136284 186556
rect 137140 186552 137204 186556
rect 137140 186496 137190 186552
rect 137190 186496 137204 186552
rect 137140 186492 137204 186496
rect 161428 186492 161492 186556
rect 201908 186492 201972 186556
rect 151308 186356 151372 186420
rect 151860 186356 151924 186420
rect 153516 186356 153580 186420
rect 162164 186356 162228 186420
rect 164004 186356 164068 186420
rect 164924 186356 164988 186420
rect 169892 186356 169956 186420
rect 170996 186356 171060 186420
rect 136036 186220 136100 186284
rect 139164 186280 139228 186284
rect 139164 186224 139214 186280
rect 139214 186224 139228 186280
rect 139164 186220 139228 186224
rect 139532 186220 139596 186284
rect 140268 186220 140332 186284
rect 146892 186220 146956 186284
rect 148180 186220 148244 186284
rect 153332 186280 153396 186284
rect 153332 186224 153346 186280
rect 153346 186224 153396 186280
rect 153332 186220 153396 186224
rect 154068 186220 154132 186284
rect 155908 186220 155972 186284
rect 158116 186220 158180 186284
rect 160140 186220 160204 186284
rect 162532 186280 162596 186284
rect 162532 186224 162546 186280
rect 162546 186224 162596 186280
rect 162532 186220 162596 186224
rect 163268 186220 163332 186284
rect 164740 186220 164804 186284
rect 170996 186220 171060 186284
rect 174308 186220 174372 186284
rect 176516 186220 176580 186284
rect 176884 186220 176948 186284
rect 133092 186084 133156 186148
rect 134564 186084 134628 186148
rect 149284 186084 149348 186148
rect 162900 186084 162964 186148
rect 173388 186084 173452 186148
rect 125364 185948 125428 186012
rect 173204 185948 173268 186012
rect 136956 185812 137020 185876
rect 142660 185812 142724 185876
rect 169156 185872 169220 185876
rect 169156 185816 169206 185872
rect 169206 185816 169220 185872
rect 169156 185812 169220 185816
rect 175964 185812 176028 185876
rect 119844 185676 119908 185740
rect 133460 185676 133524 185740
rect 134932 185676 134996 185740
rect 147076 185676 147140 185740
rect 166028 185736 166092 185740
rect 166028 185680 166042 185736
rect 166042 185680 166092 185736
rect 166028 185676 166092 185680
rect 166212 185676 166276 185740
rect 167316 185676 167380 185740
rect 169156 185676 169220 185740
rect 172284 185736 172348 185740
rect 172284 185680 172298 185736
rect 172298 185680 172348 185736
rect 172284 185676 172348 185680
rect 200620 185676 200684 185740
rect 131620 185540 131684 185604
rect 132908 185540 132972 185604
rect 134380 185540 134444 185604
rect 134564 185540 134628 185604
rect 137692 185540 137756 185604
rect 140636 185600 140700 185604
rect 140636 185544 140650 185600
rect 140650 185544 140700 185600
rect 140636 185540 140700 185544
rect 141004 185540 141068 185604
rect 143028 185600 143092 185604
rect 143028 185544 143042 185600
rect 143042 185544 143092 185600
rect 143028 185540 143092 185544
rect 149836 185600 149900 185604
rect 149836 185544 149886 185600
rect 149886 185544 149900 185600
rect 149836 185540 149900 185544
rect 151492 185600 151556 185604
rect 151492 185544 151506 185600
rect 151506 185544 151556 185600
rect 151492 185540 151556 185544
rect 152228 185600 152292 185604
rect 152228 185544 152278 185600
rect 152278 185544 152292 185600
rect 152228 185540 152292 185544
rect 152596 185600 152660 185604
rect 152596 185544 152610 185600
rect 152610 185544 152660 185600
rect 152596 185540 152660 185544
rect 153700 185540 153764 185604
rect 155540 185540 155604 185604
rect 156828 185540 156892 185604
rect 157196 185540 157260 185604
rect 160692 185540 160756 185604
rect 165844 185540 165908 185604
rect 167500 185600 167564 185604
rect 167500 185544 167550 185600
rect 167550 185544 167564 185600
rect 167500 185540 167564 185544
rect 168052 185600 168116 185604
rect 168052 185544 168066 185600
rect 168066 185544 168116 185600
rect 168052 185540 168116 185544
rect 168604 185540 168668 185604
rect 171548 185540 171612 185604
rect 172100 185600 172164 185604
rect 172100 185544 172114 185600
rect 172114 185544 172164 185600
rect 172100 185540 172164 185544
rect 173020 185540 173084 185604
rect 197860 185540 197924 185604
rect 134748 185404 134812 185468
rect 142108 185404 142172 185468
rect 145236 185404 145300 185468
rect 200804 185404 200868 185468
rect 133828 185268 133892 185332
rect 143764 185268 143828 185332
rect 166764 185268 166828 185332
rect 197676 185268 197740 185332
rect 133276 185192 133340 185196
rect 133276 185136 133290 185192
rect 133290 185136 133340 185192
rect 133276 185132 133340 185136
rect 197308 185132 197372 185196
rect 170812 184860 170876 184924
rect 148732 183364 148796 183428
rect 136220 183092 136284 183156
rect 147076 181868 147140 181932
rect 147444 181732 147508 181796
rect 175596 180780 175660 180844
rect 166580 180236 166644 180300
rect 168788 179964 168852 180028
rect 159036 179420 159100 179484
rect 140084 179284 140148 179348
rect 146524 179284 146588 179348
rect 145604 179012 145668 179076
rect 148916 178468 148980 178532
rect 165292 178468 165356 178532
rect 161060 177924 161124 177988
rect 138428 177168 138492 177172
rect 138428 177112 138442 177168
rect 138442 177112 138492 177168
rect 138428 177108 138492 177112
rect 177068 176564 177132 176628
rect 138980 174992 139044 174996
rect 138980 174936 139030 174992
rect 139030 174936 139044 174992
rect 138980 174932 139044 174936
rect 197492 174524 197556 174588
rect 201540 173496 201604 173500
rect 201540 173440 201554 173496
rect 201554 173440 201604 173496
rect 201540 173436 201604 173440
rect 161428 171124 161492 171188
rect 142108 171048 142172 171052
rect 142108 170992 142122 171048
rect 142122 170992 142172 171048
rect 142108 170988 142172 170992
rect 161428 170988 161492 171052
rect 142108 161604 142172 161668
rect 161428 161468 161492 161532
rect 142108 161392 142172 161396
rect 142108 161336 142122 161392
rect 142122 161336 142172 161392
rect 142108 161332 142172 161336
rect 161428 161332 161492 161396
rect 185348 152628 185412 152692
rect 185164 152492 185228 152556
rect 145236 152356 145300 152420
rect 142108 151948 142172 152012
rect 161428 151812 161492 151876
rect 142108 151736 142172 151740
rect 142108 151680 142122 151736
rect 142122 151680 142172 151736
rect 142108 151676 142172 151680
rect 161428 151676 161492 151740
rect 181116 150316 181180 150380
rect 183876 150180 183940 150244
rect 203012 150044 203076 150108
rect 203196 149908 203260 149972
rect 182772 149772 182836 149836
rect 187372 149636 187436 149700
rect 187004 149152 187068 149156
rect 187004 149096 187018 149152
rect 187018 149096 187068 149152
rect 187004 149092 187068 149096
rect 143764 148412 143828 148476
rect 191604 148412 191668 148476
rect 188292 148276 188356 148340
rect 196572 147732 196636 147796
rect 199332 147732 199396 147796
rect 142476 147596 142540 147660
rect 193628 147596 193692 147660
rect 189396 147460 189460 147524
rect 192156 147324 192220 147388
rect 198964 147188 199028 147252
rect 183140 147052 183204 147116
rect 142292 146916 142356 146980
rect 181300 146916 181364 146980
rect 112852 145828 112916 145892
rect 194732 145828 194796 145892
rect 111196 145692 111260 145756
rect 120580 145556 120644 145620
rect 119660 144876 119724 144940
rect 115612 144740 115676 144804
rect 182956 144740 183020 144804
rect 116900 144604 116964 144668
rect 191972 144604 192036 144668
rect 114140 144468 114204 144532
rect 191788 144468 191852 144532
rect 117084 144332 117148 144396
rect 194548 144332 194612 144396
rect 118188 144196 118252 144260
rect 190500 144196 190564 144260
rect 115796 144060 115860 144124
rect 188108 144060 188172 144124
rect 113588 143924 113652 143988
rect 190500 143516 190564 143580
rect 111380 143380 111444 143444
rect 111564 143244 111628 143308
rect 121132 143108 121196 143172
rect 113956 142564 114020 142628
rect 142292 142292 142356 142356
rect 161612 142292 161676 142356
rect 189028 142156 189092 142220
rect 188844 142020 188908 142084
rect 142660 141884 142724 141948
rect 118372 141748 118436 141812
rect 117084 141612 117148 141676
rect 141372 141672 141436 141676
rect 141372 141616 141422 141672
rect 141422 141616 141436 141672
rect 141372 141612 141436 141616
rect 177620 141612 177684 141676
rect 120948 141476 121012 141540
rect 193444 141476 193508 141540
rect 118556 141340 118620 141404
rect 141556 141264 141620 141268
rect 141556 141208 141570 141264
rect 141570 141208 141620 141264
rect 141556 141204 141620 141208
rect 177252 141204 177316 141268
rect 189580 141204 189644 141268
rect 188108 141068 188172 141132
rect 192340 141204 192404 141268
rect 116532 140796 116596 140860
rect 186820 140796 186884 140860
rect 190868 140796 190932 140860
rect 120764 140660 120828 140724
rect 193260 140660 193324 140724
rect 193444 140660 193508 140724
rect 117820 140524 117884 140588
rect 193260 140584 193324 140588
rect 193260 140528 193274 140584
rect 193274 140528 193324 140584
rect 193260 140524 193324 140528
rect 108252 140388 108316 140452
rect 127756 140252 127820 140316
rect 113036 139980 113100 140044
rect 173940 140116 174004 140180
rect 186084 140252 186148 140316
rect 178724 140116 178788 140180
rect 179828 139980 179892 140044
rect 183324 139980 183388 140044
rect 184796 140040 184860 140044
rect 184796 139984 184810 140040
rect 184810 139984 184860 140040
rect 184796 139980 184860 139984
rect 119292 139844 119356 139908
rect 186084 139844 186148 139908
rect 173940 139708 174004 139772
rect 180012 139708 180076 139772
rect 180196 139436 180260 139500
rect 122052 139300 122116 139364
rect 126468 139300 126532 139364
rect 129596 139360 129660 139364
rect 129596 139304 129646 139360
rect 129646 139304 129660 139360
rect 129596 139300 129660 139304
rect 120028 139164 120092 139228
rect 120948 139028 121012 139092
rect 150940 139300 151004 139364
rect 118556 138620 118620 138684
rect 154804 139300 154868 139364
rect 155356 139300 155420 139364
rect 159220 139300 159284 139364
rect 159956 139360 160020 139364
rect 159956 139304 160006 139360
rect 160006 139304 160020 139360
rect 159956 139300 160020 139304
rect 195100 139436 195164 139500
rect 183324 138892 183388 138956
rect 184796 138484 184860 138548
rect 187004 138136 187068 138140
rect 187004 138080 187054 138136
rect 187054 138080 187068 138136
rect 187004 138076 187068 138080
rect 122788 138000 122852 138004
rect 122788 137944 122802 138000
rect 122802 137944 122852 138000
rect 122788 137940 122852 137944
rect 186084 137396 186148 137460
rect 189028 137260 189092 137324
rect 119660 130324 119724 130388
rect 120028 130324 120092 130388
rect 122788 128480 122852 128484
rect 122788 128424 122802 128480
rect 122802 128424 122852 128480
rect 122788 128420 122852 128424
rect 122788 122904 122852 122908
rect 122788 122848 122802 122904
rect 122802 122848 122852 122904
rect 122788 122844 122852 122848
rect 122788 122768 122852 122772
rect 122788 122712 122802 122768
rect 122802 122712 122852 122768
rect 122788 122708 122852 122712
rect 191052 114412 191116 114476
rect 122788 113324 122852 113388
rect 122788 112916 122852 112980
rect 122788 103592 122852 103596
rect 122788 103536 122802 103592
rect 122802 103536 122852 103592
rect 122788 103532 122852 103536
rect 122788 103260 122852 103324
rect 119476 96596 119540 96660
rect 122788 93936 122852 93940
rect 122788 93880 122802 93936
rect 122802 93880 122852 93936
rect 122788 93876 122852 93880
rect 122788 93604 122852 93668
rect 122788 89720 122852 89724
rect 122788 89664 122802 89720
rect 122802 89664 122852 89720
rect 122788 89660 122852 89664
rect 119292 84220 119356 84284
rect 119660 83404 119724 83468
rect 120028 83404 120092 83468
rect 127572 81908 127636 81972
rect 145788 81908 145852 81972
rect 160692 81908 160756 81972
rect 161244 81908 161308 81972
rect 185348 81908 185412 81972
rect 122236 81364 122300 81428
rect 140820 81364 140884 81428
rect 141740 81364 141804 81428
rect 130700 81228 130764 81292
rect 143028 81228 143092 81292
rect 172468 81228 172532 81292
rect 130516 81092 130580 81156
rect 143396 81092 143460 81156
rect 171916 81092 171980 81156
rect 122972 80956 123036 81020
rect 143212 80956 143276 81020
rect 145420 80956 145484 81020
rect 147628 80956 147692 81020
rect 155908 80956 155972 81020
rect 187188 81016 187252 81020
rect 187188 80960 187202 81016
rect 187202 80960 187252 81016
rect 187188 80956 187252 80960
rect 126652 80820 126716 80884
rect 146524 80820 146588 80884
rect 148364 80820 148428 80884
rect 161428 80820 161492 80884
rect 122420 80548 122484 80612
rect 146708 80684 146772 80748
rect 154436 80684 154500 80748
rect 180012 80820 180076 80884
rect 177252 80684 177316 80748
rect 178356 80744 178420 80748
rect 178356 80688 178406 80744
rect 178406 80688 178420 80744
rect 178356 80684 178420 80688
rect 133092 80548 133156 80612
rect 147444 80548 147508 80612
rect 133460 80412 133524 80476
rect 138612 80412 138676 80476
rect 147260 80412 147324 80476
rect 149468 80412 149532 80476
rect 159220 80548 159284 80612
rect 122788 80336 122852 80340
rect 122788 80280 122838 80336
rect 122838 80280 122852 80336
rect 122788 80276 122852 80280
rect 140820 80276 140884 80340
rect 141924 80276 141988 80340
rect 138612 80140 138676 80204
rect 161796 80412 161860 80476
rect 150940 80276 151004 80340
rect 151676 80276 151740 80340
rect 158852 80276 158916 80340
rect 178540 80412 178604 80476
rect 131620 79868 131684 79932
rect 134932 80004 134996 80068
rect 135116 80004 135180 80068
rect 126468 79732 126532 79796
rect 133460 79868 133524 79932
rect 134196 79868 134260 79932
rect 134748 79868 134812 79932
rect 135484 79868 135548 79932
rect 136404 79868 136468 79932
rect 136956 79928 137020 79932
rect 136956 79872 136960 79928
rect 136960 79872 137016 79928
rect 137016 79872 137020 79928
rect 136956 79868 137020 79872
rect 137876 80004 137940 80068
rect 137508 79868 137572 79932
rect 138060 79868 138124 79932
rect 138796 80004 138860 80068
rect 140268 80004 140332 80068
rect 140452 80004 140516 80068
rect 151860 80004 151924 80068
rect 138980 79928 139044 79932
rect 138980 79872 138984 79928
rect 138984 79872 139040 79928
rect 139040 79872 139044 79928
rect 138980 79868 139044 79872
rect 139532 79928 139596 79932
rect 139532 79872 139536 79928
rect 139536 79872 139592 79928
rect 139592 79872 139596 79928
rect 139532 79868 139596 79872
rect 139900 79868 139964 79932
rect 140636 79928 140700 79932
rect 140636 79872 140640 79928
rect 140640 79872 140696 79928
rect 140696 79872 140700 79928
rect 140636 79868 140700 79872
rect 141556 79868 141620 79932
rect 141740 79928 141804 79932
rect 141740 79872 141744 79928
rect 141744 79872 141800 79928
rect 141800 79872 141804 79928
rect 141740 79868 141804 79872
rect 133828 79732 133892 79796
rect 134380 79792 134444 79796
rect 134380 79736 134394 79792
rect 134394 79736 134444 79792
rect 134380 79732 134444 79736
rect 135668 79732 135732 79796
rect 143212 79868 143276 79932
rect 143948 79928 144012 79932
rect 143948 79872 143952 79928
rect 143952 79872 144008 79928
rect 144008 79872 144012 79928
rect 143948 79868 144012 79872
rect 145420 79868 145484 79932
rect 146524 79868 146588 79932
rect 146892 79868 146956 79932
rect 147444 79868 147508 79932
rect 147812 79868 147876 79932
rect 149100 79868 149164 79932
rect 120764 79596 120828 79660
rect 132908 79596 132972 79660
rect 138428 79732 138492 79796
rect 138796 79792 138860 79796
rect 138796 79736 138846 79792
rect 138846 79736 138860 79792
rect 138796 79732 138860 79736
rect 140084 79732 140148 79796
rect 140820 79732 140884 79796
rect 144132 79732 144196 79796
rect 145788 79792 145852 79796
rect 145788 79736 145838 79792
rect 145838 79736 145852 79792
rect 145788 79732 145852 79736
rect 146708 79732 146772 79796
rect 147260 79732 147324 79796
rect 147996 79792 148060 79796
rect 147996 79736 148000 79792
rect 148000 79736 148056 79792
rect 148056 79736 148060 79792
rect 147996 79732 148060 79736
rect 149836 79868 149900 79932
rect 149652 79732 149716 79796
rect 151124 79906 151128 79932
rect 151128 79906 151184 79932
rect 151184 79906 151188 79932
rect 151124 79868 151188 79906
rect 151492 79868 151556 79932
rect 151676 79928 151740 79932
rect 151676 79872 151680 79928
rect 151680 79872 151736 79928
rect 151736 79872 151740 79928
rect 151676 79868 151740 79872
rect 152228 79928 152292 79932
rect 152228 79872 152232 79928
rect 152232 79872 152288 79928
rect 152288 79872 152292 79928
rect 152228 79868 152292 79872
rect 154068 80004 154132 80068
rect 157196 80004 157260 80068
rect 154068 79868 154132 79932
rect 154436 79868 154500 79932
rect 154620 79868 154684 79932
rect 151308 79732 151372 79796
rect 151676 79732 151740 79796
rect 152044 79792 152108 79796
rect 152044 79736 152048 79792
rect 152048 79736 152104 79792
rect 152104 79736 152108 79792
rect 152044 79732 152108 79736
rect 152596 79732 152660 79796
rect 133644 79596 133708 79660
rect 135852 79596 135916 79660
rect 136036 79596 136100 79660
rect 137140 79656 137204 79660
rect 137140 79600 137154 79656
rect 137154 79600 137204 79656
rect 137140 79596 137204 79600
rect 137692 79596 137756 79660
rect 152412 79596 152476 79660
rect 153516 79596 153580 79660
rect 154068 79596 154132 79660
rect 155172 79868 155236 79932
rect 155540 79868 155604 79932
rect 173204 80276 173268 80340
rect 183692 80336 183756 80340
rect 190868 80548 190932 80612
rect 183692 80280 183742 80336
rect 183742 80280 183756 80336
rect 183692 80276 183756 80280
rect 162164 80004 162228 80068
rect 163268 80004 163332 80068
rect 155908 79928 155972 79932
rect 155908 79872 155912 79928
rect 155912 79872 155968 79928
rect 155968 79872 155972 79928
rect 155908 79868 155972 79872
rect 156460 79868 156524 79932
rect 157196 79868 157260 79932
rect 155356 79656 155420 79660
rect 155356 79600 155406 79656
rect 155406 79600 155420 79656
rect 155356 79596 155420 79600
rect 157012 79732 157076 79796
rect 158300 79868 158364 79932
rect 158116 79732 158180 79796
rect 159036 79732 159100 79796
rect 156828 79596 156892 79660
rect 158484 79596 158548 79660
rect 160140 79868 160204 79932
rect 160876 79868 160940 79932
rect 161244 79868 161308 79932
rect 161980 79906 161984 79932
rect 161984 79906 162040 79932
rect 162040 79906 162044 79932
rect 161980 79868 162044 79906
rect 159772 79656 159836 79660
rect 159772 79600 159822 79656
rect 159822 79600 159836 79656
rect 159772 79596 159836 79600
rect 138244 79460 138308 79524
rect 147076 79520 147140 79524
rect 147076 79464 147126 79520
rect 147126 79464 147140 79520
rect 147076 79460 147140 79464
rect 147444 79520 147508 79524
rect 147444 79464 147458 79520
rect 147458 79464 147508 79520
rect 147444 79460 147508 79464
rect 147628 79520 147692 79524
rect 147628 79464 147678 79520
rect 147678 79464 147692 79520
rect 147628 79460 147692 79464
rect 148180 79520 148244 79524
rect 148180 79464 148194 79520
rect 148194 79464 148244 79520
rect 148180 79460 148244 79464
rect 148548 79460 148612 79524
rect 149284 79460 149348 79524
rect 153884 79460 153948 79524
rect 159220 79460 159284 79524
rect 160876 79732 160940 79796
rect 161428 79732 161492 79796
rect 160508 79596 160572 79660
rect 161060 79460 161124 79524
rect 163452 79868 163516 79932
rect 166948 80140 167012 80204
rect 169156 80140 169220 80204
rect 169892 80140 169956 80204
rect 164556 79868 164620 79932
rect 164740 79868 164804 79932
rect 165292 79868 165356 79932
rect 166212 79868 166276 79932
rect 167684 79868 167748 79932
rect 168236 79906 168240 79932
rect 168240 79906 168296 79932
rect 168296 79906 168300 79932
rect 168236 79868 168300 79906
rect 168788 79868 168852 79932
rect 170812 80004 170876 80068
rect 169708 79906 169712 79932
rect 169712 79906 169768 79932
rect 169768 79906 169772 79932
rect 169708 79868 169772 79906
rect 171364 79906 171368 79932
rect 171368 79906 171424 79932
rect 171424 79906 171428 79932
rect 171364 79868 171428 79906
rect 171732 79868 171796 79932
rect 171916 79868 171980 79932
rect 173756 80004 173820 80068
rect 197676 80004 197740 80068
rect 172468 79868 172532 79932
rect 174308 79868 174372 79932
rect 175044 79868 175108 79932
rect 175412 79928 175476 79932
rect 175412 79872 175416 79928
rect 175416 79872 175472 79928
rect 175472 79872 175476 79928
rect 175412 79868 175476 79872
rect 175780 79868 175844 79932
rect 176148 79868 176212 79932
rect 164004 79732 164068 79796
rect 166028 79792 166092 79796
rect 166028 79736 166032 79792
rect 166032 79736 166088 79792
rect 166088 79736 166092 79792
rect 166028 79732 166092 79736
rect 166396 79732 166460 79796
rect 167500 79732 167564 79796
rect 169340 79732 169404 79796
rect 161796 79656 161860 79660
rect 161796 79600 161846 79656
rect 161846 79600 161860 79656
rect 161796 79596 161860 79600
rect 162348 79596 162412 79660
rect 163636 79596 163700 79660
rect 164924 79596 164988 79660
rect 167684 79596 167748 79660
rect 168972 79596 169036 79660
rect 169524 79656 169588 79660
rect 169524 79600 169538 79656
rect 169538 79600 169588 79656
rect 169524 79596 169588 79600
rect 170076 79596 170140 79660
rect 170996 79732 171060 79796
rect 171548 79732 171612 79796
rect 172100 79792 172164 79796
rect 172100 79736 172114 79792
rect 172114 79736 172164 79792
rect 172100 79732 172164 79736
rect 172836 79732 172900 79796
rect 175044 79732 175108 79796
rect 175918 79792 175982 79796
rect 175918 79736 175922 79792
rect 175922 79736 175978 79792
rect 175978 79736 175982 79792
rect 175918 79732 175982 79736
rect 176148 79792 176212 79796
rect 176148 79736 176152 79792
rect 176152 79736 176208 79792
rect 176208 79736 176212 79792
rect 176148 79732 176212 79736
rect 176516 79732 176580 79796
rect 170628 79596 170692 79660
rect 176884 79868 176948 79932
rect 177620 79928 177684 79932
rect 177620 79872 177634 79928
rect 177634 79872 177684 79928
rect 177620 79868 177684 79872
rect 197860 79868 197924 79932
rect 177068 79732 177132 79796
rect 162532 79460 162596 79524
rect 162900 79460 162964 79524
rect 177068 79596 177132 79660
rect 178172 79792 178236 79796
rect 178172 79736 178222 79792
rect 178222 79736 178236 79792
rect 178172 79732 178236 79736
rect 178540 79596 178604 79660
rect 132356 79324 132420 79388
rect 152780 79384 152844 79388
rect 152780 79328 152830 79384
rect 152830 79328 152844 79384
rect 152780 79324 152844 79328
rect 153700 79324 153764 79388
rect 154804 79324 154868 79388
rect 155724 79384 155788 79388
rect 155724 79328 155738 79384
rect 155738 79328 155788 79384
rect 155724 79324 155788 79328
rect 157748 79324 157812 79388
rect 157932 79324 157996 79388
rect 161612 79324 161676 79388
rect 125364 79188 125428 79252
rect 148916 79188 148980 79252
rect 129596 79052 129660 79116
rect 151124 79052 151188 79116
rect 151308 79112 151372 79116
rect 152044 79188 152108 79252
rect 164740 79188 164804 79252
rect 165292 79188 165356 79252
rect 166580 79188 166644 79252
rect 167316 79248 167380 79252
rect 167316 79192 167330 79248
rect 167330 79192 167380 79248
rect 167316 79188 167380 79192
rect 168052 79188 168116 79252
rect 168236 79248 168300 79252
rect 168236 79192 168250 79248
rect 168250 79192 168300 79248
rect 168236 79188 168300 79192
rect 168604 79188 168668 79252
rect 171732 79188 171796 79252
rect 172284 79384 172348 79388
rect 172284 79328 172334 79384
rect 172334 79328 172348 79384
rect 172284 79324 172348 79328
rect 173020 79384 173084 79388
rect 173020 79328 173034 79384
rect 173034 79328 173084 79384
rect 173020 79324 173084 79328
rect 174492 79384 174556 79388
rect 174492 79328 174506 79384
rect 174506 79328 174556 79384
rect 174492 79324 174556 79328
rect 176148 79324 176212 79388
rect 177252 79324 177316 79388
rect 191052 79324 191116 79388
rect 172284 79188 172348 79252
rect 189212 79188 189276 79252
rect 151308 79056 151358 79112
rect 151358 79056 151372 79112
rect 151308 79052 151372 79056
rect 166580 79052 166644 79116
rect 190500 79052 190564 79116
rect 122604 78916 122668 78980
rect 138060 78916 138124 78980
rect 139164 78976 139228 78980
rect 139164 78920 139214 78976
rect 139214 78920 139228 78976
rect 139164 78916 139228 78920
rect 140636 78916 140700 78980
rect 141372 78916 141436 78980
rect 142476 78976 142540 78980
rect 142476 78920 142490 78976
rect 142490 78920 142540 78976
rect 142476 78916 142540 78920
rect 143396 78916 143460 78980
rect 149836 78916 149900 78980
rect 154620 78916 154684 78980
rect 158300 78916 158364 78980
rect 159956 78916 160020 78980
rect 173204 78916 173268 78980
rect 173572 78916 173636 78980
rect 203196 78916 203260 78980
rect 122052 78780 122116 78844
rect 158116 78780 158180 78844
rect 160692 78780 160756 78844
rect 171916 78780 171980 78844
rect 172652 78780 172716 78844
rect 174492 78780 174556 78844
rect 130884 78644 130948 78708
rect 151308 78704 151372 78708
rect 151308 78648 151322 78704
rect 151322 78648 151372 78704
rect 151308 78644 151372 78648
rect 156460 78644 156524 78708
rect 163452 78644 163516 78708
rect 165844 78644 165908 78708
rect 166396 78644 166460 78708
rect 174676 78644 174740 78708
rect 175780 78644 175844 78708
rect 175964 78644 176028 78708
rect 130332 78568 130396 78572
rect 130332 78512 130382 78568
rect 130382 78512 130396 78568
rect 130332 78508 130396 78512
rect 133460 78508 133524 78572
rect 134564 78508 134628 78572
rect 136220 78568 136284 78572
rect 136220 78512 136234 78568
rect 136234 78512 136284 78568
rect 136220 78508 136284 78512
rect 136588 78508 136652 78572
rect 136956 78568 137020 78572
rect 136956 78512 136970 78568
rect 136970 78512 137020 78568
rect 136956 78508 137020 78512
rect 138060 78568 138124 78572
rect 138060 78512 138074 78568
rect 138074 78512 138124 78568
rect 138060 78508 138124 78512
rect 141004 78508 141068 78572
rect 143028 78508 143092 78572
rect 151492 78508 151556 78572
rect 156644 78508 156708 78572
rect 158300 78508 158364 78572
rect 161060 78568 161124 78572
rect 161060 78512 161110 78568
rect 161110 78512 161124 78568
rect 161060 78508 161124 78512
rect 162716 78568 162780 78572
rect 162716 78512 162766 78568
rect 162766 78512 162780 78568
rect 162716 78508 162780 78512
rect 184980 78508 185044 78572
rect 186820 78508 186884 78572
rect 187372 78568 187436 78572
rect 187372 78512 187422 78568
rect 187422 78512 187436 78568
rect 187372 78508 187436 78512
rect 193628 78568 193692 78572
rect 193628 78512 193642 78568
rect 193642 78512 193692 78568
rect 193628 78508 193692 78512
rect 125180 78372 125244 78436
rect 141740 78432 141804 78436
rect 141740 78376 141754 78432
rect 141754 78376 141804 78432
rect 141740 78372 141804 78376
rect 143212 78372 143276 78436
rect 165476 78432 165540 78436
rect 165476 78376 165526 78432
rect 165526 78376 165540 78432
rect 165476 78372 165540 78376
rect 171364 78372 171428 78436
rect 126836 78236 126900 78300
rect 138612 78296 138676 78300
rect 138612 78240 138626 78296
rect 138626 78240 138676 78296
rect 138612 78236 138676 78240
rect 148180 78236 148244 78300
rect 150020 78236 150084 78300
rect 124076 78100 124140 78164
rect 155172 78160 155236 78164
rect 155172 78104 155186 78160
rect 155186 78104 155236 78160
rect 155172 78100 155236 78104
rect 127388 77964 127452 78028
rect 148732 77964 148796 78028
rect 164556 78236 164620 78300
rect 164004 78100 164068 78164
rect 167868 78100 167932 78164
rect 170812 78100 170876 78164
rect 173756 77964 173820 78028
rect 119844 77828 119908 77892
rect 133276 77888 133340 77892
rect 133276 77832 133290 77888
rect 133290 77832 133340 77888
rect 133276 77828 133340 77832
rect 134748 77828 134812 77892
rect 136036 77828 136100 77892
rect 137876 77828 137940 77892
rect 138980 77828 139044 77892
rect 139716 77828 139780 77892
rect 140084 77888 140148 77892
rect 140084 77832 140098 77888
rect 140098 77832 140148 77888
rect 140084 77828 140148 77832
rect 140820 77828 140884 77892
rect 147076 77828 147140 77892
rect 147996 77828 148060 77892
rect 149100 77828 149164 77892
rect 160324 77828 160388 77892
rect 176332 77828 176396 77892
rect 124812 77692 124876 77756
rect 142292 77752 142356 77756
rect 142292 77696 142342 77752
rect 142342 77696 142356 77752
rect 142292 77692 142356 77696
rect 145052 77692 145116 77756
rect 146892 77692 146956 77756
rect 147812 77692 147876 77756
rect 149284 77692 149348 77756
rect 165476 77692 165540 77756
rect 172468 77692 172532 77756
rect 131988 77556 132052 77620
rect 136404 77556 136468 77620
rect 137508 77616 137572 77620
rect 137508 77560 137558 77616
rect 137558 77560 137572 77616
rect 137508 77556 137572 77560
rect 137692 77420 137756 77484
rect 124996 77284 125060 77348
rect 145604 77556 145668 77620
rect 157012 77556 157076 77620
rect 163636 77556 163700 77620
rect 164556 77556 164620 77620
rect 173940 77556 174004 77620
rect 138244 77420 138308 77484
rect 147996 77420 148060 77484
rect 148364 77420 148428 77484
rect 154068 77420 154132 77484
rect 165108 77420 165172 77484
rect 170812 77480 170876 77484
rect 170812 77424 170862 77480
rect 170862 77424 170876 77480
rect 170812 77420 170876 77424
rect 144316 77284 144380 77348
rect 154436 77344 154500 77348
rect 154436 77288 154486 77344
rect 154486 77288 154500 77344
rect 154436 77284 154500 77288
rect 170444 77344 170508 77348
rect 170444 77288 170494 77344
rect 170494 77288 170508 77344
rect 170444 77284 170508 77288
rect 170996 77284 171060 77348
rect 146892 77148 146956 77212
rect 178724 77148 178788 77212
rect 148364 77012 148428 77076
rect 181484 77012 181548 77076
rect 193444 76876 193508 76940
rect 192156 76740 192220 76804
rect 135484 76468 135548 76532
rect 189396 76468 189460 76532
rect 193260 76332 193324 76396
rect 175412 76196 175476 76260
rect 172100 76120 172164 76124
rect 172100 76064 172150 76120
rect 172150 76064 172164 76120
rect 172100 76060 172164 76064
rect 173572 76060 173636 76124
rect 157932 75924 157996 75988
rect 169340 75984 169404 75988
rect 169340 75928 169390 75984
rect 169390 75928 169404 75984
rect 169340 75924 169404 75928
rect 171916 75924 171980 75988
rect 117084 75788 117148 75852
rect 174860 75788 174924 75852
rect 147076 75652 147140 75716
rect 176516 75712 176580 75716
rect 176516 75656 176566 75712
rect 176566 75656 176580 75712
rect 176516 75652 176580 75656
rect 148916 75516 148980 75580
rect 203012 75516 203076 75580
rect 196388 75380 196452 75444
rect 119844 75108 119908 75172
rect 159036 74972 159100 75036
rect 154252 74564 154316 74628
rect 120580 74428 120644 74492
rect 156460 74428 156524 74492
rect 143948 74352 144012 74356
rect 143948 74296 143962 74352
rect 143962 74296 144012 74352
rect 143948 74292 144012 74296
rect 181116 74292 181180 74356
rect 161244 74216 161308 74220
rect 161244 74160 161258 74216
rect 161258 74160 161308 74216
rect 161244 74156 161308 74160
rect 198964 74156 199028 74220
rect 144132 74020 144196 74084
rect 135668 73884 135732 73948
rect 149652 73884 149716 73948
rect 135300 73748 135364 73812
rect 152964 73748 153028 73812
rect 167684 73748 167748 73812
rect 173756 73748 173820 73812
rect 166764 73612 166828 73676
rect 152596 73476 152660 73540
rect 168052 73476 168116 73540
rect 168052 73340 168116 73404
rect 121316 73068 121380 73132
rect 179644 73128 179708 73132
rect 179644 73072 179694 73128
rect 179694 73072 179708 73128
rect 179644 73068 179708 73072
rect 180932 73068 180996 73132
rect 152596 72932 152660 72996
rect 183876 72932 183940 72996
rect 149284 72796 149348 72860
rect 149836 72796 149900 72860
rect 183140 72796 183204 72860
rect 142292 72524 142356 72588
rect 179828 72660 179892 72724
rect 185164 72524 185228 72588
rect 169708 72388 169772 72452
rect 158852 71844 158916 71908
rect 149100 71708 149164 71772
rect 162532 71768 162596 71772
rect 162532 71712 162546 71768
rect 162546 71712 162596 71768
rect 162532 71708 162596 71712
rect 120028 71572 120092 71636
rect 118556 71436 118620 71500
rect 152412 71436 152476 71500
rect 145052 71300 145116 71364
rect 166948 71300 167012 71364
rect 145604 71164 145668 71228
rect 148916 71028 148980 71092
rect 144316 70484 144380 70548
rect 195100 70408 195164 70412
rect 195100 70352 195150 70408
rect 195150 70352 195164 70408
rect 195100 70348 195164 70352
rect 191604 70212 191668 70276
rect 166948 70076 167012 70140
rect 200804 69532 200868 69596
rect 169156 68988 169220 69052
rect 120948 68852 121012 68916
rect 200988 68852 201052 68916
rect 144500 68776 144564 68780
rect 144500 68720 144550 68776
rect 144550 68720 144564 68776
rect 144500 68716 144564 68720
rect 150020 68716 150084 68780
rect 179460 68716 179524 68780
rect 148180 68580 148244 68644
rect 144684 68444 144748 68508
rect 140820 68308 140884 68372
rect 188292 68776 188356 68780
rect 188292 68720 188306 68776
rect 188306 68720 188356 68776
rect 188292 68716 188356 68720
rect 131620 68172 131684 68236
rect 147076 68172 147140 68236
rect 160876 67688 160940 67692
rect 160876 67632 160926 67688
rect 160926 67632 160940 67688
rect 160876 67628 160940 67632
rect 138612 67492 138676 67556
rect 161244 67492 161308 67556
rect 151308 67356 151372 67420
rect 182588 67356 182652 67420
rect 148364 67220 148428 67284
rect 137508 66948 137572 67012
rect 133828 66812 133892 66876
rect 146892 66812 146956 66876
rect 176148 66676 176212 66740
rect 200620 66812 200684 66876
rect 139900 66132 139964 66196
rect 187924 66132 187988 66196
rect 188108 66192 188172 66196
rect 188108 66136 188122 66192
rect 188122 66136 188172 66192
rect 188108 66132 188172 66136
rect 139716 65996 139780 66060
rect 161980 65996 162044 66060
rect 187924 65588 187988 65652
rect 133092 65452 133156 65516
rect 188108 65044 188172 65108
rect 197492 65104 197556 65108
rect 197492 65048 197542 65104
rect 197542 65048 197556 65104
rect 197492 65044 197556 65048
rect 135852 64772 135916 64836
rect 152964 64772 153028 64836
rect 174676 64636 174740 64700
rect 201724 64636 201788 64700
rect 171916 64500 171980 64564
rect 197308 64500 197372 64564
rect 201724 64092 201788 64156
rect 139532 63412 139596 63476
rect 157932 63412 157996 63476
rect 138428 63276 138492 63340
rect 165108 63004 165172 63068
rect 172100 62868 172164 62932
rect 196572 62868 196636 62932
rect 176332 62732 176396 62796
rect 201908 62732 201972 62796
rect 151492 62052 151556 62116
rect 183692 62052 183756 62116
rect 187740 61916 187804 61980
rect 156828 61780 156892 61844
rect 151676 61236 151740 61300
rect 180564 61236 180628 61300
rect 138244 60556 138308 60620
rect 155724 60556 155788 60620
rect 158116 60420 158180 60484
rect 173572 60284 173636 60348
rect 198964 60284 199028 60348
rect 147260 59876 147324 59940
rect 198964 59876 199028 59940
rect 140084 59196 140148 59260
rect 160692 59196 160756 59260
rect 158300 59060 158364 59124
rect 174860 58924 174924 58988
rect 138060 57836 138124 57900
rect 157012 57836 157076 57900
rect 165292 57700 165356 57764
rect 175044 57564 175108 57628
rect 201540 57564 201604 57628
rect 202828 57564 202892 57628
rect 202828 57156 202892 57220
rect 163268 56476 163332 56540
rect 149836 56340 149900 56404
rect 157196 56204 157260 56268
rect 167684 55932 167748 55996
rect 170444 55796 170508 55860
rect 136588 55116 136652 55180
rect 160876 55116 160940 55180
rect 113772 55040 113836 55044
rect 113772 54984 113822 55040
rect 113822 54984 113836 55040
rect 113772 54980 113836 54984
rect 158484 54980 158548 55044
rect 148180 54844 148244 54908
rect 165476 54436 165540 54500
rect 196204 54436 196268 54500
rect 166580 53756 166644 53820
rect 162532 53620 162596 53684
rect 154252 53484 154316 53548
rect 182772 53484 182836 53548
rect 158852 53348 158916 53412
rect 134196 52396 134260 52460
rect 170628 52396 170692 52460
rect 169340 52260 169404 52324
rect 203012 52260 203076 52324
rect 204116 52260 204180 52324
rect 161244 52124 161308 52188
rect 161060 51988 161124 52052
rect 204116 51852 204180 51916
rect 159036 50900 159100 50964
rect 166764 50764 166828 50828
rect 163452 50628 163516 50692
rect 177068 50220 177132 50284
rect 135668 49540 135732 49604
rect 167868 49540 167932 49604
rect 170812 49404 170876 49468
rect 198780 49404 198844 49468
rect 175964 49268 176028 49332
rect 198780 48996 198844 49060
rect 135484 48180 135548 48244
rect 162716 48180 162780 48244
rect 196020 48180 196084 48244
rect 173756 48044 173820 48108
rect 196020 47636 196084 47700
rect 147444 47500 147508 47564
rect 135300 46820 135364 46884
rect 169524 46820 169588 46884
rect 170996 46684 171060 46748
rect 192340 45596 192404 45660
rect 163636 45460 163700 45524
rect 148916 45052 148980 45116
rect 152596 44916 152660 44980
rect 116532 44236 116596 44300
rect 168052 44100 168116 44164
rect 154436 43964 154500 44028
rect 187004 43964 187068 44028
rect 187004 43556 187068 43620
rect 172284 42740 172348 42804
rect 145604 37844 145668 37908
rect 133644 33764 133708 33828
rect 144684 33764 144748 33828
rect 117820 31724 117884 31788
rect 189580 31724 189644 31788
rect 149652 30908 149716 30972
rect 152412 28188 152476 28252
rect 144500 26828 144564 26892
rect 108252 19348 108316 19412
rect 145420 17172 145484 17236
rect 144132 15812 144196 15876
rect 144316 11596 144380 11660
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 682954 -8106 711002
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 -8106 682954
rect -8726 682634 -8106 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 -8106 682634
rect -8726 646954 -8106 682398
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 -8106 646954
rect -8726 646634 -8106 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 -8106 646634
rect -8726 610954 -8106 646398
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 -8106 610954
rect -8726 610634 -8106 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 -8106 610634
rect -8726 574954 -8106 610398
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 -8106 574954
rect -8726 574634 -8106 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 -8106 574634
rect -8726 538954 -8106 574398
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 -8106 538954
rect -8726 538634 -8106 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 -8106 538634
rect -8726 502954 -8106 538398
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 -8106 502954
rect -8726 502634 -8106 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 -8106 502634
rect -8726 466954 -8106 502398
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 -8106 466954
rect -8726 466634 -8106 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 -8106 466634
rect -8726 430954 -8106 466398
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 -8106 430954
rect -8726 430634 -8106 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 -8106 430634
rect -8726 394954 -8106 430398
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 -8106 394954
rect -8726 394634 -8106 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 -8106 394634
rect -8726 358954 -8106 394398
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 -8106 358954
rect -8726 358634 -8106 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 -8106 358634
rect -8726 322954 -8106 358398
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 -8106 322954
rect -8726 322634 -8106 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 -8106 322634
rect -8726 286954 -8106 322398
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 -8106 286954
rect -8726 286634 -8106 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 -8106 286634
rect -8726 250954 -8106 286398
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 -8106 250954
rect -8726 250634 -8106 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 -8106 250634
rect -8726 214954 -8106 250398
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 -8106 214954
rect -8726 214634 -8106 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 -8106 214634
rect -8726 178954 -8106 214398
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 -8106 178954
rect -8726 178634 -8106 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 -8106 178634
rect -8726 142954 -8106 178398
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 -8106 142954
rect -8726 142634 -8106 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 -8106 142634
rect -8726 106954 -8106 142398
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 -8106 106954
rect -8726 106634 -8106 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 -8106 106634
rect -8726 70954 -8106 106398
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 -8106 70954
rect -8726 70634 -8106 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 -8106 70634
rect -8726 34954 -8106 70398
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 -8106 34954
rect -8726 34634 -8106 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 -8106 34634
rect -8726 -7066 -8106 34398
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 678454 -7146 710042
rect -7766 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 -7146 678454
rect -7766 678134 -7146 678218
rect -7766 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 -7146 678134
rect -7766 642454 -7146 677898
rect -7766 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 -7146 642454
rect -7766 642134 -7146 642218
rect -7766 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 -7146 642134
rect -7766 606454 -7146 641898
rect -7766 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 -7146 606454
rect -7766 606134 -7146 606218
rect -7766 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 -7146 606134
rect -7766 570454 -7146 605898
rect -7766 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 -7146 570454
rect -7766 570134 -7146 570218
rect -7766 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 -7146 570134
rect -7766 534454 -7146 569898
rect -7766 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 -7146 534454
rect -7766 534134 -7146 534218
rect -7766 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 -7146 534134
rect -7766 498454 -7146 533898
rect -7766 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 -7146 498454
rect -7766 498134 -7146 498218
rect -7766 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 -7146 498134
rect -7766 462454 -7146 497898
rect -7766 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 -7146 462454
rect -7766 462134 -7146 462218
rect -7766 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 -7146 462134
rect -7766 426454 -7146 461898
rect -7766 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 -7146 426454
rect -7766 426134 -7146 426218
rect -7766 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 -7146 426134
rect -7766 390454 -7146 425898
rect -7766 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 -7146 390454
rect -7766 390134 -7146 390218
rect -7766 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 -7146 390134
rect -7766 354454 -7146 389898
rect -7766 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 -7146 354454
rect -7766 354134 -7146 354218
rect -7766 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 -7146 354134
rect -7766 318454 -7146 353898
rect -7766 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 -7146 318454
rect -7766 318134 -7146 318218
rect -7766 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 -7146 318134
rect -7766 282454 -7146 317898
rect -7766 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 -7146 282454
rect -7766 282134 -7146 282218
rect -7766 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 -7146 282134
rect -7766 246454 -7146 281898
rect -7766 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 -7146 246454
rect -7766 246134 -7146 246218
rect -7766 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 -7146 246134
rect -7766 210454 -7146 245898
rect -7766 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 -7146 210454
rect -7766 210134 -7146 210218
rect -7766 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 -7146 210134
rect -7766 174454 -7146 209898
rect -7766 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 -7146 174454
rect -7766 174134 -7146 174218
rect -7766 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 -7146 174134
rect -7766 138454 -7146 173898
rect -7766 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 -7146 138454
rect -7766 138134 -7146 138218
rect -7766 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 -7146 138134
rect -7766 102454 -7146 137898
rect -7766 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 -7146 102454
rect -7766 102134 -7146 102218
rect -7766 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 -7146 102134
rect -7766 66454 -7146 101898
rect -7766 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 -7146 66454
rect -7766 66134 -7146 66218
rect -7766 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 -7146 66134
rect -7766 30454 -7146 65898
rect -7766 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 -7146 30454
rect -7766 30134 -7146 30218
rect -7766 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 -7146 30134
rect -7766 -6106 -7146 29898
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 673954 -6186 709082
rect -6806 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 -6186 673954
rect -6806 673634 -6186 673718
rect -6806 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 -6186 673634
rect -6806 637954 -6186 673398
rect -6806 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 -6186 637954
rect -6806 637634 -6186 637718
rect -6806 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 -6186 637634
rect -6806 601954 -6186 637398
rect -6806 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 -6186 601954
rect -6806 601634 -6186 601718
rect -6806 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 -6186 601634
rect -6806 565954 -6186 601398
rect -6806 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 -6186 565954
rect -6806 565634 -6186 565718
rect -6806 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 -6186 565634
rect -6806 529954 -6186 565398
rect -6806 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 -6186 529954
rect -6806 529634 -6186 529718
rect -6806 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 -6186 529634
rect -6806 493954 -6186 529398
rect -6806 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 -6186 493954
rect -6806 493634 -6186 493718
rect -6806 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 -6186 493634
rect -6806 457954 -6186 493398
rect -6806 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 -6186 457954
rect -6806 457634 -6186 457718
rect -6806 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 -6186 457634
rect -6806 421954 -6186 457398
rect -6806 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 -6186 421954
rect -6806 421634 -6186 421718
rect -6806 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 -6186 421634
rect -6806 385954 -6186 421398
rect -6806 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 -6186 385954
rect -6806 385634 -6186 385718
rect -6806 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 -6186 385634
rect -6806 349954 -6186 385398
rect -6806 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 -6186 349954
rect -6806 349634 -6186 349718
rect -6806 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 -6186 349634
rect -6806 313954 -6186 349398
rect -6806 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 -6186 313954
rect -6806 313634 -6186 313718
rect -6806 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 -6186 313634
rect -6806 277954 -6186 313398
rect -6806 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 -6186 277954
rect -6806 277634 -6186 277718
rect -6806 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 -6186 277634
rect -6806 241954 -6186 277398
rect -6806 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 -6186 241954
rect -6806 241634 -6186 241718
rect -6806 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 -6186 241634
rect -6806 205954 -6186 241398
rect -6806 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 -6186 205954
rect -6806 205634 -6186 205718
rect -6806 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 -6186 205634
rect -6806 169954 -6186 205398
rect -6806 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 -6186 169954
rect -6806 169634 -6186 169718
rect -6806 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 -6186 169634
rect -6806 133954 -6186 169398
rect -6806 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 -6186 133954
rect -6806 133634 -6186 133718
rect -6806 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 -6186 133634
rect -6806 97954 -6186 133398
rect -6806 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 -6186 97954
rect -6806 97634 -6186 97718
rect -6806 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 -6186 97634
rect -6806 61954 -6186 97398
rect -6806 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 -6186 61954
rect -6806 61634 -6186 61718
rect -6806 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 -6186 61634
rect -6806 25954 -6186 61398
rect -6806 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 -6186 25954
rect -6806 25634 -6186 25718
rect -6806 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 -6186 25634
rect -6806 -5146 -6186 25398
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 669454 -5226 708122
rect -5846 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 -5226 669454
rect -5846 669134 -5226 669218
rect -5846 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 -5226 669134
rect -5846 633454 -5226 668898
rect -5846 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 -5226 633454
rect -5846 633134 -5226 633218
rect -5846 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 -5226 633134
rect -5846 597454 -5226 632898
rect -5846 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 -5226 597454
rect -5846 597134 -5226 597218
rect -5846 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 -5226 597134
rect -5846 561454 -5226 596898
rect -5846 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 -5226 561454
rect -5846 561134 -5226 561218
rect -5846 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 -5226 561134
rect -5846 525454 -5226 560898
rect -5846 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 -5226 525454
rect -5846 525134 -5226 525218
rect -5846 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 -5226 525134
rect -5846 489454 -5226 524898
rect -5846 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 -5226 489454
rect -5846 489134 -5226 489218
rect -5846 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 -5226 489134
rect -5846 453454 -5226 488898
rect -5846 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 -5226 453454
rect -5846 453134 -5226 453218
rect -5846 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 -5226 453134
rect -5846 417454 -5226 452898
rect -5846 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 -5226 417454
rect -5846 417134 -5226 417218
rect -5846 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 -5226 417134
rect -5846 381454 -5226 416898
rect -5846 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 -5226 381454
rect -5846 381134 -5226 381218
rect -5846 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 -5226 381134
rect -5846 345454 -5226 380898
rect -5846 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 -5226 345454
rect -5846 345134 -5226 345218
rect -5846 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 -5226 345134
rect -5846 309454 -5226 344898
rect -5846 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 -5226 309454
rect -5846 309134 -5226 309218
rect -5846 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 -5226 309134
rect -5846 273454 -5226 308898
rect -5846 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 -5226 273454
rect -5846 273134 -5226 273218
rect -5846 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 -5226 273134
rect -5846 237454 -5226 272898
rect -5846 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 -5226 237454
rect -5846 237134 -5226 237218
rect -5846 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 -5226 237134
rect -5846 201454 -5226 236898
rect -5846 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 -5226 201454
rect -5846 201134 -5226 201218
rect -5846 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 -5226 201134
rect -5846 165454 -5226 200898
rect -5846 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 -5226 165454
rect -5846 165134 -5226 165218
rect -5846 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 -5226 165134
rect -5846 129454 -5226 164898
rect -5846 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 -5226 129454
rect -5846 129134 -5226 129218
rect -5846 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 -5226 129134
rect -5846 93454 -5226 128898
rect -5846 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 -5226 93454
rect -5846 93134 -5226 93218
rect -5846 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 -5226 93134
rect -5846 57454 -5226 92898
rect -5846 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 -5226 57454
rect -5846 57134 -5226 57218
rect -5846 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 -5226 57134
rect -5846 21454 -5226 56898
rect -5846 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 -5226 21454
rect -5846 21134 -5226 21218
rect -5846 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 -5226 21134
rect -5846 -4186 -5226 20898
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 700954 -4266 707162
rect -4886 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 -4266 700954
rect -4886 700634 -4266 700718
rect -4886 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 -4266 700634
rect -4886 664954 -4266 700398
rect -4886 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 -4266 664954
rect -4886 664634 -4266 664718
rect -4886 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 -4266 664634
rect -4886 628954 -4266 664398
rect -4886 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 -4266 628954
rect -4886 628634 -4266 628718
rect -4886 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 -4266 628634
rect -4886 592954 -4266 628398
rect -4886 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 -4266 592954
rect -4886 592634 -4266 592718
rect -4886 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 -4266 592634
rect -4886 556954 -4266 592398
rect -4886 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 -4266 556954
rect -4886 556634 -4266 556718
rect -4886 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 -4266 556634
rect -4886 520954 -4266 556398
rect -4886 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 -4266 520954
rect -4886 520634 -4266 520718
rect -4886 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 -4266 520634
rect -4886 484954 -4266 520398
rect -4886 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 -4266 484954
rect -4886 484634 -4266 484718
rect -4886 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 -4266 484634
rect -4886 448954 -4266 484398
rect -4886 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 -4266 448954
rect -4886 448634 -4266 448718
rect -4886 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 -4266 448634
rect -4886 412954 -4266 448398
rect -4886 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 -4266 412954
rect -4886 412634 -4266 412718
rect -4886 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 -4266 412634
rect -4886 376954 -4266 412398
rect -4886 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 -4266 376954
rect -4886 376634 -4266 376718
rect -4886 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 -4266 376634
rect -4886 340954 -4266 376398
rect -4886 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 -4266 340954
rect -4886 340634 -4266 340718
rect -4886 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 -4266 340634
rect -4886 304954 -4266 340398
rect -4886 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 -4266 304954
rect -4886 304634 -4266 304718
rect -4886 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 -4266 304634
rect -4886 268954 -4266 304398
rect -4886 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 -4266 268954
rect -4886 268634 -4266 268718
rect -4886 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 -4266 268634
rect -4886 232954 -4266 268398
rect -4886 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 -4266 232954
rect -4886 232634 -4266 232718
rect -4886 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 -4266 232634
rect -4886 196954 -4266 232398
rect -4886 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 -4266 196954
rect -4886 196634 -4266 196718
rect -4886 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 -4266 196634
rect -4886 160954 -4266 196398
rect -4886 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 -4266 160954
rect -4886 160634 -4266 160718
rect -4886 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 -4266 160634
rect -4886 124954 -4266 160398
rect -4886 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 -4266 124954
rect -4886 124634 -4266 124718
rect -4886 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 -4266 124634
rect -4886 88954 -4266 124398
rect -4886 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 -4266 88954
rect -4886 88634 -4266 88718
rect -4886 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 -4266 88634
rect -4886 52954 -4266 88398
rect -4886 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 -4266 52954
rect -4886 52634 -4266 52718
rect -4886 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 -4266 52634
rect -4886 16954 -4266 52398
rect -4886 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 -4266 16954
rect -4886 16634 -4266 16718
rect -4886 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 -4266 16634
rect -4886 -3226 -4266 16398
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 696454 -3306 706202
rect -3926 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 -3306 696454
rect -3926 696134 -3306 696218
rect -3926 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 -3306 696134
rect -3926 660454 -3306 695898
rect -3926 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 -3306 660454
rect -3926 660134 -3306 660218
rect -3926 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 -3306 660134
rect -3926 624454 -3306 659898
rect -3926 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 -3306 624454
rect -3926 624134 -3306 624218
rect -3926 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 -3306 624134
rect -3926 588454 -3306 623898
rect -3926 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 -3306 588454
rect -3926 588134 -3306 588218
rect -3926 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 -3306 588134
rect -3926 552454 -3306 587898
rect -3926 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 -3306 552454
rect -3926 552134 -3306 552218
rect -3926 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 -3306 552134
rect -3926 516454 -3306 551898
rect -3926 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 -3306 516454
rect -3926 516134 -3306 516218
rect -3926 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 -3306 516134
rect -3926 480454 -3306 515898
rect -3926 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 -3306 480454
rect -3926 480134 -3306 480218
rect -3926 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 -3306 480134
rect -3926 444454 -3306 479898
rect -3926 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 -3306 444454
rect -3926 444134 -3306 444218
rect -3926 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 -3306 444134
rect -3926 408454 -3306 443898
rect -3926 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 -3306 408454
rect -3926 408134 -3306 408218
rect -3926 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 -3306 408134
rect -3926 372454 -3306 407898
rect -3926 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 -3306 372454
rect -3926 372134 -3306 372218
rect -3926 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 -3306 372134
rect -3926 336454 -3306 371898
rect -3926 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 -3306 336454
rect -3926 336134 -3306 336218
rect -3926 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 -3306 336134
rect -3926 300454 -3306 335898
rect -3926 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 -3306 300454
rect -3926 300134 -3306 300218
rect -3926 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 -3306 300134
rect -3926 264454 -3306 299898
rect -3926 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 -3306 264454
rect -3926 264134 -3306 264218
rect -3926 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 -3306 264134
rect -3926 228454 -3306 263898
rect -3926 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 -3306 228454
rect -3926 228134 -3306 228218
rect -3926 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 -3306 228134
rect -3926 192454 -3306 227898
rect -3926 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 -3306 192454
rect -3926 192134 -3306 192218
rect -3926 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 -3306 192134
rect -3926 156454 -3306 191898
rect -3926 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 -3306 156454
rect -3926 156134 -3306 156218
rect -3926 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 -3306 156134
rect -3926 120454 -3306 155898
rect -3926 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 -3306 120454
rect -3926 120134 -3306 120218
rect -3926 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 -3306 120134
rect -3926 84454 -3306 119898
rect -3926 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 -3306 84454
rect -3926 84134 -3306 84218
rect -3926 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 -3306 84134
rect -3926 48454 -3306 83898
rect -3926 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 -3306 48454
rect -3926 48134 -3306 48218
rect -3926 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 -3306 48134
rect -3926 12454 -3306 47898
rect -3926 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 -3306 12454
rect -3926 12134 -3306 12218
rect -3926 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 -3306 12134
rect -3926 -2266 -3306 11898
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 691954 -2346 705242
rect -2966 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 -2346 691954
rect -2966 691634 -2346 691718
rect -2966 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 -2346 691634
rect -2966 655954 -2346 691398
rect -2966 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 -2346 655954
rect -2966 655634 -2346 655718
rect -2966 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 -2346 655634
rect -2966 619954 -2346 655398
rect -2966 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 -2346 619954
rect -2966 619634 -2346 619718
rect -2966 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 -2346 619634
rect -2966 583954 -2346 619398
rect -2966 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 -2346 583954
rect -2966 583634 -2346 583718
rect -2966 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 -2346 583634
rect -2966 547954 -2346 583398
rect -2966 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 -2346 547954
rect -2966 547634 -2346 547718
rect -2966 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 -2346 547634
rect -2966 511954 -2346 547398
rect -2966 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 -2346 511954
rect -2966 511634 -2346 511718
rect -2966 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 -2346 511634
rect -2966 475954 -2346 511398
rect -2966 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 -2346 475954
rect -2966 475634 -2346 475718
rect -2966 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 -2346 475634
rect -2966 439954 -2346 475398
rect -2966 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 -2346 439954
rect -2966 439634 -2346 439718
rect -2966 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 -2346 439634
rect -2966 403954 -2346 439398
rect -2966 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 -2346 403954
rect -2966 403634 -2346 403718
rect -2966 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 -2346 403634
rect -2966 367954 -2346 403398
rect -2966 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 -2346 367954
rect -2966 367634 -2346 367718
rect -2966 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 -2346 367634
rect -2966 331954 -2346 367398
rect -2966 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 -2346 331954
rect -2966 331634 -2346 331718
rect -2966 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 -2346 331634
rect -2966 295954 -2346 331398
rect -2966 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 -2346 295954
rect -2966 295634 -2346 295718
rect -2966 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 -2346 295634
rect -2966 259954 -2346 295398
rect -2966 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 -2346 259954
rect -2966 259634 -2346 259718
rect -2966 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 -2346 259634
rect -2966 223954 -2346 259398
rect -2966 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 -2346 223954
rect -2966 223634 -2346 223718
rect -2966 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 -2346 223634
rect -2966 187954 -2346 223398
rect -2966 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 -2346 187954
rect -2966 187634 -2346 187718
rect -2966 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 -2346 187634
rect -2966 151954 -2346 187398
rect -2966 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 -2346 151954
rect -2966 151634 -2346 151718
rect -2966 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 -2346 151634
rect -2966 115954 -2346 151398
rect -2966 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 -2346 115954
rect -2966 115634 -2346 115718
rect -2966 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 -2346 115634
rect -2966 79954 -2346 115398
rect -2966 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 -2346 79954
rect -2966 79634 -2346 79718
rect -2966 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 -2346 79634
rect -2966 43954 -2346 79398
rect -2966 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 -2346 43954
rect -2966 43634 -2346 43718
rect -2966 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 -2346 43634
rect -2966 7954 -2346 43398
rect -2966 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 -2346 7954
rect -2966 7634 -2346 7718
rect -2966 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 -2346 7634
rect -2966 -1306 -2346 7398
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 711590
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 1794 -7654 2414 -902
rect 6294 705798 6914 711590
rect 6294 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 6914 705798
rect 6294 705478 6914 705562
rect 6294 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 6914 705478
rect 6294 691954 6914 705242
rect 6294 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 6914 691954
rect 6294 691634 6914 691718
rect 6294 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 6914 691634
rect 6294 655954 6914 691398
rect 6294 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 6914 655954
rect 6294 655634 6914 655718
rect 6294 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 6914 655634
rect 6294 619954 6914 655398
rect 6294 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 6914 619954
rect 6294 619634 6914 619718
rect 6294 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 6914 619634
rect 6294 583954 6914 619398
rect 6294 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 6914 583954
rect 6294 583634 6914 583718
rect 6294 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 6914 583634
rect 6294 547954 6914 583398
rect 6294 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 6914 547954
rect 6294 547634 6914 547718
rect 6294 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 6914 547634
rect 6294 511954 6914 547398
rect 6294 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 6914 511954
rect 6294 511634 6914 511718
rect 6294 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 6914 511634
rect 6294 475954 6914 511398
rect 6294 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 6914 475954
rect 6294 475634 6914 475718
rect 6294 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 6914 475634
rect 6294 439954 6914 475398
rect 6294 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 6914 439954
rect 6294 439634 6914 439718
rect 6294 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 6914 439634
rect 6294 403954 6914 439398
rect 6294 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 6914 403954
rect 6294 403634 6914 403718
rect 6294 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 6914 403634
rect 6294 367954 6914 403398
rect 6294 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 6914 367954
rect 6294 367634 6914 367718
rect 6294 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 6914 367634
rect 6294 331954 6914 367398
rect 6294 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 6914 331954
rect 6294 331634 6914 331718
rect 6294 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 6914 331634
rect 6294 295954 6914 331398
rect 6294 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 6914 295954
rect 6294 295634 6914 295718
rect 6294 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 6914 295634
rect 6294 259954 6914 295398
rect 6294 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 6914 259954
rect 6294 259634 6914 259718
rect 6294 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 6914 259634
rect 6294 223954 6914 259398
rect 6294 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 6914 223954
rect 6294 223634 6914 223718
rect 6294 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 6914 223634
rect 6294 187954 6914 223398
rect 6294 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 6914 187954
rect 6294 187634 6914 187718
rect 6294 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 6914 187634
rect 6294 151954 6914 187398
rect 6294 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 6914 151954
rect 6294 151634 6914 151718
rect 6294 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 6914 151634
rect 6294 115954 6914 151398
rect 6294 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 6914 115954
rect 6294 115634 6914 115718
rect 6294 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 6914 115634
rect 6294 79954 6914 115398
rect 6294 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 6914 79954
rect 6294 79634 6914 79718
rect 6294 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 6914 79634
rect 6294 43954 6914 79398
rect 6294 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 6914 43954
rect 6294 43634 6914 43718
rect 6294 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 6914 43634
rect 6294 7954 6914 43398
rect 6294 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 6914 7954
rect 6294 7634 6914 7718
rect 6294 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 6914 7634
rect 6294 -1306 6914 7398
rect 6294 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 6914 -1306
rect 6294 -1626 6914 -1542
rect 6294 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 6914 -1626
rect 6294 -7654 6914 -1862
rect 10794 706758 11414 711590
rect 10794 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 11414 706758
rect 10794 706438 11414 706522
rect 10794 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 11414 706438
rect 10794 696454 11414 706202
rect 10794 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 11414 696454
rect 10794 696134 11414 696218
rect 10794 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 11414 696134
rect 10794 660454 11414 695898
rect 10794 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 11414 660454
rect 10794 660134 11414 660218
rect 10794 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 11414 660134
rect 10794 624454 11414 659898
rect 10794 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 11414 624454
rect 10794 624134 11414 624218
rect 10794 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 11414 624134
rect 10794 588454 11414 623898
rect 10794 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 11414 588454
rect 10794 588134 11414 588218
rect 10794 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 11414 588134
rect 10794 552454 11414 587898
rect 10794 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 11414 552454
rect 10794 552134 11414 552218
rect 10794 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 11414 552134
rect 10794 516454 11414 551898
rect 10794 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 11414 516454
rect 10794 516134 11414 516218
rect 10794 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 11414 516134
rect 10794 480454 11414 515898
rect 10794 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 11414 480454
rect 10794 480134 11414 480218
rect 10794 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 11414 480134
rect 10794 444454 11414 479898
rect 10794 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 11414 444454
rect 10794 444134 11414 444218
rect 10794 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 11414 444134
rect 10794 408454 11414 443898
rect 10794 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 11414 408454
rect 10794 408134 11414 408218
rect 10794 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 11414 408134
rect 10794 372454 11414 407898
rect 10794 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 11414 372454
rect 10794 372134 11414 372218
rect 10794 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 11414 372134
rect 10794 336454 11414 371898
rect 10794 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 11414 336454
rect 10794 336134 11414 336218
rect 10794 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 11414 336134
rect 10794 300454 11414 335898
rect 10794 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 11414 300454
rect 10794 300134 11414 300218
rect 10794 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 11414 300134
rect 10794 264454 11414 299898
rect 10794 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 11414 264454
rect 10794 264134 11414 264218
rect 10794 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 11414 264134
rect 10794 228454 11414 263898
rect 10794 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 11414 228454
rect 10794 228134 11414 228218
rect 10794 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 11414 228134
rect 10794 192454 11414 227898
rect 10794 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 11414 192454
rect 10794 192134 11414 192218
rect 10794 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 11414 192134
rect 10794 156454 11414 191898
rect 10794 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 11414 156454
rect 10794 156134 11414 156218
rect 10794 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 11414 156134
rect 10794 120454 11414 155898
rect 10794 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 11414 120454
rect 10794 120134 11414 120218
rect 10794 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 11414 120134
rect 10794 84454 11414 119898
rect 10794 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 11414 84454
rect 10794 84134 11414 84218
rect 10794 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 11414 84134
rect 10794 48454 11414 83898
rect 10794 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 11414 48454
rect 10794 48134 11414 48218
rect 10794 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 11414 48134
rect 10794 12454 11414 47898
rect 10794 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 11414 12454
rect 10794 12134 11414 12218
rect 10794 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 11414 12134
rect 10794 -2266 11414 11898
rect 10794 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 11414 -2266
rect 10794 -2586 11414 -2502
rect 10794 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 11414 -2586
rect 10794 -7654 11414 -2822
rect 15294 707718 15914 711590
rect 15294 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 15914 707718
rect 15294 707398 15914 707482
rect 15294 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 15914 707398
rect 15294 700954 15914 707162
rect 15294 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 15914 700954
rect 15294 700634 15914 700718
rect 15294 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 15914 700634
rect 15294 664954 15914 700398
rect 15294 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 15914 664954
rect 15294 664634 15914 664718
rect 15294 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 15914 664634
rect 15294 628954 15914 664398
rect 15294 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 15914 628954
rect 15294 628634 15914 628718
rect 15294 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 15914 628634
rect 15294 592954 15914 628398
rect 15294 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 15914 592954
rect 15294 592634 15914 592718
rect 15294 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 15914 592634
rect 15294 556954 15914 592398
rect 15294 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 15914 556954
rect 15294 556634 15914 556718
rect 15294 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 15914 556634
rect 15294 520954 15914 556398
rect 15294 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 15914 520954
rect 15294 520634 15914 520718
rect 15294 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 15914 520634
rect 15294 484954 15914 520398
rect 15294 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 15914 484954
rect 15294 484634 15914 484718
rect 15294 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 15914 484634
rect 15294 448954 15914 484398
rect 15294 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 15914 448954
rect 15294 448634 15914 448718
rect 15294 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 15914 448634
rect 15294 412954 15914 448398
rect 15294 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 15914 412954
rect 15294 412634 15914 412718
rect 15294 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 15914 412634
rect 15294 376954 15914 412398
rect 15294 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 15914 376954
rect 15294 376634 15914 376718
rect 15294 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 15914 376634
rect 15294 340954 15914 376398
rect 15294 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 15914 340954
rect 15294 340634 15914 340718
rect 15294 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 15914 340634
rect 15294 304954 15914 340398
rect 15294 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 15914 304954
rect 15294 304634 15914 304718
rect 15294 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 15914 304634
rect 15294 268954 15914 304398
rect 15294 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 15914 268954
rect 15294 268634 15914 268718
rect 15294 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 15914 268634
rect 15294 232954 15914 268398
rect 15294 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 15914 232954
rect 15294 232634 15914 232718
rect 15294 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 15914 232634
rect 15294 196954 15914 232398
rect 15294 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 15914 196954
rect 15294 196634 15914 196718
rect 15294 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 15914 196634
rect 15294 160954 15914 196398
rect 15294 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 15914 160954
rect 15294 160634 15914 160718
rect 15294 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 15914 160634
rect 15294 124954 15914 160398
rect 15294 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 15914 124954
rect 15294 124634 15914 124718
rect 15294 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 15914 124634
rect 15294 88954 15914 124398
rect 15294 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 15914 88954
rect 15294 88634 15914 88718
rect 15294 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 15914 88634
rect 15294 52954 15914 88398
rect 15294 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 15914 52954
rect 15294 52634 15914 52718
rect 15294 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 15914 52634
rect 15294 16954 15914 52398
rect 15294 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 15914 16954
rect 15294 16634 15914 16718
rect 15294 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 15914 16634
rect 15294 -3226 15914 16398
rect 15294 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 15914 -3226
rect 15294 -3546 15914 -3462
rect 15294 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 15914 -3546
rect 15294 -7654 15914 -3782
rect 19794 708678 20414 711590
rect 19794 708442 19826 708678
rect 20062 708442 20146 708678
rect 20382 708442 20414 708678
rect 19794 708358 20414 708442
rect 19794 708122 19826 708358
rect 20062 708122 20146 708358
rect 20382 708122 20414 708358
rect 19794 669454 20414 708122
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -4186 20414 20898
rect 19794 -4422 19826 -4186
rect 20062 -4422 20146 -4186
rect 20382 -4422 20414 -4186
rect 19794 -4506 20414 -4422
rect 19794 -4742 19826 -4506
rect 20062 -4742 20146 -4506
rect 20382 -4742 20414 -4506
rect 19794 -7654 20414 -4742
rect 24294 709638 24914 711590
rect 24294 709402 24326 709638
rect 24562 709402 24646 709638
rect 24882 709402 24914 709638
rect 24294 709318 24914 709402
rect 24294 709082 24326 709318
rect 24562 709082 24646 709318
rect 24882 709082 24914 709318
rect 24294 673954 24914 709082
rect 24294 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 24914 673954
rect 24294 673634 24914 673718
rect 24294 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 24914 673634
rect 24294 637954 24914 673398
rect 24294 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 24914 637954
rect 24294 637634 24914 637718
rect 24294 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 24914 637634
rect 24294 601954 24914 637398
rect 24294 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 24914 601954
rect 24294 601634 24914 601718
rect 24294 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 24914 601634
rect 24294 565954 24914 601398
rect 24294 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 24914 565954
rect 24294 565634 24914 565718
rect 24294 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 24914 565634
rect 24294 529954 24914 565398
rect 24294 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 24914 529954
rect 24294 529634 24914 529718
rect 24294 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 24914 529634
rect 24294 493954 24914 529398
rect 24294 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 24914 493954
rect 24294 493634 24914 493718
rect 24294 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 24914 493634
rect 24294 457954 24914 493398
rect 24294 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 24914 457954
rect 24294 457634 24914 457718
rect 24294 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 24914 457634
rect 24294 421954 24914 457398
rect 24294 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 24914 421954
rect 24294 421634 24914 421718
rect 24294 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 24914 421634
rect 24294 385954 24914 421398
rect 24294 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 24914 385954
rect 24294 385634 24914 385718
rect 24294 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 24914 385634
rect 24294 349954 24914 385398
rect 24294 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 24914 349954
rect 24294 349634 24914 349718
rect 24294 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 24914 349634
rect 24294 313954 24914 349398
rect 24294 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 24914 313954
rect 24294 313634 24914 313718
rect 24294 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 24914 313634
rect 24294 277954 24914 313398
rect 24294 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 24914 277954
rect 24294 277634 24914 277718
rect 24294 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 24914 277634
rect 24294 241954 24914 277398
rect 24294 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241718 24914 241954
rect 24294 241634 24914 241718
rect 24294 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241398 24914 241634
rect 24294 205954 24914 241398
rect 24294 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 24914 205954
rect 24294 205634 24914 205718
rect 24294 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 24914 205634
rect 24294 169954 24914 205398
rect 24294 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 24914 169954
rect 24294 169634 24914 169718
rect 24294 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 24914 169634
rect 24294 133954 24914 169398
rect 24294 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 24914 133954
rect 24294 133634 24914 133718
rect 24294 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 24914 133634
rect 24294 97954 24914 133398
rect 24294 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 24914 97954
rect 24294 97634 24914 97718
rect 24294 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 24914 97634
rect 24294 61954 24914 97398
rect 24294 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 24914 61954
rect 24294 61634 24914 61718
rect 24294 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 24914 61634
rect 24294 25954 24914 61398
rect 24294 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 24914 25954
rect 24294 25634 24914 25718
rect 24294 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 24914 25634
rect 24294 -5146 24914 25398
rect 24294 -5382 24326 -5146
rect 24562 -5382 24646 -5146
rect 24882 -5382 24914 -5146
rect 24294 -5466 24914 -5382
rect 24294 -5702 24326 -5466
rect 24562 -5702 24646 -5466
rect 24882 -5702 24914 -5466
rect 24294 -7654 24914 -5702
rect 28794 710598 29414 711590
rect 28794 710362 28826 710598
rect 29062 710362 29146 710598
rect 29382 710362 29414 710598
rect 28794 710278 29414 710362
rect 28794 710042 28826 710278
rect 29062 710042 29146 710278
rect 29382 710042 29414 710278
rect 28794 678454 29414 710042
rect 28794 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 29414 678454
rect 28794 678134 29414 678218
rect 28794 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 29414 678134
rect 28794 642454 29414 677898
rect 28794 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 29414 642454
rect 28794 642134 29414 642218
rect 28794 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 29414 642134
rect 28794 606454 29414 641898
rect 28794 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 29414 606454
rect 28794 606134 29414 606218
rect 28794 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 29414 606134
rect 28794 570454 29414 605898
rect 28794 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 29414 570454
rect 28794 570134 29414 570218
rect 28794 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 29414 570134
rect 28794 534454 29414 569898
rect 28794 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 29414 534454
rect 28794 534134 29414 534218
rect 28794 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 29414 534134
rect 28794 498454 29414 533898
rect 28794 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 29414 498454
rect 28794 498134 29414 498218
rect 28794 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 29414 498134
rect 28794 462454 29414 497898
rect 28794 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 29414 462454
rect 28794 462134 29414 462218
rect 28794 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 29414 462134
rect 28794 426454 29414 461898
rect 28794 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 29414 426454
rect 28794 426134 29414 426218
rect 28794 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 29414 426134
rect 28794 390454 29414 425898
rect 28794 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 29414 390454
rect 28794 390134 29414 390218
rect 28794 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 29414 390134
rect 28794 354454 29414 389898
rect 28794 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 29414 354454
rect 28794 354134 29414 354218
rect 28794 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 29414 354134
rect 28794 318454 29414 353898
rect 28794 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 29414 318454
rect 28794 318134 29414 318218
rect 28794 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 29414 318134
rect 28794 282454 29414 317898
rect 28794 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 29414 282454
rect 28794 282134 29414 282218
rect 28794 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 29414 282134
rect 28794 246454 29414 281898
rect 28794 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246218 29414 246454
rect 28794 246134 29414 246218
rect 28794 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 245898 29414 246134
rect 28794 210454 29414 245898
rect 28794 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 29414 210454
rect 28794 210134 29414 210218
rect 28794 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 29414 210134
rect 28794 174454 29414 209898
rect 28794 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 29414 174454
rect 28794 174134 29414 174218
rect 28794 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 29414 174134
rect 28794 138454 29414 173898
rect 28794 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 29414 138454
rect 28794 138134 29414 138218
rect 28794 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 29414 138134
rect 28794 102454 29414 137898
rect 28794 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 29414 102454
rect 28794 102134 29414 102218
rect 28794 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 29414 102134
rect 28794 66454 29414 101898
rect 28794 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 29414 66454
rect 28794 66134 29414 66218
rect 28794 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 29414 66134
rect 28794 30454 29414 65898
rect 28794 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 29414 30454
rect 28794 30134 29414 30218
rect 28794 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 29414 30134
rect 28794 -6106 29414 29898
rect 28794 -6342 28826 -6106
rect 29062 -6342 29146 -6106
rect 29382 -6342 29414 -6106
rect 28794 -6426 29414 -6342
rect 28794 -6662 28826 -6426
rect 29062 -6662 29146 -6426
rect 29382 -6662 29414 -6426
rect 28794 -7654 29414 -6662
rect 33294 711558 33914 711590
rect 33294 711322 33326 711558
rect 33562 711322 33646 711558
rect 33882 711322 33914 711558
rect 33294 711238 33914 711322
rect 33294 711002 33326 711238
rect 33562 711002 33646 711238
rect 33882 711002 33914 711238
rect 33294 682954 33914 711002
rect 33294 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 33914 682954
rect 33294 682634 33914 682718
rect 33294 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 33914 682634
rect 33294 646954 33914 682398
rect 33294 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 33914 646954
rect 33294 646634 33914 646718
rect 33294 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 33914 646634
rect 33294 610954 33914 646398
rect 33294 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 33914 610954
rect 33294 610634 33914 610718
rect 33294 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 33914 610634
rect 33294 574954 33914 610398
rect 33294 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 33914 574954
rect 33294 574634 33914 574718
rect 33294 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 33914 574634
rect 33294 538954 33914 574398
rect 33294 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 33914 538954
rect 33294 538634 33914 538718
rect 33294 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 33914 538634
rect 33294 502954 33914 538398
rect 33294 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 33914 502954
rect 33294 502634 33914 502718
rect 33294 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 33914 502634
rect 33294 466954 33914 502398
rect 33294 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 33914 466954
rect 33294 466634 33914 466718
rect 33294 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 33914 466634
rect 33294 430954 33914 466398
rect 33294 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 33914 430954
rect 33294 430634 33914 430718
rect 33294 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 33914 430634
rect 33294 394954 33914 430398
rect 33294 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 33914 394954
rect 33294 394634 33914 394718
rect 33294 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 33914 394634
rect 33294 358954 33914 394398
rect 33294 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 33914 358954
rect 33294 358634 33914 358718
rect 33294 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 33914 358634
rect 33294 322954 33914 358398
rect 33294 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 33914 322954
rect 33294 322634 33914 322718
rect 33294 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 33914 322634
rect 33294 286954 33914 322398
rect 33294 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 33914 286954
rect 33294 286634 33914 286718
rect 33294 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 33914 286634
rect 33294 250954 33914 286398
rect 33294 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 33914 250954
rect 33294 250634 33914 250718
rect 33294 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 33914 250634
rect 33294 214954 33914 250398
rect 33294 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 33914 214954
rect 33294 214634 33914 214718
rect 33294 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 33914 214634
rect 33294 178954 33914 214398
rect 33294 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 33914 178954
rect 33294 178634 33914 178718
rect 33294 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 33914 178634
rect 33294 142954 33914 178398
rect 33294 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 33914 142954
rect 33294 142634 33914 142718
rect 33294 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 33914 142634
rect 33294 106954 33914 142398
rect 33294 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 33914 106954
rect 33294 106634 33914 106718
rect 33294 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 33914 106634
rect 33294 70954 33914 106398
rect 33294 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 33914 70954
rect 33294 70634 33914 70718
rect 33294 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 33914 70634
rect 33294 34954 33914 70398
rect 33294 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 33914 34954
rect 33294 34634 33914 34718
rect 33294 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 33914 34634
rect 33294 -7066 33914 34398
rect 33294 -7302 33326 -7066
rect 33562 -7302 33646 -7066
rect 33882 -7302 33914 -7066
rect 33294 -7386 33914 -7302
rect 33294 -7622 33326 -7386
rect 33562 -7622 33646 -7386
rect 33882 -7622 33914 -7386
rect 33294 -7654 33914 -7622
rect 37794 704838 38414 711590
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -7654 38414 -902
rect 42294 705798 42914 711590
rect 42294 705562 42326 705798
rect 42562 705562 42646 705798
rect 42882 705562 42914 705798
rect 42294 705478 42914 705562
rect 42294 705242 42326 705478
rect 42562 705242 42646 705478
rect 42882 705242 42914 705478
rect 42294 691954 42914 705242
rect 42294 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 42914 691954
rect 42294 691634 42914 691718
rect 42294 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 42914 691634
rect 42294 655954 42914 691398
rect 42294 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 42914 655954
rect 42294 655634 42914 655718
rect 42294 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 42914 655634
rect 42294 619954 42914 655398
rect 42294 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 42914 619954
rect 42294 619634 42914 619718
rect 42294 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 42914 619634
rect 42294 583954 42914 619398
rect 42294 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 42914 583954
rect 42294 583634 42914 583718
rect 42294 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 42914 583634
rect 42294 547954 42914 583398
rect 42294 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 42914 547954
rect 42294 547634 42914 547718
rect 42294 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 42914 547634
rect 42294 511954 42914 547398
rect 42294 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 42914 511954
rect 42294 511634 42914 511718
rect 42294 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 42914 511634
rect 42294 475954 42914 511398
rect 42294 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 42914 475954
rect 42294 475634 42914 475718
rect 42294 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 42914 475634
rect 42294 439954 42914 475398
rect 42294 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 42914 439954
rect 42294 439634 42914 439718
rect 42294 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 42914 439634
rect 42294 403954 42914 439398
rect 42294 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 42914 403954
rect 42294 403634 42914 403718
rect 42294 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 42914 403634
rect 42294 367954 42914 403398
rect 42294 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 42914 367954
rect 42294 367634 42914 367718
rect 42294 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 42914 367634
rect 42294 331954 42914 367398
rect 42294 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 42914 331954
rect 42294 331634 42914 331718
rect 42294 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 42914 331634
rect 42294 295954 42914 331398
rect 42294 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 42914 295954
rect 42294 295634 42914 295718
rect 42294 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 42914 295634
rect 42294 259954 42914 295398
rect 42294 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 42914 259954
rect 42294 259634 42914 259718
rect 42294 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 42914 259634
rect 42294 223954 42914 259398
rect 42294 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 42914 223954
rect 42294 223634 42914 223718
rect 42294 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 42914 223634
rect 42294 187954 42914 223398
rect 42294 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 42914 187954
rect 42294 187634 42914 187718
rect 42294 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 42914 187634
rect 42294 151954 42914 187398
rect 42294 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 42914 151954
rect 42294 151634 42914 151718
rect 42294 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 42914 151634
rect 42294 115954 42914 151398
rect 42294 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 42914 115954
rect 42294 115634 42914 115718
rect 42294 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 42914 115634
rect 42294 79954 42914 115398
rect 42294 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 42914 79954
rect 42294 79634 42914 79718
rect 42294 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 42914 79634
rect 42294 43954 42914 79398
rect 42294 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 42914 43954
rect 42294 43634 42914 43718
rect 42294 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 42914 43634
rect 42294 7954 42914 43398
rect 42294 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 42914 7954
rect 42294 7634 42914 7718
rect 42294 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 42914 7634
rect 42294 -1306 42914 7398
rect 42294 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 42914 -1306
rect 42294 -1626 42914 -1542
rect 42294 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 42914 -1626
rect 42294 -7654 42914 -1862
rect 46794 706758 47414 711590
rect 46794 706522 46826 706758
rect 47062 706522 47146 706758
rect 47382 706522 47414 706758
rect 46794 706438 47414 706522
rect 46794 706202 46826 706438
rect 47062 706202 47146 706438
rect 47382 706202 47414 706438
rect 46794 696454 47414 706202
rect 46794 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 47414 696454
rect 46794 696134 47414 696218
rect 46794 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 47414 696134
rect 46794 660454 47414 695898
rect 46794 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 47414 660454
rect 46794 660134 47414 660218
rect 46794 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 47414 660134
rect 46794 624454 47414 659898
rect 46794 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 47414 624454
rect 46794 624134 47414 624218
rect 46794 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 47414 624134
rect 46794 588454 47414 623898
rect 46794 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 47414 588454
rect 46794 588134 47414 588218
rect 46794 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 47414 588134
rect 46794 552454 47414 587898
rect 46794 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 47414 552454
rect 46794 552134 47414 552218
rect 46794 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 47414 552134
rect 46794 516454 47414 551898
rect 46794 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 47414 516454
rect 46794 516134 47414 516218
rect 46794 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 47414 516134
rect 46794 480454 47414 515898
rect 46794 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 47414 480454
rect 46794 480134 47414 480218
rect 46794 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 47414 480134
rect 46794 444454 47414 479898
rect 46794 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 47414 444454
rect 46794 444134 47414 444218
rect 46794 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 47414 444134
rect 46794 408454 47414 443898
rect 46794 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 47414 408454
rect 46794 408134 47414 408218
rect 46794 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 47414 408134
rect 46794 372454 47414 407898
rect 46794 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 47414 372454
rect 46794 372134 47414 372218
rect 46794 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 47414 372134
rect 46794 336454 47414 371898
rect 46794 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 47414 336454
rect 46794 336134 47414 336218
rect 46794 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 47414 336134
rect 46794 300454 47414 335898
rect 46794 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 47414 300454
rect 46794 300134 47414 300218
rect 46794 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 47414 300134
rect 46794 264454 47414 299898
rect 46794 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 47414 264454
rect 46794 264134 47414 264218
rect 46794 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 47414 264134
rect 46794 228454 47414 263898
rect 46794 228218 46826 228454
rect 47062 228218 47146 228454
rect 47382 228218 47414 228454
rect 46794 228134 47414 228218
rect 46794 227898 46826 228134
rect 47062 227898 47146 228134
rect 47382 227898 47414 228134
rect 46794 192454 47414 227898
rect 46794 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 47414 192454
rect 46794 192134 47414 192218
rect 46794 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 47414 192134
rect 46794 156454 47414 191898
rect 46794 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 47414 156454
rect 46794 156134 47414 156218
rect 46794 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 47414 156134
rect 46794 120454 47414 155898
rect 46794 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 47414 120454
rect 46794 120134 47414 120218
rect 46794 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 47414 120134
rect 46794 84454 47414 119898
rect 46794 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 47414 84454
rect 46794 84134 47414 84218
rect 46794 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 47414 84134
rect 46794 48454 47414 83898
rect 46794 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 47414 48454
rect 46794 48134 47414 48218
rect 46794 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 47414 48134
rect 46794 12454 47414 47898
rect 46794 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 47414 12454
rect 46794 12134 47414 12218
rect 46794 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 47414 12134
rect 46794 -2266 47414 11898
rect 46794 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 47414 -2266
rect 46794 -2586 47414 -2502
rect 46794 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 47414 -2586
rect 46794 -7654 47414 -2822
rect 51294 707718 51914 711590
rect 51294 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 51914 707718
rect 51294 707398 51914 707482
rect 51294 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 51914 707398
rect 51294 700954 51914 707162
rect 51294 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 51914 700954
rect 51294 700634 51914 700718
rect 51294 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 51914 700634
rect 51294 664954 51914 700398
rect 51294 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 51914 664954
rect 51294 664634 51914 664718
rect 51294 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 51914 664634
rect 51294 628954 51914 664398
rect 51294 628718 51326 628954
rect 51562 628718 51646 628954
rect 51882 628718 51914 628954
rect 51294 628634 51914 628718
rect 51294 628398 51326 628634
rect 51562 628398 51646 628634
rect 51882 628398 51914 628634
rect 51294 592954 51914 628398
rect 51294 592718 51326 592954
rect 51562 592718 51646 592954
rect 51882 592718 51914 592954
rect 51294 592634 51914 592718
rect 51294 592398 51326 592634
rect 51562 592398 51646 592634
rect 51882 592398 51914 592634
rect 51294 556954 51914 592398
rect 51294 556718 51326 556954
rect 51562 556718 51646 556954
rect 51882 556718 51914 556954
rect 51294 556634 51914 556718
rect 51294 556398 51326 556634
rect 51562 556398 51646 556634
rect 51882 556398 51914 556634
rect 51294 520954 51914 556398
rect 51294 520718 51326 520954
rect 51562 520718 51646 520954
rect 51882 520718 51914 520954
rect 51294 520634 51914 520718
rect 51294 520398 51326 520634
rect 51562 520398 51646 520634
rect 51882 520398 51914 520634
rect 51294 484954 51914 520398
rect 51294 484718 51326 484954
rect 51562 484718 51646 484954
rect 51882 484718 51914 484954
rect 51294 484634 51914 484718
rect 51294 484398 51326 484634
rect 51562 484398 51646 484634
rect 51882 484398 51914 484634
rect 51294 448954 51914 484398
rect 51294 448718 51326 448954
rect 51562 448718 51646 448954
rect 51882 448718 51914 448954
rect 51294 448634 51914 448718
rect 51294 448398 51326 448634
rect 51562 448398 51646 448634
rect 51882 448398 51914 448634
rect 51294 412954 51914 448398
rect 51294 412718 51326 412954
rect 51562 412718 51646 412954
rect 51882 412718 51914 412954
rect 51294 412634 51914 412718
rect 51294 412398 51326 412634
rect 51562 412398 51646 412634
rect 51882 412398 51914 412634
rect 51294 376954 51914 412398
rect 51294 376718 51326 376954
rect 51562 376718 51646 376954
rect 51882 376718 51914 376954
rect 51294 376634 51914 376718
rect 51294 376398 51326 376634
rect 51562 376398 51646 376634
rect 51882 376398 51914 376634
rect 51294 340954 51914 376398
rect 51294 340718 51326 340954
rect 51562 340718 51646 340954
rect 51882 340718 51914 340954
rect 51294 340634 51914 340718
rect 51294 340398 51326 340634
rect 51562 340398 51646 340634
rect 51882 340398 51914 340634
rect 51294 304954 51914 340398
rect 51294 304718 51326 304954
rect 51562 304718 51646 304954
rect 51882 304718 51914 304954
rect 51294 304634 51914 304718
rect 51294 304398 51326 304634
rect 51562 304398 51646 304634
rect 51882 304398 51914 304634
rect 51294 268954 51914 304398
rect 51294 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 51914 268954
rect 51294 268634 51914 268718
rect 51294 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 51914 268634
rect 51294 232954 51914 268398
rect 51294 232718 51326 232954
rect 51562 232718 51646 232954
rect 51882 232718 51914 232954
rect 51294 232634 51914 232718
rect 51294 232398 51326 232634
rect 51562 232398 51646 232634
rect 51882 232398 51914 232634
rect 51294 196954 51914 232398
rect 51294 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 51914 196954
rect 51294 196634 51914 196718
rect 51294 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 51914 196634
rect 51294 160954 51914 196398
rect 51294 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 51914 160954
rect 51294 160634 51914 160718
rect 51294 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 51914 160634
rect 51294 124954 51914 160398
rect 51294 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 51914 124954
rect 51294 124634 51914 124718
rect 51294 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 51914 124634
rect 51294 88954 51914 124398
rect 51294 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 51914 88954
rect 51294 88634 51914 88718
rect 51294 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 51914 88634
rect 51294 52954 51914 88398
rect 51294 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 51914 52954
rect 51294 52634 51914 52718
rect 51294 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 51914 52634
rect 51294 16954 51914 52398
rect 51294 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 51914 16954
rect 51294 16634 51914 16718
rect 51294 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 51914 16634
rect 51294 -3226 51914 16398
rect 51294 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 51914 -3226
rect 51294 -3546 51914 -3462
rect 51294 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 51914 -3546
rect 51294 -7654 51914 -3782
rect 55794 708678 56414 711590
rect 55794 708442 55826 708678
rect 56062 708442 56146 708678
rect 56382 708442 56414 708678
rect 55794 708358 56414 708442
rect 55794 708122 55826 708358
rect 56062 708122 56146 708358
rect 56382 708122 56414 708358
rect 55794 669454 56414 708122
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -4186 56414 20898
rect 55794 -4422 55826 -4186
rect 56062 -4422 56146 -4186
rect 56382 -4422 56414 -4186
rect 55794 -4506 56414 -4422
rect 55794 -4742 55826 -4506
rect 56062 -4742 56146 -4506
rect 56382 -4742 56414 -4506
rect 55794 -7654 56414 -4742
rect 60294 709638 60914 711590
rect 60294 709402 60326 709638
rect 60562 709402 60646 709638
rect 60882 709402 60914 709638
rect 60294 709318 60914 709402
rect 60294 709082 60326 709318
rect 60562 709082 60646 709318
rect 60882 709082 60914 709318
rect 60294 673954 60914 709082
rect 60294 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 60914 673954
rect 60294 673634 60914 673718
rect 60294 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 60914 673634
rect 60294 637954 60914 673398
rect 60294 637718 60326 637954
rect 60562 637718 60646 637954
rect 60882 637718 60914 637954
rect 60294 637634 60914 637718
rect 60294 637398 60326 637634
rect 60562 637398 60646 637634
rect 60882 637398 60914 637634
rect 60294 601954 60914 637398
rect 60294 601718 60326 601954
rect 60562 601718 60646 601954
rect 60882 601718 60914 601954
rect 60294 601634 60914 601718
rect 60294 601398 60326 601634
rect 60562 601398 60646 601634
rect 60882 601398 60914 601634
rect 60294 565954 60914 601398
rect 60294 565718 60326 565954
rect 60562 565718 60646 565954
rect 60882 565718 60914 565954
rect 60294 565634 60914 565718
rect 60294 565398 60326 565634
rect 60562 565398 60646 565634
rect 60882 565398 60914 565634
rect 60294 529954 60914 565398
rect 60294 529718 60326 529954
rect 60562 529718 60646 529954
rect 60882 529718 60914 529954
rect 60294 529634 60914 529718
rect 60294 529398 60326 529634
rect 60562 529398 60646 529634
rect 60882 529398 60914 529634
rect 60294 493954 60914 529398
rect 60294 493718 60326 493954
rect 60562 493718 60646 493954
rect 60882 493718 60914 493954
rect 60294 493634 60914 493718
rect 60294 493398 60326 493634
rect 60562 493398 60646 493634
rect 60882 493398 60914 493634
rect 60294 457954 60914 493398
rect 60294 457718 60326 457954
rect 60562 457718 60646 457954
rect 60882 457718 60914 457954
rect 60294 457634 60914 457718
rect 60294 457398 60326 457634
rect 60562 457398 60646 457634
rect 60882 457398 60914 457634
rect 60294 421954 60914 457398
rect 60294 421718 60326 421954
rect 60562 421718 60646 421954
rect 60882 421718 60914 421954
rect 60294 421634 60914 421718
rect 60294 421398 60326 421634
rect 60562 421398 60646 421634
rect 60882 421398 60914 421634
rect 60294 385954 60914 421398
rect 60294 385718 60326 385954
rect 60562 385718 60646 385954
rect 60882 385718 60914 385954
rect 60294 385634 60914 385718
rect 60294 385398 60326 385634
rect 60562 385398 60646 385634
rect 60882 385398 60914 385634
rect 60294 349954 60914 385398
rect 60294 349718 60326 349954
rect 60562 349718 60646 349954
rect 60882 349718 60914 349954
rect 60294 349634 60914 349718
rect 60294 349398 60326 349634
rect 60562 349398 60646 349634
rect 60882 349398 60914 349634
rect 60294 313954 60914 349398
rect 60294 313718 60326 313954
rect 60562 313718 60646 313954
rect 60882 313718 60914 313954
rect 60294 313634 60914 313718
rect 60294 313398 60326 313634
rect 60562 313398 60646 313634
rect 60882 313398 60914 313634
rect 60294 277954 60914 313398
rect 60294 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 60914 277954
rect 60294 277634 60914 277718
rect 60294 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 60914 277634
rect 60294 241954 60914 277398
rect 60294 241718 60326 241954
rect 60562 241718 60646 241954
rect 60882 241718 60914 241954
rect 60294 241634 60914 241718
rect 60294 241398 60326 241634
rect 60562 241398 60646 241634
rect 60882 241398 60914 241634
rect 60294 205954 60914 241398
rect 60294 205718 60326 205954
rect 60562 205718 60646 205954
rect 60882 205718 60914 205954
rect 60294 205634 60914 205718
rect 60294 205398 60326 205634
rect 60562 205398 60646 205634
rect 60882 205398 60914 205634
rect 60294 169954 60914 205398
rect 60294 169718 60326 169954
rect 60562 169718 60646 169954
rect 60882 169718 60914 169954
rect 60294 169634 60914 169718
rect 60294 169398 60326 169634
rect 60562 169398 60646 169634
rect 60882 169398 60914 169634
rect 60294 133954 60914 169398
rect 60294 133718 60326 133954
rect 60562 133718 60646 133954
rect 60882 133718 60914 133954
rect 60294 133634 60914 133718
rect 60294 133398 60326 133634
rect 60562 133398 60646 133634
rect 60882 133398 60914 133634
rect 60294 97954 60914 133398
rect 60294 97718 60326 97954
rect 60562 97718 60646 97954
rect 60882 97718 60914 97954
rect 60294 97634 60914 97718
rect 60294 97398 60326 97634
rect 60562 97398 60646 97634
rect 60882 97398 60914 97634
rect 60294 61954 60914 97398
rect 60294 61718 60326 61954
rect 60562 61718 60646 61954
rect 60882 61718 60914 61954
rect 60294 61634 60914 61718
rect 60294 61398 60326 61634
rect 60562 61398 60646 61634
rect 60882 61398 60914 61634
rect 60294 25954 60914 61398
rect 60294 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 60914 25954
rect 60294 25634 60914 25718
rect 60294 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 60914 25634
rect 60294 -5146 60914 25398
rect 60294 -5382 60326 -5146
rect 60562 -5382 60646 -5146
rect 60882 -5382 60914 -5146
rect 60294 -5466 60914 -5382
rect 60294 -5702 60326 -5466
rect 60562 -5702 60646 -5466
rect 60882 -5702 60914 -5466
rect 60294 -7654 60914 -5702
rect 64794 710598 65414 711590
rect 64794 710362 64826 710598
rect 65062 710362 65146 710598
rect 65382 710362 65414 710598
rect 64794 710278 65414 710362
rect 64794 710042 64826 710278
rect 65062 710042 65146 710278
rect 65382 710042 65414 710278
rect 64794 678454 65414 710042
rect 64794 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 65414 678454
rect 64794 678134 65414 678218
rect 64794 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 65414 678134
rect 64794 642454 65414 677898
rect 64794 642218 64826 642454
rect 65062 642218 65146 642454
rect 65382 642218 65414 642454
rect 64794 642134 65414 642218
rect 64794 641898 64826 642134
rect 65062 641898 65146 642134
rect 65382 641898 65414 642134
rect 64794 606454 65414 641898
rect 64794 606218 64826 606454
rect 65062 606218 65146 606454
rect 65382 606218 65414 606454
rect 64794 606134 65414 606218
rect 64794 605898 64826 606134
rect 65062 605898 65146 606134
rect 65382 605898 65414 606134
rect 64794 570454 65414 605898
rect 64794 570218 64826 570454
rect 65062 570218 65146 570454
rect 65382 570218 65414 570454
rect 64794 570134 65414 570218
rect 64794 569898 64826 570134
rect 65062 569898 65146 570134
rect 65382 569898 65414 570134
rect 64794 534454 65414 569898
rect 64794 534218 64826 534454
rect 65062 534218 65146 534454
rect 65382 534218 65414 534454
rect 64794 534134 65414 534218
rect 64794 533898 64826 534134
rect 65062 533898 65146 534134
rect 65382 533898 65414 534134
rect 64794 498454 65414 533898
rect 64794 498218 64826 498454
rect 65062 498218 65146 498454
rect 65382 498218 65414 498454
rect 64794 498134 65414 498218
rect 64794 497898 64826 498134
rect 65062 497898 65146 498134
rect 65382 497898 65414 498134
rect 64794 462454 65414 497898
rect 64794 462218 64826 462454
rect 65062 462218 65146 462454
rect 65382 462218 65414 462454
rect 64794 462134 65414 462218
rect 64794 461898 64826 462134
rect 65062 461898 65146 462134
rect 65382 461898 65414 462134
rect 64794 426454 65414 461898
rect 64794 426218 64826 426454
rect 65062 426218 65146 426454
rect 65382 426218 65414 426454
rect 64794 426134 65414 426218
rect 64794 425898 64826 426134
rect 65062 425898 65146 426134
rect 65382 425898 65414 426134
rect 64794 390454 65414 425898
rect 64794 390218 64826 390454
rect 65062 390218 65146 390454
rect 65382 390218 65414 390454
rect 64794 390134 65414 390218
rect 64794 389898 64826 390134
rect 65062 389898 65146 390134
rect 65382 389898 65414 390134
rect 64794 354454 65414 389898
rect 64794 354218 64826 354454
rect 65062 354218 65146 354454
rect 65382 354218 65414 354454
rect 64794 354134 65414 354218
rect 64794 353898 64826 354134
rect 65062 353898 65146 354134
rect 65382 353898 65414 354134
rect 64794 318454 65414 353898
rect 64794 318218 64826 318454
rect 65062 318218 65146 318454
rect 65382 318218 65414 318454
rect 64794 318134 65414 318218
rect 64794 317898 64826 318134
rect 65062 317898 65146 318134
rect 65382 317898 65414 318134
rect 64794 282454 65414 317898
rect 64794 282218 64826 282454
rect 65062 282218 65146 282454
rect 65382 282218 65414 282454
rect 64794 282134 65414 282218
rect 64794 281898 64826 282134
rect 65062 281898 65146 282134
rect 65382 281898 65414 282134
rect 64794 246454 65414 281898
rect 64794 246218 64826 246454
rect 65062 246218 65146 246454
rect 65382 246218 65414 246454
rect 64794 246134 65414 246218
rect 64794 245898 64826 246134
rect 65062 245898 65146 246134
rect 65382 245898 65414 246134
rect 64794 210454 65414 245898
rect 64794 210218 64826 210454
rect 65062 210218 65146 210454
rect 65382 210218 65414 210454
rect 64794 210134 65414 210218
rect 64794 209898 64826 210134
rect 65062 209898 65146 210134
rect 65382 209898 65414 210134
rect 64794 174454 65414 209898
rect 64794 174218 64826 174454
rect 65062 174218 65146 174454
rect 65382 174218 65414 174454
rect 64794 174134 65414 174218
rect 64794 173898 64826 174134
rect 65062 173898 65146 174134
rect 65382 173898 65414 174134
rect 64794 138454 65414 173898
rect 64794 138218 64826 138454
rect 65062 138218 65146 138454
rect 65382 138218 65414 138454
rect 64794 138134 65414 138218
rect 64794 137898 64826 138134
rect 65062 137898 65146 138134
rect 65382 137898 65414 138134
rect 64794 102454 65414 137898
rect 64794 102218 64826 102454
rect 65062 102218 65146 102454
rect 65382 102218 65414 102454
rect 64794 102134 65414 102218
rect 64794 101898 64826 102134
rect 65062 101898 65146 102134
rect 65382 101898 65414 102134
rect 64794 66454 65414 101898
rect 64794 66218 64826 66454
rect 65062 66218 65146 66454
rect 65382 66218 65414 66454
rect 64794 66134 65414 66218
rect 64794 65898 64826 66134
rect 65062 65898 65146 66134
rect 65382 65898 65414 66134
rect 64794 30454 65414 65898
rect 64794 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 65414 30454
rect 64794 30134 65414 30218
rect 64794 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 65414 30134
rect 64794 -6106 65414 29898
rect 64794 -6342 64826 -6106
rect 65062 -6342 65146 -6106
rect 65382 -6342 65414 -6106
rect 64794 -6426 65414 -6342
rect 64794 -6662 64826 -6426
rect 65062 -6662 65146 -6426
rect 65382 -6662 65414 -6426
rect 64794 -7654 65414 -6662
rect 69294 711558 69914 711590
rect 69294 711322 69326 711558
rect 69562 711322 69646 711558
rect 69882 711322 69914 711558
rect 69294 711238 69914 711322
rect 69294 711002 69326 711238
rect 69562 711002 69646 711238
rect 69882 711002 69914 711238
rect 69294 682954 69914 711002
rect 69294 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 69914 682954
rect 69294 682634 69914 682718
rect 69294 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 69914 682634
rect 69294 646954 69914 682398
rect 69294 646718 69326 646954
rect 69562 646718 69646 646954
rect 69882 646718 69914 646954
rect 69294 646634 69914 646718
rect 69294 646398 69326 646634
rect 69562 646398 69646 646634
rect 69882 646398 69914 646634
rect 69294 610954 69914 646398
rect 69294 610718 69326 610954
rect 69562 610718 69646 610954
rect 69882 610718 69914 610954
rect 69294 610634 69914 610718
rect 69294 610398 69326 610634
rect 69562 610398 69646 610634
rect 69882 610398 69914 610634
rect 69294 574954 69914 610398
rect 69294 574718 69326 574954
rect 69562 574718 69646 574954
rect 69882 574718 69914 574954
rect 69294 574634 69914 574718
rect 69294 574398 69326 574634
rect 69562 574398 69646 574634
rect 69882 574398 69914 574634
rect 69294 538954 69914 574398
rect 69294 538718 69326 538954
rect 69562 538718 69646 538954
rect 69882 538718 69914 538954
rect 69294 538634 69914 538718
rect 69294 538398 69326 538634
rect 69562 538398 69646 538634
rect 69882 538398 69914 538634
rect 69294 502954 69914 538398
rect 69294 502718 69326 502954
rect 69562 502718 69646 502954
rect 69882 502718 69914 502954
rect 69294 502634 69914 502718
rect 69294 502398 69326 502634
rect 69562 502398 69646 502634
rect 69882 502398 69914 502634
rect 69294 466954 69914 502398
rect 69294 466718 69326 466954
rect 69562 466718 69646 466954
rect 69882 466718 69914 466954
rect 69294 466634 69914 466718
rect 69294 466398 69326 466634
rect 69562 466398 69646 466634
rect 69882 466398 69914 466634
rect 69294 430954 69914 466398
rect 69294 430718 69326 430954
rect 69562 430718 69646 430954
rect 69882 430718 69914 430954
rect 69294 430634 69914 430718
rect 69294 430398 69326 430634
rect 69562 430398 69646 430634
rect 69882 430398 69914 430634
rect 69294 394954 69914 430398
rect 69294 394718 69326 394954
rect 69562 394718 69646 394954
rect 69882 394718 69914 394954
rect 69294 394634 69914 394718
rect 69294 394398 69326 394634
rect 69562 394398 69646 394634
rect 69882 394398 69914 394634
rect 69294 358954 69914 394398
rect 69294 358718 69326 358954
rect 69562 358718 69646 358954
rect 69882 358718 69914 358954
rect 69294 358634 69914 358718
rect 69294 358398 69326 358634
rect 69562 358398 69646 358634
rect 69882 358398 69914 358634
rect 69294 322954 69914 358398
rect 69294 322718 69326 322954
rect 69562 322718 69646 322954
rect 69882 322718 69914 322954
rect 69294 322634 69914 322718
rect 69294 322398 69326 322634
rect 69562 322398 69646 322634
rect 69882 322398 69914 322634
rect 69294 286954 69914 322398
rect 69294 286718 69326 286954
rect 69562 286718 69646 286954
rect 69882 286718 69914 286954
rect 69294 286634 69914 286718
rect 69294 286398 69326 286634
rect 69562 286398 69646 286634
rect 69882 286398 69914 286634
rect 69294 250954 69914 286398
rect 69294 250718 69326 250954
rect 69562 250718 69646 250954
rect 69882 250718 69914 250954
rect 69294 250634 69914 250718
rect 69294 250398 69326 250634
rect 69562 250398 69646 250634
rect 69882 250398 69914 250634
rect 69294 214954 69914 250398
rect 69294 214718 69326 214954
rect 69562 214718 69646 214954
rect 69882 214718 69914 214954
rect 69294 214634 69914 214718
rect 69294 214398 69326 214634
rect 69562 214398 69646 214634
rect 69882 214398 69914 214634
rect 69294 178954 69914 214398
rect 69294 178718 69326 178954
rect 69562 178718 69646 178954
rect 69882 178718 69914 178954
rect 69294 178634 69914 178718
rect 69294 178398 69326 178634
rect 69562 178398 69646 178634
rect 69882 178398 69914 178634
rect 69294 142954 69914 178398
rect 69294 142718 69326 142954
rect 69562 142718 69646 142954
rect 69882 142718 69914 142954
rect 69294 142634 69914 142718
rect 69294 142398 69326 142634
rect 69562 142398 69646 142634
rect 69882 142398 69914 142634
rect 69294 106954 69914 142398
rect 69294 106718 69326 106954
rect 69562 106718 69646 106954
rect 69882 106718 69914 106954
rect 69294 106634 69914 106718
rect 69294 106398 69326 106634
rect 69562 106398 69646 106634
rect 69882 106398 69914 106634
rect 69294 70954 69914 106398
rect 69294 70718 69326 70954
rect 69562 70718 69646 70954
rect 69882 70718 69914 70954
rect 69294 70634 69914 70718
rect 69294 70398 69326 70634
rect 69562 70398 69646 70634
rect 69882 70398 69914 70634
rect 69294 34954 69914 70398
rect 69294 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 69914 34954
rect 69294 34634 69914 34718
rect 69294 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 69914 34634
rect 69294 -7066 69914 34398
rect 69294 -7302 69326 -7066
rect 69562 -7302 69646 -7066
rect 69882 -7302 69914 -7066
rect 69294 -7386 69914 -7302
rect 69294 -7622 69326 -7386
rect 69562 -7622 69646 -7386
rect 69882 -7622 69914 -7386
rect 69294 -7654 69914 -7622
rect 73794 704838 74414 711590
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 579454 74414 614898
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 73794 543454 74414 578898
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 73794 507454 74414 542898
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 435454 74414 470898
rect 73794 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 74414 435454
rect 73794 435134 74414 435218
rect 73794 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 74414 435134
rect 73794 399454 74414 434898
rect 73794 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 74414 399454
rect 73794 399134 74414 399218
rect 73794 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 74414 399134
rect 73794 363454 74414 398898
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 327454 74414 362898
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 73794 291454 74414 326898
rect 73794 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 74414 291454
rect 73794 291134 74414 291218
rect 73794 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 74414 291134
rect 73794 255454 74414 290898
rect 73794 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 74414 255454
rect 73794 255134 74414 255218
rect 73794 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 74414 255134
rect 73794 219454 74414 254898
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 73794 183454 74414 218898
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 147454 74414 182898
rect 73794 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 74414 147454
rect 73794 147134 74414 147218
rect 73794 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 74414 147134
rect 73794 111454 74414 146898
rect 73794 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 74414 111454
rect 73794 111134 74414 111218
rect 73794 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 74414 111134
rect 73794 75454 74414 110898
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -7654 74414 -902
rect 78294 705798 78914 711590
rect 78294 705562 78326 705798
rect 78562 705562 78646 705798
rect 78882 705562 78914 705798
rect 78294 705478 78914 705562
rect 78294 705242 78326 705478
rect 78562 705242 78646 705478
rect 78882 705242 78914 705478
rect 78294 691954 78914 705242
rect 78294 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 78914 691954
rect 78294 691634 78914 691718
rect 78294 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 78914 691634
rect 78294 655954 78914 691398
rect 78294 655718 78326 655954
rect 78562 655718 78646 655954
rect 78882 655718 78914 655954
rect 78294 655634 78914 655718
rect 78294 655398 78326 655634
rect 78562 655398 78646 655634
rect 78882 655398 78914 655634
rect 78294 619954 78914 655398
rect 78294 619718 78326 619954
rect 78562 619718 78646 619954
rect 78882 619718 78914 619954
rect 78294 619634 78914 619718
rect 78294 619398 78326 619634
rect 78562 619398 78646 619634
rect 78882 619398 78914 619634
rect 78294 583954 78914 619398
rect 78294 583718 78326 583954
rect 78562 583718 78646 583954
rect 78882 583718 78914 583954
rect 78294 583634 78914 583718
rect 78294 583398 78326 583634
rect 78562 583398 78646 583634
rect 78882 583398 78914 583634
rect 78294 547954 78914 583398
rect 78294 547718 78326 547954
rect 78562 547718 78646 547954
rect 78882 547718 78914 547954
rect 78294 547634 78914 547718
rect 78294 547398 78326 547634
rect 78562 547398 78646 547634
rect 78882 547398 78914 547634
rect 78294 511954 78914 547398
rect 78294 511718 78326 511954
rect 78562 511718 78646 511954
rect 78882 511718 78914 511954
rect 78294 511634 78914 511718
rect 78294 511398 78326 511634
rect 78562 511398 78646 511634
rect 78882 511398 78914 511634
rect 78294 475954 78914 511398
rect 78294 475718 78326 475954
rect 78562 475718 78646 475954
rect 78882 475718 78914 475954
rect 78294 475634 78914 475718
rect 78294 475398 78326 475634
rect 78562 475398 78646 475634
rect 78882 475398 78914 475634
rect 78294 439954 78914 475398
rect 78294 439718 78326 439954
rect 78562 439718 78646 439954
rect 78882 439718 78914 439954
rect 78294 439634 78914 439718
rect 78294 439398 78326 439634
rect 78562 439398 78646 439634
rect 78882 439398 78914 439634
rect 78294 403954 78914 439398
rect 78294 403718 78326 403954
rect 78562 403718 78646 403954
rect 78882 403718 78914 403954
rect 78294 403634 78914 403718
rect 78294 403398 78326 403634
rect 78562 403398 78646 403634
rect 78882 403398 78914 403634
rect 78294 367954 78914 403398
rect 78294 367718 78326 367954
rect 78562 367718 78646 367954
rect 78882 367718 78914 367954
rect 78294 367634 78914 367718
rect 78294 367398 78326 367634
rect 78562 367398 78646 367634
rect 78882 367398 78914 367634
rect 78294 331954 78914 367398
rect 78294 331718 78326 331954
rect 78562 331718 78646 331954
rect 78882 331718 78914 331954
rect 78294 331634 78914 331718
rect 78294 331398 78326 331634
rect 78562 331398 78646 331634
rect 78882 331398 78914 331634
rect 78294 295954 78914 331398
rect 78294 295718 78326 295954
rect 78562 295718 78646 295954
rect 78882 295718 78914 295954
rect 78294 295634 78914 295718
rect 78294 295398 78326 295634
rect 78562 295398 78646 295634
rect 78882 295398 78914 295634
rect 78294 259954 78914 295398
rect 78294 259718 78326 259954
rect 78562 259718 78646 259954
rect 78882 259718 78914 259954
rect 78294 259634 78914 259718
rect 78294 259398 78326 259634
rect 78562 259398 78646 259634
rect 78882 259398 78914 259634
rect 78294 223954 78914 259398
rect 78294 223718 78326 223954
rect 78562 223718 78646 223954
rect 78882 223718 78914 223954
rect 78294 223634 78914 223718
rect 78294 223398 78326 223634
rect 78562 223398 78646 223634
rect 78882 223398 78914 223634
rect 78294 187954 78914 223398
rect 78294 187718 78326 187954
rect 78562 187718 78646 187954
rect 78882 187718 78914 187954
rect 78294 187634 78914 187718
rect 78294 187398 78326 187634
rect 78562 187398 78646 187634
rect 78882 187398 78914 187634
rect 78294 151954 78914 187398
rect 78294 151718 78326 151954
rect 78562 151718 78646 151954
rect 78882 151718 78914 151954
rect 78294 151634 78914 151718
rect 78294 151398 78326 151634
rect 78562 151398 78646 151634
rect 78882 151398 78914 151634
rect 78294 115954 78914 151398
rect 78294 115718 78326 115954
rect 78562 115718 78646 115954
rect 78882 115718 78914 115954
rect 78294 115634 78914 115718
rect 78294 115398 78326 115634
rect 78562 115398 78646 115634
rect 78882 115398 78914 115634
rect 78294 79954 78914 115398
rect 78294 79718 78326 79954
rect 78562 79718 78646 79954
rect 78882 79718 78914 79954
rect 78294 79634 78914 79718
rect 78294 79398 78326 79634
rect 78562 79398 78646 79634
rect 78882 79398 78914 79634
rect 78294 43954 78914 79398
rect 78294 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 78914 43954
rect 78294 43634 78914 43718
rect 78294 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 78914 43634
rect 78294 7954 78914 43398
rect 78294 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 78914 7954
rect 78294 7634 78914 7718
rect 78294 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 78914 7634
rect 78294 -1306 78914 7398
rect 78294 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 78914 -1306
rect 78294 -1626 78914 -1542
rect 78294 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 78914 -1626
rect 78294 -7654 78914 -1862
rect 82794 706758 83414 711590
rect 82794 706522 82826 706758
rect 83062 706522 83146 706758
rect 83382 706522 83414 706758
rect 82794 706438 83414 706522
rect 82794 706202 82826 706438
rect 83062 706202 83146 706438
rect 83382 706202 83414 706438
rect 82794 696454 83414 706202
rect 82794 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 83414 696454
rect 82794 696134 83414 696218
rect 82794 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 83414 696134
rect 82794 660454 83414 695898
rect 82794 660218 82826 660454
rect 83062 660218 83146 660454
rect 83382 660218 83414 660454
rect 82794 660134 83414 660218
rect 82794 659898 82826 660134
rect 83062 659898 83146 660134
rect 83382 659898 83414 660134
rect 82794 624454 83414 659898
rect 82794 624218 82826 624454
rect 83062 624218 83146 624454
rect 83382 624218 83414 624454
rect 82794 624134 83414 624218
rect 82794 623898 82826 624134
rect 83062 623898 83146 624134
rect 83382 623898 83414 624134
rect 82794 588454 83414 623898
rect 82794 588218 82826 588454
rect 83062 588218 83146 588454
rect 83382 588218 83414 588454
rect 82794 588134 83414 588218
rect 82794 587898 82826 588134
rect 83062 587898 83146 588134
rect 83382 587898 83414 588134
rect 82794 552454 83414 587898
rect 82794 552218 82826 552454
rect 83062 552218 83146 552454
rect 83382 552218 83414 552454
rect 82794 552134 83414 552218
rect 82794 551898 82826 552134
rect 83062 551898 83146 552134
rect 83382 551898 83414 552134
rect 82794 516454 83414 551898
rect 82794 516218 82826 516454
rect 83062 516218 83146 516454
rect 83382 516218 83414 516454
rect 82794 516134 83414 516218
rect 82794 515898 82826 516134
rect 83062 515898 83146 516134
rect 83382 515898 83414 516134
rect 82794 480454 83414 515898
rect 82794 480218 82826 480454
rect 83062 480218 83146 480454
rect 83382 480218 83414 480454
rect 82794 480134 83414 480218
rect 82794 479898 82826 480134
rect 83062 479898 83146 480134
rect 83382 479898 83414 480134
rect 82794 444454 83414 479898
rect 82794 444218 82826 444454
rect 83062 444218 83146 444454
rect 83382 444218 83414 444454
rect 82794 444134 83414 444218
rect 82794 443898 82826 444134
rect 83062 443898 83146 444134
rect 83382 443898 83414 444134
rect 82794 408454 83414 443898
rect 82794 408218 82826 408454
rect 83062 408218 83146 408454
rect 83382 408218 83414 408454
rect 82794 408134 83414 408218
rect 82794 407898 82826 408134
rect 83062 407898 83146 408134
rect 83382 407898 83414 408134
rect 82794 372454 83414 407898
rect 82794 372218 82826 372454
rect 83062 372218 83146 372454
rect 83382 372218 83414 372454
rect 82794 372134 83414 372218
rect 82794 371898 82826 372134
rect 83062 371898 83146 372134
rect 83382 371898 83414 372134
rect 82794 336454 83414 371898
rect 82794 336218 82826 336454
rect 83062 336218 83146 336454
rect 83382 336218 83414 336454
rect 82794 336134 83414 336218
rect 82794 335898 82826 336134
rect 83062 335898 83146 336134
rect 83382 335898 83414 336134
rect 82794 300454 83414 335898
rect 82794 300218 82826 300454
rect 83062 300218 83146 300454
rect 83382 300218 83414 300454
rect 82794 300134 83414 300218
rect 82794 299898 82826 300134
rect 83062 299898 83146 300134
rect 83382 299898 83414 300134
rect 82794 264454 83414 299898
rect 82794 264218 82826 264454
rect 83062 264218 83146 264454
rect 83382 264218 83414 264454
rect 82794 264134 83414 264218
rect 82794 263898 82826 264134
rect 83062 263898 83146 264134
rect 83382 263898 83414 264134
rect 82794 228454 83414 263898
rect 82794 228218 82826 228454
rect 83062 228218 83146 228454
rect 83382 228218 83414 228454
rect 82794 228134 83414 228218
rect 82794 227898 82826 228134
rect 83062 227898 83146 228134
rect 83382 227898 83414 228134
rect 82794 192454 83414 227898
rect 82794 192218 82826 192454
rect 83062 192218 83146 192454
rect 83382 192218 83414 192454
rect 82794 192134 83414 192218
rect 82794 191898 82826 192134
rect 83062 191898 83146 192134
rect 83382 191898 83414 192134
rect 82794 156454 83414 191898
rect 82794 156218 82826 156454
rect 83062 156218 83146 156454
rect 83382 156218 83414 156454
rect 82794 156134 83414 156218
rect 82794 155898 82826 156134
rect 83062 155898 83146 156134
rect 83382 155898 83414 156134
rect 82794 120454 83414 155898
rect 82794 120218 82826 120454
rect 83062 120218 83146 120454
rect 83382 120218 83414 120454
rect 82794 120134 83414 120218
rect 82794 119898 82826 120134
rect 83062 119898 83146 120134
rect 83382 119898 83414 120134
rect 82794 84454 83414 119898
rect 82794 84218 82826 84454
rect 83062 84218 83146 84454
rect 83382 84218 83414 84454
rect 82794 84134 83414 84218
rect 82794 83898 82826 84134
rect 83062 83898 83146 84134
rect 83382 83898 83414 84134
rect 82794 48454 83414 83898
rect 82794 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 83414 48454
rect 82794 48134 83414 48218
rect 82794 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 83414 48134
rect 82794 12454 83414 47898
rect 82794 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 83414 12454
rect 82794 12134 83414 12218
rect 82794 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 83414 12134
rect 82794 -2266 83414 11898
rect 82794 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 83414 -2266
rect 82794 -2586 83414 -2502
rect 82794 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 83414 -2586
rect 82794 -7654 83414 -2822
rect 87294 707718 87914 711590
rect 87294 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 87914 707718
rect 87294 707398 87914 707482
rect 87294 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 87914 707398
rect 87294 700954 87914 707162
rect 87294 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 87914 700954
rect 87294 700634 87914 700718
rect 87294 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 87914 700634
rect 87294 664954 87914 700398
rect 87294 664718 87326 664954
rect 87562 664718 87646 664954
rect 87882 664718 87914 664954
rect 87294 664634 87914 664718
rect 87294 664398 87326 664634
rect 87562 664398 87646 664634
rect 87882 664398 87914 664634
rect 87294 628954 87914 664398
rect 87294 628718 87326 628954
rect 87562 628718 87646 628954
rect 87882 628718 87914 628954
rect 87294 628634 87914 628718
rect 87294 628398 87326 628634
rect 87562 628398 87646 628634
rect 87882 628398 87914 628634
rect 87294 592954 87914 628398
rect 87294 592718 87326 592954
rect 87562 592718 87646 592954
rect 87882 592718 87914 592954
rect 87294 592634 87914 592718
rect 87294 592398 87326 592634
rect 87562 592398 87646 592634
rect 87882 592398 87914 592634
rect 87294 556954 87914 592398
rect 87294 556718 87326 556954
rect 87562 556718 87646 556954
rect 87882 556718 87914 556954
rect 87294 556634 87914 556718
rect 87294 556398 87326 556634
rect 87562 556398 87646 556634
rect 87882 556398 87914 556634
rect 87294 520954 87914 556398
rect 87294 520718 87326 520954
rect 87562 520718 87646 520954
rect 87882 520718 87914 520954
rect 87294 520634 87914 520718
rect 87294 520398 87326 520634
rect 87562 520398 87646 520634
rect 87882 520398 87914 520634
rect 87294 484954 87914 520398
rect 87294 484718 87326 484954
rect 87562 484718 87646 484954
rect 87882 484718 87914 484954
rect 87294 484634 87914 484718
rect 87294 484398 87326 484634
rect 87562 484398 87646 484634
rect 87882 484398 87914 484634
rect 87294 448954 87914 484398
rect 87294 448718 87326 448954
rect 87562 448718 87646 448954
rect 87882 448718 87914 448954
rect 87294 448634 87914 448718
rect 87294 448398 87326 448634
rect 87562 448398 87646 448634
rect 87882 448398 87914 448634
rect 87294 412954 87914 448398
rect 87294 412718 87326 412954
rect 87562 412718 87646 412954
rect 87882 412718 87914 412954
rect 87294 412634 87914 412718
rect 87294 412398 87326 412634
rect 87562 412398 87646 412634
rect 87882 412398 87914 412634
rect 87294 376954 87914 412398
rect 87294 376718 87326 376954
rect 87562 376718 87646 376954
rect 87882 376718 87914 376954
rect 87294 376634 87914 376718
rect 87294 376398 87326 376634
rect 87562 376398 87646 376634
rect 87882 376398 87914 376634
rect 87294 340954 87914 376398
rect 87294 340718 87326 340954
rect 87562 340718 87646 340954
rect 87882 340718 87914 340954
rect 87294 340634 87914 340718
rect 87294 340398 87326 340634
rect 87562 340398 87646 340634
rect 87882 340398 87914 340634
rect 87294 304954 87914 340398
rect 87294 304718 87326 304954
rect 87562 304718 87646 304954
rect 87882 304718 87914 304954
rect 87294 304634 87914 304718
rect 87294 304398 87326 304634
rect 87562 304398 87646 304634
rect 87882 304398 87914 304634
rect 87294 268954 87914 304398
rect 87294 268718 87326 268954
rect 87562 268718 87646 268954
rect 87882 268718 87914 268954
rect 87294 268634 87914 268718
rect 87294 268398 87326 268634
rect 87562 268398 87646 268634
rect 87882 268398 87914 268634
rect 87294 232954 87914 268398
rect 87294 232718 87326 232954
rect 87562 232718 87646 232954
rect 87882 232718 87914 232954
rect 87294 232634 87914 232718
rect 87294 232398 87326 232634
rect 87562 232398 87646 232634
rect 87882 232398 87914 232634
rect 87294 196954 87914 232398
rect 87294 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 87914 196954
rect 87294 196634 87914 196718
rect 87294 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 87914 196634
rect 87294 160954 87914 196398
rect 87294 160718 87326 160954
rect 87562 160718 87646 160954
rect 87882 160718 87914 160954
rect 87294 160634 87914 160718
rect 87294 160398 87326 160634
rect 87562 160398 87646 160634
rect 87882 160398 87914 160634
rect 87294 124954 87914 160398
rect 87294 124718 87326 124954
rect 87562 124718 87646 124954
rect 87882 124718 87914 124954
rect 87294 124634 87914 124718
rect 87294 124398 87326 124634
rect 87562 124398 87646 124634
rect 87882 124398 87914 124634
rect 87294 88954 87914 124398
rect 87294 88718 87326 88954
rect 87562 88718 87646 88954
rect 87882 88718 87914 88954
rect 87294 88634 87914 88718
rect 87294 88398 87326 88634
rect 87562 88398 87646 88634
rect 87882 88398 87914 88634
rect 87294 52954 87914 88398
rect 87294 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 87914 52954
rect 87294 52634 87914 52718
rect 87294 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 87914 52634
rect 87294 16954 87914 52398
rect 87294 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 87914 16954
rect 87294 16634 87914 16718
rect 87294 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 87914 16634
rect 87294 -3226 87914 16398
rect 87294 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 87914 -3226
rect 87294 -3546 87914 -3462
rect 87294 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 87914 -3546
rect 87294 -7654 87914 -3782
rect 91794 708678 92414 711590
rect 91794 708442 91826 708678
rect 92062 708442 92146 708678
rect 92382 708442 92414 708678
rect 91794 708358 92414 708442
rect 91794 708122 91826 708358
rect 92062 708122 92146 708358
rect 92382 708122 92414 708358
rect 91794 669454 92414 708122
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 561454 92414 596898
rect 91794 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 92414 561454
rect 91794 561134 92414 561218
rect 91794 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 92414 561134
rect 91794 525454 92414 560898
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 489454 92414 524898
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 91794 453454 92414 488898
rect 91794 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 92414 453454
rect 91794 453134 92414 453218
rect 91794 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 92414 453134
rect 91794 417454 92414 452898
rect 91794 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 92414 417454
rect 91794 417134 92414 417218
rect 91794 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 92414 417134
rect 91794 381454 92414 416898
rect 91794 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 92414 381454
rect 91794 381134 92414 381218
rect 91794 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 92414 381134
rect 91794 345454 92414 380898
rect 91794 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 92414 345454
rect 91794 345134 92414 345218
rect 91794 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 92414 345134
rect 91794 309454 92414 344898
rect 91794 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 92414 309454
rect 91794 309134 92414 309218
rect 91794 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 92414 309134
rect 91794 273454 92414 308898
rect 91794 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 92414 273454
rect 91794 273134 92414 273218
rect 91794 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 92414 273134
rect 91794 237454 92414 272898
rect 91794 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 92414 237454
rect 91794 237134 92414 237218
rect 91794 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 92414 237134
rect 91794 201454 92414 236898
rect 91794 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 92414 201454
rect 91794 201134 92414 201218
rect 91794 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 92414 201134
rect 91794 165454 92414 200898
rect 91794 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 92414 165454
rect 91794 165134 92414 165218
rect 91794 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 92414 165134
rect 91794 129454 92414 164898
rect 91794 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 92414 129454
rect 91794 129134 92414 129218
rect 91794 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 92414 129134
rect 91794 93454 92414 128898
rect 91794 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 92414 93454
rect 91794 93134 92414 93218
rect 91794 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 92414 93134
rect 91794 57454 92414 92898
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -4186 92414 20898
rect 91794 -4422 91826 -4186
rect 92062 -4422 92146 -4186
rect 92382 -4422 92414 -4186
rect 91794 -4506 92414 -4422
rect 91794 -4742 91826 -4506
rect 92062 -4742 92146 -4506
rect 92382 -4742 92414 -4506
rect 91794 -7654 92414 -4742
rect 96294 709638 96914 711590
rect 96294 709402 96326 709638
rect 96562 709402 96646 709638
rect 96882 709402 96914 709638
rect 96294 709318 96914 709402
rect 96294 709082 96326 709318
rect 96562 709082 96646 709318
rect 96882 709082 96914 709318
rect 96294 673954 96914 709082
rect 96294 673718 96326 673954
rect 96562 673718 96646 673954
rect 96882 673718 96914 673954
rect 96294 673634 96914 673718
rect 96294 673398 96326 673634
rect 96562 673398 96646 673634
rect 96882 673398 96914 673634
rect 96294 637954 96914 673398
rect 96294 637718 96326 637954
rect 96562 637718 96646 637954
rect 96882 637718 96914 637954
rect 96294 637634 96914 637718
rect 96294 637398 96326 637634
rect 96562 637398 96646 637634
rect 96882 637398 96914 637634
rect 96294 601954 96914 637398
rect 96294 601718 96326 601954
rect 96562 601718 96646 601954
rect 96882 601718 96914 601954
rect 96294 601634 96914 601718
rect 96294 601398 96326 601634
rect 96562 601398 96646 601634
rect 96882 601398 96914 601634
rect 96294 565954 96914 601398
rect 96294 565718 96326 565954
rect 96562 565718 96646 565954
rect 96882 565718 96914 565954
rect 96294 565634 96914 565718
rect 96294 565398 96326 565634
rect 96562 565398 96646 565634
rect 96882 565398 96914 565634
rect 96294 529954 96914 565398
rect 96294 529718 96326 529954
rect 96562 529718 96646 529954
rect 96882 529718 96914 529954
rect 96294 529634 96914 529718
rect 96294 529398 96326 529634
rect 96562 529398 96646 529634
rect 96882 529398 96914 529634
rect 96294 493954 96914 529398
rect 96294 493718 96326 493954
rect 96562 493718 96646 493954
rect 96882 493718 96914 493954
rect 96294 493634 96914 493718
rect 96294 493398 96326 493634
rect 96562 493398 96646 493634
rect 96882 493398 96914 493634
rect 96294 457954 96914 493398
rect 96294 457718 96326 457954
rect 96562 457718 96646 457954
rect 96882 457718 96914 457954
rect 96294 457634 96914 457718
rect 96294 457398 96326 457634
rect 96562 457398 96646 457634
rect 96882 457398 96914 457634
rect 96294 421954 96914 457398
rect 96294 421718 96326 421954
rect 96562 421718 96646 421954
rect 96882 421718 96914 421954
rect 96294 421634 96914 421718
rect 96294 421398 96326 421634
rect 96562 421398 96646 421634
rect 96882 421398 96914 421634
rect 96294 385954 96914 421398
rect 96294 385718 96326 385954
rect 96562 385718 96646 385954
rect 96882 385718 96914 385954
rect 96294 385634 96914 385718
rect 96294 385398 96326 385634
rect 96562 385398 96646 385634
rect 96882 385398 96914 385634
rect 96294 349954 96914 385398
rect 96294 349718 96326 349954
rect 96562 349718 96646 349954
rect 96882 349718 96914 349954
rect 96294 349634 96914 349718
rect 96294 349398 96326 349634
rect 96562 349398 96646 349634
rect 96882 349398 96914 349634
rect 96294 313954 96914 349398
rect 96294 313718 96326 313954
rect 96562 313718 96646 313954
rect 96882 313718 96914 313954
rect 96294 313634 96914 313718
rect 96294 313398 96326 313634
rect 96562 313398 96646 313634
rect 96882 313398 96914 313634
rect 96294 277954 96914 313398
rect 96294 277718 96326 277954
rect 96562 277718 96646 277954
rect 96882 277718 96914 277954
rect 96294 277634 96914 277718
rect 96294 277398 96326 277634
rect 96562 277398 96646 277634
rect 96882 277398 96914 277634
rect 96294 241954 96914 277398
rect 96294 241718 96326 241954
rect 96562 241718 96646 241954
rect 96882 241718 96914 241954
rect 96294 241634 96914 241718
rect 96294 241398 96326 241634
rect 96562 241398 96646 241634
rect 96882 241398 96914 241634
rect 96294 205954 96914 241398
rect 96294 205718 96326 205954
rect 96562 205718 96646 205954
rect 96882 205718 96914 205954
rect 96294 205634 96914 205718
rect 96294 205398 96326 205634
rect 96562 205398 96646 205634
rect 96882 205398 96914 205634
rect 96294 169954 96914 205398
rect 96294 169718 96326 169954
rect 96562 169718 96646 169954
rect 96882 169718 96914 169954
rect 96294 169634 96914 169718
rect 96294 169398 96326 169634
rect 96562 169398 96646 169634
rect 96882 169398 96914 169634
rect 96294 133954 96914 169398
rect 96294 133718 96326 133954
rect 96562 133718 96646 133954
rect 96882 133718 96914 133954
rect 96294 133634 96914 133718
rect 96294 133398 96326 133634
rect 96562 133398 96646 133634
rect 96882 133398 96914 133634
rect 96294 97954 96914 133398
rect 96294 97718 96326 97954
rect 96562 97718 96646 97954
rect 96882 97718 96914 97954
rect 96294 97634 96914 97718
rect 96294 97398 96326 97634
rect 96562 97398 96646 97634
rect 96882 97398 96914 97634
rect 96294 61954 96914 97398
rect 96294 61718 96326 61954
rect 96562 61718 96646 61954
rect 96882 61718 96914 61954
rect 96294 61634 96914 61718
rect 96294 61398 96326 61634
rect 96562 61398 96646 61634
rect 96882 61398 96914 61634
rect 96294 25954 96914 61398
rect 96294 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 96914 25954
rect 96294 25634 96914 25718
rect 96294 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 96914 25634
rect 96294 -5146 96914 25398
rect 96294 -5382 96326 -5146
rect 96562 -5382 96646 -5146
rect 96882 -5382 96914 -5146
rect 96294 -5466 96914 -5382
rect 96294 -5702 96326 -5466
rect 96562 -5702 96646 -5466
rect 96882 -5702 96914 -5466
rect 96294 -7654 96914 -5702
rect 100794 710598 101414 711590
rect 100794 710362 100826 710598
rect 101062 710362 101146 710598
rect 101382 710362 101414 710598
rect 100794 710278 101414 710362
rect 100794 710042 100826 710278
rect 101062 710042 101146 710278
rect 101382 710042 101414 710278
rect 100794 678454 101414 710042
rect 100794 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 101414 678454
rect 100794 678134 101414 678218
rect 100794 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 101414 678134
rect 100794 642454 101414 677898
rect 100794 642218 100826 642454
rect 101062 642218 101146 642454
rect 101382 642218 101414 642454
rect 100794 642134 101414 642218
rect 100794 641898 100826 642134
rect 101062 641898 101146 642134
rect 101382 641898 101414 642134
rect 100794 606454 101414 641898
rect 100794 606218 100826 606454
rect 101062 606218 101146 606454
rect 101382 606218 101414 606454
rect 100794 606134 101414 606218
rect 100794 605898 100826 606134
rect 101062 605898 101146 606134
rect 101382 605898 101414 606134
rect 100794 570454 101414 605898
rect 100794 570218 100826 570454
rect 101062 570218 101146 570454
rect 101382 570218 101414 570454
rect 100794 570134 101414 570218
rect 100794 569898 100826 570134
rect 101062 569898 101146 570134
rect 101382 569898 101414 570134
rect 100794 534454 101414 569898
rect 100794 534218 100826 534454
rect 101062 534218 101146 534454
rect 101382 534218 101414 534454
rect 100794 534134 101414 534218
rect 100794 533898 100826 534134
rect 101062 533898 101146 534134
rect 101382 533898 101414 534134
rect 100794 498454 101414 533898
rect 100794 498218 100826 498454
rect 101062 498218 101146 498454
rect 101382 498218 101414 498454
rect 100794 498134 101414 498218
rect 100794 497898 100826 498134
rect 101062 497898 101146 498134
rect 101382 497898 101414 498134
rect 100794 462454 101414 497898
rect 100794 462218 100826 462454
rect 101062 462218 101146 462454
rect 101382 462218 101414 462454
rect 100794 462134 101414 462218
rect 100794 461898 100826 462134
rect 101062 461898 101146 462134
rect 101382 461898 101414 462134
rect 100794 426454 101414 461898
rect 100794 426218 100826 426454
rect 101062 426218 101146 426454
rect 101382 426218 101414 426454
rect 100794 426134 101414 426218
rect 100794 425898 100826 426134
rect 101062 425898 101146 426134
rect 101382 425898 101414 426134
rect 100794 390454 101414 425898
rect 100794 390218 100826 390454
rect 101062 390218 101146 390454
rect 101382 390218 101414 390454
rect 100794 390134 101414 390218
rect 100794 389898 100826 390134
rect 101062 389898 101146 390134
rect 101382 389898 101414 390134
rect 100794 354454 101414 389898
rect 100794 354218 100826 354454
rect 101062 354218 101146 354454
rect 101382 354218 101414 354454
rect 100794 354134 101414 354218
rect 100794 353898 100826 354134
rect 101062 353898 101146 354134
rect 101382 353898 101414 354134
rect 100794 318454 101414 353898
rect 100794 318218 100826 318454
rect 101062 318218 101146 318454
rect 101382 318218 101414 318454
rect 100794 318134 101414 318218
rect 100794 317898 100826 318134
rect 101062 317898 101146 318134
rect 101382 317898 101414 318134
rect 100794 282454 101414 317898
rect 100794 282218 100826 282454
rect 101062 282218 101146 282454
rect 101382 282218 101414 282454
rect 100794 282134 101414 282218
rect 100794 281898 100826 282134
rect 101062 281898 101146 282134
rect 101382 281898 101414 282134
rect 100794 246454 101414 281898
rect 100794 246218 100826 246454
rect 101062 246218 101146 246454
rect 101382 246218 101414 246454
rect 100794 246134 101414 246218
rect 100794 245898 100826 246134
rect 101062 245898 101146 246134
rect 101382 245898 101414 246134
rect 100794 210454 101414 245898
rect 100794 210218 100826 210454
rect 101062 210218 101146 210454
rect 101382 210218 101414 210454
rect 100794 210134 101414 210218
rect 100794 209898 100826 210134
rect 101062 209898 101146 210134
rect 101382 209898 101414 210134
rect 100794 174454 101414 209898
rect 100794 174218 100826 174454
rect 101062 174218 101146 174454
rect 101382 174218 101414 174454
rect 100794 174134 101414 174218
rect 100794 173898 100826 174134
rect 101062 173898 101146 174134
rect 101382 173898 101414 174134
rect 100794 138454 101414 173898
rect 100794 138218 100826 138454
rect 101062 138218 101146 138454
rect 101382 138218 101414 138454
rect 100794 138134 101414 138218
rect 100794 137898 100826 138134
rect 101062 137898 101146 138134
rect 101382 137898 101414 138134
rect 100794 102454 101414 137898
rect 100794 102218 100826 102454
rect 101062 102218 101146 102454
rect 101382 102218 101414 102454
rect 100794 102134 101414 102218
rect 100794 101898 100826 102134
rect 101062 101898 101146 102134
rect 101382 101898 101414 102134
rect 100794 66454 101414 101898
rect 100794 66218 100826 66454
rect 101062 66218 101146 66454
rect 101382 66218 101414 66454
rect 100794 66134 101414 66218
rect 100794 65898 100826 66134
rect 101062 65898 101146 66134
rect 101382 65898 101414 66134
rect 100794 30454 101414 65898
rect 100794 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 101414 30454
rect 100794 30134 101414 30218
rect 100794 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 101414 30134
rect 100794 -6106 101414 29898
rect 100794 -6342 100826 -6106
rect 101062 -6342 101146 -6106
rect 101382 -6342 101414 -6106
rect 100794 -6426 101414 -6342
rect 100794 -6662 100826 -6426
rect 101062 -6662 101146 -6426
rect 101382 -6662 101414 -6426
rect 100794 -7654 101414 -6662
rect 105294 711558 105914 711590
rect 105294 711322 105326 711558
rect 105562 711322 105646 711558
rect 105882 711322 105914 711558
rect 105294 711238 105914 711322
rect 105294 711002 105326 711238
rect 105562 711002 105646 711238
rect 105882 711002 105914 711238
rect 105294 682954 105914 711002
rect 105294 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 105914 682954
rect 105294 682634 105914 682718
rect 105294 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 105914 682634
rect 105294 646954 105914 682398
rect 105294 646718 105326 646954
rect 105562 646718 105646 646954
rect 105882 646718 105914 646954
rect 105294 646634 105914 646718
rect 105294 646398 105326 646634
rect 105562 646398 105646 646634
rect 105882 646398 105914 646634
rect 105294 610954 105914 646398
rect 105294 610718 105326 610954
rect 105562 610718 105646 610954
rect 105882 610718 105914 610954
rect 105294 610634 105914 610718
rect 105294 610398 105326 610634
rect 105562 610398 105646 610634
rect 105882 610398 105914 610634
rect 105294 574954 105914 610398
rect 105294 574718 105326 574954
rect 105562 574718 105646 574954
rect 105882 574718 105914 574954
rect 105294 574634 105914 574718
rect 105294 574398 105326 574634
rect 105562 574398 105646 574634
rect 105882 574398 105914 574634
rect 105294 538954 105914 574398
rect 105294 538718 105326 538954
rect 105562 538718 105646 538954
rect 105882 538718 105914 538954
rect 105294 538634 105914 538718
rect 105294 538398 105326 538634
rect 105562 538398 105646 538634
rect 105882 538398 105914 538634
rect 105294 502954 105914 538398
rect 105294 502718 105326 502954
rect 105562 502718 105646 502954
rect 105882 502718 105914 502954
rect 105294 502634 105914 502718
rect 105294 502398 105326 502634
rect 105562 502398 105646 502634
rect 105882 502398 105914 502634
rect 105294 466954 105914 502398
rect 105294 466718 105326 466954
rect 105562 466718 105646 466954
rect 105882 466718 105914 466954
rect 105294 466634 105914 466718
rect 105294 466398 105326 466634
rect 105562 466398 105646 466634
rect 105882 466398 105914 466634
rect 105294 430954 105914 466398
rect 105294 430718 105326 430954
rect 105562 430718 105646 430954
rect 105882 430718 105914 430954
rect 105294 430634 105914 430718
rect 105294 430398 105326 430634
rect 105562 430398 105646 430634
rect 105882 430398 105914 430634
rect 105294 394954 105914 430398
rect 105294 394718 105326 394954
rect 105562 394718 105646 394954
rect 105882 394718 105914 394954
rect 105294 394634 105914 394718
rect 105294 394398 105326 394634
rect 105562 394398 105646 394634
rect 105882 394398 105914 394634
rect 105294 358954 105914 394398
rect 105294 358718 105326 358954
rect 105562 358718 105646 358954
rect 105882 358718 105914 358954
rect 105294 358634 105914 358718
rect 105294 358398 105326 358634
rect 105562 358398 105646 358634
rect 105882 358398 105914 358634
rect 105294 322954 105914 358398
rect 105294 322718 105326 322954
rect 105562 322718 105646 322954
rect 105882 322718 105914 322954
rect 105294 322634 105914 322718
rect 105294 322398 105326 322634
rect 105562 322398 105646 322634
rect 105882 322398 105914 322634
rect 105294 286954 105914 322398
rect 105294 286718 105326 286954
rect 105562 286718 105646 286954
rect 105882 286718 105914 286954
rect 105294 286634 105914 286718
rect 105294 286398 105326 286634
rect 105562 286398 105646 286634
rect 105882 286398 105914 286634
rect 105294 250954 105914 286398
rect 105294 250718 105326 250954
rect 105562 250718 105646 250954
rect 105882 250718 105914 250954
rect 105294 250634 105914 250718
rect 105294 250398 105326 250634
rect 105562 250398 105646 250634
rect 105882 250398 105914 250634
rect 105294 214954 105914 250398
rect 105294 214718 105326 214954
rect 105562 214718 105646 214954
rect 105882 214718 105914 214954
rect 105294 214634 105914 214718
rect 105294 214398 105326 214634
rect 105562 214398 105646 214634
rect 105882 214398 105914 214634
rect 105294 178954 105914 214398
rect 105294 178718 105326 178954
rect 105562 178718 105646 178954
rect 105882 178718 105914 178954
rect 105294 178634 105914 178718
rect 105294 178398 105326 178634
rect 105562 178398 105646 178634
rect 105882 178398 105914 178634
rect 105294 142954 105914 178398
rect 105294 142718 105326 142954
rect 105562 142718 105646 142954
rect 105882 142718 105914 142954
rect 105294 142634 105914 142718
rect 105294 142398 105326 142634
rect 105562 142398 105646 142634
rect 105882 142398 105914 142634
rect 105294 106954 105914 142398
rect 109794 704838 110414 711590
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 543454 110414 578898
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 109794 471454 110414 506898
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 435454 110414 470898
rect 109794 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 110414 435454
rect 109794 435134 110414 435218
rect 109794 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 110414 435134
rect 109794 399454 110414 434898
rect 109794 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 110414 399454
rect 109794 399134 110414 399218
rect 109794 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 110414 399134
rect 109794 363454 110414 398898
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 327454 110414 362898
rect 109794 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 110414 327454
rect 109794 327134 110414 327218
rect 109794 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 110414 327134
rect 109794 291454 110414 326898
rect 109794 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 110414 291454
rect 109794 291134 110414 291218
rect 109794 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 110414 291134
rect 109794 255454 110414 290898
rect 114294 705798 114914 711590
rect 114294 705562 114326 705798
rect 114562 705562 114646 705798
rect 114882 705562 114914 705798
rect 114294 705478 114914 705562
rect 114294 705242 114326 705478
rect 114562 705242 114646 705478
rect 114882 705242 114914 705478
rect 114294 691954 114914 705242
rect 114294 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 114914 691954
rect 114294 691634 114914 691718
rect 114294 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 114914 691634
rect 114294 655954 114914 691398
rect 114294 655718 114326 655954
rect 114562 655718 114646 655954
rect 114882 655718 114914 655954
rect 114294 655634 114914 655718
rect 114294 655398 114326 655634
rect 114562 655398 114646 655634
rect 114882 655398 114914 655634
rect 114294 619954 114914 655398
rect 114294 619718 114326 619954
rect 114562 619718 114646 619954
rect 114882 619718 114914 619954
rect 114294 619634 114914 619718
rect 114294 619398 114326 619634
rect 114562 619398 114646 619634
rect 114882 619398 114914 619634
rect 114294 583954 114914 619398
rect 114294 583718 114326 583954
rect 114562 583718 114646 583954
rect 114882 583718 114914 583954
rect 114294 583634 114914 583718
rect 114294 583398 114326 583634
rect 114562 583398 114646 583634
rect 114882 583398 114914 583634
rect 114294 547954 114914 583398
rect 114294 547718 114326 547954
rect 114562 547718 114646 547954
rect 114882 547718 114914 547954
rect 114294 547634 114914 547718
rect 114294 547398 114326 547634
rect 114562 547398 114646 547634
rect 114882 547398 114914 547634
rect 114294 511954 114914 547398
rect 114294 511718 114326 511954
rect 114562 511718 114646 511954
rect 114882 511718 114914 511954
rect 114294 511634 114914 511718
rect 114294 511398 114326 511634
rect 114562 511398 114646 511634
rect 114882 511398 114914 511634
rect 114294 475954 114914 511398
rect 114294 475718 114326 475954
rect 114562 475718 114646 475954
rect 114882 475718 114914 475954
rect 114294 475634 114914 475718
rect 114294 475398 114326 475634
rect 114562 475398 114646 475634
rect 114882 475398 114914 475634
rect 114294 439954 114914 475398
rect 114294 439718 114326 439954
rect 114562 439718 114646 439954
rect 114882 439718 114914 439954
rect 114294 439634 114914 439718
rect 114294 439398 114326 439634
rect 114562 439398 114646 439634
rect 114882 439398 114914 439634
rect 114294 403954 114914 439398
rect 114294 403718 114326 403954
rect 114562 403718 114646 403954
rect 114882 403718 114914 403954
rect 114294 403634 114914 403718
rect 114294 403398 114326 403634
rect 114562 403398 114646 403634
rect 114882 403398 114914 403634
rect 114294 367954 114914 403398
rect 114294 367718 114326 367954
rect 114562 367718 114646 367954
rect 114882 367718 114914 367954
rect 114294 367634 114914 367718
rect 114294 367398 114326 367634
rect 114562 367398 114646 367634
rect 114882 367398 114914 367634
rect 114294 331954 114914 367398
rect 114294 331718 114326 331954
rect 114562 331718 114646 331954
rect 114882 331718 114914 331954
rect 114294 331634 114914 331718
rect 114294 331398 114326 331634
rect 114562 331398 114646 331634
rect 114882 331398 114914 331634
rect 114294 295954 114914 331398
rect 114294 295718 114326 295954
rect 114562 295718 114646 295954
rect 114882 295718 114914 295954
rect 114294 295634 114914 295718
rect 114294 295398 114326 295634
rect 114562 295398 114646 295634
rect 114882 295398 114914 295634
rect 113035 265028 113101 265029
rect 113035 264964 113036 265028
rect 113100 264964 113101 265028
rect 113035 264963 113101 264964
rect 112851 262716 112917 262717
rect 112851 262652 112852 262716
rect 112916 262652 112917 262716
rect 112851 262651 112917 262652
rect 111563 262580 111629 262581
rect 111563 262516 111564 262580
rect 111628 262516 111629 262580
rect 111563 262515 111629 262516
rect 111379 262308 111445 262309
rect 111379 262244 111380 262308
rect 111444 262244 111445 262308
rect 111379 262243 111445 262244
rect 111195 260948 111261 260949
rect 111195 260884 111196 260948
rect 111260 260884 111261 260948
rect 111195 260883 111261 260884
rect 109794 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 110414 255454
rect 109794 255134 110414 255218
rect 109794 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 110414 255134
rect 109794 219454 110414 254898
rect 109794 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 110414 219454
rect 109794 219134 110414 219218
rect 109794 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 110414 219134
rect 109794 183454 110414 218898
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 109794 147454 110414 182898
rect 109794 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 110414 147454
rect 109794 147134 110414 147218
rect 109794 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 110414 147134
rect 108251 140452 108317 140453
rect 108251 140388 108252 140452
rect 108316 140388 108317 140452
rect 108251 140387 108317 140388
rect 105294 106718 105326 106954
rect 105562 106718 105646 106954
rect 105882 106718 105914 106954
rect 105294 106634 105914 106718
rect 105294 106398 105326 106634
rect 105562 106398 105646 106634
rect 105882 106398 105914 106634
rect 105294 70954 105914 106398
rect 105294 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 105914 70954
rect 105294 70634 105914 70718
rect 105294 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 105914 70634
rect 105294 34954 105914 70398
rect 105294 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 105914 34954
rect 105294 34634 105914 34718
rect 105294 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 105914 34634
rect 105294 -7066 105914 34398
rect 108254 19413 108314 140387
rect 109794 111454 110414 146898
rect 111198 145757 111258 260883
rect 111195 145756 111261 145757
rect 111195 145692 111196 145756
rect 111260 145692 111261 145756
rect 111195 145691 111261 145692
rect 111382 143445 111442 262243
rect 111379 143444 111445 143445
rect 111379 143380 111380 143444
rect 111444 143380 111445 143444
rect 111379 143379 111445 143380
rect 111566 143309 111626 262515
rect 112854 145893 112914 262651
rect 112851 145892 112917 145893
rect 112851 145828 112852 145892
rect 112916 145828 112917 145892
rect 112851 145827 112917 145828
rect 111563 143308 111629 143309
rect 111563 143244 111564 143308
rect 111628 143244 111629 143308
rect 111563 143243 111629 143244
rect 113038 140045 113098 264963
rect 114139 262444 114205 262445
rect 114139 262380 114140 262444
rect 114204 262380 114205 262444
rect 114139 262379 114205 262380
rect 113587 260404 113653 260405
rect 113587 260340 113588 260404
rect 113652 260340 113653 260404
rect 113587 260339 113653 260340
rect 113590 143989 113650 260339
rect 113955 259724 114021 259725
rect 113955 259660 113956 259724
rect 114020 259660 114021 259724
rect 113955 259659 114021 259660
rect 113771 189684 113837 189685
rect 113771 189620 113772 189684
rect 113836 189620 113837 189684
rect 113771 189619 113837 189620
rect 113587 143988 113653 143989
rect 113587 143924 113588 143988
rect 113652 143924 113653 143988
rect 113587 143923 113653 143924
rect 113035 140044 113101 140045
rect 113035 139980 113036 140044
rect 113100 139980 113101 140044
rect 113035 139979 113101 139980
rect 109794 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 110414 111454
rect 109794 111134 110414 111218
rect 109794 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 110414 111134
rect 109794 75454 110414 110898
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 113774 55045 113834 189619
rect 113958 142629 114018 259659
rect 114142 144533 114202 262379
rect 114294 259954 114914 295398
rect 118794 706758 119414 711590
rect 118794 706522 118826 706758
rect 119062 706522 119146 706758
rect 119382 706522 119414 706758
rect 118794 706438 119414 706522
rect 118794 706202 118826 706438
rect 119062 706202 119146 706438
rect 119382 706202 119414 706438
rect 118794 696454 119414 706202
rect 118794 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 119414 696454
rect 118794 696134 119414 696218
rect 118794 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 119414 696134
rect 118794 660454 119414 695898
rect 118794 660218 118826 660454
rect 119062 660218 119146 660454
rect 119382 660218 119414 660454
rect 118794 660134 119414 660218
rect 118794 659898 118826 660134
rect 119062 659898 119146 660134
rect 119382 659898 119414 660134
rect 118794 624454 119414 659898
rect 118794 624218 118826 624454
rect 119062 624218 119146 624454
rect 119382 624218 119414 624454
rect 118794 624134 119414 624218
rect 118794 623898 118826 624134
rect 119062 623898 119146 624134
rect 119382 623898 119414 624134
rect 118794 588454 119414 623898
rect 118794 588218 118826 588454
rect 119062 588218 119146 588454
rect 119382 588218 119414 588454
rect 118794 588134 119414 588218
rect 118794 587898 118826 588134
rect 119062 587898 119146 588134
rect 119382 587898 119414 588134
rect 118794 552454 119414 587898
rect 118794 552218 118826 552454
rect 119062 552218 119146 552454
rect 119382 552218 119414 552454
rect 118794 552134 119414 552218
rect 118794 551898 118826 552134
rect 119062 551898 119146 552134
rect 119382 551898 119414 552134
rect 118794 516454 119414 551898
rect 118794 516218 118826 516454
rect 119062 516218 119146 516454
rect 119382 516218 119414 516454
rect 118794 516134 119414 516218
rect 118794 515898 118826 516134
rect 119062 515898 119146 516134
rect 119382 515898 119414 516134
rect 118794 480454 119414 515898
rect 118794 480218 118826 480454
rect 119062 480218 119146 480454
rect 119382 480218 119414 480454
rect 118794 480134 119414 480218
rect 118794 479898 118826 480134
rect 119062 479898 119146 480134
rect 119382 479898 119414 480134
rect 118794 444454 119414 479898
rect 118794 444218 118826 444454
rect 119062 444218 119146 444454
rect 119382 444218 119414 444454
rect 118794 444134 119414 444218
rect 118794 443898 118826 444134
rect 119062 443898 119146 444134
rect 119382 443898 119414 444134
rect 118794 408454 119414 443898
rect 118794 408218 118826 408454
rect 119062 408218 119146 408454
rect 119382 408218 119414 408454
rect 118794 408134 119414 408218
rect 118794 407898 118826 408134
rect 119062 407898 119146 408134
rect 119382 407898 119414 408134
rect 118794 372454 119414 407898
rect 118794 372218 118826 372454
rect 119062 372218 119146 372454
rect 119382 372218 119414 372454
rect 118794 372134 119414 372218
rect 118794 371898 118826 372134
rect 119062 371898 119146 372134
rect 119382 371898 119414 372134
rect 118794 336454 119414 371898
rect 118794 336218 118826 336454
rect 119062 336218 119146 336454
rect 119382 336218 119414 336454
rect 118794 336134 119414 336218
rect 118794 335898 118826 336134
rect 119062 335898 119146 336134
rect 119382 335898 119414 336134
rect 118794 300454 119414 335898
rect 118794 300218 118826 300454
rect 119062 300218 119146 300454
rect 119382 300218 119414 300454
rect 118794 300134 119414 300218
rect 118794 299898 118826 300134
rect 119062 299898 119146 300134
rect 119382 299898 119414 300134
rect 118794 264454 119414 299898
rect 118794 264218 118826 264454
rect 119062 264218 119146 264454
rect 119382 264218 119414 264454
rect 118794 264134 119414 264218
rect 118794 263898 118826 264134
rect 119062 263898 119146 264134
rect 119382 263898 119414 264134
rect 118555 263668 118621 263669
rect 118555 263604 118556 263668
rect 118620 263604 118621 263668
rect 118555 263603 118621 263604
rect 115795 262852 115861 262853
rect 115795 262788 115796 262852
rect 115860 262788 115861 262852
rect 115795 262787 115861 262788
rect 115611 260132 115677 260133
rect 115611 260068 115612 260132
rect 115676 260068 115677 260132
rect 115611 260067 115677 260068
rect 114294 259718 114326 259954
rect 114562 259718 114646 259954
rect 114882 259718 114914 259954
rect 114294 259634 114914 259718
rect 114294 259398 114326 259634
rect 114562 259398 114646 259634
rect 114882 259398 114914 259634
rect 114294 223954 114914 259398
rect 114294 223718 114326 223954
rect 114562 223718 114646 223954
rect 114882 223718 114914 223954
rect 114294 223634 114914 223718
rect 114294 223398 114326 223634
rect 114562 223398 114646 223634
rect 114882 223398 114914 223634
rect 114294 187954 114914 223398
rect 114294 187718 114326 187954
rect 114562 187718 114646 187954
rect 114882 187718 114914 187954
rect 114294 187634 114914 187718
rect 114294 187398 114326 187634
rect 114562 187398 114646 187634
rect 114882 187398 114914 187634
rect 114294 151954 114914 187398
rect 114294 151718 114326 151954
rect 114562 151718 114646 151954
rect 114882 151718 114914 151954
rect 114294 151634 114914 151718
rect 114294 151398 114326 151634
rect 114562 151398 114646 151634
rect 114882 151398 114914 151634
rect 114139 144532 114205 144533
rect 114139 144468 114140 144532
rect 114204 144468 114205 144532
rect 114139 144467 114205 144468
rect 113955 142628 114021 142629
rect 113955 142564 113956 142628
rect 114020 142564 114021 142628
rect 113955 142563 114021 142564
rect 114294 115954 114914 151398
rect 115614 144805 115674 260067
rect 115611 144804 115677 144805
rect 115611 144740 115612 144804
rect 115676 144740 115677 144804
rect 115611 144739 115677 144740
rect 115798 144125 115858 262787
rect 118371 260268 118437 260269
rect 118371 260204 118372 260268
rect 118436 260204 118437 260268
rect 118371 260203 118437 260204
rect 116899 259996 116965 259997
rect 116899 259932 116900 259996
rect 116964 259932 116965 259996
rect 116899 259931 116965 259932
rect 116902 144669 116962 259931
rect 117083 259860 117149 259861
rect 117083 259796 117084 259860
rect 117148 259796 117149 259860
rect 117083 259795 117149 259796
rect 116899 144668 116965 144669
rect 116899 144604 116900 144668
rect 116964 144604 116965 144668
rect 116899 144603 116965 144604
rect 117086 144397 117146 259795
rect 118187 259588 118253 259589
rect 118187 259524 118188 259588
rect 118252 259524 118253 259588
rect 118187 259523 118253 259524
rect 117083 144396 117149 144397
rect 117083 144332 117084 144396
rect 117148 144332 117149 144396
rect 117083 144331 117149 144332
rect 118190 144261 118250 259523
rect 118187 144260 118253 144261
rect 118187 144196 118188 144260
rect 118252 144196 118253 144260
rect 118187 144195 118253 144196
rect 115795 144124 115861 144125
rect 115795 144060 115796 144124
rect 115860 144060 115861 144124
rect 115795 144059 115861 144060
rect 118374 141813 118434 260203
rect 118371 141812 118437 141813
rect 118371 141748 118372 141812
rect 118436 141748 118437 141812
rect 118371 141747 118437 141748
rect 117083 141676 117149 141677
rect 117083 141612 117084 141676
rect 117148 141612 117149 141676
rect 117083 141611 117149 141612
rect 116531 140860 116597 140861
rect 116531 140796 116532 140860
rect 116596 140796 116597 140860
rect 116531 140795 116597 140796
rect 114294 115718 114326 115954
rect 114562 115718 114646 115954
rect 114882 115718 114914 115954
rect 114294 115634 114914 115718
rect 114294 115398 114326 115634
rect 114562 115398 114646 115634
rect 114882 115398 114914 115634
rect 114294 79954 114914 115398
rect 114294 79718 114326 79954
rect 114562 79718 114646 79954
rect 114882 79718 114914 79954
rect 114294 79634 114914 79718
rect 114294 79398 114326 79634
rect 114562 79398 114646 79634
rect 114882 79398 114914 79634
rect 113771 55044 113837 55045
rect 113771 54980 113772 55044
rect 113836 54980 113837 55044
rect 113771 54979 113837 54980
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 108251 19412 108317 19413
rect 108251 19348 108252 19412
rect 108316 19348 108317 19412
rect 108251 19347 108317 19348
rect 105294 -7302 105326 -7066
rect 105562 -7302 105646 -7066
rect 105882 -7302 105914 -7066
rect 105294 -7386 105914 -7302
rect 105294 -7622 105326 -7386
rect 105562 -7622 105646 -7386
rect 105882 -7622 105914 -7386
rect 105294 -7654 105914 -7622
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -7654 110414 -902
rect 114294 43954 114914 79398
rect 116534 44301 116594 140795
rect 117086 75853 117146 141611
rect 118558 141405 118618 263603
rect 118794 262000 119414 263898
rect 123294 707718 123914 711590
rect 123294 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 123914 707718
rect 123294 707398 123914 707482
rect 123294 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 123914 707398
rect 123294 700954 123914 707162
rect 123294 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 123914 700954
rect 123294 700634 123914 700718
rect 123294 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 123914 700634
rect 123294 664954 123914 700398
rect 123294 664718 123326 664954
rect 123562 664718 123646 664954
rect 123882 664718 123914 664954
rect 123294 664634 123914 664718
rect 123294 664398 123326 664634
rect 123562 664398 123646 664634
rect 123882 664398 123914 664634
rect 123294 628954 123914 664398
rect 123294 628718 123326 628954
rect 123562 628718 123646 628954
rect 123882 628718 123914 628954
rect 123294 628634 123914 628718
rect 123294 628398 123326 628634
rect 123562 628398 123646 628634
rect 123882 628398 123914 628634
rect 123294 592954 123914 628398
rect 123294 592718 123326 592954
rect 123562 592718 123646 592954
rect 123882 592718 123914 592954
rect 123294 592634 123914 592718
rect 123294 592398 123326 592634
rect 123562 592398 123646 592634
rect 123882 592398 123914 592634
rect 123294 556954 123914 592398
rect 123294 556718 123326 556954
rect 123562 556718 123646 556954
rect 123882 556718 123914 556954
rect 123294 556634 123914 556718
rect 123294 556398 123326 556634
rect 123562 556398 123646 556634
rect 123882 556398 123914 556634
rect 123294 520954 123914 556398
rect 123294 520718 123326 520954
rect 123562 520718 123646 520954
rect 123882 520718 123914 520954
rect 123294 520634 123914 520718
rect 123294 520398 123326 520634
rect 123562 520398 123646 520634
rect 123882 520398 123914 520634
rect 123294 484954 123914 520398
rect 123294 484718 123326 484954
rect 123562 484718 123646 484954
rect 123882 484718 123914 484954
rect 123294 484634 123914 484718
rect 123294 484398 123326 484634
rect 123562 484398 123646 484634
rect 123882 484398 123914 484634
rect 123294 448954 123914 484398
rect 123294 448718 123326 448954
rect 123562 448718 123646 448954
rect 123882 448718 123914 448954
rect 123294 448634 123914 448718
rect 123294 448398 123326 448634
rect 123562 448398 123646 448634
rect 123882 448398 123914 448634
rect 123294 412954 123914 448398
rect 123294 412718 123326 412954
rect 123562 412718 123646 412954
rect 123882 412718 123914 412954
rect 123294 412634 123914 412718
rect 123294 412398 123326 412634
rect 123562 412398 123646 412634
rect 123882 412398 123914 412634
rect 123294 376954 123914 412398
rect 123294 376718 123326 376954
rect 123562 376718 123646 376954
rect 123882 376718 123914 376954
rect 123294 376634 123914 376718
rect 123294 376398 123326 376634
rect 123562 376398 123646 376634
rect 123882 376398 123914 376634
rect 123294 340954 123914 376398
rect 123294 340718 123326 340954
rect 123562 340718 123646 340954
rect 123882 340718 123914 340954
rect 123294 340634 123914 340718
rect 123294 340398 123326 340634
rect 123562 340398 123646 340634
rect 123882 340398 123914 340634
rect 123294 304954 123914 340398
rect 123294 304718 123326 304954
rect 123562 304718 123646 304954
rect 123882 304718 123914 304954
rect 123294 304634 123914 304718
rect 123294 304398 123326 304634
rect 123562 304398 123646 304634
rect 123882 304398 123914 304634
rect 123294 268954 123914 304398
rect 123294 268718 123326 268954
rect 123562 268718 123646 268954
rect 123882 268718 123914 268954
rect 123294 268634 123914 268718
rect 123294 268398 123326 268634
rect 123562 268398 123646 268634
rect 123882 268398 123914 268634
rect 121131 263804 121197 263805
rect 121131 263740 121132 263804
rect 121196 263740 121197 263804
rect 121131 263739 121197 263740
rect 120947 260540 121013 260541
rect 120947 260476 120948 260540
rect 121012 260476 121013 260540
rect 120947 260475 121013 260476
rect 118794 192454 119414 198000
rect 118794 192218 118826 192454
rect 119062 192218 119146 192454
rect 119382 192218 119414 192454
rect 118794 192134 119414 192218
rect 118794 191898 118826 192134
rect 119062 191898 119146 192134
rect 119382 191898 119414 192134
rect 118794 156454 119414 191898
rect 119843 185740 119909 185741
rect 119843 185676 119844 185740
rect 119908 185676 119909 185740
rect 119843 185675 119909 185676
rect 118794 156218 118826 156454
rect 119062 156218 119146 156454
rect 119382 156218 119414 156454
rect 118794 156134 119414 156218
rect 118794 155898 118826 156134
rect 119062 155898 119146 156134
rect 119382 155898 119414 156134
rect 118794 142000 119414 155898
rect 119659 144940 119725 144941
rect 119659 144876 119660 144940
rect 119724 144876 119725 144940
rect 119659 144875 119725 144876
rect 118555 141404 118621 141405
rect 118555 141340 118556 141404
rect 118620 141340 118621 141404
rect 118555 141339 118621 141340
rect 117819 140588 117885 140589
rect 117819 140524 117820 140588
rect 117884 140524 117885 140588
rect 117819 140523 117885 140524
rect 117083 75852 117149 75853
rect 117083 75788 117084 75852
rect 117148 75788 117149 75852
rect 117083 75787 117149 75788
rect 116531 44300 116597 44301
rect 116531 44236 116532 44300
rect 116596 44236 116597 44300
rect 116531 44235 116597 44236
rect 114294 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 114914 43954
rect 114294 43634 114914 43718
rect 114294 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 114914 43634
rect 114294 7954 114914 43398
rect 117822 31789 117882 140523
rect 119291 139908 119357 139909
rect 119291 139844 119292 139908
rect 119356 139844 119357 139908
rect 119291 139843 119357 139844
rect 118555 138684 118621 138685
rect 118555 138620 118556 138684
rect 118620 138620 118621 138684
rect 118555 138619 118621 138620
rect 118558 71501 118618 138619
rect 119294 84285 119354 139843
rect 119662 138030 119722 144875
rect 119478 137970 119722 138030
rect 119478 96661 119538 137970
rect 119659 130388 119725 130389
rect 119659 130324 119660 130388
rect 119724 130324 119725 130388
rect 119659 130323 119725 130324
rect 119475 96660 119541 96661
rect 119475 96596 119476 96660
rect 119540 96596 119541 96660
rect 119475 96595 119541 96596
rect 119291 84284 119357 84285
rect 119291 84220 119292 84284
rect 119356 84220 119357 84284
rect 119291 84219 119357 84220
rect 119662 83469 119722 130323
rect 119659 83468 119725 83469
rect 119659 83404 119660 83468
rect 119724 83404 119725 83468
rect 119659 83403 119725 83404
rect 118555 71500 118621 71501
rect 118555 71436 118556 71500
rect 118620 71436 118621 71500
rect 118555 71435 118621 71436
rect 118794 48454 119414 78000
rect 119846 77893 119906 185675
rect 120579 145620 120645 145621
rect 120579 145556 120580 145620
rect 120644 145556 120645 145620
rect 120579 145555 120645 145556
rect 120027 139228 120093 139229
rect 120027 139164 120028 139228
rect 120092 139164 120093 139228
rect 120027 139163 120093 139164
rect 120030 130389 120090 139163
rect 120027 130388 120093 130389
rect 120027 130324 120028 130388
rect 120092 130324 120093 130388
rect 120027 130323 120093 130324
rect 120027 83468 120093 83469
rect 120027 83404 120028 83468
rect 120092 83404 120093 83468
rect 120027 83403 120093 83404
rect 119843 77892 119909 77893
rect 119843 77828 119844 77892
rect 119908 77828 119909 77892
rect 119843 77827 119909 77828
rect 119846 75173 119906 77827
rect 119843 75172 119909 75173
rect 119843 75108 119844 75172
rect 119908 75108 119909 75172
rect 119843 75107 119909 75108
rect 120030 71637 120090 83403
rect 120582 74493 120642 145555
rect 120950 141541 121010 260475
rect 121134 143173 121194 263739
rect 123294 262000 123914 268398
rect 127794 708678 128414 711590
rect 127794 708442 127826 708678
rect 128062 708442 128146 708678
rect 128382 708442 128414 708678
rect 127794 708358 128414 708442
rect 127794 708122 127826 708358
rect 128062 708122 128146 708358
rect 128382 708122 128414 708358
rect 127794 669454 128414 708122
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 525454 128414 560898
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 127794 489454 128414 524898
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 127794 453454 128414 488898
rect 127794 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 128414 453454
rect 127794 453134 128414 453218
rect 127794 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 128414 453134
rect 127794 417454 128414 452898
rect 127794 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 128414 417454
rect 127794 417134 128414 417218
rect 127794 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 128414 417134
rect 127794 381454 128414 416898
rect 127794 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 128414 381454
rect 127794 381134 128414 381218
rect 127794 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 128414 381134
rect 127794 345454 128414 380898
rect 127794 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 128414 345454
rect 127794 345134 128414 345218
rect 127794 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 128414 345134
rect 127794 309454 128414 344898
rect 127794 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 128414 309454
rect 127794 309134 128414 309218
rect 127794 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 128414 309134
rect 127794 273454 128414 308898
rect 127794 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 128414 273454
rect 127794 273134 128414 273218
rect 127794 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 128414 273134
rect 127794 262000 128414 272898
rect 132294 709638 132914 711590
rect 132294 709402 132326 709638
rect 132562 709402 132646 709638
rect 132882 709402 132914 709638
rect 132294 709318 132914 709402
rect 132294 709082 132326 709318
rect 132562 709082 132646 709318
rect 132882 709082 132914 709318
rect 132294 673954 132914 709082
rect 132294 673718 132326 673954
rect 132562 673718 132646 673954
rect 132882 673718 132914 673954
rect 132294 673634 132914 673718
rect 132294 673398 132326 673634
rect 132562 673398 132646 673634
rect 132882 673398 132914 673634
rect 132294 637954 132914 673398
rect 132294 637718 132326 637954
rect 132562 637718 132646 637954
rect 132882 637718 132914 637954
rect 132294 637634 132914 637718
rect 132294 637398 132326 637634
rect 132562 637398 132646 637634
rect 132882 637398 132914 637634
rect 132294 601954 132914 637398
rect 132294 601718 132326 601954
rect 132562 601718 132646 601954
rect 132882 601718 132914 601954
rect 132294 601634 132914 601718
rect 132294 601398 132326 601634
rect 132562 601398 132646 601634
rect 132882 601398 132914 601634
rect 132294 565954 132914 601398
rect 132294 565718 132326 565954
rect 132562 565718 132646 565954
rect 132882 565718 132914 565954
rect 132294 565634 132914 565718
rect 132294 565398 132326 565634
rect 132562 565398 132646 565634
rect 132882 565398 132914 565634
rect 132294 529954 132914 565398
rect 132294 529718 132326 529954
rect 132562 529718 132646 529954
rect 132882 529718 132914 529954
rect 132294 529634 132914 529718
rect 132294 529398 132326 529634
rect 132562 529398 132646 529634
rect 132882 529398 132914 529634
rect 132294 493954 132914 529398
rect 132294 493718 132326 493954
rect 132562 493718 132646 493954
rect 132882 493718 132914 493954
rect 132294 493634 132914 493718
rect 132294 493398 132326 493634
rect 132562 493398 132646 493634
rect 132882 493398 132914 493634
rect 132294 457954 132914 493398
rect 132294 457718 132326 457954
rect 132562 457718 132646 457954
rect 132882 457718 132914 457954
rect 132294 457634 132914 457718
rect 132294 457398 132326 457634
rect 132562 457398 132646 457634
rect 132882 457398 132914 457634
rect 132294 421954 132914 457398
rect 132294 421718 132326 421954
rect 132562 421718 132646 421954
rect 132882 421718 132914 421954
rect 132294 421634 132914 421718
rect 132294 421398 132326 421634
rect 132562 421398 132646 421634
rect 132882 421398 132914 421634
rect 132294 385954 132914 421398
rect 132294 385718 132326 385954
rect 132562 385718 132646 385954
rect 132882 385718 132914 385954
rect 132294 385634 132914 385718
rect 132294 385398 132326 385634
rect 132562 385398 132646 385634
rect 132882 385398 132914 385634
rect 132294 349954 132914 385398
rect 132294 349718 132326 349954
rect 132562 349718 132646 349954
rect 132882 349718 132914 349954
rect 132294 349634 132914 349718
rect 132294 349398 132326 349634
rect 132562 349398 132646 349634
rect 132882 349398 132914 349634
rect 132294 313954 132914 349398
rect 132294 313718 132326 313954
rect 132562 313718 132646 313954
rect 132882 313718 132914 313954
rect 132294 313634 132914 313718
rect 132294 313398 132326 313634
rect 132562 313398 132646 313634
rect 132882 313398 132914 313634
rect 132294 277954 132914 313398
rect 132294 277718 132326 277954
rect 132562 277718 132646 277954
rect 132882 277718 132914 277954
rect 132294 277634 132914 277718
rect 132294 277398 132326 277634
rect 132562 277398 132646 277634
rect 132882 277398 132914 277634
rect 132294 262000 132914 277398
rect 136794 710598 137414 711590
rect 136794 710362 136826 710598
rect 137062 710362 137146 710598
rect 137382 710362 137414 710598
rect 136794 710278 137414 710362
rect 136794 710042 136826 710278
rect 137062 710042 137146 710278
rect 137382 710042 137414 710278
rect 136794 678454 137414 710042
rect 136794 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 137414 678454
rect 136794 678134 137414 678218
rect 136794 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 137414 678134
rect 136794 642454 137414 677898
rect 136794 642218 136826 642454
rect 137062 642218 137146 642454
rect 137382 642218 137414 642454
rect 136794 642134 137414 642218
rect 136794 641898 136826 642134
rect 137062 641898 137146 642134
rect 137382 641898 137414 642134
rect 136794 606454 137414 641898
rect 136794 606218 136826 606454
rect 137062 606218 137146 606454
rect 137382 606218 137414 606454
rect 136794 606134 137414 606218
rect 136794 605898 136826 606134
rect 137062 605898 137146 606134
rect 137382 605898 137414 606134
rect 136794 570454 137414 605898
rect 136794 570218 136826 570454
rect 137062 570218 137146 570454
rect 137382 570218 137414 570454
rect 136794 570134 137414 570218
rect 136794 569898 136826 570134
rect 137062 569898 137146 570134
rect 137382 569898 137414 570134
rect 136794 534454 137414 569898
rect 136794 534218 136826 534454
rect 137062 534218 137146 534454
rect 137382 534218 137414 534454
rect 136794 534134 137414 534218
rect 136794 533898 136826 534134
rect 137062 533898 137146 534134
rect 137382 533898 137414 534134
rect 136794 498454 137414 533898
rect 136794 498218 136826 498454
rect 137062 498218 137146 498454
rect 137382 498218 137414 498454
rect 136794 498134 137414 498218
rect 136794 497898 136826 498134
rect 137062 497898 137146 498134
rect 137382 497898 137414 498134
rect 136794 462454 137414 497898
rect 136794 462218 136826 462454
rect 137062 462218 137146 462454
rect 137382 462218 137414 462454
rect 136794 462134 137414 462218
rect 136794 461898 136826 462134
rect 137062 461898 137146 462134
rect 137382 461898 137414 462134
rect 136794 426454 137414 461898
rect 136794 426218 136826 426454
rect 137062 426218 137146 426454
rect 137382 426218 137414 426454
rect 136794 426134 137414 426218
rect 136794 425898 136826 426134
rect 137062 425898 137146 426134
rect 137382 425898 137414 426134
rect 136794 390454 137414 425898
rect 136794 390218 136826 390454
rect 137062 390218 137146 390454
rect 137382 390218 137414 390454
rect 136794 390134 137414 390218
rect 136794 389898 136826 390134
rect 137062 389898 137146 390134
rect 137382 389898 137414 390134
rect 136794 354454 137414 389898
rect 136794 354218 136826 354454
rect 137062 354218 137146 354454
rect 137382 354218 137414 354454
rect 136794 354134 137414 354218
rect 136794 353898 136826 354134
rect 137062 353898 137146 354134
rect 137382 353898 137414 354134
rect 136794 318454 137414 353898
rect 136794 318218 136826 318454
rect 137062 318218 137146 318454
rect 137382 318218 137414 318454
rect 136794 318134 137414 318218
rect 136794 317898 136826 318134
rect 137062 317898 137146 318134
rect 137382 317898 137414 318134
rect 136794 282454 137414 317898
rect 136794 282218 136826 282454
rect 137062 282218 137146 282454
rect 137382 282218 137414 282454
rect 136794 282134 137414 282218
rect 136794 281898 136826 282134
rect 137062 281898 137146 282134
rect 137382 281898 137414 282134
rect 136794 262000 137414 281898
rect 141294 711558 141914 711590
rect 141294 711322 141326 711558
rect 141562 711322 141646 711558
rect 141882 711322 141914 711558
rect 141294 711238 141914 711322
rect 141294 711002 141326 711238
rect 141562 711002 141646 711238
rect 141882 711002 141914 711238
rect 141294 682954 141914 711002
rect 141294 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 141914 682954
rect 141294 682634 141914 682718
rect 141294 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 141914 682634
rect 141294 646954 141914 682398
rect 141294 646718 141326 646954
rect 141562 646718 141646 646954
rect 141882 646718 141914 646954
rect 141294 646634 141914 646718
rect 141294 646398 141326 646634
rect 141562 646398 141646 646634
rect 141882 646398 141914 646634
rect 141294 610954 141914 646398
rect 141294 610718 141326 610954
rect 141562 610718 141646 610954
rect 141882 610718 141914 610954
rect 141294 610634 141914 610718
rect 141294 610398 141326 610634
rect 141562 610398 141646 610634
rect 141882 610398 141914 610634
rect 141294 574954 141914 610398
rect 141294 574718 141326 574954
rect 141562 574718 141646 574954
rect 141882 574718 141914 574954
rect 141294 574634 141914 574718
rect 141294 574398 141326 574634
rect 141562 574398 141646 574634
rect 141882 574398 141914 574634
rect 141294 538954 141914 574398
rect 141294 538718 141326 538954
rect 141562 538718 141646 538954
rect 141882 538718 141914 538954
rect 141294 538634 141914 538718
rect 141294 538398 141326 538634
rect 141562 538398 141646 538634
rect 141882 538398 141914 538634
rect 141294 502954 141914 538398
rect 141294 502718 141326 502954
rect 141562 502718 141646 502954
rect 141882 502718 141914 502954
rect 141294 502634 141914 502718
rect 141294 502398 141326 502634
rect 141562 502398 141646 502634
rect 141882 502398 141914 502634
rect 141294 466954 141914 502398
rect 141294 466718 141326 466954
rect 141562 466718 141646 466954
rect 141882 466718 141914 466954
rect 141294 466634 141914 466718
rect 141294 466398 141326 466634
rect 141562 466398 141646 466634
rect 141882 466398 141914 466634
rect 141294 430954 141914 466398
rect 141294 430718 141326 430954
rect 141562 430718 141646 430954
rect 141882 430718 141914 430954
rect 141294 430634 141914 430718
rect 141294 430398 141326 430634
rect 141562 430398 141646 430634
rect 141882 430398 141914 430634
rect 141294 394954 141914 430398
rect 141294 394718 141326 394954
rect 141562 394718 141646 394954
rect 141882 394718 141914 394954
rect 141294 394634 141914 394718
rect 141294 394398 141326 394634
rect 141562 394398 141646 394634
rect 141882 394398 141914 394634
rect 141294 358954 141914 394398
rect 141294 358718 141326 358954
rect 141562 358718 141646 358954
rect 141882 358718 141914 358954
rect 141294 358634 141914 358718
rect 141294 358398 141326 358634
rect 141562 358398 141646 358634
rect 141882 358398 141914 358634
rect 141294 322954 141914 358398
rect 141294 322718 141326 322954
rect 141562 322718 141646 322954
rect 141882 322718 141914 322954
rect 141294 322634 141914 322718
rect 141294 322398 141326 322634
rect 141562 322398 141646 322634
rect 141882 322398 141914 322634
rect 141294 286954 141914 322398
rect 141294 286718 141326 286954
rect 141562 286718 141646 286954
rect 141882 286718 141914 286954
rect 141294 286634 141914 286718
rect 141294 286398 141326 286634
rect 141562 286398 141646 286634
rect 141882 286398 141914 286634
rect 141294 262000 141914 286398
rect 145794 704838 146414 711590
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 363454 146414 398898
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 327454 146414 362898
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 145794 291454 146414 326898
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 262000 146414 290898
rect 150294 705798 150914 711590
rect 150294 705562 150326 705798
rect 150562 705562 150646 705798
rect 150882 705562 150914 705798
rect 150294 705478 150914 705562
rect 150294 705242 150326 705478
rect 150562 705242 150646 705478
rect 150882 705242 150914 705478
rect 150294 691954 150914 705242
rect 150294 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 150914 691954
rect 150294 691634 150914 691718
rect 150294 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 150914 691634
rect 150294 655954 150914 691398
rect 150294 655718 150326 655954
rect 150562 655718 150646 655954
rect 150882 655718 150914 655954
rect 150294 655634 150914 655718
rect 150294 655398 150326 655634
rect 150562 655398 150646 655634
rect 150882 655398 150914 655634
rect 150294 619954 150914 655398
rect 150294 619718 150326 619954
rect 150562 619718 150646 619954
rect 150882 619718 150914 619954
rect 150294 619634 150914 619718
rect 150294 619398 150326 619634
rect 150562 619398 150646 619634
rect 150882 619398 150914 619634
rect 150294 583954 150914 619398
rect 150294 583718 150326 583954
rect 150562 583718 150646 583954
rect 150882 583718 150914 583954
rect 150294 583634 150914 583718
rect 150294 583398 150326 583634
rect 150562 583398 150646 583634
rect 150882 583398 150914 583634
rect 150294 547954 150914 583398
rect 150294 547718 150326 547954
rect 150562 547718 150646 547954
rect 150882 547718 150914 547954
rect 150294 547634 150914 547718
rect 150294 547398 150326 547634
rect 150562 547398 150646 547634
rect 150882 547398 150914 547634
rect 150294 511954 150914 547398
rect 150294 511718 150326 511954
rect 150562 511718 150646 511954
rect 150882 511718 150914 511954
rect 150294 511634 150914 511718
rect 150294 511398 150326 511634
rect 150562 511398 150646 511634
rect 150882 511398 150914 511634
rect 150294 475954 150914 511398
rect 150294 475718 150326 475954
rect 150562 475718 150646 475954
rect 150882 475718 150914 475954
rect 150294 475634 150914 475718
rect 150294 475398 150326 475634
rect 150562 475398 150646 475634
rect 150882 475398 150914 475634
rect 150294 439954 150914 475398
rect 150294 439718 150326 439954
rect 150562 439718 150646 439954
rect 150882 439718 150914 439954
rect 150294 439634 150914 439718
rect 150294 439398 150326 439634
rect 150562 439398 150646 439634
rect 150882 439398 150914 439634
rect 150294 403954 150914 439398
rect 150294 403718 150326 403954
rect 150562 403718 150646 403954
rect 150882 403718 150914 403954
rect 150294 403634 150914 403718
rect 150294 403398 150326 403634
rect 150562 403398 150646 403634
rect 150882 403398 150914 403634
rect 150294 367954 150914 403398
rect 150294 367718 150326 367954
rect 150562 367718 150646 367954
rect 150882 367718 150914 367954
rect 150294 367634 150914 367718
rect 150294 367398 150326 367634
rect 150562 367398 150646 367634
rect 150882 367398 150914 367634
rect 150294 331954 150914 367398
rect 150294 331718 150326 331954
rect 150562 331718 150646 331954
rect 150882 331718 150914 331954
rect 150294 331634 150914 331718
rect 150294 331398 150326 331634
rect 150562 331398 150646 331634
rect 150882 331398 150914 331634
rect 150294 295954 150914 331398
rect 150294 295718 150326 295954
rect 150562 295718 150646 295954
rect 150882 295718 150914 295954
rect 150294 295634 150914 295718
rect 150294 295398 150326 295634
rect 150562 295398 150646 295634
rect 150882 295398 150914 295634
rect 150294 262000 150914 295398
rect 154794 706758 155414 711590
rect 154794 706522 154826 706758
rect 155062 706522 155146 706758
rect 155382 706522 155414 706758
rect 154794 706438 155414 706522
rect 154794 706202 154826 706438
rect 155062 706202 155146 706438
rect 155382 706202 155414 706438
rect 154794 696454 155414 706202
rect 154794 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 155414 696454
rect 154794 696134 155414 696218
rect 154794 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 155414 696134
rect 154794 660454 155414 695898
rect 154794 660218 154826 660454
rect 155062 660218 155146 660454
rect 155382 660218 155414 660454
rect 154794 660134 155414 660218
rect 154794 659898 154826 660134
rect 155062 659898 155146 660134
rect 155382 659898 155414 660134
rect 154794 624454 155414 659898
rect 154794 624218 154826 624454
rect 155062 624218 155146 624454
rect 155382 624218 155414 624454
rect 154794 624134 155414 624218
rect 154794 623898 154826 624134
rect 155062 623898 155146 624134
rect 155382 623898 155414 624134
rect 154794 588454 155414 623898
rect 154794 588218 154826 588454
rect 155062 588218 155146 588454
rect 155382 588218 155414 588454
rect 154794 588134 155414 588218
rect 154794 587898 154826 588134
rect 155062 587898 155146 588134
rect 155382 587898 155414 588134
rect 154794 552454 155414 587898
rect 154794 552218 154826 552454
rect 155062 552218 155146 552454
rect 155382 552218 155414 552454
rect 154794 552134 155414 552218
rect 154794 551898 154826 552134
rect 155062 551898 155146 552134
rect 155382 551898 155414 552134
rect 154794 516454 155414 551898
rect 154794 516218 154826 516454
rect 155062 516218 155146 516454
rect 155382 516218 155414 516454
rect 154794 516134 155414 516218
rect 154794 515898 154826 516134
rect 155062 515898 155146 516134
rect 155382 515898 155414 516134
rect 154794 480454 155414 515898
rect 154794 480218 154826 480454
rect 155062 480218 155146 480454
rect 155382 480218 155414 480454
rect 154794 480134 155414 480218
rect 154794 479898 154826 480134
rect 155062 479898 155146 480134
rect 155382 479898 155414 480134
rect 154794 444454 155414 479898
rect 154794 444218 154826 444454
rect 155062 444218 155146 444454
rect 155382 444218 155414 444454
rect 154794 444134 155414 444218
rect 154794 443898 154826 444134
rect 155062 443898 155146 444134
rect 155382 443898 155414 444134
rect 154794 408454 155414 443898
rect 154794 408218 154826 408454
rect 155062 408218 155146 408454
rect 155382 408218 155414 408454
rect 154794 408134 155414 408218
rect 154794 407898 154826 408134
rect 155062 407898 155146 408134
rect 155382 407898 155414 408134
rect 154794 372454 155414 407898
rect 154794 372218 154826 372454
rect 155062 372218 155146 372454
rect 155382 372218 155414 372454
rect 154794 372134 155414 372218
rect 154794 371898 154826 372134
rect 155062 371898 155146 372134
rect 155382 371898 155414 372134
rect 154794 336454 155414 371898
rect 154794 336218 154826 336454
rect 155062 336218 155146 336454
rect 155382 336218 155414 336454
rect 154794 336134 155414 336218
rect 154794 335898 154826 336134
rect 155062 335898 155146 336134
rect 155382 335898 155414 336134
rect 154794 300454 155414 335898
rect 154794 300218 154826 300454
rect 155062 300218 155146 300454
rect 155382 300218 155414 300454
rect 154794 300134 155414 300218
rect 154794 299898 154826 300134
rect 155062 299898 155146 300134
rect 155382 299898 155414 300134
rect 154794 264454 155414 299898
rect 154794 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 155414 264454
rect 154794 264134 155414 264218
rect 154794 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 155414 264134
rect 154794 262000 155414 263898
rect 159294 707718 159914 711590
rect 159294 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 159914 707718
rect 159294 707398 159914 707482
rect 159294 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 159914 707398
rect 159294 700954 159914 707162
rect 159294 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 159914 700954
rect 159294 700634 159914 700718
rect 159294 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 159914 700634
rect 159294 664954 159914 700398
rect 159294 664718 159326 664954
rect 159562 664718 159646 664954
rect 159882 664718 159914 664954
rect 159294 664634 159914 664718
rect 159294 664398 159326 664634
rect 159562 664398 159646 664634
rect 159882 664398 159914 664634
rect 159294 628954 159914 664398
rect 159294 628718 159326 628954
rect 159562 628718 159646 628954
rect 159882 628718 159914 628954
rect 159294 628634 159914 628718
rect 159294 628398 159326 628634
rect 159562 628398 159646 628634
rect 159882 628398 159914 628634
rect 159294 592954 159914 628398
rect 159294 592718 159326 592954
rect 159562 592718 159646 592954
rect 159882 592718 159914 592954
rect 159294 592634 159914 592718
rect 159294 592398 159326 592634
rect 159562 592398 159646 592634
rect 159882 592398 159914 592634
rect 159294 556954 159914 592398
rect 159294 556718 159326 556954
rect 159562 556718 159646 556954
rect 159882 556718 159914 556954
rect 159294 556634 159914 556718
rect 159294 556398 159326 556634
rect 159562 556398 159646 556634
rect 159882 556398 159914 556634
rect 159294 520954 159914 556398
rect 159294 520718 159326 520954
rect 159562 520718 159646 520954
rect 159882 520718 159914 520954
rect 159294 520634 159914 520718
rect 159294 520398 159326 520634
rect 159562 520398 159646 520634
rect 159882 520398 159914 520634
rect 159294 484954 159914 520398
rect 159294 484718 159326 484954
rect 159562 484718 159646 484954
rect 159882 484718 159914 484954
rect 159294 484634 159914 484718
rect 159294 484398 159326 484634
rect 159562 484398 159646 484634
rect 159882 484398 159914 484634
rect 159294 448954 159914 484398
rect 159294 448718 159326 448954
rect 159562 448718 159646 448954
rect 159882 448718 159914 448954
rect 159294 448634 159914 448718
rect 159294 448398 159326 448634
rect 159562 448398 159646 448634
rect 159882 448398 159914 448634
rect 159294 412954 159914 448398
rect 159294 412718 159326 412954
rect 159562 412718 159646 412954
rect 159882 412718 159914 412954
rect 159294 412634 159914 412718
rect 159294 412398 159326 412634
rect 159562 412398 159646 412634
rect 159882 412398 159914 412634
rect 159294 376954 159914 412398
rect 159294 376718 159326 376954
rect 159562 376718 159646 376954
rect 159882 376718 159914 376954
rect 159294 376634 159914 376718
rect 159294 376398 159326 376634
rect 159562 376398 159646 376634
rect 159882 376398 159914 376634
rect 159294 340954 159914 376398
rect 159294 340718 159326 340954
rect 159562 340718 159646 340954
rect 159882 340718 159914 340954
rect 159294 340634 159914 340718
rect 159294 340398 159326 340634
rect 159562 340398 159646 340634
rect 159882 340398 159914 340634
rect 159294 304954 159914 340398
rect 159294 304718 159326 304954
rect 159562 304718 159646 304954
rect 159882 304718 159914 304954
rect 159294 304634 159914 304718
rect 159294 304398 159326 304634
rect 159562 304398 159646 304634
rect 159882 304398 159914 304634
rect 159294 268954 159914 304398
rect 159294 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 159914 268954
rect 159294 268634 159914 268718
rect 159294 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 159914 268634
rect 159294 262000 159914 268398
rect 163794 708678 164414 711590
rect 163794 708442 163826 708678
rect 164062 708442 164146 708678
rect 164382 708442 164414 708678
rect 163794 708358 164414 708442
rect 163794 708122 163826 708358
rect 164062 708122 164146 708358
rect 164382 708122 164414 708358
rect 163794 669454 164414 708122
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 525454 164414 560898
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 163794 489454 164414 524898
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 453454 164414 488898
rect 163794 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 164414 453454
rect 163794 453134 164414 453218
rect 163794 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 164414 453134
rect 163794 417454 164414 452898
rect 163794 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 164414 417454
rect 163794 417134 164414 417218
rect 163794 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 164414 417134
rect 163794 381454 164414 416898
rect 163794 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 164414 381454
rect 163794 381134 164414 381218
rect 163794 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 164414 381134
rect 163794 345454 164414 380898
rect 163794 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 164414 345454
rect 163794 345134 164414 345218
rect 163794 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 164414 345134
rect 163794 309454 164414 344898
rect 163794 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 164414 309454
rect 163794 309134 164414 309218
rect 163794 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 164414 309134
rect 163794 273454 164414 308898
rect 163794 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 164414 273454
rect 163794 273134 164414 273218
rect 163794 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 164414 273134
rect 163794 262000 164414 272898
rect 168294 709638 168914 711590
rect 168294 709402 168326 709638
rect 168562 709402 168646 709638
rect 168882 709402 168914 709638
rect 168294 709318 168914 709402
rect 168294 709082 168326 709318
rect 168562 709082 168646 709318
rect 168882 709082 168914 709318
rect 168294 673954 168914 709082
rect 168294 673718 168326 673954
rect 168562 673718 168646 673954
rect 168882 673718 168914 673954
rect 168294 673634 168914 673718
rect 168294 673398 168326 673634
rect 168562 673398 168646 673634
rect 168882 673398 168914 673634
rect 168294 637954 168914 673398
rect 168294 637718 168326 637954
rect 168562 637718 168646 637954
rect 168882 637718 168914 637954
rect 168294 637634 168914 637718
rect 168294 637398 168326 637634
rect 168562 637398 168646 637634
rect 168882 637398 168914 637634
rect 168294 601954 168914 637398
rect 168294 601718 168326 601954
rect 168562 601718 168646 601954
rect 168882 601718 168914 601954
rect 168294 601634 168914 601718
rect 168294 601398 168326 601634
rect 168562 601398 168646 601634
rect 168882 601398 168914 601634
rect 168294 565954 168914 601398
rect 168294 565718 168326 565954
rect 168562 565718 168646 565954
rect 168882 565718 168914 565954
rect 168294 565634 168914 565718
rect 168294 565398 168326 565634
rect 168562 565398 168646 565634
rect 168882 565398 168914 565634
rect 168294 529954 168914 565398
rect 168294 529718 168326 529954
rect 168562 529718 168646 529954
rect 168882 529718 168914 529954
rect 168294 529634 168914 529718
rect 168294 529398 168326 529634
rect 168562 529398 168646 529634
rect 168882 529398 168914 529634
rect 168294 493954 168914 529398
rect 168294 493718 168326 493954
rect 168562 493718 168646 493954
rect 168882 493718 168914 493954
rect 168294 493634 168914 493718
rect 168294 493398 168326 493634
rect 168562 493398 168646 493634
rect 168882 493398 168914 493634
rect 168294 457954 168914 493398
rect 168294 457718 168326 457954
rect 168562 457718 168646 457954
rect 168882 457718 168914 457954
rect 168294 457634 168914 457718
rect 168294 457398 168326 457634
rect 168562 457398 168646 457634
rect 168882 457398 168914 457634
rect 168294 421954 168914 457398
rect 168294 421718 168326 421954
rect 168562 421718 168646 421954
rect 168882 421718 168914 421954
rect 168294 421634 168914 421718
rect 168294 421398 168326 421634
rect 168562 421398 168646 421634
rect 168882 421398 168914 421634
rect 168294 385954 168914 421398
rect 168294 385718 168326 385954
rect 168562 385718 168646 385954
rect 168882 385718 168914 385954
rect 168294 385634 168914 385718
rect 168294 385398 168326 385634
rect 168562 385398 168646 385634
rect 168882 385398 168914 385634
rect 168294 349954 168914 385398
rect 168294 349718 168326 349954
rect 168562 349718 168646 349954
rect 168882 349718 168914 349954
rect 168294 349634 168914 349718
rect 168294 349398 168326 349634
rect 168562 349398 168646 349634
rect 168882 349398 168914 349634
rect 168294 313954 168914 349398
rect 168294 313718 168326 313954
rect 168562 313718 168646 313954
rect 168882 313718 168914 313954
rect 168294 313634 168914 313718
rect 168294 313398 168326 313634
rect 168562 313398 168646 313634
rect 168882 313398 168914 313634
rect 168294 277954 168914 313398
rect 168294 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 168914 277954
rect 168294 277634 168914 277718
rect 168294 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 168914 277634
rect 168294 262000 168914 277398
rect 172794 710598 173414 711590
rect 172794 710362 172826 710598
rect 173062 710362 173146 710598
rect 173382 710362 173414 710598
rect 172794 710278 173414 710362
rect 172794 710042 172826 710278
rect 173062 710042 173146 710278
rect 173382 710042 173414 710278
rect 172794 678454 173414 710042
rect 172794 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 173414 678454
rect 172794 678134 173414 678218
rect 172794 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 173414 678134
rect 172794 642454 173414 677898
rect 172794 642218 172826 642454
rect 173062 642218 173146 642454
rect 173382 642218 173414 642454
rect 172794 642134 173414 642218
rect 172794 641898 172826 642134
rect 173062 641898 173146 642134
rect 173382 641898 173414 642134
rect 172794 606454 173414 641898
rect 172794 606218 172826 606454
rect 173062 606218 173146 606454
rect 173382 606218 173414 606454
rect 172794 606134 173414 606218
rect 172794 605898 172826 606134
rect 173062 605898 173146 606134
rect 173382 605898 173414 606134
rect 172794 570454 173414 605898
rect 172794 570218 172826 570454
rect 173062 570218 173146 570454
rect 173382 570218 173414 570454
rect 172794 570134 173414 570218
rect 172794 569898 172826 570134
rect 173062 569898 173146 570134
rect 173382 569898 173414 570134
rect 172794 534454 173414 569898
rect 172794 534218 172826 534454
rect 173062 534218 173146 534454
rect 173382 534218 173414 534454
rect 172794 534134 173414 534218
rect 172794 533898 172826 534134
rect 173062 533898 173146 534134
rect 173382 533898 173414 534134
rect 172794 498454 173414 533898
rect 172794 498218 172826 498454
rect 173062 498218 173146 498454
rect 173382 498218 173414 498454
rect 172794 498134 173414 498218
rect 172794 497898 172826 498134
rect 173062 497898 173146 498134
rect 173382 497898 173414 498134
rect 172794 462454 173414 497898
rect 172794 462218 172826 462454
rect 173062 462218 173146 462454
rect 173382 462218 173414 462454
rect 172794 462134 173414 462218
rect 172794 461898 172826 462134
rect 173062 461898 173146 462134
rect 173382 461898 173414 462134
rect 172794 426454 173414 461898
rect 172794 426218 172826 426454
rect 173062 426218 173146 426454
rect 173382 426218 173414 426454
rect 172794 426134 173414 426218
rect 172794 425898 172826 426134
rect 173062 425898 173146 426134
rect 173382 425898 173414 426134
rect 172794 390454 173414 425898
rect 172794 390218 172826 390454
rect 173062 390218 173146 390454
rect 173382 390218 173414 390454
rect 172794 390134 173414 390218
rect 172794 389898 172826 390134
rect 173062 389898 173146 390134
rect 173382 389898 173414 390134
rect 172794 354454 173414 389898
rect 172794 354218 172826 354454
rect 173062 354218 173146 354454
rect 173382 354218 173414 354454
rect 172794 354134 173414 354218
rect 172794 353898 172826 354134
rect 173062 353898 173146 354134
rect 173382 353898 173414 354134
rect 172794 318454 173414 353898
rect 172794 318218 172826 318454
rect 173062 318218 173146 318454
rect 173382 318218 173414 318454
rect 172794 318134 173414 318218
rect 172794 317898 172826 318134
rect 173062 317898 173146 318134
rect 173382 317898 173414 318134
rect 172794 282454 173414 317898
rect 172794 282218 172826 282454
rect 173062 282218 173146 282454
rect 173382 282218 173414 282454
rect 172794 282134 173414 282218
rect 172794 281898 172826 282134
rect 173062 281898 173146 282134
rect 173382 281898 173414 282134
rect 172794 262000 173414 281898
rect 177294 711558 177914 711590
rect 177294 711322 177326 711558
rect 177562 711322 177646 711558
rect 177882 711322 177914 711558
rect 177294 711238 177914 711322
rect 177294 711002 177326 711238
rect 177562 711002 177646 711238
rect 177882 711002 177914 711238
rect 177294 682954 177914 711002
rect 177294 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 177914 682954
rect 177294 682634 177914 682718
rect 177294 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 177914 682634
rect 177294 646954 177914 682398
rect 177294 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 177914 646954
rect 177294 646634 177914 646718
rect 177294 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 177914 646634
rect 177294 610954 177914 646398
rect 177294 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 177914 610954
rect 177294 610634 177914 610718
rect 177294 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 177914 610634
rect 177294 574954 177914 610398
rect 177294 574718 177326 574954
rect 177562 574718 177646 574954
rect 177882 574718 177914 574954
rect 177294 574634 177914 574718
rect 177294 574398 177326 574634
rect 177562 574398 177646 574634
rect 177882 574398 177914 574634
rect 177294 538954 177914 574398
rect 177294 538718 177326 538954
rect 177562 538718 177646 538954
rect 177882 538718 177914 538954
rect 177294 538634 177914 538718
rect 177294 538398 177326 538634
rect 177562 538398 177646 538634
rect 177882 538398 177914 538634
rect 177294 502954 177914 538398
rect 177294 502718 177326 502954
rect 177562 502718 177646 502954
rect 177882 502718 177914 502954
rect 177294 502634 177914 502718
rect 177294 502398 177326 502634
rect 177562 502398 177646 502634
rect 177882 502398 177914 502634
rect 177294 466954 177914 502398
rect 177294 466718 177326 466954
rect 177562 466718 177646 466954
rect 177882 466718 177914 466954
rect 177294 466634 177914 466718
rect 177294 466398 177326 466634
rect 177562 466398 177646 466634
rect 177882 466398 177914 466634
rect 177294 430954 177914 466398
rect 177294 430718 177326 430954
rect 177562 430718 177646 430954
rect 177882 430718 177914 430954
rect 177294 430634 177914 430718
rect 177294 430398 177326 430634
rect 177562 430398 177646 430634
rect 177882 430398 177914 430634
rect 177294 394954 177914 430398
rect 177294 394718 177326 394954
rect 177562 394718 177646 394954
rect 177882 394718 177914 394954
rect 177294 394634 177914 394718
rect 177294 394398 177326 394634
rect 177562 394398 177646 394634
rect 177882 394398 177914 394634
rect 177294 358954 177914 394398
rect 177294 358718 177326 358954
rect 177562 358718 177646 358954
rect 177882 358718 177914 358954
rect 177294 358634 177914 358718
rect 177294 358398 177326 358634
rect 177562 358398 177646 358634
rect 177882 358398 177914 358634
rect 177294 322954 177914 358398
rect 177294 322718 177326 322954
rect 177562 322718 177646 322954
rect 177882 322718 177914 322954
rect 177294 322634 177914 322718
rect 177294 322398 177326 322634
rect 177562 322398 177646 322634
rect 177882 322398 177914 322634
rect 177294 286954 177914 322398
rect 177294 286718 177326 286954
rect 177562 286718 177646 286954
rect 177882 286718 177914 286954
rect 177294 286634 177914 286718
rect 177294 286398 177326 286634
rect 177562 286398 177646 286634
rect 177882 286398 177914 286634
rect 177294 262000 177914 286398
rect 181794 704838 182414 711590
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181794 363454 182414 398898
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 181794 291454 182414 326898
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181794 262000 182414 290898
rect 186294 705798 186914 711590
rect 186294 705562 186326 705798
rect 186562 705562 186646 705798
rect 186882 705562 186914 705798
rect 186294 705478 186914 705562
rect 186294 705242 186326 705478
rect 186562 705242 186646 705478
rect 186882 705242 186914 705478
rect 186294 691954 186914 705242
rect 186294 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 186914 691954
rect 186294 691634 186914 691718
rect 186294 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 186914 691634
rect 186294 655954 186914 691398
rect 186294 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 186914 655954
rect 186294 655634 186914 655718
rect 186294 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 186914 655634
rect 186294 619954 186914 655398
rect 186294 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 186914 619954
rect 186294 619634 186914 619718
rect 186294 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 186914 619634
rect 186294 583954 186914 619398
rect 186294 583718 186326 583954
rect 186562 583718 186646 583954
rect 186882 583718 186914 583954
rect 186294 583634 186914 583718
rect 186294 583398 186326 583634
rect 186562 583398 186646 583634
rect 186882 583398 186914 583634
rect 186294 547954 186914 583398
rect 186294 547718 186326 547954
rect 186562 547718 186646 547954
rect 186882 547718 186914 547954
rect 186294 547634 186914 547718
rect 186294 547398 186326 547634
rect 186562 547398 186646 547634
rect 186882 547398 186914 547634
rect 186294 511954 186914 547398
rect 186294 511718 186326 511954
rect 186562 511718 186646 511954
rect 186882 511718 186914 511954
rect 186294 511634 186914 511718
rect 186294 511398 186326 511634
rect 186562 511398 186646 511634
rect 186882 511398 186914 511634
rect 186294 475954 186914 511398
rect 186294 475718 186326 475954
rect 186562 475718 186646 475954
rect 186882 475718 186914 475954
rect 186294 475634 186914 475718
rect 186294 475398 186326 475634
rect 186562 475398 186646 475634
rect 186882 475398 186914 475634
rect 186294 439954 186914 475398
rect 186294 439718 186326 439954
rect 186562 439718 186646 439954
rect 186882 439718 186914 439954
rect 186294 439634 186914 439718
rect 186294 439398 186326 439634
rect 186562 439398 186646 439634
rect 186882 439398 186914 439634
rect 186294 403954 186914 439398
rect 186294 403718 186326 403954
rect 186562 403718 186646 403954
rect 186882 403718 186914 403954
rect 186294 403634 186914 403718
rect 186294 403398 186326 403634
rect 186562 403398 186646 403634
rect 186882 403398 186914 403634
rect 186294 367954 186914 403398
rect 186294 367718 186326 367954
rect 186562 367718 186646 367954
rect 186882 367718 186914 367954
rect 186294 367634 186914 367718
rect 186294 367398 186326 367634
rect 186562 367398 186646 367634
rect 186882 367398 186914 367634
rect 186294 331954 186914 367398
rect 186294 331718 186326 331954
rect 186562 331718 186646 331954
rect 186882 331718 186914 331954
rect 186294 331634 186914 331718
rect 186294 331398 186326 331634
rect 186562 331398 186646 331634
rect 186882 331398 186914 331634
rect 186294 295954 186914 331398
rect 186294 295718 186326 295954
rect 186562 295718 186646 295954
rect 186882 295718 186914 295954
rect 186294 295634 186914 295718
rect 186294 295398 186326 295634
rect 186562 295398 186646 295634
rect 186882 295398 186914 295634
rect 186294 262000 186914 295398
rect 190794 706758 191414 711590
rect 190794 706522 190826 706758
rect 191062 706522 191146 706758
rect 191382 706522 191414 706758
rect 190794 706438 191414 706522
rect 190794 706202 190826 706438
rect 191062 706202 191146 706438
rect 191382 706202 191414 706438
rect 190794 696454 191414 706202
rect 190794 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 191414 696454
rect 190794 696134 191414 696218
rect 190794 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 191414 696134
rect 190794 660454 191414 695898
rect 190794 660218 190826 660454
rect 191062 660218 191146 660454
rect 191382 660218 191414 660454
rect 190794 660134 191414 660218
rect 190794 659898 190826 660134
rect 191062 659898 191146 660134
rect 191382 659898 191414 660134
rect 190794 624454 191414 659898
rect 190794 624218 190826 624454
rect 191062 624218 191146 624454
rect 191382 624218 191414 624454
rect 190794 624134 191414 624218
rect 190794 623898 190826 624134
rect 191062 623898 191146 624134
rect 191382 623898 191414 624134
rect 190794 588454 191414 623898
rect 190794 588218 190826 588454
rect 191062 588218 191146 588454
rect 191382 588218 191414 588454
rect 190794 588134 191414 588218
rect 190794 587898 190826 588134
rect 191062 587898 191146 588134
rect 191382 587898 191414 588134
rect 190794 552454 191414 587898
rect 190794 552218 190826 552454
rect 191062 552218 191146 552454
rect 191382 552218 191414 552454
rect 190794 552134 191414 552218
rect 190794 551898 190826 552134
rect 191062 551898 191146 552134
rect 191382 551898 191414 552134
rect 190794 516454 191414 551898
rect 190794 516218 190826 516454
rect 191062 516218 191146 516454
rect 191382 516218 191414 516454
rect 190794 516134 191414 516218
rect 190794 515898 190826 516134
rect 191062 515898 191146 516134
rect 191382 515898 191414 516134
rect 190794 480454 191414 515898
rect 190794 480218 190826 480454
rect 191062 480218 191146 480454
rect 191382 480218 191414 480454
rect 190794 480134 191414 480218
rect 190794 479898 190826 480134
rect 191062 479898 191146 480134
rect 191382 479898 191414 480134
rect 190794 444454 191414 479898
rect 190794 444218 190826 444454
rect 191062 444218 191146 444454
rect 191382 444218 191414 444454
rect 190794 444134 191414 444218
rect 190794 443898 190826 444134
rect 191062 443898 191146 444134
rect 191382 443898 191414 444134
rect 190794 408454 191414 443898
rect 190794 408218 190826 408454
rect 191062 408218 191146 408454
rect 191382 408218 191414 408454
rect 190794 408134 191414 408218
rect 190794 407898 190826 408134
rect 191062 407898 191146 408134
rect 191382 407898 191414 408134
rect 190794 372454 191414 407898
rect 190794 372218 190826 372454
rect 191062 372218 191146 372454
rect 191382 372218 191414 372454
rect 190794 372134 191414 372218
rect 190794 371898 190826 372134
rect 191062 371898 191146 372134
rect 191382 371898 191414 372134
rect 190794 336454 191414 371898
rect 190794 336218 190826 336454
rect 191062 336218 191146 336454
rect 191382 336218 191414 336454
rect 190794 336134 191414 336218
rect 190794 335898 190826 336134
rect 191062 335898 191146 336134
rect 191382 335898 191414 336134
rect 190794 300454 191414 335898
rect 190794 300218 190826 300454
rect 191062 300218 191146 300454
rect 191382 300218 191414 300454
rect 190794 300134 191414 300218
rect 190794 299898 190826 300134
rect 191062 299898 191146 300134
rect 191382 299898 191414 300134
rect 189027 276044 189093 276045
rect 189027 275980 189028 276044
rect 189092 275980 189093 276044
rect 189027 275979 189093 275980
rect 187003 271148 187069 271149
rect 187003 271084 187004 271148
rect 187068 271084 187069 271148
rect 187003 271083 187069 271084
rect 187006 270605 187066 271083
rect 187003 270604 187069 270605
rect 187003 270540 187004 270604
rect 187068 270540 187069 270604
rect 187003 270539 187069 270540
rect 185347 259588 185413 259589
rect 185347 259524 185348 259588
rect 185412 259524 185413 259588
rect 185347 259523 185413 259524
rect 186083 259588 186149 259589
rect 186083 259524 186084 259588
rect 186148 259524 186149 259588
rect 186083 259523 186149 259524
rect 124208 255454 124528 255486
rect 124208 255218 124250 255454
rect 124486 255218 124528 255454
rect 124208 255134 124528 255218
rect 124208 254898 124250 255134
rect 124486 254898 124528 255134
rect 124208 254866 124528 254898
rect 154928 255454 155248 255486
rect 154928 255218 154970 255454
rect 155206 255218 155248 255454
rect 154928 255134 155248 255218
rect 154928 254898 154970 255134
rect 155206 254898 155248 255134
rect 154928 254866 155248 254898
rect 139568 223954 139888 223986
rect 139568 223718 139610 223954
rect 139846 223718 139888 223954
rect 139568 223634 139888 223718
rect 139568 223398 139610 223634
rect 139846 223398 139888 223634
rect 139568 223366 139888 223398
rect 170288 223954 170608 223986
rect 170288 223718 170330 223954
rect 170566 223718 170608 223954
rect 170288 223634 170608 223718
rect 170288 223398 170330 223634
rect 170566 223398 170608 223634
rect 170288 223366 170608 223398
rect 124208 219454 124528 219486
rect 124208 219218 124250 219454
rect 124486 219218 124528 219454
rect 124208 219134 124528 219218
rect 124208 218898 124250 219134
rect 124486 218898 124528 219134
rect 124208 218866 124528 218898
rect 154928 219454 155248 219486
rect 154928 219218 154970 219454
rect 155206 219218 155248 219454
rect 154928 219134 155248 219218
rect 154928 218898 154970 219134
rect 155206 218898 155248 219134
rect 154928 218866 155248 218898
rect 185350 201789 185410 259523
rect 185648 255454 185968 255486
rect 185648 255218 185690 255454
rect 185926 255218 185968 255454
rect 185648 255134 185968 255218
rect 185648 254898 185690 255134
rect 185926 254898 185968 255134
rect 185648 254866 185968 254898
rect 186086 222210 186146 259523
rect 186086 222150 186514 222210
rect 185648 219454 185968 219486
rect 185648 219218 185690 219454
rect 185926 219218 185968 219454
rect 185648 219134 185968 219218
rect 185648 218898 185690 219134
rect 185926 218898 185968 219134
rect 185648 218866 185968 218898
rect 186454 210357 186514 222150
rect 186451 210356 186517 210357
rect 186451 210292 186452 210356
rect 186516 210292 186517 210356
rect 186451 210291 186517 210292
rect 186083 202876 186149 202877
rect 186083 202812 186084 202876
rect 186148 202812 186149 202876
rect 186083 202811 186149 202812
rect 185347 201788 185413 201789
rect 185347 201724 185348 201788
rect 185412 201724 185413 201788
rect 185347 201723 185413 201724
rect 157195 200700 157261 200701
rect 157195 200636 157196 200700
rect 157260 200636 157261 200700
rect 157195 200635 157261 200636
rect 179827 200700 179893 200701
rect 179827 200636 179828 200700
rect 179892 200636 179893 200700
rect 179827 200635 179893 200636
rect 137875 200292 137941 200293
rect 137875 200228 137876 200292
rect 137940 200228 137941 200292
rect 137875 200227 137941 200228
rect 136403 200156 136469 200157
rect 136403 200092 136404 200156
rect 136468 200092 136469 200156
rect 136403 200091 136469 200092
rect 137507 200156 137573 200157
rect 137507 200092 137508 200156
rect 137572 200092 137573 200156
rect 137507 200091 137573 200092
rect 132723 199884 132789 199885
rect 132723 199820 132724 199884
rect 132788 199820 132789 199884
rect 132723 199819 132789 199820
rect 133091 199884 133157 199885
rect 133091 199820 133092 199884
rect 133156 199820 133157 199884
rect 133091 199819 133157 199820
rect 133459 199884 133525 199885
rect 133459 199820 133460 199884
rect 133524 199820 133525 199884
rect 133459 199819 133525 199820
rect 134195 199884 134261 199885
rect 134195 199820 134196 199884
rect 134260 199820 134261 199884
rect 134195 199819 134261 199820
rect 134379 199884 134445 199885
rect 134379 199820 134380 199884
rect 134444 199820 134445 199884
rect 134379 199819 134445 199820
rect 134747 199884 134813 199885
rect 134747 199820 134748 199884
rect 134812 199820 134813 199884
rect 134747 199819 134813 199820
rect 135115 199884 135181 199885
rect 135115 199820 135116 199884
rect 135180 199820 135181 199884
rect 135115 199819 135181 199820
rect 135483 199884 135549 199885
rect 135483 199820 135484 199884
rect 135548 199820 135549 199884
rect 135483 199819 135549 199820
rect 135851 199884 135917 199885
rect 135851 199820 135852 199884
rect 135916 199820 135917 199884
rect 135851 199819 135917 199820
rect 121315 197300 121381 197301
rect 121315 197236 121316 197300
rect 121380 197236 121381 197300
rect 121315 197235 121381 197236
rect 121131 143172 121197 143173
rect 121131 143108 121132 143172
rect 121196 143108 121197 143172
rect 121131 143107 121197 143108
rect 120947 141540 121013 141541
rect 120947 141476 120948 141540
rect 121012 141476 121013 141540
rect 120947 141475 121013 141476
rect 120763 140724 120829 140725
rect 120763 140660 120764 140724
rect 120828 140660 120829 140724
rect 120763 140659 120829 140660
rect 120766 79661 120826 140659
rect 120947 139092 121013 139093
rect 120947 139028 120948 139092
rect 121012 139028 121013 139092
rect 120947 139027 121013 139028
rect 120763 79660 120829 79661
rect 120763 79596 120764 79660
rect 120828 79596 120829 79660
rect 120763 79595 120829 79596
rect 120579 74492 120645 74493
rect 120579 74428 120580 74492
rect 120644 74428 120645 74492
rect 120579 74427 120645 74428
rect 120027 71636 120093 71637
rect 120027 71572 120028 71636
rect 120092 71572 120093 71636
rect 120027 71571 120093 71572
rect 120950 68917 121010 139027
rect 121318 73133 121378 197235
rect 123294 196954 123914 198000
rect 132726 197981 132786 199819
rect 133094 199613 133154 199819
rect 133091 199612 133157 199613
rect 133091 199548 133092 199612
rect 133156 199548 133157 199612
rect 133091 199547 133157 199548
rect 133462 197981 133522 199819
rect 134198 199341 134258 199819
rect 134195 199340 134261 199341
rect 134195 199276 134196 199340
rect 134260 199276 134261 199340
rect 134195 199275 134261 199276
rect 133827 198388 133893 198389
rect 133827 198324 133828 198388
rect 133892 198324 133893 198388
rect 133827 198323 133893 198324
rect 134195 198388 134261 198389
rect 134195 198324 134196 198388
rect 134260 198324 134261 198388
rect 134195 198323 134261 198324
rect 132723 197980 132789 197981
rect 132723 197916 132724 197980
rect 132788 197916 132789 197980
rect 132723 197915 132789 197916
rect 133459 197980 133525 197981
rect 133459 197916 133460 197980
rect 133524 197916 133525 197980
rect 133459 197915 133525 197916
rect 132355 197844 132421 197845
rect 132355 197780 132356 197844
rect 132420 197780 132421 197844
rect 132355 197779 132421 197780
rect 123294 196718 123326 196954
rect 123562 196718 123646 196954
rect 123882 196718 123914 196954
rect 123294 196634 123914 196718
rect 123294 196398 123326 196634
rect 123562 196398 123646 196634
rect 123882 196398 123914 196634
rect 122971 192268 123037 192269
rect 122971 192204 122972 192268
rect 123036 192204 123037 192268
rect 122971 192203 123037 192204
rect 122235 191316 122301 191317
rect 122235 191252 122236 191316
rect 122300 191252 122301 191316
rect 122235 191251 122301 191252
rect 122051 139364 122117 139365
rect 122051 139300 122052 139364
rect 122116 139300 122117 139364
rect 122051 139299 122117 139300
rect 122054 78845 122114 139299
rect 122238 81429 122298 191251
rect 122603 189956 122669 189957
rect 122603 189892 122604 189956
rect 122668 189892 122669 189956
rect 122603 189891 122669 189892
rect 122419 186692 122485 186693
rect 122419 186628 122420 186692
rect 122484 186628 122485 186692
rect 122419 186627 122485 186628
rect 122235 81428 122301 81429
rect 122235 81364 122236 81428
rect 122300 81364 122301 81428
rect 122235 81363 122301 81364
rect 122422 80613 122482 186627
rect 122419 80612 122485 80613
rect 122419 80548 122420 80612
rect 122484 80548 122485 80612
rect 122419 80547 122485 80548
rect 122606 78981 122666 189891
rect 122787 138004 122853 138005
rect 122787 137940 122788 138004
rect 122852 137940 122853 138004
rect 122787 137939 122853 137940
rect 122790 128485 122850 137939
rect 122787 128484 122853 128485
rect 122787 128420 122788 128484
rect 122852 128420 122853 128484
rect 122787 128419 122853 128420
rect 122787 122908 122853 122909
rect 122787 122844 122788 122908
rect 122852 122844 122853 122908
rect 122787 122843 122853 122844
rect 122790 122773 122850 122843
rect 122787 122772 122853 122773
rect 122787 122708 122788 122772
rect 122852 122708 122853 122772
rect 122787 122707 122853 122708
rect 122787 113388 122853 113389
rect 122787 113324 122788 113388
rect 122852 113324 122853 113388
rect 122787 113323 122853 113324
rect 122790 112981 122850 113323
rect 122787 112980 122853 112981
rect 122787 112916 122788 112980
rect 122852 112916 122853 112980
rect 122787 112915 122853 112916
rect 122787 103596 122853 103597
rect 122787 103532 122788 103596
rect 122852 103532 122853 103596
rect 122787 103531 122853 103532
rect 122790 103325 122850 103531
rect 122787 103324 122853 103325
rect 122787 103260 122788 103324
rect 122852 103260 122853 103324
rect 122787 103259 122853 103260
rect 122787 93940 122853 93941
rect 122787 93876 122788 93940
rect 122852 93876 122853 93940
rect 122787 93875 122853 93876
rect 122790 93669 122850 93875
rect 122787 93668 122853 93669
rect 122787 93604 122788 93668
rect 122852 93604 122853 93668
rect 122787 93603 122853 93604
rect 122787 89724 122853 89725
rect 122787 89660 122788 89724
rect 122852 89660 122853 89724
rect 122787 89659 122853 89660
rect 122790 80341 122850 89659
rect 122974 81021 123034 192203
rect 123294 160954 123914 196398
rect 130331 194308 130397 194309
rect 130331 194244 130332 194308
rect 130396 194244 130397 194308
rect 130331 194243 130397 194244
rect 127571 193764 127637 193765
rect 127571 193700 127572 193764
rect 127636 193700 127637 193764
rect 127571 193699 127637 193700
rect 124995 192948 125061 192949
rect 124995 192884 124996 192948
rect 125060 192884 125061 192948
rect 124995 192883 125061 192884
rect 124811 191860 124877 191861
rect 124811 191796 124812 191860
rect 124876 191796 124877 191860
rect 124811 191795 124877 191796
rect 124075 191180 124141 191181
rect 124075 191116 124076 191180
rect 124140 191116 124141 191180
rect 124075 191115 124141 191116
rect 123294 160718 123326 160954
rect 123562 160718 123646 160954
rect 123882 160718 123914 160954
rect 123294 160634 123914 160718
rect 123294 160398 123326 160634
rect 123562 160398 123646 160634
rect 123882 160398 123914 160634
rect 123294 142000 123914 160398
rect 122971 81020 123037 81021
rect 122971 80956 122972 81020
rect 123036 80956 123037 81020
rect 122971 80955 123037 80956
rect 122787 80340 122853 80341
rect 122787 80276 122788 80340
rect 122852 80276 122853 80340
rect 122787 80275 122853 80276
rect 122603 78980 122669 78981
rect 122603 78916 122604 78980
rect 122668 78916 122669 78980
rect 122603 78915 122669 78916
rect 122051 78844 122117 78845
rect 122051 78780 122052 78844
rect 122116 78780 122117 78844
rect 122051 78779 122117 78780
rect 124078 78165 124138 191115
rect 124208 111454 124528 111486
rect 124208 111218 124250 111454
rect 124486 111218 124528 111454
rect 124208 111134 124528 111218
rect 124208 110898 124250 111134
rect 124486 110898 124528 111134
rect 124208 110866 124528 110898
rect 124075 78164 124141 78165
rect 124075 78100 124076 78164
rect 124140 78100 124141 78164
rect 124075 78099 124141 78100
rect 121315 73132 121381 73133
rect 121315 73068 121316 73132
rect 121380 73068 121381 73132
rect 121315 73067 121381 73068
rect 120947 68916 121013 68917
rect 120947 68852 120948 68916
rect 121012 68852 121013 68916
rect 120947 68851 121013 68852
rect 118794 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 119414 48454
rect 118794 48134 119414 48218
rect 118794 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 119414 48134
rect 117819 31788 117885 31789
rect 117819 31724 117820 31788
rect 117884 31724 117885 31788
rect 117819 31723 117885 31724
rect 114294 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 114914 7954
rect 114294 7634 114914 7718
rect 114294 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 114914 7634
rect 114294 -1306 114914 7398
rect 114294 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 114914 -1306
rect 114294 -1626 114914 -1542
rect 114294 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 114914 -1626
rect 114294 -7654 114914 -1862
rect 118794 12454 119414 47898
rect 118794 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 119414 12454
rect 118794 12134 119414 12218
rect 118794 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 119414 12134
rect 118794 -2266 119414 11898
rect 118794 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 119414 -2266
rect 118794 -2586 119414 -2502
rect 118794 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 119414 -2586
rect 118794 -7654 119414 -2822
rect 123294 52954 123914 78000
rect 124814 77757 124874 191795
rect 124811 77756 124877 77757
rect 124811 77692 124812 77756
rect 124876 77692 124877 77756
rect 124811 77691 124877 77692
rect 124998 77349 125058 192883
rect 126835 191452 126901 191453
rect 126835 191388 126836 191452
rect 126900 191388 126901 191452
rect 126835 191387 126901 191388
rect 125179 190364 125245 190365
rect 125179 190300 125180 190364
rect 125244 190300 125245 190364
rect 125179 190299 125245 190300
rect 125182 78437 125242 190299
rect 126651 187372 126717 187373
rect 126651 187308 126652 187372
rect 126716 187308 126717 187372
rect 126651 187307 126717 187308
rect 125363 186012 125429 186013
rect 125363 185948 125364 186012
rect 125428 185948 125429 186012
rect 125363 185947 125429 185948
rect 125366 79253 125426 185947
rect 126467 139364 126533 139365
rect 126467 139300 126468 139364
rect 126532 139300 126533 139364
rect 126467 139299 126533 139300
rect 126470 79797 126530 139299
rect 126654 80885 126714 187307
rect 126651 80884 126717 80885
rect 126651 80820 126652 80884
rect 126716 80820 126717 80884
rect 126651 80819 126717 80820
rect 126467 79796 126533 79797
rect 126467 79732 126468 79796
rect 126532 79732 126533 79796
rect 126467 79731 126533 79732
rect 125363 79252 125429 79253
rect 125363 79188 125364 79252
rect 125428 79188 125429 79252
rect 125363 79187 125429 79188
rect 125179 78436 125245 78437
rect 125179 78372 125180 78436
rect 125244 78372 125245 78436
rect 125179 78371 125245 78372
rect 126838 78301 126898 191387
rect 127387 187236 127453 187237
rect 127387 187172 127388 187236
rect 127452 187172 127453 187236
rect 127387 187171 127453 187172
rect 126835 78300 126901 78301
rect 126835 78236 126836 78300
rect 126900 78236 126901 78300
rect 126835 78235 126901 78236
rect 127390 78029 127450 187171
rect 127574 81973 127634 193699
rect 127755 192132 127821 192133
rect 127755 192068 127756 192132
rect 127820 192068 127821 192132
rect 127755 192067 127821 192068
rect 127758 140317 127818 192067
rect 127755 140316 127821 140317
rect 127755 140252 127756 140316
rect 127820 140252 127821 140316
rect 127755 140251 127821 140252
rect 129595 139364 129661 139365
rect 129595 139300 129596 139364
rect 129660 139300 129661 139364
rect 129595 139299 129661 139300
rect 127571 81972 127637 81973
rect 127571 81908 127572 81972
rect 127636 81908 127637 81972
rect 127571 81907 127637 81908
rect 129598 79117 129658 139299
rect 129595 79116 129661 79117
rect 129595 79052 129596 79116
rect 129660 79052 129661 79116
rect 129595 79051 129661 79052
rect 130334 78573 130394 194243
rect 131987 190908 132053 190909
rect 131987 190844 131988 190908
rect 132052 190844 132053 190908
rect 131987 190843 132053 190844
rect 130883 190772 130949 190773
rect 130883 190708 130884 190772
rect 130948 190708 130949 190772
rect 130883 190707 130949 190708
rect 130699 190636 130765 190637
rect 130699 190572 130700 190636
rect 130764 190572 130765 190636
rect 130699 190571 130765 190572
rect 130515 190500 130581 190501
rect 130515 190436 130516 190500
rect 130580 190436 130581 190500
rect 130515 190435 130581 190436
rect 130518 81157 130578 190435
rect 130702 81293 130762 190571
rect 130699 81292 130765 81293
rect 130699 81228 130700 81292
rect 130764 81228 130765 81292
rect 130699 81227 130765 81228
rect 130515 81156 130581 81157
rect 130515 81092 130516 81156
rect 130580 81092 130581 81156
rect 130515 81091 130581 81092
rect 130886 78709 130946 190707
rect 131619 185604 131685 185605
rect 131619 185540 131620 185604
rect 131684 185540 131685 185604
rect 131619 185539 131685 185540
rect 131622 79933 131682 185539
rect 131619 79932 131685 79933
rect 131619 79868 131620 79932
rect 131684 79868 131685 79932
rect 131619 79867 131685 79868
rect 130883 78708 130949 78709
rect 130883 78644 130884 78708
rect 130948 78644 130949 78708
rect 130883 78643 130949 78644
rect 130331 78572 130397 78573
rect 130331 78508 130332 78572
rect 130396 78508 130397 78572
rect 130331 78507 130397 78508
rect 127387 78028 127453 78029
rect 127387 77964 127388 78028
rect 127452 77964 127453 78028
rect 127387 77963 127453 77964
rect 124995 77348 125061 77349
rect 124995 77284 124996 77348
rect 125060 77284 125061 77348
rect 124995 77283 125061 77284
rect 123294 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 123914 52954
rect 123294 52634 123914 52718
rect 123294 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 123914 52634
rect 123294 16954 123914 52398
rect 123294 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 123914 16954
rect 123294 16634 123914 16718
rect 123294 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 123914 16634
rect 123294 -3226 123914 16398
rect 123294 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 123914 -3226
rect 123294 -3546 123914 -3462
rect 123294 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 123914 -3546
rect 123294 -7654 123914 -3782
rect 127794 57454 128414 78000
rect 131622 68237 131682 79867
rect 131990 77621 132050 190843
rect 132358 79389 132418 197779
rect 133091 186148 133157 186149
rect 133091 186084 133092 186148
rect 133156 186084 133157 186148
rect 133091 186083 133157 186084
rect 132907 185604 132973 185605
rect 132907 185540 132908 185604
rect 132972 185540 132973 185604
rect 132907 185539 132973 185540
rect 132910 79661 132970 185539
rect 133094 80613 133154 186083
rect 133459 185740 133525 185741
rect 133459 185676 133460 185740
rect 133524 185676 133525 185740
rect 133459 185675 133525 185676
rect 133275 185196 133341 185197
rect 133275 185132 133276 185196
rect 133340 185132 133341 185196
rect 133275 185131 133341 185132
rect 133091 80612 133157 80613
rect 133091 80548 133092 80612
rect 133156 80548 133157 80612
rect 133091 80547 133157 80548
rect 132907 79660 132973 79661
rect 132907 79596 132908 79660
rect 132972 79596 132973 79660
rect 132907 79595 132973 79596
rect 132355 79388 132421 79389
rect 132355 79324 132356 79388
rect 132420 79324 132421 79388
rect 132355 79323 132421 79324
rect 131987 77620 132053 77621
rect 131987 77556 131988 77620
rect 132052 77556 132053 77620
rect 131987 77555 132053 77556
rect 131619 68236 131685 68237
rect 131619 68172 131620 68236
rect 131684 68172 131685 68236
rect 131619 68171 131685 68172
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -4186 128414 20898
rect 127794 -4422 127826 -4186
rect 128062 -4422 128146 -4186
rect 128382 -4422 128414 -4186
rect 127794 -4506 128414 -4422
rect 127794 -4742 127826 -4506
rect 128062 -4742 128146 -4506
rect 128382 -4742 128414 -4506
rect 127794 -7654 128414 -4742
rect 132294 61954 132914 78000
rect 133094 65517 133154 80547
rect 133278 77893 133338 185131
rect 133462 80477 133522 185675
rect 133830 185333 133890 198323
rect 133827 185332 133893 185333
rect 133827 185268 133828 185332
rect 133892 185268 133893 185332
rect 133827 185267 133893 185268
rect 134198 89730 134258 198323
rect 134382 197709 134442 199819
rect 134750 197845 134810 199819
rect 135118 198389 135178 199819
rect 135486 199341 135546 199819
rect 135483 199340 135549 199341
rect 135483 199276 135484 199340
rect 135548 199276 135549 199340
rect 135483 199275 135549 199276
rect 135483 199204 135549 199205
rect 135483 199140 135484 199204
rect 135548 199140 135549 199204
rect 135483 199139 135549 199140
rect 135115 198388 135181 198389
rect 135115 198324 135116 198388
rect 135180 198324 135181 198388
rect 135115 198323 135181 198324
rect 134563 197844 134629 197845
rect 134563 197780 134564 197844
rect 134628 197780 134629 197844
rect 134563 197779 134629 197780
rect 134747 197844 134813 197845
rect 134747 197780 134748 197844
rect 134812 197780 134813 197844
rect 134747 197779 134813 197780
rect 135115 197844 135181 197845
rect 135115 197780 135116 197844
rect 135180 197780 135181 197844
rect 135115 197779 135181 197780
rect 134379 197708 134445 197709
rect 134379 197644 134380 197708
rect 134444 197644 134445 197708
rect 134379 197643 134445 197644
rect 134379 197572 134445 197573
rect 134379 197508 134380 197572
rect 134444 197508 134445 197572
rect 134379 197507 134445 197508
rect 134382 185605 134442 197507
rect 134566 186149 134626 197779
rect 135118 195125 135178 197779
rect 135115 195124 135181 195125
rect 135115 195060 135116 195124
rect 135180 195060 135181 195124
rect 135115 195059 135181 195060
rect 134563 186148 134629 186149
rect 134563 186084 134564 186148
rect 134628 186084 134629 186148
rect 134563 186083 134629 186084
rect 134931 185740 134997 185741
rect 134931 185676 134932 185740
rect 134996 185676 134997 185740
rect 134931 185675 134997 185676
rect 134379 185604 134445 185605
rect 134379 185540 134380 185604
rect 134444 185540 134445 185604
rect 134379 185539 134445 185540
rect 134563 185604 134629 185605
rect 134563 185540 134564 185604
rect 134628 185540 134629 185604
rect 134563 185539 134629 185540
rect 134198 89670 134442 89730
rect 133459 80476 133525 80477
rect 133459 80412 133460 80476
rect 133524 80412 133525 80476
rect 133459 80411 133525 80412
rect 133459 79932 133525 79933
rect 133459 79868 133460 79932
rect 133524 79868 133525 79932
rect 133459 79867 133525 79868
rect 134195 79932 134261 79933
rect 134195 79868 134196 79932
rect 134260 79868 134261 79932
rect 134195 79867 134261 79868
rect 133462 78573 133522 79867
rect 133827 79796 133893 79797
rect 133827 79732 133828 79796
rect 133892 79732 133893 79796
rect 133827 79731 133893 79732
rect 133643 79660 133709 79661
rect 133643 79596 133644 79660
rect 133708 79596 133709 79660
rect 133643 79595 133709 79596
rect 133459 78572 133525 78573
rect 133459 78508 133460 78572
rect 133524 78508 133525 78572
rect 133459 78507 133525 78508
rect 133275 77892 133341 77893
rect 133275 77828 133276 77892
rect 133340 77828 133341 77892
rect 133275 77827 133341 77828
rect 133091 65516 133157 65517
rect 133091 65452 133092 65516
rect 133156 65452 133157 65516
rect 133091 65451 133157 65452
rect 132294 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 132914 61954
rect 132294 61634 132914 61718
rect 132294 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 132914 61634
rect 132294 25954 132914 61398
rect 133646 33829 133706 79595
rect 133830 66877 133890 79731
rect 133827 66876 133893 66877
rect 133827 66812 133828 66876
rect 133892 66812 133893 66876
rect 133827 66811 133893 66812
rect 134198 52461 134258 79867
rect 134382 79797 134442 89670
rect 134379 79796 134445 79797
rect 134379 79732 134380 79796
rect 134444 79732 134445 79796
rect 134379 79731 134445 79732
rect 134566 78573 134626 185539
rect 134747 185468 134813 185469
rect 134747 185404 134748 185468
rect 134812 185404 134813 185468
rect 134747 185403 134813 185404
rect 134750 79933 134810 185403
rect 134934 80069 134994 185675
rect 135486 85590 135546 199139
rect 135854 197981 135914 199819
rect 136406 199613 136466 200091
rect 136955 199884 137021 199885
rect 136955 199820 136956 199884
rect 137020 199820 137021 199884
rect 136955 199819 137021 199820
rect 137139 199884 137205 199885
rect 137139 199820 137140 199884
rect 137204 199820 137205 199884
rect 137139 199819 137205 199820
rect 136403 199612 136469 199613
rect 136403 199548 136404 199612
rect 136468 199548 136469 199612
rect 136403 199547 136469 199548
rect 136219 198388 136285 198389
rect 136219 198324 136220 198388
rect 136284 198324 136285 198388
rect 136219 198323 136285 198324
rect 135851 197980 135917 197981
rect 135851 197916 135852 197980
rect 135916 197916 135917 197980
rect 135851 197915 135917 197916
rect 135851 197844 135917 197845
rect 135851 197780 135852 197844
rect 135916 197780 135917 197844
rect 135851 197779 135917 197780
rect 135118 85530 135546 85590
rect 135118 80069 135178 85530
rect 135854 84210 135914 197779
rect 136222 186557 136282 198323
rect 136219 186556 136285 186557
rect 136219 186492 136220 186556
rect 136284 186492 136285 186556
rect 136219 186491 136285 186492
rect 136035 186284 136101 186285
rect 136035 186220 136036 186284
rect 136100 186220 136101 186284
rect 136035 186219 136101 186220
rect 135670 84150 135914 84210
rect 134931 80068 134997 80069
rect 134931 80004 134932 80068
rect 134996 80004 134997 80068
rect 134931 80003 134997 80004
rect 135115 80068 135181 80069
rect 135115 80004 135116 80068
rect 135180 80004 135181 80068
rect 135115 80003 135181 80004
rect 134747 79932 134813 79933
rect 134747 79868 134748 79932
rect 134812 79868 134813 79932
rect 134747 79867 134813 79868
rect 135483 79932 135549 79933
rect 135483 79868 135484 79932
rect 135548 79868 135549 79932
rect 135483 79867 135549 79868
rect 134563 78572 134629 78573
rect 134563 78508 134564 78572
rect 134628 78508 134629 78572
rect 134563 78507 134629 78508
rect 134750 77893 134810 79867
rect 135486 79522 135546 79867
rect 135670 79797 135730 84150
rect 135667 79796 135733 79797
rect 135667 79732 135668 79796
rect 135732 79732 135733 79796
rect 136038 79794 136098 186219
rect 136958 185877 137018 199819
rect 137142 197981 137202 199819
rect 137139 197980 137205 197981
rect 137139 197916 137140 197980
rect 137204 197916 137205 197980
rect 137139 197915 137205 197916
rect 137139 186556 137205 186557
rect 137139 186492 137140 186556
rect 137204 186492 137205 186556
rect 137139 186491 137205 186492
rect 136955 185876 137021 185877
rect 136955 185812 136956 185876
rect 137020 185812 137021 185876
rect 136955 185811 137021 185812
rect 136219 183156 136285 183157
rect 136219 183092 136220 183156
rect 136284 183092 136285 183156
rect 136219 183091 136285 183092
rect 135667 79731 135733 79732
rect 135854 79734 136098 79794
rect 135854 79661 135914 79734
rect 135851 79660 135917 79661
rect 135851 79596 135852 79660
rect 135916 79596 135917 79660
rect 135851 79595 135917 79596
rect 136035 79660 136101 79661
rect 136035 79596 136036 79660
rect 136100 79596 136101 79660
rect 136035 79595 136101 79596
rect 135486 79462 135914 79522
rect 134747 77892 134813 77893
rect 134747 77828 134748 77892
rect 134812 77828 134813 77892
rect 134747 77827 134813 77828
rect 135483 76532 135549 76533
rect 135483 76468 135484 76532
rect 135548 76468 135549 76532
rect 135483 76467 135549 76468
rect 135299 73812 135365 73813
rect 135299 73748 135300 73812
rect 135364 73748 135365 73812
rect 135299 73747 135365 73748
rect 134195 52460 134261 52461
rect 134195 52396 134196 52460
rect 134260 52396 134261 52460
rect 134195 52395 134261 52396
rect 135302 46885 135362 73747
rect 135486 48245 135546 76467
rect 135667 73948 135733 73949
rect 135667 73884 135668 73948
rect 135732 73884 135733 73948
rect 135667 73883 135733 73884
rect 135670 49605 135730 73883
rect 135854 64837 135914 79462
rect 136038 77893 136098 79595
rect 136222 78573 136282 183091
rect 136403 79932 136469 79933
rect 136403 79868 136404 79932
rect 136468 79868 136469 79932
rect 136403 79867 136469 79868
rect 136955 79932 137021 79933
rect 136955 79868 136956 79932
rect 137020 79868 137021 79932
rect 136955 79867 137021 79868
rect 136219 78572 136285 78573
rect 136219 78508 136220 78572
rect 136284 78508 136285 78572
rect 136219 78507 136285 78508
rect 136035 77892 136101 77893
rect 136035 77828 136036 77892
rect 136100 77828 136101 77892
rect 136035 77827 136101 77828
rect 136406 77621 136466 79867
rect 136958 78573 137018 79867
rect 137142 79661 137202 186491
rect 137510 79933 137570 200091
rect 137691 199884 137757 199885
rect 137691 199820 137692 199884
rect 137756 199820 137757 199884
rect 137691 199819 137757 199820
rect 137694 186690 137754 199819
rect 137878 199613 137938 200227
rect 139531 200156 139597 200157
rect 139531 200092 139532 200156
rect 139596 200092 139597 200156
rect 139531 200091 139597 200092
rect 140819 200156 140885 200157
rect 140819 200092 140820 200156
rect 140884 200092 140885 200156
rect 140819 200091 140885 200092
rect 145419 200156 145485 200157
rect 145419 200092 145420 200156
rect 145484 200092 145485 200156
rect 145419 200091 145485 200092
rect 138059 199884 138125 199885
rect 138059 199820 138060 199884
rect 138124 199820 138125 199884
rect 138059 199819 138125 199820
rect 138611 199884 138677 199885
rect 138611 199820 138612 199884
rect 138676 199820 138677 199884
rect 138611 199819 138677 199820
rect 138795 199884 138861 199885
rect 138795 199820 138796 199884
rect 138860 199820 138861 199884
rect 138795 199819 138861 199820
rect 139347 199884 139413 199885
rect 139347 199820 139348 199884
rect 139412 199820 139413 199884
rect 139347 199819 139413 199820
rect 137875 199612 137941 199613
rect 137875 199548 137876 199612
rect 137940 199548 137941 199612
rect 137875 199547 137941 199548
rect 138062 192405 138122 199819
rect 138059 192404 138125 192405
rect 138059 192340 138060 192404
rect 138124 192340 138125 192404
rect 138059 192339 138125 192340
rect 137694 186630 137938 186690
rect 137691 185604 137757 185605
rect 137691 185540 137692 185604
rect 137756 185540 137757 185604
rect 137691 185539 137757 185540
rect 137507 79932 137573 79933
rect 137507 79868 137508 79932
rect 137572 79868 137573 79932
rect 137507 79867 137573 79868
rect 137694 79661 137754 185539
rect 137878 80069 137938 186630
rect 138427 177172 138493 177173
rect 138427 177108 138428 177172
rect 138492 177108 138493 177172
rect 138427 177107 138493 177108
rect 137875 80068 137941 80069
rect 137875 80004 137876 80068
rect 137940 80004 137941 80068
rect 137875 80003 137941 80004
rect 138059 79932 138125 79933
rect 138059 79930 138060 79932
rect 137878 79870 138060 79930
rect 137139 79660 137205 79661
rect 137139 79596 137140 79660
rect 137204 79596 137205 79660
rect 137139 79595 137205 79596
rect 137691 79660 137757 79661
rect 137691 79596 137692 79660
rect 137756 79596 137757 79660
rect 137691 79595 137757 79596
rect 136587 78572 136653 78573
rect 136587 78508 136588 78572
rect 136652 78508 136653 78572
rect 136587 78507 136653 78508
rect 136955 78572 137021 78573
rect 136955 78508 136956 78572
rect 137020 78508 137021 78572
rect 136955 78507 137021 78508
rect 136403 77620 136469 77621
rect 136403 77556 136404 77620
rect 136468 77556 136469 77620
rect 136403 77555 136469 77556
rect 135851 64836 135917 64837
rect 135851 64772 135852 64836
rect 135916 64772 135917 64836
rect 135851 64771 135917 64772
rect 136590 55181 136650 78507
rect 136794 66454 137414 78000
rect 137507 77620 137573 77621
rect 137507 77556 137508 77620
rect 137572 77556 137573 77620
rect 137507 77555 137573 77556
rect 137510 67013 137570 77555
rect 137694 77485 137754 79595
rect 137878 77893 137938 79870
rect 138059 79868 138060 79870
rect 138124 79868 138125 79932
rect 138430 79930 138490 177107
rect 138614 86970 138674 199819
rect 138798 194853 138858 199819
rect 139350 196893 139410 199819
rect 139347 196892 139413 196893
rect 139347 196828 139348 196892
rect 139412 196828 139413 196892
rect 139347 196827 139413 196828
rect 138795 194852 138861 194853
rect 138795 194788 138796 194852
rect 138860 194788 138861 194852
rect 138795 194787 138861 194788
rect 139534 186285 139594 200091
rect 139715 199884 139781 199885
rect 139715 199820 139716 199884
rect 139780 199820 139781 199884
rect 139715 199819 139781 199820
rect 140083 199884 140149 199885
rect 140083 199820 140084 199884
rect 140148 199820 140149 199884
rect 140083 199819 140149 199820
rect 140451 199884 140517 199885
rect 140451 199820 140452 199884
rect 140516 199820 140517 199884
rect 140451 199819 140517 199820
rect 139718 189821 139778 199819
rect 140086 199205 140146 199819
rect 140083 199204 140149 199205
rect 140083 199140 140084 199204
rect 140148 199140 140149 199204
rect 140083 199139 140149 199140
rect 140454 198525 140514 199819
rect 140451 198524 140517 198525
rect 140451 198460 140452 198524
rect 140516 198460 140517 198524
rect 140451 198459 140517 198460
rect 140451 198116 140517 198117
rect 140451 198052 140452 198116
rect 140516 198052 140517 198116
rect 140451 198051 140517 198052
rect 139715 189820 139781 189821
rect 139715 189756 139716 189820
rect 139780 189756 139781 189820
rect 139715 189755 139781 189756
rect 139163 186284 139229 186285
rect 139163 186220 139164 186284
rect 139228 186220 139229 186284
rect 139163 186219 139229 186220
rect 139531 186284 139597 186285
rect 139531 186220 139532 186284
rect 139596 186220 139597 186284
rect 139531 186219 139597 186220
rect 140267 186284 140333 186285
rect 140267 186220 140268 186284
rect 140332 186220 140333 186284
rect 140267 186219 140333 186220
rect 138979 174996 139045 174997
rect 138979 174932 138980 174996
rect 139044 174932 139045 174996
rect 138979 174931 139045 174932
rect 138614 86910 138858 86970
rect 138611 80476 138677 80477
rect 138611 80412 138612 80476
rect 138676 80412 138677 80476
rect 138611 80411 138677 80412
rect 138614 80205 138674 80411
rect 138611 80204 138677 80205
rect 138611 80140 138612 80204
rect 138676 80140 138677 80204
rect 138611 80139 138677 80140
rect 138798 80069 138858 86910
rect 138795 80068 138861 80069
rect 138795 80004 138796 80068
rect 138860 80004 138861 80068
rect 138795 80003 138861 80004
rect 138982 79933 139042 174931
rect 138979 79932 139045 79933
rect 138430 79870 138858 79930
rect 138059 79867 138125 79868
rect 138798 79797 138858 79870
rect 138979 79868 138980 79932
rect 139044 79868 139045 79932
rect 138979 79867 139045 79868
rect 138427 79796 138493 79797
rect 138427 79732 138428 79796
rect 138492 79732 138493 79796
rect 138427 79731 138493 79732
rect 138795 79796 138861 79797
rect 138795 79732 138796 79796
rect 138860 79732 138861 79796
rect 138795 79731 138861 79732
rect 138243 79524 138309 79525
rect 138243 79460 138244 79524
rect 138308 79460 138309 79524
rect 138243 79459 138309 79460
rect 138246 79250 138306 79459
rect 138062 79190 138306 79250
rect 138062 78981 138122 79190
rect 138059 78980 138125 78981
rect 138059 78916 138060 78980
rect 138124 78916 138125 78980
rect 138059 78915 138125 78916
rect 138059 78572 138125 78573
rect 138059 78508 138060 78572
rect 138124 78508 138125 78572
rect 138059 78507 138125 78508
rect 137875 77892 137941 77893
rect 137875 77828 137876 77892
rect 137940 77828 137941 77892
rect 137875 77827 137941 77828
rect 137691 77484 137757 77485
rect 137691 77420 137692 77484
rect 137756 77420 137757 77484
rect 137691 77419 137757 77420
rect 137507 67012 137573 67013
rect 137507 66948 137508 67012
rect 137572 66948 137573 67012
rect 137507 66947 137573 66948
rect 136794 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 137414 66454
rect 136794 66134 137414 66218
rect 136794 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 137414 66134
rect 136587 55180 136653 55181
rect 136587 55116 136588 55180
rect 136652 55116 136653 55180
rect 136587 55115 136653 55116
rect 135667 49604 135733 49605
rect 135667 49540 135668 49604
rect 135732 49540 135733 49604
rect 135667 49539 135733 49540
rect 135483 48244 135549 48245
rect 135483 48180 135484 48244
rect 135548 48180 135549 48244
rect 135483 48179 135549 48180
rect 135299 46884 135365 46885
rect 135299 46820 135300 46884
rect 135364 46820 135365 46884
rect 135299 46819 135365 46820
rect 133643 33828 133709 33829
rect 133643 33764 133644 33828
rect 133708 33764 133709 33828
rect 133643 33763 133709 33764
rect 132294 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 132914 25954
rect 132294 25634 132914 25718
rect 132294 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 132914 25634
rect 132294 -5146 132914 25398
rect 132294 -5382 132326 -5146
rect 132562 -5382 132646 -5146
rect 132882 -5382 132914 -5146
rect 132294 -5466 132914 -5382
rect 132294 -5702 132326 -5466
rect 132562 -5702 132646 -5466
rect 132882 -5702 132914 -5466
rect 132294 -7654 132914 -5702
rect 136794 30454 137414 65898
rect 138062 57901 138122 78507
rect 138243 77484 138309 77485
rect 138243 77420 138244 77484
rect 138308 77420 138309 77484
rect 138243 77419 138309 77420
rect 138246 60621 138306 77419
rect 138430 63341 138490 79731
rect 138611 78300 138677 78301
rect 138611 78236 138612 78300
rect 138676 78236 138677 78300
rect 138611 78235 138677 78236
rect 138614 67557 138674 78235
rect 138982 77893 139042 79867
rect 139166 78981 139226 186219
rect 140083 179348 140149 179349
rect 140083 179284 140084 179348
rect 140148 179284 140149 179348
rect 140083 179283 140149 179284
rect 139568 115954 139888 115986
rect 139568 115718 139610 115954
rect 139846 115718 139888 115954
rect 139568 115634 139888 115718
rect 139568 115398 139610 115634
rect 139846 115398 139888 115634
rect 139568 115366 139888 115398
rect 139531 79932 139597 79933
rect 139531 79868 139532 79932
rect 139596 79868 139597 79932
rect 139531 79867 139597 79868
rect 139899 79932 139965 79933
rect 139899 79868 139900 79932
rect 139964 79868 139965 79932
rect 139899 79867 139965 79868
rect 139163 78980 139229 78981
rect 139163 78916 139164 78980
rect 139228 78916 139229 78980
rect 139163 78915 139229 78916
rect 138979 77892 139045 77893
rect 138979 77828 138980 77892
rect 139044 77828 139045 77892
rect 138979 77827 139045 77828
rect 138611 67556 138677 67557
rect 138611 67492 138612 67556
rect 138676 67492 138677 67556
rect 138611 67491 138677 67492
rect 139534 63477 139594 79867
rect 139715 77892 139781 77893
rect 139715 77828 139716 77892
rect 139780 77828 139781 77892
rect 139715 77827 139781 77828
rect 139718 66061 139778 77827
rect 139902 66197 139962 79867
rect 140086 79797 140146 179283
rect 140270 80069 140330 186219
rect 140454 80069 140514 198051
rect 140635 185604 140701 185605
rect 140635 185540 140636 185604
rect 140700 185540 140701 185604
rect 140635 185539 140701 185540
rect 140267 80068 140333 80069
rect 140267 80004 140268 80068
rect 140332 80004 140333 80068
rect 140267 80003 140333 80004
rect 140451 80068 140517 80069
rect 140451 80004 140452 80068
rect 140516 80004 140517 80068
rect 140451 80003 140517 80004
rect 140638 79933 140698 185539
rect 140822 81429 140882 200091
rect 141003 199884 141069 199885
rect 141003 199820 141004 199884
rect 141068 199820 141069 199884
rect 141003 199819 141069 199820
rect 141187 199884 141253 199885
rect 141187 199820 141188 199884
rect 141252 199820 141253 199884
rect 141187 199819 141253 199820
rect 142475 199884 142541 199885
rect 142475 199820 142476 199884
rect 142540 199820 142541 199884
rect 142475 199819 142541 199820
rect 143027 199884 143093 199885
rect 143027 199820 143028 199884
rect 143092 199820 143093 199884
rect 143027 199819 143093 199820
rect 144683 199884 144749 199885
rect 144683 199820 144684 199884
rect 144748 199820 144749 199884
rect 144683 199819 144749 199820
rect 145051 199884 145117 199885
rect 145051 199820 145052 199884
rect 145116 199820 145117 199884
rect 145051 199819 145117 199820
rect 141006 195397 141066 199819
rect 141190 198389 141250 199819
rect 141187 198388 141253 198389
rect 141187 198324 141188 198388
rect 141252 198324 141253 198388
rect 141187 198323 141253 198324
rect 142478 198117 142538 199819
rect 142659 199748 142725 199749
rect 142659 199684 142660 199748
rect 142724 199684 142725 199748
rect 142659 199683 142725 199684
rect 142662 198253 142722 199683
rect 142659 198252 142725 198253
rect 142659 198188 142660 198252
rect 142724 198188 142725 198252
rect 142659 198187 142725 198188
rect 142291 198116 142357 198117
rect 142291 198052 142292 198116
rect 142356 198052 142357 198116
rect 142291 198051 142357 198052
rect 142475 198116 142541 198117
rect 142475 198052 142476 198116
rect 142540 198052 142541 198116
rect 142475 198051 142541 198052
rect 141003 195396 141069 195397
rect 141003 195332 141004 195396
rect 141068 195332 141069 195396
rect 141003 195331 141069 195332
rect 141003 185604 141069 185605
rect 141003 185540 141004 185604
rect 141068 185540 141069 185604
rect 141003 185539 141069 185540
rect 140819 81428 140885 81429
rect 140819 81364 140820 81428
rect 140884 81364 140885 81428
rect 140819 81363 140885 81364
rect 140819 80340 140885 80341
rect 140819 80276 140820 80340
rect 140884 80276 140885 80340
rect 140819 80275 140885 80276
rect 140635 79932 140701 79933
rect 140635 79868 140636 79932
rect 140700 79868 140701 79932
rect 140635 79867 140701 79868
rect 140083 79796 140149 79797
rect 140083 79732 140084 79796
rect 140148 79732 140149 79796
rect 140083 79731 140149 79732
rect 140638 78981 140698 79867
rect 140822 79797 140882 80275
rect 140819 79796 140885 79797
rect 140819 79732 140820 79796
rect 140884 79732 140885 79796
rect 140819 79731 140885 79732
rect 140635 78980 140701 78981
rect 140635 78916 140636 78980
rect 140700 78916 140701 78980
rect 140635 78915 140701 78916
rect 141006 78573 141066 185539
rect 141294 178954 141914 198000
rect 142107 185468 142173 185469
rect 142107 185404 142108 185468
rect 142172 185404 142173 185468
rect 142107 185403 142173 185404
rect 141294 178718 141326 178954
rect 141562 178718 141646 178954
rect 141882 178718 141914 178954
rect 141294 178634 141914 178718
rect 141294 178398 141326 178634
rect 141562 178398 141646 178634
rect 141882 178398 141914 178634
rect 141294 142954 141914 178398
rect 142110 171053 142170 185403
rect 142107 171052 142173 171053
rect 142107 170988 142108 171052
rect 142172 170988 142173 171052
rect 142107 170987 142173 170988
rect 142107 161668 142173 161669
rect 142107 161604 142108 161668
rect 142172 161604 142173 161668
rect 142107 161603 142173 161604
rect 142110 161397 142170 161603
rect 142107 161396 142173 161397
rect 142107 161332 142108 161396
rect 142172 161332 142173 161396
rect 142107 161331 142173 161332
rect 142107 152012 142173 152013
rect 142107 151948 142108 152012
rect 142172 151948 142173 152012
rect 142107 151947 142173 151948
rect 142110 151741 142170 151947
rect 142107 151740 142173 151741
rect 142107 151676 142108 151740
rect 142172 151676 142173 151740
rect 142107 151675 142173 151676
rect 142294 146981 142354 198051
rect 142659 185876 142725 185877
rect 142659 185812 142660 185876
rect 142724 185812 142725 185876
rect 142659 185811 142725 185812
rect 142475 147660 142541 147661
rect 142475 147596 142476 147660
rect 142540 147596 142541 147660
rect 142475 147595 142541 147596
rect 142291 146980 142357 146981
rect 142291 146916 142292 146980
rect 142356 146916 142357 146980
rect 142291 146915 142357 146916
rect 141294 142718 141326 142954
rect 141562 142718 141646 142954
rect 141882 142718 141914 142954
rect 141294 142634 141914 142718
rect 141294 142398 141326 142634
rect 141562 142398 141646 142634
rect 141882 142398 141914 142634
rect 141294 142000 141914 142398
rect 142291 142356 142357 142357
rect 142291 142292 142292 142356
rect 142356 142292 142357 142356
rect 142291 142291 142357 142292
rect 142294 142170 142354 142291
rect 142110 142110 142354 142170
rect 142110 141810 142170 142110
rect 141926 141750 142170 141810
rect 141371 141676 141437 141677
rect 141371 141612 141372 141676
rect 141436 141612 141437 141676
rect 141371 141611 141437 141612
rect 141374 78981 141434 141611
rect 141555 141268 141621 141269
rect 141555 141204 141556 141268
rect 141620 141204 141621 141268
rect 141555 141203 141621 141204
rect 141558 79933 141618 141203
rect 141926 89730 141986 141750
rect 141926 89670 142170 89730
rect 142110 84210 142170 89670
rect 141926 84150 142170 84210
rect 141739 81428 141805 81429
rect 141739 81364 141740 81428
rect 141804 81364 141805 81428
rect 141739 81363 141805 81364
rect 141742 79933 141802 81363
rect 141926 80341 141986 84150
rect 141923 80340 141989 80341
rect 141923 80276 141924 80340
rect 141988 80276 141989 80340
rect 141923 80275 141989 80276
rect 141555 79932 141621 79933
rect 141555 79868 141556 79932
rect 141620 79868 141621 79932
rect 141555 79867 141621 79868
rect 141739 79932 141805 79933
rect 141739 79868 141740 79932
rect 141804 79868 141805 79932
rect 141739 79867 141805 79868
rect 141371 78980 141437 78981
rect 141371 78916 141372 78980
rect 141436 78916 141437 78980
rect 141371 78915 141437 78916
rect 141003 78572 141069 78573
rect 141003 78508 141004 78572
rect 141068 78508 141069 78572
rect 141003 78507 141069 78508
rect 141742 78437 141802 79867
rect 142478 78981 142538 147595
rect 142662 141949 142722 185811
rect 143030 185605 143090 199819
rect 144686 195805 144746 199819
rect 145054 199205 145114 199819
rect 145051 199204 145117 199205
rect 145051 199140 145052 199204
rect 145116 199140 145117 199204
rect 145051 199139 145117 199140
rect 144683 195804 144749 195805
rect 144683 195740 144684 195804
rect 144748 195740 144749 195804
rect 144683 195739 144749 195740
rect 144315 190092 144381 190093
rect 144315 190028 144316 190092
rect 144380 190028 144381 190092
rect 144315 190027 144381 190028
rect 143027 185604 143093 185605
rect 143027 185540 143028 185604
rect 143092 185540 143093 185604
rect 143027 185539 143093 185540
rect 143763 185332 143829 185333
rect 143763 185268 143764 185332
rect 143828 185268 143829 185332
rect 143763 185267 143829 185268
rect 143766 148477 143826 185267
rect 143763 148476 143829 148477
rect 143763 148412 143764 148476
rect 143828 148412 143829 148476
rect 143763 148411 143829 148412
rect 142659 141948 142725 141949
rect 142659 141884 142660 141948
rect 142724 141884 142725 141948
rect 142659 141883 142725 141884
rect 143027 81292 143093 81293
rect 143027 81228 143028 81292
rect 143092 81228 143093 81292
rect 143027 81227 143093 81228
rect 142475 78980 142541 78981
rect 142475 78916 142476 78980
rect 142540 78916 142541 78980
rect 142475 78915 142541 78916
rect 143030 78573 143090 81227
rect 143395 81156 143461 81157
rect 143395 81092 143396 81156
rect 143460 81092 143461 81156
rect 143395 81091 143461 81092
rect 143211 81020 143277 81021
rect 143211 80956 143212 81020
rect 143276 80956 143277 81020
rect 143211 80955 143277 80956
rect 143214 79933 143274 80955
rect 143211 79932 143277 79933
rect 143211 79868 143212 79932
rect 143276 79868 143277 79932
rect 143211 79867 143277 79868
rect 143027 78572 143093 78573
rect 143027 78508 143028 78572
rect 143092 78508 143093 78572
rect 143027 78507 143093 78508
rect 143214 78437 143274 79867
rect 143398 78981 143458 81091
rect 143947 79932 144013 79933
rect 143947 79868 143948 79932
rect 144012 79868 144013 79932
rect 143947 79867 144013 79868
rect 143395 78980 143461 78981
rect 143395 78916 143396 78980
rect 143460 78916 143461 78980
rect 143395 78915 143461 78916
rect 141739 78436 141805 78437
rect 141739 78372 141740 78436
rect 141804 78372 141805 78436
rect 141739 78371 141805 78372
rect 143211 78436 143277 78437
rect 143211 78372 143212 78436
rect 143276 78372 143277 78436
rect 143211 78371 143277 78372
rect 140083 77892 140149 77893
rect 140083 77828 140084 77892
rect 140148 77828 140149 77892
rect 140083 77827 140149 77828
rect 140819 77892 140885 77893
rect 140819 77828 140820 77892
rect 140884 77828 140885 77892
rect 140819 77827 140885 77828
rect 139899 66196 139965 66197
rect 139899 66132 139900 66196
rect 139964 66132 139965 66196
rect 139899 66131 139965 66132
rect 139715 66060 139781 66061
rect 139715 65996 139716 66060
rect 139780 65996 139781 66060
rect 139715 65995 139781 65996
rect 139531 63476 139597 63477
rect 139531 63412 139532 63476
rect 139596 63412 139597 63476
rect 139531 63411 139597 63412
rect 138427 63340 138493 63341
rect 138427 63276 138428 63340
rect 138492 63276 138493 63340
rect 138427 63275 138493 63276
rect 138243 60620 138309 60621
rect 138243 60556 138244 60620
rect 138308 60556 138309 60620
rect 138243 60555 138309 60556
rect 140086 59261 140146 77827
rect 140822 68373 140882 77827
rect 141294 70954 141914 78000
rect 142291 77756 142357 77757
rect 142291 77692 142292 77756
rect 142356 77692 142357 77756
rect 142291 77691 142357 77692
rect 142294 72589 142354 77691
rect 143950 74357 144010 79867
rect 144131 79796 144197 79797
rect 144131 79732 144132 79796
rect 144196 79732 144197 79796
rect 144131 79731 144197 79732
rect 143947 74356 144013 74357
rect 143947 74292 143948 74356
rect 144012 74292 144013 74356
rect 143947 74291 144013 74292
rect 144134 74085 144194 79731
rect 144318 77349 144378 190027
rect 145235 185468 145301 185469
rect 145235 185404 145236 185468
rect 145300 185404 145301 185468
rect 145235 185403 145301 185404
rect 145238 152421 145298 185403
rect 145235 152420 145301 152421
rect 145235 152356 145236 152420
rect 145300 152356 145301 152420
rect 145235 152355 145301 152356
rect 145422 81021 145482 200091
rect 146523 199884 146589 199885
rect 146523 199820 146524 199884
rect 146588 199820 146589 199884
rect 146523 199819 146589 199820
rect 146707 199884 146773 199885
rect 146707 199820 146708 199884
rect 146772 199820 146773 199884
rect 146707 199819 146773 199820
rect 147075 199884 147141 199885
rect 147075 199820 147076 199884
rect 147140 199820 147141 199884
rect 147075 199819 147141 199820
rect 148179 199884 148245 199885
rect 148179 199820 148180 199884
rect 148244 199820 148245 199884
rect 148179 199819 148245 199820
rect 149283 199884 149349 199885
rect 149283 199820 149284 199884
rect 149348 199820 149349 199884
rect 149283 199819 149349 199820
rect 149651 199884 149717 199885
rect 149651 199820 149652 199884
rect 149716 199820 149717 199884
rect 149651 199819 149717 199820
rect 150939 199884 151005 199885
rect 150939 199820 150940 199884
rect 151004 199820 151005 199884
rect 152595 199884 152661 199885
rect 152595 199882 152596 199884
rect 150939 199819 151005 199820
rect 152414 199822 152596 199882
rect 145794 183454 146414 198000
rect 145794 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 146414 183454
rect 145794 183134 146414 183218
rect 145794 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 146414 183134
rect 145603 179076 145669 179077
rect 145603 179012 145604 179076
rect 145668 179012 145669 179076
rect 145603 179011 145669 179012
rect 145419 81020 145485 81021
rect 145419 80956 145420 81020
rect 145484 80956 145485 81020
rect 145419 80955 145485 80956
rect 145419 79932 145485 79933
rect 145419 79868 145420 79932
rect 145484 79868 145485 79932
rect 145419 79867 145485 79868
rect 145051 77756 145117 77757
rect 145051 77692 145052 77756
rect 145116 77692 145117 77756
rect 145051 77691 145117 77692
rect 144315 77348 144381 77349
rect 144315 77284 144316 77348
rect 144380 77284 144381 77348
rect 144315 77283 144381 77284
rect 144131 74084 144197 74085
rect 144131 74020 144132 74084
rect 144196 74020 144197 74084
rect 144131 74019 144197 74020
rect 142291 72588 142357 72589
rect 142291 72524 142292 72588
rect 142356 72524 142357 72588
rect 142291 72523 142357 72524
rect 141294 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 141914 70954
rect 141294 70634 141914 70718
rect 141294 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 141914 70634
rect 140819 68372 140885 68373
rect 140819 68308 140820 68372
rect 140884 68308 140885 68372
rect 140819 68307 140885 68308
rect 140083 59260 140149 59261
rect 140083 59196 140084 59260
rect 140148 59196 140149 59260
rect 140083 59195 140149 59196
rect 138059 57900 138125 57901
rect 138059 57836 138060 57900
rect 138124 57836 138125 57900
rect 138059 57835 138125 57836
rect 136794 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 137414 30454
rect 136794 30134 137414 30218
rect 136794 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 137414 30134
rect 136794 -6106 137414 29898
rect 136794 -6342 136826 -6106
rect 137062 -6342 137146 -6106
rect 137382 -6342 137414 -6106
rect 136794 -6426 137414 -6342
rect 136794 -6662 136826 -6426
rect 137062 -6662 137146 -6426
rect 137382 -6662 137414 -6426
rect 136794 -7654 137414 -6662
rect 141294 34954 141914 70398
rect 141294 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 141914 34954
rect 141294 34634 141914 34718
rect 141294 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 141914 34634
rect 141294 -7066 141914 34398
rect 144134 15877 144194 74019
rect 145054 71365 145114 77691
rect 145422 74550 145482 79867
rect 145606 77621 145666 179011
rect 145794 147454 146414 182898
rect 146526 179349 146586 199819
rect 146710 187373 146770 199819
rect 146891 199748 146957 199749
rect 146891 199684 146892 199748
rect 146956 199684 146957 199748
rect 146891 199683 146957 199684
rect 146894 199341 146954 199683
rect 146891 199340 146957 199341
rect 146891 199276 146892 199340
rect 146956 199276 146957 199340
rect 146891 199275 146957 199276
rect 146707 187372 146773 187373
rect 146707 187308 146708 187372
rect 146772 187308 146773 187372
rect 146707 187307 146773 187308
rect 146891 186284 146957 186285
rect 146891 186220 146892 186284
rect 146956 186220 146957 186284
rect 146891 186219 146957 186220
rect 146523 179348 146589 179349
rect 146523 179284 146524 179348
rect 146588 179284 146589 179348
rect 146523 179283 146589 179284
rect 145794 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 146414 147454
rect 145794 147134 146414 147218
rect 145794 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 146414 147134
rect 145794 142000 146414 146898
rect 145787 81972 145853 81973
rect 145787 81908 145788 81972
rect 145852 81908 145853 81972
rect 145787 81907 145853 81908
rect 145790 79797 145850 81907
rect 146523 80884 146589 80885
rect 146523 80820 146524 80884
rect 146588 80820 146589 80884
rect 146523 80819 146589 80820
rect 146526 79933 146586 80819
rect 146707 80748 146773 80749
rect 146707 80684 146708 80748
rect 146772 80684 146773 80748
rect 146707 80683 146773 80684
rect 146523 79932 146589 79933
rect 146523 79868 146524 79932
rect 146588 79868 146589 79932
rect 146523 79867 146589 79868
rect 146710 79797 146770 80683
rect 146894 79933 146954 186219
rect 147078 185741 147138 199819
rect 148182 198525 148242 199819
rect 148179 198524 148245 198525
rect 148179 198460 148180 198524
rect 148244 198460 148245 198524
rect 148179 198459 148245 198460
rect 149286 191181 149346 199819
rect 149467 192676 149533 192677
rect 149467 192612 149468 192676
rect 149532 192612 149533 192676
rect 149467 192611 149533 192612
rect 149283 191180 149349 191181
rect 149283 191116 149284 191180
rect 149348 191116 149349 191180
rect 149283 191115 149349 191116
rect 148547 186692 148613 186693
rect 148547 186628 148548 186692
rect 148612 186628 148613 186692
rect 148547 186627 148613 186628
rect 148179 186284 148245 186285
rect 148179 186220 148180 186284
rect 148244 186220 148245 186284
rect 148179 186219 148245 186220
rect 147075 185740 147141 185741
rect 147075 185676 147076 185740
rect 147140 185676 147141 185740
rect 147075 185675 147141 185676
rect 147075 181932 147141 181933
rect 147075 181868 147076 181932
rect 147140 181868 147141 181932
rect 147075 181867 147141 181868
rect 146891 79932 146957 79933
rect 146891 79868 146892 79932
rect 146956 79868 146957 79932
rect 146891 79867 146957 79868
rect 145787 79796 145853 79797
rect 145787 79732 145788 79796
rect 145852 79732 145853 79796
rect 145787 79731 145853 79732
rect 146707 79796 146773 79797
rect 146707 79732 146708 79796
rect 146772 79732 146773 79796
rect 146707 79731 146773 79732
rect 147078 79525 147138 181867
rect 147443 181796 147509 181797
rect 147443 181732 147444 181796
rect 147508 181732 147509 181796
rect 147443 181731 147509 181732
rect 147446 80613 147506 181731
rect 147627 81020 147693 81021
rect 147627 80956 147628 81020
rect 147692 80956 147693 81020
rect 147627 80955 147693 80956
rect 147443 80612 147509 80613
rect 147443 80548 147444 80612
rect 147508 80548 147509 80612
rect 147443 80547 147509 80548
rect 147259 80476 147325 80477
rect 147259 80412 147260 80476
rect 147324 80412 147325 80476
rect 147259 80411 147325 80412
rect 147262 79797 147322 80411
rect 147443 79932 147509 79933
rect 147443 79868 147444 79932
rect 147508 79868 147509 79932
rect 147443 79867 147509 79868
rect 147259 79796 147325 79797
rect 147259 79732 147260 79796
rect 147324 79732 147325 79796
rect 147259 79731 147325 79732
rect 147075 79524 147141 79525
rect 147075 79460 147076 79524
rect 147140 79460 147141 79524
rect 147075 79459 147141 79460
rect 145603 77620 145669 77621
rect 145603 77556 145604 77620
rect 145668 77556 145669 77620
rect 145603 77555 145669 77556
rect 145794 75454 146414 78000
rect 147075 77892 147141 77893
rect 147075 77828 147076 77892
rect 147140 77828 147141 77892
rect 147075 77827 147141 77828
rect 146891 77756 146957 77757
rect 146891 77692 146892 77756
rect 146956 77692 146957 77756
rect 146891 77691 146957 77692
rect 146894 77213 146954 77691
rect 146891 77212 146957 77213
rect 146891 77148 146892 77212
rect 146956 77148 146957 77212
rect 146891 77147 146957 77148
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145422 74490 145666 74550
rect 145051 71364 145117 71365
rect 145051 71300 145052 71364
rect 145116 71300 145117 71364
rect 145051 71299 145117 71300
rect 144315 70548 144381 70549
rect 144315 70484 144316 70548
rect 144380 70484 144381 70548
rect 144315 70483 144381 70484
rect 144131 15876 144197 15877
rect 144131 15812 144132 15876
rect 144196 15812 144197 15876
rect 144131 15811 144197 15812
rect 144318 11661 144378 70483
rect 144499 68780 144565 68781
rect 144499 68716 144500 68780
rect 144564 68716 144565 68780
rect 144499 68715 144565 68716
rect 144502 26893 144562 68715
rect 144683 68508 144749 68509
rect 144683 68444 144684 68508
rect 144748 68444 144749 68508
rect 144683 68443 144749 68444
rect 144686 33829 144746 68443
rect 145054 64890 145114 71299
rect 145606 71229 145666 74490
rect 145603 71228 145669 71229
rect 145603 71164 145604 71228
rect 145668 71164 145669 71228
rect 145603 71163 145669 71164
rect 145054 64830 145482 64890
rect 144683 33828 144749 33829
rect 144683 33764 144684 33828
rect 144748 33764 144749 33828
rect 144683 33763 144749 33764
rect 144499 26892 144565 26893
rect 144499 26828 144500 26892
rect 144564 26828 144565 26892
rect 144499 26827 144565 26828
rect 145422 17237 145482 64830
rect 145606 37909 145666 71163
rect 145794 39454 146414 74898
rect 146894 66877 146954 77147
rect 147078 75717 147138 77827
rect 147075 75716 147141 75717
rect 147075 75652 147076 75716
rect 147140 75652 147141 75716
rect 147075 75651 147141 75652
rect 147078 68237 147138 75651
rect 147075 68236 147141 68237
rect 147075 68172 147076 68236
rect 147140 68172 147141 68236
rect 147075 68171 147141 68172
rect 146891 66876 146957 66877
rect 146891 66812 146892 66876
rect 146956 66812 146957 66876
rect 146891 66811 146957 66812
rect 147262 59941 147322 79731
rect 147446 79525 147506 79867
rect 147630 79525 147690 80955
rect 147811 79932 147877 79933
rect 147811 79868 147812 79932
rect 147876 79868 147877 79932
rect 147811 79867 147877 79868
rect 147443 79524 147509 79525
rect 147443 79460 147444 79524
rect 147508 79460 147509 79524
rect 147443 79459 147509 79460
rect 147627 79524 147693 79525
rect 147627 79460 147628 79524
rect 147692 79460 147693 79524
rect 147627 79459 147693 79460
rect 147259 59940 147325 59941
rect 147259 59876 147260 59940
rect 147324 59876 147325 59940
rect 147259 59875 147325 59876
rect 147446 47565 147506 79459
rect 147814 77757 147874 79867
rect 147995 79796 148061 79797
rect 147995 79732 147996 79796
rect 148060 79732 148061 79796
rect 147995 79731 148061 79732
rect 147998 77893 148058 79731
rect 148182 79525 148242 186219
rect 148550 89730 148610 186627
rect 149283 186148 149349 186149
rect 149283 186084 149284 186148
rect 149348 186084 149349 186148
rect 149283 186083 149349 186084
rect 148731 183428 148797 183429
rect 148731 183364 148732 183428
rect 148796 183364 148797 183428
rect 148731 183363 148797 183364
rect 148366 89670 148610 89730
rect 148366 80885 148426 89670
rect 148363 80884 148429 80885
rect 148363 80820 148364 80884
rect 148428 80820 148429 80884
rect 148363 80819 148429 80820
rect 148179 79524 148245 79525
rect 148179 79460 148180 79524
rect 148244 79460 148245 79524
rect 148179 79459 148245 79460
rect 148547 79524 148613 79525
rect 148547 79460 148548 79524
rect 148612 79460 148613 79524
rect 148547 79459 148613 79460
rect 148179 78300 148245 78301
rect 148179 78236 148180 78300
rect 148244 78236 148245 78300
rect 148179 78235 148245 78236
rect 147995 77892 148061 77893
rect 147995 77828 147996 77892
rect 148060 77828 148061 77892
rect 147995 77827 148061 77828
rect 147811 77756 147877 77757
rect 147811 77692 147812 77756
rect 147876 77692 147877 77756
rect 147811 77691 147877 77692
rect 147998 77485 148058 77827
rect 147995 77484 148061 77485
rect 147995 77420 147996 77484
rect 148060 77420 148061 77484
rect 147995 77419 148061 77420
rect 148182 68645 148242 78235
rect 148363 77484 148429 77485
rect 148363 77420 148364 77484
rect 148428 77420 148429 77484
rect 148363 77419 148429 77420
rect 148366 77077 148426 77419
rect 148363 77076 148429 77077
rect 148363 77012 148364 77076
rect 148428 77012 148429 77076
rect 148363 77011 148429 77012
rect 148179 68644 148245 68645
rect 148179 68580 148180 68644
rect 148244 68580 148245 68644
rect 148179 68579 148245 68580
rect 148182 54909 148242 68579
rect 148366 67285 148426 77011
rect 148550 70410 148610 79459
rect 148734 78029 148794 183363
rect 148915 178532 148981 178533
rect 148915 178468 148916 178532
rect 148980 178468 148981 178532
rect 148915 178467 148981 178468
rect 148918 79253 148978 178467
rect 149099 79932 149165 79933
rect 149099 79868 149100 79932
rect 149164 79868 149165 79932
rect 149099 79867 149165 79868
rect 148915 79252 148981 79253
rect 148915 79188 148916 79252
rect 148980 79188 148981 79252
rect 148915 79187 148981 79188
rect 148731 78028 148797 78029
rect 148731 77964 148732 78028
rect 148796 77964 148797 78028
rect 149102 78026 149162 79867
rect 149286 79525 149346 186083
rect 149470 80477 149530 192611
rect 149467 80476 149533 80477
rect 149467 80412 149468 80476
rect 149532 80412 149533 80476
rect 149467 80411 149533 80412
rect 149654 79797 149714 199819
rect 150942 199205 151002 199819
rect 151123 199748 151189 199749
rect 151123 199684 151124 199748
rect 151188 199684 151189 199748
rect 151123 199683 151189 199684
rect 150939 199204 151005 199205
rect 150939 199140 150940 199204
rect 151004 199140 151005 199204
rect 150939 199139 151005 199140
rect 150294 187954 150914 198000
rect 150294 187718 150326 187954
rect 150562 187718 150646 187954
rect 150882 187718 150914 187954
rect 150294 187634 150914 187718
rect 150294 187398 150326 187634
rect 150562 187398 150646 187634
rect 150882 187398 150914 187634
rect 149835 185604 149901 185605
rect 149835 185540 149836 185604
rect 149900 185540 149901 185604
rect 149835 185539 149901 185540
rect 149838 79933 149898 185539
rect 150294 151954 150914 187398
rect 150294 151718 150326 151954
rect 150562 151718 150646 151954
rect 150882 151718 150914 151954
rect 150294 151634 150914 151718
rect 150294 151398 150326 151634
rect 150562 151398 150646 151634
rect 150882 151398 150914 151634
rect 150294 142000 150914 151398
rect 150939 139364 151005 139365
rect 150939 139300 150940 139364
rect 151004 139300 151005 139364
rect 150939 139299 151005 139300
rect 150942 80341 151002 139299
rect 150939 80340 151005 80341
rect 150939 80276 150940 80340
rect 151004 80276 151005 80340
rect 150939 80275 151005 80276
rect 151126 79933 151186 199683
rect 151307 186420 151373 186421
rect 151307 186356 151308 186420
rect 151372 186356 151373 186420
rect 151307 186355 151373 186356
rect 151859 186420 151925 186421
rect 151859 186356 151860 186420
rect 151924 186356 151925 186420
rect 151859 186355 151925 186356
rect 149835 79932 149901 79933
rect 149835 79868 149836 79932
rect 149900 79868 149901 79932
rect 149835 79867 149901 79868
rect 151123 79932 151189 79933
rect 151123 79868 151124 79932
rect 151188 79868 151189 79932
rect 151123 79867 151189 79868
rect 149651 79796 149717 79797
rect 149651 79732 149652 79796
rect 149716 79732 149717 79796
rect 149651 79731 149717 79732
rect 149283 79524 149349 79525
rect 149283 79460 149284 79524
rect 149348 79460 149349 79524
rect 149283 79459 149349 79460
rect 148731 77963 148797 77964
rect 148918 77966 149162 78026
rect 148918 75581 148978 77966
rect 149099 77892 149165 77893
rect 149099 77828 149100 77892
rect 149164 77828 149165 77892
rect 149099 77827 149165 77828
rect 148915 75580 148981 75581
rect 148915 75516 148916 75580
rect 148980 75516 148981 75580
rect 148915 75515 148981 75516
rect 148918 71093 148978 75515
rect 149102 71773 149162 77827
rect 149283 77756 149349 77757
rect 149283 77692 149284 77756
rect 149348 77692 149349 77756
rect 149283 77691 149349 77692
rect 149286 72861 149346 77691
rect 149654 73949 149714 79731
rect 149838 78981 149898 79867
rect 151126 79117 151186 79867
rect 151310 79797 151370 186355
rect 151491 185604 151557 185605
rect 151491 185540 151492 185604
rect 151556 185540 151557 185604
rect 151491 185539 151557 185540
rect 151494 79933 151554 185539
rect 151675 80340 151741 80341
rect 151675 80276 151676 80340
rect 151740 80276 151741 80340
rect 151675 80275 151741 80276
rect 151678 79933 151738 80275
rect 151862 80069 151922 186355
rect 152227 185604 152293 185605
rect 152227 185540 152228 185604
rect 152292 185540 152293 185604
rect 152227 185539 152293 185540
rect 151859 80068 151925 80069
rect 151859 80004 151860 80068
rect 151924 80004 151925 80068
rect 151859 80003 151925 80004
rect 152230 79933 152290 185539
rect 151491 79932 151557 79933
rect 151491 79868 151492 79932
rect 151556 79868 151557 79932
rect 151491 79867 151557 79868
rect 151675 79932 151741 79933
rect 151675 79868 151676 79932
rect 151740 79868 151741 79932
rect 151675 79867 151741 79868
rect 152227 79932 152293 79933
rect 152227 79868 152228 79932
rect 152292 79868 152293 79932
rect 152227 79867 152293 79868
rect 151307 79796 151373 79797
rect 151307 79732 151308 79796
rect 151372 79732 151373 79796
rect 151307 79731 151373 79732
rect 151675 79796 151741 79797
rect 151675 79732 151676 79796
rect 151740 79732 151741 79796
rect 151675 79731 151741 79732
rect 152043 79796 152109 79797
rect 152043 79732 152044 79796
rect 152108 79732 152109 79796
rect 152043 79731 152109 79732
rect 151310 79117 151370 79731
rect 151123 79116 151189 79117
rect 151123 79052 151124 79116
rect 151188 79052 151189 79116
rect 151123 79051 151189 79052
rect 151307 79116 151373 79117
rect 151307 79052 151308 79116
rect 151372 79052 151373 79116
rect 151307 79051 151373 79052
rect 149835 78980 149901 78981
rect 149835 78916 149836 78980
rect 149900 78916 149901 78980
rect 149835 78915 149901 78916
rect 151307 78708 151373 78709
rect 151307 78644 151308 78708
rect 151372 78644 151373 78708
rect 151307 78643 151373 78644
rect 150019 78300 150085 78301
rect 150019 78236 150020 78300
rect 150084 78236 150085 78300
rect 150019 78235 150085 78236
rect 149651 73948 149717 73949
rect 149651 73884 149652 73948
rect 149716 73884 149717 73948
rect 149651 73883 149717 73884
rect 149283 72860 149349 72861
rect 149283 72796 149284 72860
rect 149348 72796 149349 72860
rect 149283 72795 149349 72796
rect 149835 72860 149901 72861
rect 149835 72796 149836 72860
rect 149900 72796 149901 72860
rect 149835 72795 149901 72796
rect 149099 71772 149165 71773
rect 149099 71708 149100 71772
rect 149164 71708 149165 71772
rect 149099 71707 149165 71708
rect 148915 71092 148981 71093
rect 148915 71028 148916 71092
rect 148980 71028 148981 71092
rect 148915 71027 148981 71028
rect 148550 70350 148978 70410
rect 148363 67284 148429 67285
rect 148363 67220 148364 67284
rect 148428 67220 148429 67284
rect 148363 67219 148429 67220
rect 148179 54908 148245 54909
rect 148179 54844 148180 54908
rect 148244 54844 148245 54908
rect 148179 54843 148245 54844
rect 147443 47564 147509 47565
rect 147443 47500 147444 47564
rect 147508 47500 147509 47564
rect 147443 47499 147509 47500
rect 148918 45117 148978 70350
rect 149102 64890 149162 71707
rect 149102 64830 149714 64890
rect 148915 45116 148981 45117
rect 148915 45052 148916 45116
rect 148980 45052 148981 45116
rect 148915 45051 148981 45052
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145603 37908 145669 37909
rect 145603 37844 145604 37908
rect 145668 37844 145669 37908
rect 145603 37843 145669 37844
rect 145419 17236 145485 17237
rect 145419 17172 145420 17236
rect 145484 17172 145485 17236
rect 145419 17171 145485 17172
rect 144315 11660 144381 11661
rect 144315 11596 144316 11660
rect 144380 11596 144381 11660
rect 144315 11595 144381 11596
rect 141294 -7302 141326 -7066
rect 141562 -7302 141646 -7066
rect 141882 -7302 141914 -7066
rect 141294 -7386 141914 -7302
rect 141294 -7622 141326 -7386
rect 141562 -7622 141646 -7386
rect 141882 -7622 141914 -7386
rect 141294 -7654 141914 -7622
rect 145794 3454 146414 38898
rect 149654 30973 149714 64830
rect 149838 56405 149898 72795
rect 150022 68781 150082 78235
rect 150019 68780 150085 68781
rect 150019 68716 150020 68780
rect 150084 68716 150085 68780
rect 150019 68715 150085 68716
rect 149835 56404 149901 56405
rect 149835 56340 149836 56404
rect 149900 56340 149901 56404
rect 149835 56339 149901 56340
rect 150294 43954 150914 78000
rect 151310 67421 151370 78643
rect 151491 78572 151557 78573
rect 151491 78508 151492 78572
rect 151556 78508 151557 78572
rect 151491 78507 151557 78508
rect 151307 67420 151373 67421
rect 151307 67356 151308 67420
rect 151372 67356 151373 67420
rect 151307 67355 151373 67356
rect 151494 62117 151554 78507
rect 151491 62116 151557 62117
rect 151491 62052 151492 62116
rect 151556 62052 151557 62116
rect 151491 62051 151557 62052
rect 151678 61301 151738 79731
rect 152046 79253 152106 79731
rect 152414 79661 152474 199822
rect 152595 199820 152596 199822
rect 152660 199820 152661 199884
rect 152595 199819 152661 199820
rect 153331 199884 153397 199885
rect 153331 199820 153332 199884
rect 153396 199820 153397 199884
rect 154067 199884 154133 199885
rect 154067 199882 154068 199884
rect 153331 199819 153397 199820
rect 153886 199822 154068 199882
rect 153334 186285 153394 199819
rect 153515 186420 153581 186421
rect 153515 186356 153516 186420
rect 153580 186356 153581 186420
rect 153515 186355 153581 186356
rect 153331 186284 153397 186285
rect 153331 186220 153332 186284
rect 153396 186220 153397 186284
rect 153331 186219 153397 186220
rect 152595 185604 152661 185605
rect 152595 185540 152596 185604
rect 152660 185540 152661 185604
rect 152595 185539 152661 185540
rect 152598 89730 152658 185539
rect 152598 89670 152842 89730
rect 152595 79796 152661 79797
rect 152595 79732 152596 79796
rect 152660 79732 152661 79796
rect 152595 79731 152661 79732
rect 152411 79660 152477 79661
rect 152411 79596 152412 79660
rect 152476 79596 152477 79660
rect 152411 79595 152477 79596
rect 152043 79252 152109 79253
rect 152043 79188 152044 79252
rect 152108 79188 152109 79252
rect 152043 79187 152109 79188
rect 152598 77890 152658 79731
rect 152782 79389 152842 89670
rect 153518 79661 153578 186355
rect 153699 185604 153765 185605
rect 153699 185540 153700 185604
rect 153764 185540 153765 185604
rect 153699 185539 153765 185540
rect 153515 79660 153581 79661
rect 153515 79596 153516 79660
rect 153580 79596 153581 79660
rect 153515 79595 153581 79596
rect 153702 79389 153762 185539
rect 153886 79525 153946 199822
rect 154067 199820 154068 199822
rect 154132 199820 154133 199884
rect 154067 199819 154133 199820
rect 154619 199884 154685 199885
rect 154619 199820 154620 199884
rect 154684 199820 154685 199884
rect 154619 199819 154685 199820
rect 155907 199884 155973 199885
rect 155907 199820 155908 199884
rect 155972 199820 155973 199884
rect 155907 199819 155973 199820
rect 156643 199884 156709 199885
rect 156643 199820 156644 199884
rect 156708 199820 156709 199884
rect 156643 199819 156709 199820
rect 154067 186284 154133 186285
rect 154067 186220 154068 186284
rect 154132 186220 154133 186284
rect 154067 186219 154133 186220
rect 154070 80069 154130 186219
rect 154435 80748 154501 80749
rect 154435 80684 154436 80748
rect 154500 80684 154501 80748
rect 154435 80683 154501 80684
rect 154067 80068 154133 80069
rect 154067 80004 154068 80068
rect 154132 80004 154133 80068
rect 154067 80003 154133 80004
rect 154438 79933 154498 80683
rect 154622 79933 154682 199819
rect 154794 192454 155414 198000
rect 154794 192218 154826 192454
rect 155062 192218 155146 192454
rect 155382 192218 155414 192454
rect 154794 192134 155414 192218
rect 154794 191898 154826 192134
rect 155062 191898 155146 192134
rect 155382 191898 155414 192134
rect 154794 156454 155414 191898
rect 155910 186285 155970 199819
rect 156459 199748 156525 199749
rect 156459 199684 156460 199748
rect 156524 199684 156525 199748
rect 156459 199683 156525 199684
rect 155907 186284 155973 186285
rect 155907 186220 155908 186284
rect 155972 186220 155973 186284
rect 155907 186219 155973 186220
rect 155539 185604 155605 185605
rect 155539 185540 155540 185604
rect 155604 185540 155605 185604
rect 155539 185539 155605 185540
rect 154794 156218 154826 156454
rect 155062 156218 155146 156454
rect 155382 156218 155414 156454
rect 154794 156134 155414 156218
rect 154794 155898 154826 156134
rect 155062 155898 155146 156134
rect 155382 155898 155414 156134
rect 154794 142000 155414 155898
rect 154803 139364 154869 139365
rect 154803 139300 154804 139364
rect 154868 139300 154869 139364
rect 154803 139299 154869 139300
rect 155355 139364 155421 139365
rect 155355 139300 155356 139364
rect 155420 139300 155421 139364
rect 155355 139299 155421 139300
rect 154067 79932 154133 79933
rect 154067 79868 154068 79932
rect 154132 79868 154133 79932
rect 154067 79867 154133 79868
rect 154435 79932 154501 79933
rect 154435 79868 154436 79932
rect 154500 79868 154501 79932
rect 154435 79867 154501 79868
rect 154619 79932 154685 79933
rect 154619 79868 154620 79932
rect 154684 79868 154685 79932
rect 154619 79867 154685 79868
rect 154070 79661 154130 79867
rect 154067 79660 154133 79661
rect 154067 79596 154068 79660
rect 154132 79596 154133 79660
rect 154067 79595 154133 79596
rect 153883 79524 153949 79525
rect 153883 79460 153884 79524
rect 153948 79460 153949 79524
rect 153883 79459 153949 79460
rect 152779 79388 152845 79389
rect 152779 79324 152780 79388
rect 152844 79324 152845 79388
rect 152779 79323 152845 79324
rect 153699 79388 153765 79389
rect 153699 79324 153700 79388
rect 153764 79324 153765 79388
rect 153699 79323 153765 79324
rect 152414 77830 152658 77890
rect 152414 71501 152474 77830
rect 154070 77485 154130 79595
rect 154622 78981 154682 79867
rect 154806 79389 154866 139299
rect 154928 111454 155248 111486
rect 154928 111218 154970 111454
rect 155206 111218 155248 111454
rect 154928 111134 155248 111218
rect 154928 110898 154970 111134
rect 155206 110898 155248 111134
rect 154928 110866 155248 110898
rect 155171 79932 155237 79933
rect 155171 79868 155172 79932
rect 155236 79868 155237 79932
rect 155171 79867 155237 79868
rect 154803 79388 154869 79389
rect 154803 79324 154804 79388
rect 154868 79324 154869 79388
rect 154803 79323 154869 79324
rect 154619 78980 154685 78981
rect 154619 78916 154620 78980
rect 154684 78916 154685 78980
rect 154619 78915 154685 78916
rect 155174 78165 155234 79867
rect 155358 79661 155418 139299
rect 155542 89730 155602 185539
rect 155542 89670 155786 89730
rect 155539 79932 155605 79933
rect 155539 79868 155540 79932
rect 155604 79868 155605 79932
rect 155539 79867 155605 79868
rect 155355 79660 155421 79661
rect 155355 79596 155356 79660
rect 155420 79596 155421 79660
rect 155355 79595 155421 79596
rect 155171 78164 155237 78165
rect 155171 78100 155172 78164
rect 155236 78100 155237 78164
rect 155171 78099 155237 78100
rect 154067 77484 154133 77485
rect 154067 77420 154068 77484
rect 154132 77420 154133 77484
rect 154067 77419 154133 77420
rect 154435 77348 154501 77349
rect 154435 77284 154436 77348
rect 154500 77284 154501 77348
rect 154435 77283 154501 77284
rect 154251 74628 154317 74629
rect 154251 74564 154252 74628
rect 154316 74564 154317 74628
rect 154251 74563 154317 74564
rect 152963 73812 153029 73813
rect 152963 73748 152964 73812
rect 153028 73748 153029 73812
rect 152963 73747 153029 73748
rect 152595 73540 152661 73541
rect 152595 73476 152596 73540
rect 152660 73476 152661 73540
rect 152595 73475 152661 73476
rect 152598 72997 152658 73475
rect 152595 72996 152661 72997
rect 152595 72932 152596 72996
rect 152660 72932 152661 72996
rect 152595 72931 152661 72932
rect 152411 71500 152477 71501
rect 152411 71436 152412 71500
rect 152476 71436 152477 71500
rect 152411 71435 152477 71436
rect 151675 61300 151741 61301
rect 151675 61236 151676 61300
rect 151740 61236 151741 61300
rect 151675 61235 151741 61236
rect 150294 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 150914 43954
rect 150294 43634 150914 43718
rect 150294 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 150914 43634
rect 149651 30972 149717 30973
rect 149651 30908 149652 30972
rect 149716 30908 149717 30972
rect 149651 30907 149717 30908
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -7654 146414 -902
rect 150294 7954 150914 43398
rect 152414 28253 152474 71435
rect 152598 44981 152658 72931
rect 152966 64837 153026 73747
rect 152963 64836 153029 64837
rect 152963 64772 152964 64836
rect 153028 64772 153029 64836
rect 152963 64771 153029 64772
rect 154254 53549 154314 74563
rect 154251 53548 154317 53549
rect 154251 53484 154252 53548
rect 154316 53484 154317 53548
rect 154251 53483 154317 53484
rect 152595 44980 152661 44981
rect 152595 44916 152596 44980
rect 152660 44916 152661 44980
rect 152595 44915 152661 44916
rect 154438 44029 154498 77283
rect 154794 48454 155414 78000
rect 155542 73946 155602 79867
rect 155726 79389 155786 89670
rect 155907 81020 155973 81021
rect 155907 80956 155908 81020
rect 155972 80956 155973 81020
rect 155907 80955 155973 80956
rect 155910 79933 155970 80955
rect 156462 79933 156522 199683
rect 155907 79932 155973 79933
rect 155907 79868 155908 79932
rect 155972 79868 155973 79932
rect 155907 79867 155973 79868
rect 156459 79932 156525 79933
rect 156459 79868 156460 79932
rect 156524 79868 156525 79932
rect 156459 79867 156525 79868
rect 155723 79388 155789 79389
rect 155723 79324 155724 79388
rect 155788 79324 155789 79388
rect 155723 79323 155789 79324
rect 156459 78708 156525 78709
rect 156459 78644 156460 78708
rect 156524 78644 156525 78708
rect 156459 78643 156525 78644
rect 156462 74493 156522 78643
rect 156646 78573 156706 199819
rect 157198 199749 157258 200635
rect 166211 200564 166277 200565
rect 166211 200500 166212 200564
rect 166276 200500 166277 200564
rect 166211 200499 166277 200500
rect 163451 200156 163517 200157
rect 163451 200092 163452 200156
rect 163516 200092 163517 200156
rect 163451 200091 163517 200092
rect 157747 199884 157813 199885
rect 157747 199820 157748 199884
rect 157812 199820 157813 199884
rect 157747 199819 157813 199820
rect 158851 199884 158917 199885
rect 158851 199820 158852 199884
rect 158916 199820 158917 199884
rect 158851 199819 158917 199820
rect 160139 199884 160205 199885
rect 160139 199820 160140 199884
rect 160204 199820 160205 199884
rect 161059 199884 161125 199885
rect 161059 199882 161060 199884
rect 160139 199819 160205 199820
rect 160878 199822 161060 199882
rect 157195 199748 157261 199749
rect 157195 199684 157196 199748
rect 157260 199684 157261 199748
rect 157195 199683 157261 199684
rect 156827 185604 156893 185605
rect 156827 185540 156828 185604
rect 156892 185540 156893 185604
rect 156827 185539 156893 185540
rect 157195 185604 157261 185605
rect 157195 185540 157196 185604
rect 157260 185540 157261 185604
rect 157195 185539 157261 185540
rect 156830 79661 156890 185539
rect 157198 80069 157258 185539
rect 157195 80068 157261 80069
rect 157195 80004 157196 80068
rect 157260 80004 157261 80068
rect 157195 80003 157261 80004
rect 157195 79932 157261 79933
rect 157195 79868 157196 79932
rect 157260 79868 157261 79932
rect 157195 79867 157261 79868
rect 157011 79796 157077 79797
rect 157011 79732 157012 79796
rect 157076 79732 157077 79796
rect 157011 79731 157077 79732
rect 156827 79660 156893 79661
rect 156827 79596 156828 79660
rect 156892 79596 156893 79660
rect 156827 79595 156893 79596
rect 156643 78572 156709 78573
rect 156643 78508 156644 78572
rect 156708 78508 156709 78572
rect 157014 78570 157074 79731
rect 156643 78507 156709 78508
rect 156830 78510 157074 78570
rect 156459 74492 156525 74493
rect 156459 74428 156460 74492
rect 156524 74428 156525 74492
rect 156459 74427 156525 74428
rect 155542 73886 155786 73946
rect 155726 60621 155786 73886
rect 156830 61845 156890 78510
rect 157011 77620 157077 77621
rect 157011 77556 157012 77620
rect 157076 77556 157077 77620
rect 157011 77555 157077 77556
rect 156827 61844 156893 61845
rect 156827 61780 156828 61844
rect 156892 61780 156893 61844
rect 156827 61779 156893 61780
rect 155723 60620 155789 60621
rect 155723 60556 155724 60620
rect 155788 60556 155789 60620
rect 155723 60555 155789 60556
rect 157014 57901 157074 77555
rect 157011 57900 157077 57901
rect 157011 57836 157012 57900
rect 157076 57836 157077 57900
rect 157011 57835 157077 57836
rect 157198 56269 157258 79867
rect 157750 79389 157810 199819
rect 157931 199748 157997 199749
rect 157931 199684 157932 199748
rect 157996 199684 157997 199748
rect 157931 199683 157997 199684
rect 158299 199748 158365 199749
rect 158299 199684 158300 199748
rect 158364 199684 158365 199748
rect 158299 199683 158365 199684
rect 157934 79389 157994 199683
rect 158115 186284 158181 186285
rect 158115 186220 158116 186284
rect 158180 186220 158181 186284
rect 158115 186219 158181 186220
rect 158118 79797 158178 186219
rect 158302 79933 158362 199683
rect 158854 80341 158914 199819
rect 159294 196954 159914 198000
rect 159294 196718 159326 196954
rect 159562 196718 159646 196954
rect 159882 196718 159914 196954
rect 159294 196634 159914 196718
rect 159294 196398 159326 196634
rect 159562 196398 159646 196634
rect 159882 196398 159914 196634
rect 159035 179484 159101 179485
rect 159035 179420 159036 179484
rect 159100 179420 159101 179484
rect 159035 179419 159101 179420
rect 158851 80340 158917 80341
rect 158851 80276 158852 80340
rect 158916 80276 158917 80340
rect 158851 80275 158917 80276
rect 158299 79932 158365 79933
rect 158299 79868 158300 79932
rect 158364 79868 158365 79932
rect 158299 79867 158365 79868
rect 158115 79796 158181 79797
rect 158115 79732 158116 79796
rect 158180 79732 158181 79796
rect 158115 79731 158181 79732
rect 157747 79388 157813 79389
rect 157747 79324 157748 79388
rect 157812 79324 157813 79388
rect 157747 79323 157813 79324
rect 157931 79388 157997 79389
rect 157931 79324 157932 79388
rect 157996 79324 157997 79388
rect 157931 79323 157997 79324
rect 158302 78981 158362 79867
rect 159038 79797 159098 179419
rect 159294 160954 159914 196398
rect 160142 186285 160202 199819
rect 160139 186284 160205 186285
rect 160139 186220 160140 186284
rect 160204 186220 160205 186284
rect 160139 186219 160205 186220
rect 160691 185604 160757 185605
rect 160691 185540 160692 185604
rect 160756 185540 160757 185604
rect 160691 185539 160757 185540
rect 159294 160718 159326 160954
rect 159562 160718 159646 160954
rect 159882 160718 159914 160954
rect 159294 160634 159914 160718
rect 159294 160398 159326 160634
rect 159562 160398 159646 160634
rect 159882 160398 159914 160634
rect 159294 142000 159914 160398
rect 159219 139364 159285 139365
rect 159219 139300 159220 139364
rect 159284 139300 159285 139364
rect 159219 139299 159285 139300
rect 159955 139364 160021 139365
rect 159955 139300 159956 139364
rect 160020 139300 160021 139364
rect 159955 139299 160021 139300
rect 159222 93870 159282 139299
rect 159222 93810 159834 93870
rect 159219 80612 159285 80613
rect 159219 80548 159220 80612
rect 159284 80548 159285 80612
rect 159219 80547 159285 80548
rect 159035 79796 159101 79797
rect 159035 79732 159036 79796
rect 159100 79732 159101 79796
rect 159035 79731 159101 79732
rect 158483 79660 158549 79661
rect 158483 79596 158484 79660
rect 158548 79596 158549 79660
rect 158483 79595 158549 79596
rect 158299 78980 158365 78981
rect 158299 78916 158300 78980
rect 158364 78916 158365 78980
rect 158299 78915 158365 78916
rect 158115 78844 158181 78845
rect 158115 78780 158116 78844
rect 158180 78780 158181 78844
rect 158115 78779 158181 78780
rect 157931 75988 157997 75989
rect 157931 75924 157932 75988
rect 157996 75924 157997 75988
rect 157931 75923 157997 75924
rect 157934 63477 157994 75923
rect 157931 63476 157997 63477
rect 157931 63412 157932 63476
rect 157996 63412 157997 63476
rect 157931 63411 157997 63412
rect 158118 60485 158178 78779
rect 158299 78572 158365 78573
rect 158299 78508 158300 78572
rect 158364 78508 158365 78572
rect 158299 78507 158365 78508
rect 158115 60484 158181 60485
rect 158115 60420 158116 60484
rect 158180 60420 158181 60484
rect 158115 60419 158181 60420
rect 158302 59125 158362 78507
rect 158299 59124 158365 59125
rect 158299 59060 158300 59124
rect 158364 59060 158365 59124
rect 158299 59059 158365 59060
rect 157195 56268 157261 56269
rect 157195 56204 157196 56268
rect 157260 56204 157261 56268
rect 157195 56203 157261 56204
rect 158486 55045 158546 79595
rect 159222 79525 159282 80547
rect 159774 79661 159834 93810
rect 159771 79660 159837 79661
rect 159771 79596 159772 79660
rect 159836 79596 159837 79660
rect 159771 79595 159837 79596
rect 159219 79524 159285 79525
rect 159219 79460 159220 79524
rect 159284 79460 159285 79524
rect 159219 79459 159285 79460
rect 159958 78981 160018 139299
rect 160694 109050 160754 185539
rect 160510 108990 160754 109050
rect 160139 79932 160205 79933
rect 160139 79868 160140 79932
rect 160204 79930 160205 79932
rect 160204 79870 160386 79930
rect 160204 79868 160205 79870
rect 160139 79867 160205 79868
rect 159955 78980 160021 78981
rect 159955 78916 159956 78980
rect 160020 78916 160021 78980
rect 159955 78915 160021 78916
rect 159035 75036 159101 75037
rect 159035 74972 159036 75036
rect 159100 74972 159101 75036
rect 159035 74971 159101 74972
rect 158851 71908 158917 71909
rect 158851 71844 158852 71908
rect 158916 71844 158917 71908
rect 158851 71843 158917 71844
rect 158483 55044 158549 55045
rect 158483 54980 158484 55044
rect 158548 54980 158549 55044
rect 158483 54979 158549 54980
rect 158854 53413 158914 71843
rect 158851 53412 158917 53413
rect 158851 53348 158852 53412
rect 158916 53348 158917 53412
rect 158851 53347 158917 53348
rect 159038 50965 159098 74971
rect 159294 52954 159914 78000
rect 160326 77893 160386 79870
rect 160510 79661 160570 108990
rect 160691 81972 160757 81973
rect 160691 81908 160692 81972
rect 160756 81908 160757 81972
rect 160691 81907 160757 81908
rect 160507 79660 160573 79661
rect 160507 79596 160508 79660
rect 160572 79596 160573 79660
rect 160507 79595 160573 79596
rect 160694 78845 160754 81907
rect 160878 79933 160938 199822
rect 161059 199820 161060 199822
rect 161124 199820 161125 199884
rect 161059 199819 161125 199820
rect 161611 199884 161677 199885
rect 161611 199820 161612 199884
rect 161676 199820 161677 199884
rect 161611 199819 161677 199820
rect 162347 199884 162413 199885
rect 162347 199820 162348 199884
rect 162412 199820 162413 199884
rect 162347 199819 162413 199820
rect 163267 199884 163333 199885
rect 163267 199820 163268 199884
rect 163332 199820 163333 199884
rect 163267 199819 163333 199820
rect 161614 186693 161674 199819
rect 161611 186692 161677 186693
rect 161611 186628 161612 186692
rect 161676 186628 161677 186692
rect 161611 186627 161677 186628
rect 161427 186556 161493 186557
rect 161427 186492 161428 186556
rect 161492 186492 161493 186556
rect 161427 186491 161493 186492
rect 161430 185330 161490 186491
rect 162163 186420 162229 186421
rect 162163 186356 162164 186420
rect 162228 186356 162229 186420
rect 162163 186355 162229 186356
rect 161246 185270 161490 185330
rect 161059 177988 161125 177989
rect 161059 177924 161060 177988
rect 161124 177924 161125 177988
rect 161059 177923 161125 177924
rect 160875 79932 160941 79933
rect 160875 79868 160876 79932
rect 160940 79868 160941 79932
rect 160875 79867 160941 79868
rect 160875 79796 160941 79797
rect 160875 79732 160876 79796
rect 160940 79732 160941 79796
rect 160875 79731 160941 79732
rect 160691 78844 160757 78845
rect 160691 78780 160692 78844
rect 160756 78780 160757 78844
rect 160691 78779 160757 78780
rect 160323 77892 160389 77893
rect 160323 77828 160324 77892
rect 160388 77828 160389 77892
rect 160323 77827 160389 77828
rect 160878 68370 160938 79731
rect 161062 79525 161122 177923
rect 161246 81973 161306 185270
rect 161427 171188 161493 171189
rect 161427 171124 161428 171188
rect 161492 171124 161493 171188
rect 161427 171123 161493 171124
rect 161430 171053 161490 171123
rect 161427 171052 161493 171053
rect 161427 170988 161428 171052
rect 161492 170988 161493 171052
rect 161427 170987 161493 170988
rect 161427 161532 161493 161533
rect 161427 161468 161428 161532
rect 161492 161468 161493 161532
rect 161427 161467 161493 161468
rect 161430 161397 161490 161467
rect 161427 161396 161493 161397
rect 161427 161332 161428 161396
rect 161492 161332 161493 161396
rect 161427 161331 161493 161332
rect 161427 151876 161493 151877
rect 161427 151812 161428 151876
rect 161492 151812 161493 151876
rect 161427 151811 161493 151812
rect 161430 151741 161490 151811
rect 161427 151740 161493 151741
rect 161427 151676 161428 151740
rect 161492 151676 161493 151740
rect 161427 151675 161493 151676
rect 161611 142356 161677 142357
rect 161611 142292 161612 142356
rect 161676 142292 161677 142356
rect 161611 142291 161677 142292
rect 161243 81972 161309 81973
rect 161243 81908 161244 81972
rect 161308 81908 161309 81972
rect 161243 81907 161309 81908
rect 161427 80884 161493 80885
rect 161427 80820 161428 80884
rect 161492 80820 161493 80884
rect 161427 80819 161493 80820
rect 161243 79932 161309 79933
rect 161243 79868 161244 79932
rect 161308 79868 161309 79932
rect 161243 79867 161309 79868
rect 161059 79524 161125 79525
rect 161059 79460 161060 79524
rect 161124 79460 161125 79524
rect 161059 79459 161125 79460
rect 161059 78572 161125 78573
rect 161059 78508 161060 78572
rect 161124 78508 161125 78572
rect 161059 78507 161125 78508
rect 160694 68310 160938 68370
rect 160694 59261 160754 68310
rect 160875 67692 160941 67693
rect 160875 67628 160876 67692
rect 160940 67628 160941 67692
rect 160875 67627 160941 67628
rect 160691 59260 160757 59261
rect 160691 59196 160692 59260
rect 160756 59196 160757 59260
rect 160691 59195 160757 59196
rect 160878 55181 160938 67627
rect 160875 55180 160941 55181
rect 160875 55116 160876 55180
rect 160940 55116 160941 55180
rect 160875 55115 160941 55116
rect 159294 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 159914 52954
rect 159294 52634 159914 52718
rect 159294 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 159914 52634
rect 159035 50964 159101 50965
rect 159035 50900 159036 50964
rect 159100 50900 159101 50964
rect 159035 50899 159101 50900
rect 154794 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 155414 48454
rect 154794 48134 155414 48218
rect 154794 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 155414 48134
rect 154435 44028 154501 44029
rect 154435 43964 154436 44028
rect 154500 43964 154501 44028
rect 154435 43963 154501 43964
rect 152411 28252 152477 28253
rect 152411 28188 152412 28252
rect 152476 28188 152477 28252
rect 152411 28187 152477 28188
rect 150294 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 150914 7954
rect 150294 7634 150914 7718
rect 150294 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 150914 7634
rect 150294 -1306 150914 7398
rect 150294 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 150914 -1306
rect 150294 -1626 150914 -1542
rect 150294 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 150914 -1626
rect 150294 -7654 150914 -1862
rect 154794 12454 155414 47898
rect 154794 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 155414 12454
rect 154794 12134 155414 12218
rect 154794 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 155414 12134
rect 154794 -2266 155414 11898
rect 154794 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 155414 -2266
rect 154794 -2586 155414 -2502
rect 154794 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 155414 -2586
rect 154794 -7654 155414 -2822
rect 159294 16954 159914 52398
rect 161062 52053 161122 78507
rect 161246 74221 161306 79867
rect 161430 79797 161490 80819
rect 161427 79796 161493 79797
rect 161427 79732 161428 79796
rect 161492 79732 161493 79796
rect 161427 79731 161493 79732
rect 161614 79389 161674 142291
rect 161795 80476 161861 80477
rect 161795 80412 161796 80476
rect 161860 80412 161861 80476
rect 161795 80411 161861 80412
rect 161798 79661 161858 80411
rect 162166 80069 162226 186355
rect 162163 80068 162229 80069
rect 162163 80004 162164 80068
rect 162228 80004 162229 80068
rect 162163 80003 162229 80004
rect 161979 79932 162045 79933
rect 161979 79868 161980 79932
rect 162044 79868 162045 79932
rect 161979 79867 162045 79868
rect 161795 79660 161861 79661
rect 161795 79596 161796 79660
rect 161860 79596 161861 79660
rect 161795 79595 161861 79596
rect 161611 79388 161677 79389
rect 161611 79324 161612 79388
rect 161676 79324 161677 79388
rect 161611 79323 161677 79324
rect 161243 74220 161309 74221
rect 161243 74156 161244 74220
rect 161308 74156 161309 74220
rect 161243 74155 161309 74156
rect 161243 67556 161309 67557
rect 161243 67492 161244 67556
rect 161308 67492 161309 67556
rect 161243 67491 161309 67492
rect 161246 52189 161306 67491
rect 161982 66061 162042 79867
rect 162350 79661 162410 199819
rect 162899 199748 162965 199749
rect 162899 199684 162900 199748
rect 162964 199684 162965 199748
rect 162899 199683 162965 199684
rect 163083 199748 163149 199749
rect 163083 199684 163084 199748
rect 163148 199684 163149 199748
rect 163083 199683 163149 199684
rect 162902 198389 162962 199683
rect 162899 198388 162965 198389
rect 162899 198324 162900 198388
rect 162964 198324 162965 198388
rect 162899 198323 162965 198324
rect 162899 198252 162965 198253
rect 162899 198188 162900 198252
rect 162964 198188 162965 198252
rect 162899 198187 162965 198188
rect 162902 186829 162962 198187
rect 163086 198117 163146 199683
rect 163270 198117 163330 199819
rect 163454 198933 163514 200091
rect 164923 199884 164989 199885
rect 164923 199820 164924 199884
rect 164988 199820 164989 199884
rect 164923 199819 164989 199820
rect 163451 198932 163517 198933
rect 163451 198868 163452 198932
rect 163516 198868 163517 198932
rect 163451 198867 163517 198868
rect 164926 198117 164986 199819
rect 165475 199748 165541 199749
rect 165475 199684 165476 199748
rect 165540 199684 165541 199748
rect 165475 199683 165541 199684
rect 163083 198116 163149 198117
rect 163083 198052 163084 198116
rect 163148 198052 163149 198116
rect 163083 198051 163149 198052
rect 163267 198116 163333 198117
rect 163267 198052 163268 198116
rect 163332 198052 163333 198116
rect 163267 198051 163333 198052
rect 164923 198116 164989 198117
rect 164923 198052 164924 198116
rect 164988 198052 164989 198116
rect 164923 198051 164989 198052
rect 163635 186964 163701 186965
rect 163635 186900 163636 186964
rect 163700 186900 163701 186964
rect 163635 186899 163701 186900
rect 162899 186828 162965 186829
rect 162899 186764 162900 186828
rect 162964 186764 162965 186828
rect 162899 186763 162965 186764
rect 162531 186284 162597 186285
rect 162531 186220 162532 186284
rect 162596 186220 162597 186284
rect 162531 186219 162597 186220
rect 163267 186284 163333 186285
rect 163267 186220 163268 186284
rect 163332 186220 163333 186284
rect 163267 186219 163333 186220
rect 162347 79660 162413 79661
rect 162347 79596 162348 79660
rect 162412 79596 162413 79660
rect 162347 79595 162413 79596
rect 162534 79525 162594 186219
rect 162899 186148 162965 186149
rect 162899 186084 162900 186148
rect 162964 186084 162965 186148
rect 162899 186083 162965 186084
rect 162902 79525 162962 186083
rect 163270 80069 163330 186219
rect 163267 80068 163333 80069
rect 163267 80004 163268 80068
rect 163332 80004 163333 80068
rect 163267 80003 163333 80004
rect 163451 79932 163517 79933
rect 163451 79868 163452 79932
rect 163516 79868 163517 79932
rect 163451 79867 163517 79868
rect 162531 79524 162597 79525
rect 162531 79460 162532 79524
rect 162596 79460 162597 79524
rect 162531 79459 162597 79460
rect 162899 79524 162965 79525
rect 162899 79460 162900 79524
rect 162964 79460 162965 79524
rect 162899 79459 162965 79460
rect 163454 78842 163514 79867
rect 163638 79661 163698 186899
rect 164003 186420 164069 186421
rect 164003 186356 164004 186420
rect 164068 186356 164069 186420
rect 164003 186355 164069 186356
rect 164923 186420 164989 186421
rect 164923 186356 164924 186420
rect 164988 186356 164989 186420
rect 164923 186355 164989 186356
rect 164006 79797 164066 186355
rect 164739 186284 164805 186285
rect 164739 186220 164740 186284
rect 164804 186220 164805 186284
rect 164739 186219 164805 186220
rect 164742 79933 164802 186219
rect 164555 79932 164621 79933
rect 164555 79868 164556 79932
rect 164620 79868 164621 79932
rect 164555 79867 164621 79868
rect 164739 79932 164805 79933
rect 164739 79868 164740 79932
rect 164804 79868 164805 79932
rect 164739 79867 164805 79868
rect 164003 79796 164069 79797
rect 164003 79732 164004 79796
rect 164068 79732 164069 79796
rect 164003 79731 164069 79732
rect 163635 79660 163701 79661
rect 163635 79596 163636 79660
rect 163700 79596 163701 79660
rect 163635 79595 163701 79596
rect 163270 78782 163514 78842
rect 162715 78572 162781 78573
rect 162715 78508 162716 78572
rect 162780 78508 162781 78572
rect 162715 78507 162781 78508
rect 162531 71772 162597 71773
rect 162531 71708 162532 71772
rect 162596 71708 162597 71772
rect 162531 71707 162597 71708
rect 161979 66060 162045 66061
rect 161979 65996 161980 66060
rect 162044 65996 162045 66060
rect 161979 65995 162045 65996
rect 162534 53685 162594 71707
rect 162531 53684 162597 53685
rect 162531 53620 162532 53684
rect 162596 53620 162597 53684
rect 162531 53619 162597 53620
rect 161243 52188 161309 52189
rect 161243 52124 161244 52188
rect 161308 52124 161309 52188
rect 161243 52123 161309 52124
rect 161059 52052 161125 52053
rect 161059 51988 161060 52052
rect 161124 51988 161125 52052
rect 161059 51987 161125 51988
rect 162718 48245 162778 78507
rect 163270 56541 163330 78782
rect 163451 78708 163517 78709
rect 163451 78644 163452 78708
rect 163516 78644 163517 78708
rect 163451 78643 163517 78644
rect 163267 56540 163333 56541
rect 163267 56476 163268 56540
rect 163332 56476 163333 56540
rect 163267 56475 163333 56476
rect 163454 50693 163514 78643
rect 164006 78165 164066 79731
rect 164558 78301 164618 79867
rect 164742 79253 164802 79867
rect 164926 79661 164986 186355
rect 165291 178532 165357 178533
rect 165291 178468 165292 178532
rect 165356 178468 165357 178532
rect 165291 178467 165357 178468
rect 165294 79933 165354 178467
rect 165291 79932 165357 79933
rect 165291 79868 165292 79932
rect 165356 79868 165357 79932
rect 165291 79867 165357 79868
rect 164923 79660 164989 79661
rect 164923 79596 164924 79660
rect 164988 79596 164989 79660
rect 164923 79595 164989 79596
rect 164739 79252 164805 79253
rect 164739 79188 164740 79252
rect 164804 79188 164805 79252
rect 164739 79187 164805 79188
rect 165291 79252 165357 79253
rect 165291 79188 165292 79252
rect 165356 79188 165357 79252
rect 165291 79187 165357 79188
rect 164555 78300 164621 78301
rect 164555 78236 164556 78300
rect 164620 78236 164621 78300
rect 164555 78235 164621 78236
rect 164003 78164 164069 78165
rect 164003 78100 164004 78164
rect 164068 78100 164069 78164
rect 164003 78099 164069 78100
rect 163635 77620 163701 77621
rect 163635 77556 163636 77620
rect 163700 77556 163701 77620
rect 163635 77555 163701 77556
rect 163451 50692 163517 50693
rect 163451 50628 163452 50692
rect 163516 50628 163517 50692
rect 163451 50627 163517 50628
rect 162715 48244 162781 48245
rect 162715 48180 162716 48244
rect 162780 48180 162781 48244
rect 162715 48179 162781 48180
rect 163638 45525 163698 77555
rect 163794 57454 164414 78000
rect 164558 77621 164618 78235
rect 164555 77620 164621 77621
rect 164555 77556 164556 77620
rect 164620 77556 164621 77620
rect 164555 77555 164621 77556
rect 165107 77484 165173 77485
rect 165107 77420 165108 77484
rect 165172 77420 165173 77484
rect 165107 77419 165173 77420
rect 165110 63069 165170 77419
rect 165107 63068 165173 63069
rect 165107 63004 165108 63068
rect 165172 63004 165173 63068
rect 165107 63003 165173 63004
rect 165294 57765 165354 79187
rect 165478 78437 165538 199683
rect 166214 199069 166274 200499
rect 166579 200428 166645 200429
rect 166579 200364 166580 200428
rect 166644 200364 166645 200428
rect 166579 200363 166645 200364
rect 166582 199749 166642 200363
rect 169155 200156 169221 200157
rect 169155 200092 169156 200156
rect 169220 200092 169221 200156
rect 169155 200091 169221 200092
rect 166947 199884 167013 199885
rect 166947 199820 166948 199884
rect 167012 199820 167013 199884
rect 166947 199819 167013 199820
rect 167867 199884 167933 199885
rect 167867 199820 167868 199884
rect 167932 199820 167933 199884
rect 167867 199819 167933 199820
rect 168051 199884 168117 199885
rect 168051 199820 168052 199884
rect 168116 199820 168117 199884
rect 168051 199819 168117 199820
rect 168603 199884 168669 199885
rect 168603 199820 168604 199884
rect 168668 199820 168669 199884
rect 168603 199819 168669 199820
rect 166579 199748 166645 199749
rect 166579 199684 166580 199748
rect 166644 199684 166645 199748
rect 166579 199683 166645 199684
rect 166763 199748 166829 199749
rect 166763 199684 166764 199748
rect 166828 199684 166829 199748
rect 166763 199683 166829 199684
rect 166211 199068 166277 199069
rect 166211 199004 166212 199068
rect 166276 199004 166277 199068
rect 166211 199003 166277 199004
rect 166027 185740 166093 185741
rect 166027 185676 166028 185740
rect 166092 185676 166093 185740
rect 166027 185675 166093 185676
rect 166211 185740 166277 185741
rect 166211 185676 166212 185740
rect 166276 185676 166277 185740
rect 166211 185675 166277 185676
rect 165843 185604 165909 185605
rect 165843 185540 165844 185604
rect 165908 185540 165909 185604
rect 165843 185539 165909 185540
rect 165846 78709 165906 185539
rect 166030 79797 166090 185675
rect 166214 79933 166274 185675
rect 166766 185333 166826 199683
rect 166950 198117 167010 199819
rect 167499 199748 167565 199749
rect 167499 199684 167500 199748
rect 167564 199684 167565 199748
rect 167499 199683 167565 199684
rect 166947 198116 167013 198117
rect 166947 198052 166948 198116
rect 167012 198052 167013 198116
rect 166947 198051 167013 198052
rect 167502 197845 167562 199683
rect 167683 198252 167749 198253
rect 167683 198188 167684 198252
rect 167748 198188 167749 198252
rect 167683 198187 167749 198188
rect 167499 197844 167565 197845
rect 167499 197780 167500 197844
rect 167564 197780 167565 197844
rect 167499 197779 167565 197780
rect 167315 185740 167381 185741
rect 167315 185676 167316 185740
rect 167380 185676 167381 185740
rect 167315 185675 167381 185676
rect 166763 185332 166829 185333
rect 166763 185268 166764 185332
rect 166828 185268 166829 185332
rect 166763 185267 166829 185268
rect 166579 180300 166645 180301
rect 166579 180236 166580 180300
rect 166644 180236 166645 180300
rect 166579 180235 166645 180236
rect 166211 79932 166277 79933
rect 166211 79868 166212 79932
rect 166276 79868 166277 79932
rect 166211 79867 166277 79868
rect 166027 79796 166093 79797
rect 166027 79732 166028 79796
rect 166092 79732 166093 79796
rect 166027 79731 166093 79732
rect 166395 79796 166461 79797
rect 166395 79732 166396 79796
rect 166460 79732 166461 79796
rect 166395 79731 166461 79732
rect 166398 78709 166458 79731
rect 166582 79253 166642 180235
rect 166947 80204 167013 80205
rect 166947 80140 166948 80204
rect 167012 80140 167013 80204
rect 166947 80139 167013 80140
rect 166579 79252 166645 79253
rect 166579 79188 166580 79252
rect 166644 79188 166645 79252
rect 166579 79187 166645 79188
rect 166579 79116 166645 79117
rect 166579 79052 166580 79116
rect 166644 79052 166645 79116
rect 166579 79051 166645 79052
rect 165843 78708 165909 78709
rect 165843 78644 165844 78708
rect 165908 78644 165909 78708
rect 165843 78643 165909 78644
rect 166395 78708 166461 78709
rect 166395 78644 166396 78708
rect 166460 78644 166461 78708
rect 166395 78643 166461 78644
rect 165475 78436 165541 78437
rect 165475 78372 165476 78436
rect 165540 78372 165541 78436
rect 165475 78371 165541 78372
rect 165475 77756 165541 77757
rect 165475 77692 165476 77756
rect 165540 77692 165541 77756
rect 165475 77691 165541 77692
rect 165291 57764 165357 57765
rect 165291 57700 165292 57764
rect 165356 57700 165357 57764
rect 165291 57699 165357 57700
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163635 45524 163701 45525
rect 163635 45460 163636 45524
rect 163700 45460 163701 45524
rect 163635 45459 163701 45460
rect 159294 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 159914 16954
rect 159294 16634 159914 16718
rect 159294 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 159914 16634
rect 159294 -3226 159914 16398
rect 159294 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 159914 -3226
rect 159294 -3546 159914 -3462
rect 159294 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 159914 -3546
rect 159294 -7654 159914 -3782
rect 163794 21454 164414 56898
rect 165478 54501 165538 77691
rect 165475 54500 165541 54501
rect 165475 54436 165476 54500
rect 165540 54436 165541 54500
rect 165475 54435 165541 54436
rect 166582 53821 166642 79051
rect 166763 73676 166829 73677
rect 166763 73612 166764 73676
rect 166828 73612 166829 73676
rect 166763 73611 166829 73612
rect 166579 53820 166645 53821
rect 166579 53756 166580 53820
rect 166644 53756 166645 53820
rect 166579 53755 166645 53756
rect 166766 50829 166826 73611
rect 166950 71365 167010 80139
rect 167318 79253 167378 185675
rect 167499 185604 167565 185605
rect 167499 185540 167500 185604
rect 167564 185540 167565 185604
rect 167499 185539 167565 185540
rect 167502 79797 167562 185539
rect 167686 79933 167746 198187
rect 167870 198117 167930 199819
rect 168054 198117 168114 199819
rect 167867 198116 167933 198117
rect 167867 198052 167868 198116
rect 167932 198052 167933 198116
rect 167867 198051 167933 198052
rect 168051 198116 168117 198117
rect 168051 198052 168052 198116
rect 168116 198052 168117 198116
rect 168051 198051 168117 198052
rect 168606 196485 168666 199819
rect 168971 199748 169037 199749
rect 168971 199684 168972 199748
rect 169036 199684 169037 199748
rect 168971 199683 169037 199684
rect 168603 196484 168669 196485
rect 168603 196420 168604 196484
rect 168668 196420 168669 196484
rect 168603 196419 168669 196420
rect 168051 185604 168117 185605
rect 168051 185540 168052 185604
rect 168116 185540 168117 185604
rect 168051 185539 168117 185540
rect 168603 185604 168669 185605
rect 168603 185540 168604 185604
rect 168668 185540 168669 185604
rect 168603 185539 168669 185540
rect 168054 93870 168114 185539
rect 168054 93810 168298 93870
rect 168238 79933 168298 93810
rect 167683 79932 167749 79933
rect 167683 79868 167684 79932
rect 167748 79868 167749 79932
rect 167683 79867 167749 79868
rect 168235 79932 168301 79933
rect 168235 79868 168236 79932
rect 168300 79868 168301 79932
rect 168235 79867 168301 79868
rect 167499 79796 167565 79797
rect 167499 79732 167500 79796
rect 167564 79732 167565 79796
rect 167499 79731 167565 79732
rect 167686 79661 167746 79867
rect 167683 79660 167749 79661
rect 167683 79596 167684 79660
rect 167748 79596 167749 79660
rect 167683 79595 167749 79596
rect 168238 79253 168298 79867
rect 168606 79253 168666 185539
rect 168787 180028 168853 180029
rect 168787 179964 168788 180028
rect 168852 179964 168853 180028
rect 168787 179963 168853 179964
rect 168790 79933 168850 179963
rect 168787 79932 168853 79933
rect 168787 79868 168788 79932
rect 168852 79868 168853 79932
rect 168787 79867 168853 79868
rect 168974 79661 169034 199683
rect 169158 185877 169218 200091
rect 169339 199884 169405 199885
rect 169339 199820 169340 199884
rect 169404 199820 169405 199884
rect 169339 199819 169405 199820
rect 170995 199884 171061 199885
rect 170995 199820 170996 199884
rect 171060 199820 171061 199884
rect 170995 199819 171061 199820
rect 171731 199884 171797 199885
rect 171731 199820 171732 199884
rect 171796 199820 171797 199884
rect 171731 199819 171797 199820
rect 172835 199884 172901 199885
rect 172835 199820 172836 199884
rect 172900 199820 172901 199884
rect 172835 199819 172901 199820
rect 174491 199884 174557 199885
rect 174491 199820 174492 199884
rect 174556 199820 174557 199884
rect 174491 199819 174557 199820
rect 175043 199884 175109 199885
rect 175043 199820 175044 199884
rect 175108 199820 175109 199884
rect 175043 199819 175109 199820
rect 175411 199884 175477 199885
rect 175411 199820 175412 199884
rect 175476 199820 175477 199884
rect 176515 199884 176581 199885
rect 176515 199882 176516 199884
rect 175411 199819 175477 199820
rect 176150 199822 176516 199882
rect 169342 195941 169402 199819
rect 170075 199748 170141 199749
rect 170075 199684 170076 199748
rect 170140 199684 170141 199748
rect 170075 199683 170141 199684
rect 169339 195940 169405 195941
rect 169339 195876 169340 195940
rect 169404 195876 169405 195940
rect 169339 195875 169405 195876
rect 169891 186420 169957 186421
rect 169891 186356 169892 186420
rect 169956 186356 169957 186420
rect 169891 186355 169957 186356
rect 169155 185876 169221 185877
rect 169155 185812 169156 185876
rect 169220 185812 169221 185876
rect 169155 185811 169221 185812
rect 169155 185740 169221 185741
rect 169155 185676 169156 185740
rect 169220 185676 169221 185740
rect 169155 185675 169221 185676
rect 169158 89730 169218 185675
rect 169158 89670 169586 89730
rect 169155 80204 169221 80205
rect 169155 80140 169156 80204
rect 169220 80140 169221 80204
rect 169155 80139 169221 80140
rect 168971 79660 169037 79661
rect 168971 79596 168972 79660
rect 169036 79596 169037 79660
rect 168971 79595 169037 79596
rect 167315 79252 167381 79253
rect 167315 79188 167316 79252
rect 167380 79188 167381 79252
rect 167315 79187 167381 79188
rect 168051 79252 168117 79253
rect 168051 79188 168052 79252
rect 168116 79188 168117 79252
rect 168051 79187 168117 79188
rect 168235 79252 168301 79253
rect 168235 79188 168236 79252
rect 168300 79188 168301 79252
rect 168235 79187 168301 79188
rect 168603 79252 168669 79253
rect 168603 79188 168604 79252
rect 168668 79188 168669 79252
rect 168603 79187 168669 79188
rect 167867 78164 167933 78165
rect 167867 78100 167868 78164
rect 167932 78100 167933 78164
rect 167867 78099 167933 78100
rect 167683 73812 167749 73813
rect 167683 73748 167684 73812
rect 167748 73748 167749 73812
rect 167683 73747 167749 73748
rect 166947 71364 167013 71365
rect 166947 71300 166948 71364
rect 167012 71300 167013 71364
rect 166947 71299 167013 71300
rect 166950 70141 167010 71299
rect 166947 70140 167013 70141
rect 166947 70076 166948 70140
rect 167012 70076 167013 70140
rect 166947 70075 167013 70076
rect 167686 55997 167746 73747
rect 167683 55996 167749 55997
rect 167683 55932 167684 55996
rect 167748 55932 167749 55996
rect 167683 55931 167749 55932
rect 166763 50828 166829 50829
rect 166763 50764 166764 50828
rect 166828 50764 166829 50828
rect 166763 50763 166829 50764
rect 167870 49605 167930 78099
rect 168054 73541 168114 79187
rect 168051 73540 168117 73541
rect 168051 73476 168052 73540
rect 168116 73476 168117 73540
rect 168051 73475 168117 73476
rect 168051 73404 168117 73405
rect 168051 73340 168052 73404
rect 168116 73340 168117 73404
rect 168051 73339 168117 73340
rect 167867 49604 167933 49605
rect 167867 49540 167868 49604
rect 167932 49540 167933 49604
rect 167867 49539 167933 49540
rect 168054 44165 168114 73339
rect 168294 61954 168914 78000
rect 169158 69053 169218 80139
rect 169339 79796 169405 79797
rect 169339 79732 169340 79796
rect 169404 79732 169405 79796
rect 169339 79731 169405 79732
rect 169342 76122 169402 79731
rect 169526 79661 169586 89670
rect 169894 80205 169954 186355
rect 169891 80204 169957 80205
rect 169891 80140 169892 80204
rect 169956 80140 169957 80204
rect 169891 80139 169957 80140
rect 169707 79932 169773 79933
rect 169707 79868 169708 79932
rect 169772 79868 169773 79932
rect 169707 79867 169773 79868
rect 169523 79660 169589 79661
rect 169523 79596 169524 79660
rect 169588 79596 169589 79660
rect 169523 79595 169589 79596
rect 169342 76062 169586 76122
rect 169339 75988 169405 75989
rect 169339 75924 169340 75988
rect 169404 75924 169405 75988
rect 169339 75923 169405 75924
rect 169155 69052 169221 69053
rect 169155 68988 169156 69052
rect 169220 68988 169221 69052
rect 169155 68987 169221 68988
rect 168294 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 168914 61954
rect 168294 61634 168914 61718
rect 168294 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 168914 61634
rect 168051 44164 168117 44165
rect 168051 44100 168052 44164
rect 168116 44100 168117 44164
rect 168051 44099 168117 44100
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -4186 164414 20898
rect 163794 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 164414 -4186
rect 163794 -4506 164414 -4422
rect 163794 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 164414 -4506
rect 163794 -7654 164414 -4742
rect 168294 25954 168914 61398
rect 169342 52325 169402 75923
rect 169339 52324 169405 52325
rect 169339 52260 169340 52324
rect 169404 52260 169405 52324
rect 169339 52259 169405 52260
rect 169526 46885 169586 76062
rect 169710 72453 169770 79867
rect 170078 79661 170138 199683
rect 170998 186421 171058 199819
rect 170995 186420 171061 186421
rect 170995 186356 170996 186420
rect 171060 186356 171061 186420
rect 170995 186355 171061 186356
rect 170995 186284 171061 186285
rect 170995 186220 170996 186284
rect 171060 186220 171061 186284
rect 170995 186219 171061 186220
rect 170811 184924 170877 184925
rect 170811 184860 170812 184924
rect 170876 184860 170877 184924
rect 170811 184859 170877 184860
rect 170288 115954 170608 115986
rect 170288 115718 170330 115954
rect 170566 115718 170608 115954
rect 170288 115634 170608 115718
rect 170288 115398 170330 115634
rect 170566 115398 170608 115634
rect 170288 115366 170608 115398
rect 170814 80069 170874 184859
rect 170811 80068 170877 80069
rect 170811 80004 170812 80068
rect 170876 80004 170877 80068
rect 170811 80003 170877 80004
rect 170075 79660 170141 79661
rect 170075 79596 170076 79660
rect 170140 79596 170141 79660
rect 170075 79595 170141 79596
rect 170627 79660 170693 79661
rect 170627 79596 170628 79660
rect 170692 79596 170693 79660
rect 170627 79595 170693 79596
rect 170443 77348 170509 77349
rect 170443 77284 170444 77348
rect 170508 77284 170509 77348
rect 170443 77283 170509 77284
rect 169707 72452 169773 72453
rect 169707 72388 169708 72452
rect 169772 72388 169773 72452
rect 169707 72387 169773 72388
rect 170446 55861 170506 77283
rect 170443 55860 170509 55861
rect 170443 55796 170444 55860
rect 170508 55796 170509 55860
rect 170443 55795 170509 55796
rect 170630 52461 170690 79595
rect 170814 78165 170874 80003
rect 170998 79797 171058 186219
rect 171547 185604 171613 185605
rect 171547 185540 171548 185604
rect 171612 185540 171613 185604
rect 171547 185539 171613 185540
rect 171363 79932 171429 79933
rect 171363 79868 171364 79932
rect 171428 79868 171429 79932
rect 171363 79867 171429 79868
rect 170995 79796 171061 79797
rect 170995 79732 170996 79796
rect 171060 79732 171061 79796
rect 170995 79731 171061 79732
rect 171366 78437 171426 79867
rect 171550 79797 171610 185539
rect 171734 79933 171794 199819
rect 172651 199748 172717 199749
rect 172651 199684 172652 199748
rect 172716 199684 172717 199748
rect 172651 199683 172717 199684
rect 172283 185740 172349 185741
rect 172283 185676 172284 185740
rect 172348 185676 172349 185740
rect 172283 185675 172349 185676
rect 172099 185604 172165 185605
rect 172099 185540 172100 185604
rect 172164 185540 172165 185604
rect 172099 185539 172165 185540
rect 171915 81156 171981 81157
rect 171915 81092 171916 81156
rect 171980 81092 171981 81156
rect 171915 81091 171981 81092
rect 171918 79933 171978 81091
rect 171731 79932 171797 79933
rect 171731 79868 171732 79932
rect 171796 79868 171797 79932
rect 171731 79867 171797 79868
rect 171915 79932 171981 79933
rect 171915 79868 171916 79932
rect 171980 79868 171981 79932
rect 171915 79867 171981 79868
rect 171547 79796 171613 79797
rect 171547 79732 171548 79796
rect 171612 79732 171613 79796
rect 171547 79731 171613 79732
rect 171734 79253 171794 79867
rect 171731 79252 171797 79253
rect 171731 79188 171732 79252
rect 171796 79188 171797 79252
rect 171731 79187 171797 79188
rect 171918 78845 171978 79867
rect 172102 79797 172162 185539
rect 172099 79796 172165 79797
rect 172099 79732 172100 79796
rect 172164 79732 172165 79796
rect 172099 79731 172165 79732
rect 172286 79389 172346 185675
rect 172467 81292 172533 81293
rect 172467 81228 172468 81292
rect 172532 81228 172533 81292
rect 172467 81227 172533 81228
rect 172470 79933 172530 81227
rect 172467 79932 172533 79933
rect 172467 79868 172468 79932
rect 172532 79868 172533 79932
rect 172467 79867 172533 79868
rect 172283 79388 172349 79389
rect 172283 79324 172284 79388
rect 172348 79324 172349 79388
rect 172283 79323 172349 79324
rect 172283 79252 172349 79253
rect 172283 79188 172284 79252
rect 172348 79188 172349 79252
rect 172283 79187 172349 79188
rect 171915 78844 171981 78845
rect 171915 78780 171916 78844
rect 171980 78780 171981 78844
rect 171915 78779 171981 78780
rect 171363 78436 171429 78437
rect 171363 78372 171364 78436
rect 171428 78372 171429 78436
rect 171363 78371 171429 78372
rect 170811 78164 170877 78165
rect 170811 78100 170812 78164
rect 170876 78100 170877 78164
rect 170811 78099 170877 78100
rect 170811 77484 170877 77485
rect 170811 77420 170812 77484
rect 170876 77420 170877 77484
rect 170811 77419 170877 77420
rect 170627 52460 170693 52461
rect 170627 52396 170628 52460
rect 170692 52396 170693 52460
rect 170627 52395 170693 52396
rect 170814 49469 170874 77419
rect 170995 77348 171061 77349
rect 170995 77284 170996 77348
rect 171060 77284 171061 77348
rect 170995 77283 171061 77284
rect 170811 49468 170877 49469
rect 170811 49404 170812 49468
rect 170876 49404 170877 49468
rect 170811 49403 170877 49404
rect 169523 46884 169589 46885
rect 169523 46820 169524 46884
rect 169588 46820 169589 46884
rect 169523 46819 169589 46820
rect 170998 46749 171058 77283
rect 172099 76124 172165 76125
rect 172099 76060 172100 76124
rect 172164 76060 172165 76124
rect 172099 76059 172165 76060
rect 171915 75988 171981 75989
rect 171915 75924 171916 75988
rect 171980 75924 171981 75988
rect 171915 75923 171981 75924
rect 171918 64565 171978 75923
rect 171915 64564 171981 64565
rect 171915 64500 171916 64564
rect 171980 64500 171981 64564
rect 171915 64499 171981 64500
rect 172102 62933 172162 76059
rect 172099 62932 172165 62933
rect 172099 62868 172100 62932
rect 172164 62868 172165 62932
rect 172099 62867 172165 62868
rect 170995 46748 171061 46749
rect 170995 46684 170996 46748
rect 171060 46684 171061 46748
rect 170995 46683 171061 46684
rect 172286 42805 172346 79187
rect 172470 77757 172530 79867
rect 172654 78845 172714 199683
rect 172838 79797 172898 199819
rect 173387 199748 173453 199749
rect 173387 199684 173388 199748
rect 173452 199684 173453 199748
rect 173387 199683 173453 199684
rect 174123 199748 174189 199749
rect 174123 199684 174124 199748
rect 174188 199684 174189 199748
rect 174123 199683 174189 199684
rect 173390 186149 173450 199683
rect 173387 186148 173453 186149
rect 173387 186084 173388 186148
rect 173452 186084 173453 186148
rect 173387 186083 173453 186084
rect 173203 186012 173269 186013
rect 173203 185948 173204 186012
rect 173268 185948 173269 186012
rect 173203 185947 173269 185948
rect 173019 185604 173085 185605
rect 173019 185540 173020 185604
rect 173084 185540 173085 185604
rect 173019 185539 173085 185540
rect 172835 79796 172901 79797
rect 172835 79732 172836 79796
rect 172900 79732 172901 79796
rect 172835 79731 172901 79732
rect 173022 79389 173082 185539
rect 173206 93870 173266 185947
rect 173939 140180 174005 140181
rect 173939 140116 173940 140180
rect 174004 140116 174005 140180
rect 173939 140115 174005 140116
rect 173942 139773 174002 140115
rect 173939 139772 174005 139773
rect 173939 139708 173940 139772
rect 174004 139708 174005 139772
rect 173939 139707 174005 139708
rect 173206 93810 173634 93870
rect 173203 80340 173269 80341
rect 173203 80276 173204 80340
rect 173268 80276 173269 80340
rect 173203 80275 173269 80276
rect 173019 79388 173085 79389
rect 173019 79324 173020 79388
rect 173084 79324 173085 79388
rect 173019 79323 173085 79324
rect 173206 78981 173266 80275
rect 173574 78981 173634 93810
rect 174126 86970 174186 199683
rect 174307 186284 174373 186285
rect 174307 186220 174308 186284
rect 174372 186220 174373 186284
rect 174307 186219 174373 186220
rect 173942 86910 174186 86970
rect 173755 80068 173821 80069
rect 173755 80004 173756 80068
rect 173820 80004 173821 80068
rect 173755 80003 173821 80004
rect 173203 78980 173269 78981
rect 173203 78916 173204 78980
rect 173268 78916 173269 78980
rect 173203 78915 173269 78916
rect 173571 78980 173637 78981
rect 173571 78916 173572 78980
rect 173636 78916 173637 78980
rect 173571 78915 173637 78916
rect 172651 78844 172717 78845
rect 172651 78780 172652 78844
rect 172716 78780 172717 78844
rect 172651 78779 172717 78780
rect 173758 78029 173818 80003
rect 173755 78028 173821 78029
rect 172467 77756 172533 77757
rect 172467 77692 172468 77756
rect 172532 77692 172533 77756
rect 172467 77691 172533 77692
rect 172794 66454 173414 78000
rect 173755 77964 173756 78028
rect 173820 77964 173821 78028
rect 173755 77963 173821 77964
rect 173942 77621 174002 86910
rect 174310 79933 174370 186219
rect 174307 79932 174373 79933
rect 174307 79868 174308 79932
rect 174372 79868 174373 79932
rect 174307 79867 174373 79868
rect 174494 79389 174554 199819
rect 175046 79933 175106 199819
rect 175414 192677 175474 199819
rect 175595 199748 175661 199749
rect 175595 199684 175596 199748
rect 175660 199684 175661 199748
rect 175595 199683 175661 199684
rect 175779 199748 175845 199749
rect 175779 199684 175780 199748
rect 175844 199684 175845 199748
rect 175779 199683 175845 199684
rect 175411 192676 175477 192677
rect 175411 192612 175412 192676
rect 175476 192612 175477 192676
rect 175411 192611 175477 192612
rect 175598 180845 175658 199683
rect 175595 180844 175661 180845
rect 175595 180780 175596 180844
rect 175660 180780 175661 180844
rect 175595 180779 175661 180780
rect 175782 79933 175842 199683
rect 175963 185876 176029 185877
rect 175963 185812 175964 185876
rect 176028 185812 176029 185876
rect 175963 185811 176029 185812
rect 175043 79932 175109 79933
rect 175043 79868 175044 79932
rect 175108 79868 175109 79932
rect 175043 79867 175109 79868
rect 175411 79932 175477 79933
rect 175411 79868 175412 79932
rect 175476 79868 175477 79932
rect 175411 79867 175477 79868
rect 175779 79932 175845 79933
rect 175779 79868 175780 79932
rect 175844 79868 175845 79932
rect 175779 79867 175845 79868
rect 175043 79796 175109 79797
rect 175043 79732 175044 79796
rect 175108 79732 175109 79796
rect 175043 79731 175109 79732
rect 174491 79388 174557 79389
rect 174491 79324 174492 79388
rect 174556 79324 174557 79388
rect 174491 79323 174557 79324
rect 174494 78845 174554 79323
rect 174491 78844 174557 78845
rect 174491 78780 174492 78844
rect 174556 78780 174557 78844
rect 174491 78779 174557 78780
rect 174675 78708 174741 78709
rect 174675 78644 174676 78708
rect 174740 78644 174741 78708
rect 174675 78643 174741 78644
rect 173939 77620 174005 77621
rect 173939 77556 173940 77620
rect 174004 77556 174005 77620
rect 173939 77555 174005 77556
rect 173571 76124 173637 76125
rect 173571 76060 173572 76124
rect 173636 76060 173637 76124
rect 173571 76059 173637 76060
rect 172794 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 173414 66454
rect 172794 66134 173414 66218
rect 172794 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 173414 66134
rect 172283 42804 172349 42805
rect 172283 42740 172284 42804
rect 172348 42740 172349 42804
rect 172283 42739 172349 42740
rect 168294 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 168914 25954
rect 168294 25634 168914 25718
rect 168294 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 168914 25634
rect 168294 -5146 168914 25398
rect 168294 -5382 168326 -5146
rect 168562 -5382 168646 -5146
rect 168882 -5382 168914 -5146
rect 168294 -5466 168914 -5382
rect 168294 -5702 168326 -5466
rect 168562 -5702 168646 -5466
rect 168882 -5702 168914 -5466
rect 168294 -7654 168914 -5702
rect 172794 30454 173414 65898
rect 173574 60349 173634 76059
rect 173755 73812 173821 73813
rect 173755 73748 173756 73812
rect 173820 73748 173821 73812
rect 173755 73747 173821 73748
rect 173571 60348 173637 60349
rect 173571 60284 173572 60348
rect 173636 60284 173637 60348
rect 173571 60283 173637 60284
rect 173758 48109 173818 73747
rect 174678 64701 174738 78643
rect 174859 75852 174925 75853
rect 174859 75788 174860 75852
rect 174924 75788 174925 75852
rect 174859 75787 174925 75788
rect 174675 64700 174741 64701
rect 174675 64636 174676 64700
rect 174740 64636 174741 64700
rect 174675 64635 174741 64636
rect 174862 58989 174922 75787
rect 174859 58988 174925 58989
rect 174859 58924 174860 58988
rect 174924 58924 174925 58988
rect 174859 58923 174925 58924
rect 175046 57629 175106 79731
rect 175414 76261 175474 79867
rect 175782 78709 175842 79867
rect 175966 79797 176026 185811
rect 176150 79933 176210 199822
rect 176515 199820 176516 199822
rect 176580 199820 176581 199884
rect 176515 199819 176581 199820
rect 178171 199068 178237 199069
rect 178171 199004 178172 199068
rect 178236 199004 178237 199068
rect 178171 199003 178237 199004
rect 176515 186284 176581 186285
rect 176515 186220 176516 186284
rect 176580 186220 176581 186284
rect 176515 186219 176581 186220
rect 176883 186284 176949 186285
rect 176883 186220 176884 186284
rect 176948 186220 176949 186284
rect 176883 186219 176949 186220
rect 176147 79932 176213 79933
rect 176147 79868 176148 79932
rect 176212 79868 176213 79932
rect 176147 79867 176213 79868
rect 176518 79797 176578 186219
rect 176886 79933 176946 186219
rect 177294 178954 177914 198000
rect 177294 178718 177326 178954
rect 177562 178718 177646 178954
rect 177882 178718 177914 178954
rect 177294 178634 177914 178718
rect 177294 178398 177326 178634
rect 177562 178398 177646 178634
rect 177882 178398 177914 178634
rect 177067 176628 177133 176629
rect 177067 176564 177068 176628
rect 177132 176564 177133 176628
rect 177067 176563 177133 176564
rect 176883 79932 176949 79933
rect 176883 79868 176884 79932
rect 176948 79868 176949 79932
rect 176883 79867 176949 79868
rect 177070 79797 177130 176563
rect 177294 142954 177914 178398
rect 177294 142718 177326 142954
rect 177562 142718 177646 142954
rect 177882 142718 177914 142954
rect 177294 142634 177914 142718
rect 177294 142398 177326 142634
rect 177562 142398 177646 142634
rect 177882 142398 177914 142634
rect 177294 142000 177914 142398
rect 177619 141676 177685 141677
rect 177619 141612 177620 141676
rect 177684 141612 177685 141676
rect 177619 141611 177685 141612
rect 177251 141268 177317 141269
rect 177251 141204 177252 141268
rect 177316 141204 177317 141268
rect 177251 141203 177317 141204
rect 177254 80749 177314 141203
rect 177251 80748 177317 80749
rect 177251 80684 177252 80748
rect 177316 80684 177317 80748
rect 177251 80683 177317 80684
rect 175917 79796 176026 79797
rect 175917 79732 175918 79796
rect 175982 79734 176026 79796
rect 176147 79796 176213 79797
rect 175982 79732 175983 79734
rect 175917 79731 175983 79732
rect 176147 79732 176148 79796
rect 176212 79732 176213 79796
rect 176147 79731 176213 79732
rect 176515 79796 176581 79797
rect 176515 79732 176516 79796
rect 176580 79732 176581 79796
rect 176515 79731 176581 79732
rect 177067 79796 177133 79797
rect 177067 79732 177068 79796
rect 177132 79732 177133 79796
rect 177067 79731 177133 79732
rect 176150 79658 176210 79731
rect 177067 79660 177133 79661
rect 176150 79598 176578 79658
rect 176147 79388 176213 79389
rect 176147 79324 176148 79388
rect 176212 79324 176213 79388
rect 176147 79323 176213 79324
rect 175779 78708 175845 78709
rect 175779 78644 175780 78708
rect 175844 78644 175845 78708
rect 175779 78643 175845 78644
rect 175963 78708 176029 78709
rect 175963 78644 175964 78708
rect 176028 78644 176029 78708
rect 175963 78643 176029 78644
rect 175411 76260 175477 76261
rect 175411 76196 175412 76260
rect 175476 76196 175477 76260
rect 175411 76195 175477 76196
rect 175043 57628 175109 57629
rect 175043 57564 175044 57628
rect 175108 57564 175109 57628
rect 175043 57563 175109 57564
rect 175966 49333 176026 78643
rect 176150 66741 176210 79323
rect 176331 77892 176397 77893
rect 176331 77828 176332 77892
rect 176396 77828 176397 77892
rect 176331 77827 176397 77828
rect 176147 66740 176213 66741
rect 176147 66676 176148 66740
rect 176212 66676 176213 66740
rect 176147 66675 176213 66676
rect 176334 62797 176394 77827
rect 176518 75717 176578 79598
rect 177067 79596 177068 79660
rect 177132 79596 177133 79660
rect 177067 79595 177133 79596
rect 176515 75716 176581 75717
rect 176515 75652 176516 75716
rect 176580 75652 176581 75716
rect 176515 75651 176581 75652
rect 176331 62796 176397 62797
rect 176331 62732 176332 62796
rect 176396 62732 176397 62796
rect 176331 62731 176397 62732
rect 177070 50285 177130 79595
rect 177254 79389 177314 80683
rect 177622 79933 177682 141611
rect 177619 79932 177685 79933
rect 177619 79868 177620 79932
rect 177684 79868 177685 79932
rect 177619 79867 177685 79868
rect 178174 79797 178234 199003
rect 179459 197572 179525 197573
rect 179459 197508 179460 197572
rect 179524 197508 179525 197572
rect 179459 197507 179525 197508
rect 178355 193356 178421 193357
rect 178355 193292 178356 193356
rect 178420 193292 178421 193356
rect 178355 193291 178421 193292
rect 178358 80749 178418 193291
rect 178539 190500 178605 190501
rect 178539 190436 178540 190500
rect 178604 190436 178605 190500
rect 178539 190435 178605 190436
rect 178355 80748 178421 80749
rect 178355 80684 178356 80748
rect 178420 80684 178421 80748
rect 178355 80683 178421 80684
rect 178542 80477 178602 190435
rect 178723 140180 178789 140181
rect 178723 140116 178724 140180
rect 178788 140116 178789 140180
rect 178723 140115 178789 140116
rect 178539 80476 178605 80477
rect 178539 80412 178540 80476
rect 178604 80412 178605 80476
rect 178539 80411 178605 80412
rect 178171 79796 178237 79797
rect 178171 79732 178172 79796
rect 178236 79732 178237 79796
rect 178171 79731 178237 79732
rect 178542 79661 178602 80411
rect 178539 79660 178605 79661
rect 178539 79596 178540 79660
rect 178604 79596 178605 79660
rect 178539 79595 178605 79596
rect 177251 79388 177317 79389
rect 177251 79324 177252 79388
rect 177316 79324 177317 79388
rect 177251 79323 177317 79324
rect 177294 70954 177914 78000
rect 178726 77213 178786 140115
rect 178723 77212 178789 77213
rect 178723 77148 178724 77212
rect 178788 77148 178789 77212
rect 178723 77147 178789 77148
rect 177294 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 177914 70954
rect 177294 70634 177914 70718
rect 177294 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 177914 70634
rect 177067 50284 177133 50285
rect 177067 50220 177068 50284
rect 177132 50220 177133 50284
rect 177067 50219 177133 50220
rect 175963 49332 176029 49333
rect 175963 49268 175964 49332
rect 176028 49268 176029 49332
rect 175963 49267 176029 49268
rect 173755 48108 173821 48109
rect 173755 48044 173756 48108
rect 173820 48044 173821 48108
rect 173755 48043 173821 48044
rect 172794 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 173414 30454
rect 172794 30134 173414 30218
rect 172794 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 173414 30134
rect 172794 -6106 173414 29898
rect 172794 -6342 172826 -6106
rect 173062 -6342 173146 -6106
rect 173382 -6342 173414 -6106
rect 172794 -6426 173414 -6342
rect 172794 -6662 172826 -6426
rect 173062 -6662 173146 -6426
rect 173382 -6662 173414 -6426
rect 172794 -7654 173414 -6662
rect 177294 34954 177914 70398
rect 179462 68781 179522 197507
rect 179643 193084 179709 193085
rect 179643 193020 179644 193084
rect 179708 193020 179709 193084
rect 179643 193019 179709 193020
rect 179646 73133 179706 193019
rect 179830 151830 179890 200635
rect 182955 200564 183021 200565
rect 182955 200500 182956 200564
rect 183020 200500 183021 200564
rect 182955 200499 183021 200500
rect 180747 199612 180813 199613
rect 180747 199548 180748 199612
rect 180812 199548 180813 199612
rect 180747 199547 180813 199548
rect 180750 186330 180810 199547
rect 182587 199476 182653 199477
rect 182587 199412 182588 199476
rect 182652 199412 182653 199476
rect 182587 199411 182653 199412
rect 180931 192948 180997 192949
rect 180931 192884 180932 192948
rect 180996 192884 180997 192948
rect 180931 192883 180997 192884
rect 180566 186270 180810 186330
rect 179830 151770 180258 151830
rect 179827 140044 179893 140045
rect 179827 139980 179828 140044
rect 179892 139980 179893 140044
rect 179827 139979 179893 139980
rect 179643 73132 179709 73133
rect 179643 73068 179644 73132
rect 179708 73068 179709 73132
rect 179643 73067 179709 73068
rect 179830 72725 179890 139979
rect 180011 139772 180077 139773
rect 180011 139708 180012 139772
rect 180076 139708 180077 139772
rect 180011 139707 180077 139708
rect 180014 80885 180074 139707
rect 180198 139501 180258 151770
rect 180195 139500 180261 139501
rect 180195 139436 180196 139500
rect 180260 139436 180261 139500
rect 180195 139435 180261 139436
rect 180566 118710 180626 186270
rect 180566 118650 180810 118710
rect 180750 109050 180810 118650
rect 180566 108990 180810 109050
rect 180566 89730 180626 108990
rect 180566 89670 180810 89730
rect 180011 80884 180077 80885
rect 180011 80820 180012 80884
rect 180076 80820 180077 80884
rect 180011 80819 180077 80820
rect 179827 72724 179893 72725
rect 179827 72660 179828 72724
rect 179892 72660 179893 72724
rect 179827 72659 179893 72660
rect 180750 70410 180810 89670
rect 180934 73133 180994 192883
rect 181794 183454 182414 198000
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181115 150380 181181 150381
rect 181115 150316 181116 150380
rect 181180 150316 181181 150380
rect 181115 150315 181181 150316
rect 181118 74357 181178 150315
rect 181794 147454 182414 182898
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181299 146980 181365 146981
rect 181299 146916 181300 146980
rect 181364 146916 181365 146980
rect 181299 146915 181365 146916
rect 181302 93870 181362 146915
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 142000 182414 146898
rect 181302 93810 181546 93870
rect 181486 77077 181546 93810
rect 181483 77076 181549 77077
rect 181483 77012 181484 77076
rect 181548 77012 181549 77076
rect 181483 77011 181549 77012
rect 181794 75454 182414 78000
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181115 74356 181181 74357
rect 181115 74292 181116 74356
rect 181180 74292 181181 74356
rect 181115 74291 181181 74292
rect 180931 73132 180997 73133
rect 180931 73068 180932 73132
rect 180996 73068 180997 73132
rect 180931 73067 180997 73068
rect 180566 70350 180810 70410
rect 179459 68780 179525 68781
rect 179459 68716 179460 68780
rect 179524 68716 179525 68780
rect 179459 68715 179525 68716
rect 180566 61301 180626 70350
rect 180563 61300 180629 61301
rect 180563 61236 180564 61300
rect 180628 61236 180629 61300
rect 180563 61235 180629 61236
rect 177294 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 177914 34954
rect 177294 34634 177914 34718
rect 177294 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 177914 34634
rect 177294 -7066 177914 34398
rect 177294 -7302 177326 -7066
rect 177562 -7302 177646 -7066
rect 177882 -7302 177914 -7066
rect 177294 -7386 177914 -7302
rect 177294 -7622 177326 -7386
rect 177562 -7622 177646 -7386
rect 177882 -7622 177914 -7386
rect 177294 -7654 177914 -7622
rect 181794 39454 182414 74898
rect 182590 67421 182650 199411
rect 182771 149836 182837 149837
rect 182771 149772 182772 149836
rect 182836 149772 182837 149836
rect 182771 149771 182837 149772
rect 182587 67420 182653 67421
rect 182587 67356 182588 67420
rect 182652 67356 182653 67420
rect 182587 67355 182653 67356
rect 182774 53549 182834 149771
rect 182958 144805 183018 200499
rect 183507 199340 183573 199341
rect 183507 199276 183508 199340
rect 183572 199276 183573 199340
rect 183507 199275 183573 199276
rect 183139 147116 183205 147117
rect 183139 147052 183140 147116
rect 183204 147052 183205 147116
rect 183139 147051 183205 147052
rect 182955 144804 183021 144805
rect 182955 144740 182956 144804
rect 183020 144740 183021 144804
rect 182955 144739 183021 144740
rect 183142 72861 183202 147051
rect 183323 140044 183389 140045
rect 183323 139980 183324 140044
rect 183388 139980 183389 140044
rect 183323 139979 183389 139980
rect 183326 138957 183386 139979
rect 183323 138956 183389 138957
rect 183323 138892 183324 138956
rect 183388 138892 183389 138956
rect 183323 138891 183389 138892
rect 183510 73170 183570 199275
rect 183691 196892 183757 196893
rect 183691 196828 183692 196892
rect 183756 196828 183757 196892
rect 183691 196827 183757 196828
rect 183694 80341 183754 196827
rect 184979 194036 185045 194037
rect 184979 193972 184980 194036
rect 185044 193972 185045 194036
rect 184979 193971 185045 193972
rect 183875 150244 183941 150245
rect 183875 150180 183876 150244
rect 183940 150180 183941 150244
rect 183875 150179 183941 150180
rect 183878 86970 183938 150179
rect 184795 140044 184861 140045
rect 184795 139980 184796 140044
rect 184860 139980 184861 140044
rect 184795 139979 184861 139980
rect 184798 138549 184858 139979
rect 184795 138548 184861 138549
rect 184795 138484 184796 138548
rect 184860 138484 184861 138548
rect 184795 138483 184861 138484
rect 183878 86910 184122 86970
rect 183691 80340 183757 80341
rect 183691 80276 183692 80340
rect 183756 80276 183757 80340
rect 183691 80275 183757 80276
rect 184062 73170 184122 86910
rect 184982 78573 185042 193971
rect 185347 152692 185413 152693
rect 185347 152628 185348 152692
rect 185412 152628 185413 152692
rect 185347 152627 185413 152628
rect 185163 152556 185229 152557
rect 185163 152492 185164 152556
rect 185228 152492 185229 152556
rect 185163 152491 185229 152492
rect 184979 78572 185045 78573
rect 184979 78508 184980 78572
rect 185044 78508 185045 78572
rect 184979 78507 185045 78508
rect 183510 73110 183754 73170
rect 183139 72860 183205 72861
rect 183139 72796 183140 72860
rect 183204 72796 183205 72860
rect 183139 72795 183205 72796
rect 183694 62117 183754 73110
rect 183878 73110 184122 73170
rect 183878 72997 183938 73110
rect 183875 72996 183941 72997
rect 183875 72932 183876 72996
rect 183940 72932 183941 72996
rect 183875 72931 183941 72932
rect 185166 72589 185226 152491
rect 185350 81973 185410 152627
rect 186086 140317 186146 202811
rect 186294 187954 186914 198000
rect 186294 187718 186326 187954
rect 186562 187718 186646 187954
rect 186882 187718 186914 187954
rect 186294 187634 186914 187718
rect 186294 187398 186326 187634
rect 186562 187398 186646 187634
rect 186882 187398 186914 187634
rect 186294 151954 186914 187398
rect 186294 151718 186326 151954
rect 186562 151718 186646 151954
rect 186882 151718 186914 151954
rect 186294 151634 186914 151718
rect 186294 151398 186326 151634
rect 186562 151398 186646 151634
rect 186882 151398 186914 151634
rect 186294 142000 186914 151398
rect 187006 149157 187066 270539
rect 188107 262308 188173 262309
rect 188107 262244 188108 262308
rect 188172 262244 188173 262308
rect 188107 262243 188173 262244
rect 187739 196756 187805 196757
rect 187739 196692 187740 196756
rect 187804 196692 187805 196756
rect 187739 196691 187805 196692
rect 187187 195668 187253 195669
rect 187187 195604 187188 195668
rect 187252 195604 187253 195668
rect 187187 195603 187253 195604
rect 187003 149156 187069 149157
rect 187003 149092 187004 149156
rect 187068 149092 187069 149156
rect 187003 149091 187069 149092
rect 186819 140860 186885 140861
rect 186819 140796 186820 140860
rect 186884 140796 186885 140860
rect 186819 140795 186885 140796
rect 186083 140316 186149 140317
rect 186083 140252 186084 140316
rect 186148 140252 186149 140316
rect 186083 140251 186149 140252
rect 186083 139908 186149 139909
rect 186083 139844 186084 139908
rect 186148 139844 186149 139908
rect 186083 139843 186149 139844
rect 186086 137461 186146 139843
rect 186083 137460 186149 137461
rect 186083 137396 186084 137460
rect 186148 137396 186149 137460
rect 186083 137395 186149 137396
rect 185648 111454 185968 111486
rect 185648 111218 185690 111454
rect 185926 111218 185968 111454
rect 185648 111134 185968 111218
rect 185648 110898 185690 111134
rect 185926 110898 185968 111134
rect 185648 110866 185968 110898
rect 185347 81972 185413 81973
rect 185347 81908 185348 81972
rect 185412 81908 185413 81972
rect 185347 81907 185413 81908
rect 186822 78573 186882 140795
rect 187003 138140 187069 138141
rect 187003 138076 187004 138140
rect 187068 138076 187069 138140
rect 187003 138075 187069 138076
rect 186819 78572 186885 78573
rect 186819 78508 186820 78572
rect 186884 78508 186885 78572
rect 186819 78507 186885 78508
rect 185163 72588 185229 72589
rect 185163 72524 185164 72588
rect 185228 72524 185229 72588
rect 185163 72523 185229 72524
rect 183691 62116 183757 62117
rect 183691 62052 183692 62116
rect 183756 62052 183757 62116
rect 183691 62051 183757 62052
rect 182771 53548 182837 53549
rect 182771 53484 182772 53548
rect 182836 53484 182837 53548
rect 182771 53483 182837 53484
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -7654 182414 -902
rect 186294 43954 186914 78000
rect 187006 44029 187066 138075
rect 187190 81021 187250 195603
rect 187371 149700 187437 149701
rect 187371 149636 187372 149700
rect 187436 149636 187437 149700
rect 187371 149635 187437 149636
rect 187187 81020 187253 81021
rect 187187 80956 187188 81020
rect 187252 80956 187253 81020
rect 187187 80955 187253 80956
rect 187374 78573 187434 149635
rect 187371 78572 187437 78573
rect 187371 78508 187372 78572
rect 187436 78508 187437 78572
rect 187371 78507 187437 78508
rect 187742 61981 187802 196691
rect 187923 196620 187989 196621
rect 187923 196556 187924 196620
rect 187988 196556 187989 196620
rect 187923 196555 187989 196556
rect 187926 66197 187986 196555
rect 188110 144125 188170 262243
rect 188291 148340 188357 148341
rect 188291 148276 188292 148340
rect 188356 148276 188357 148340
rect 188291 148275 188357 148276
rect 188107 144124 188173 144125
rect 188107 144060 188108 144124
rect 188172 144060 188173 144124
rect 188107 144059 188173 144060
rect 188107 141132 188173 141133
rect 188107 141068 188108 141132
rect 188172 141068 188173 141132
rect 188107 141067 188173 141068
rect 188110 66197 188170 141067
rect 188294 68781 188354 148275
rect 189030 142490 189090 275979
rect 190794 264454 191414 299898
rect 195294 707718 195914 711590
rect 195294 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 195914 707718
rect 195294 707398 195914 707482
rect 195294 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 195914 707398
rect 195294 700954 195914 707162
rect 195294 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 195914 700954
rect 195294 700634 195914 700718
rect 195294 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 195914 700634
rect 195294 664954 195914 700398
rect 195294 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 195914 664954
rect 195294 664634 195914 664718
rect 195294 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 195914 664634
rect 195294 628954 195914 664398
rect 195294 628718 195326 628954
rect 195562 628718 195646 628954
rect 195882 628718 195914 628954
rect 195294 628634 195914 628718
rect 195294 628398 195326 628634
rect 195562 628398 195646 628634
rect 195882 628398 195914 628634
rect 195294 592954 195914 628398
rect 195294 592718 195326 592954
rect 195562 592718 195646 592954
rect 195882 592718 195914 592954
rect 195294 592634 195914 592718
rect 195294 592398 195326 592634
rect 195562 592398 195646 592634
rect 195882 592398 195914 592634
rect 195294 556954 195914 592398
rect 195294 556718 195326 556954
rect 195562 556718 195646 556954
rect 195882 556718 195914 556954
rect 195294 556634 195914 556718
rect 195294 556398 195326 556634
rect 195562 556398 195646 556634
rect 195882 556398 195914 556634
rect 195294 520954 195914 556398
rect 195294 520718 195326 520954
rect 195562 520718 195646 520954
rect 195882 520718 195914 520954
rect 195294 520634 195914 520718
rect 195294 520398 195326 520634
rect 195562 520398 195646 520634
rect 195882 520398 195914 520634
rect 195294 484954 195914 520398
rect 195294 484718 195326 484954
rect 195562 484718 195646 484954
rect 195882 484718 195914 484954
rect 195294 484634 195914 484718
rect 195294 484398 195326 484634
rect 195562 484398 195646 484634
rect 195882 484398 195914 484634
rect 195294 448954 195914 484398
rect 195294 448718 195326 448954
rect 195562 448718 195646 448954
rect 195882 448718 195914 448954
rect 195294 448634 195914 448718
rect 195294 448398 195326 448634
rect 195562 448398 195646 448634
rect 195882 448398 195914 448634
rect 195294 412954 195914 448398
rect 195294 412718 195326 412954
rect 195562 412718 195646 412954
rect 195882 412718 195914 412954
rect 195294 412634 195914 412718
rect 195294 412398 195326 412634
rect 195562 412398 195646 412634
rect 195882 412398 195914 412634
rect 195294 376954 195914 412398
rect 195294 376718 195326 376954
rect 195562 376718 195646 376954
rect 195882 376718 195914 376954
rect 195294 376634 195914 376718
rect 195294 376398 195326 376634
rect 195562 376398 195646 376634
rect 195882 376398 195914 376634
rect 195294 340954 195914 376398
rect 195294 340718 195326 340954
rect 195562 340718 195646 340954
rect 195882 340718 195914 340954
rect 195294 340634 195914 340718
rect 195294 340398 195326 340634
rect 195562 340398 195646 340634
rect 195882 340398 195914 340634
rect 195294 304954 195914 340398
rect 195294 304718 195326 304954
rect 195562 304718 195646 304954
rect 195882 304718 195914 304954
rect 195294 304634 195914 304718
rect 195294 304398 195326 304634
rect 195562 304398 195646 304634
rect 195882 304398 195914 304634
rect 195294 268954 195914 304398
rect 195294 268718 195326 268954
rect 195562 268718 195646 268954
rect 195882 268718 195914 268954
rect 195294 268634 195914 268718
rect 195294 268398 195326 268634
rect 195562 268398 195646 268634
rect 195882 268398 195914 268634
rect 193259 265300 193325 265301
rect 193259 265236 193260 265300
rect 193324 265236 193325 265300
rect 193259 265235 193325 265236
rect 190794 264218 190826 264454
rect 191062 264218 191146 264454
rect 191382 264218 191414 264454
rect 190794 264134 191414 264218
rect 190794 263898 190826 264134
rect 191062 263898 191146 264134
rect 191382 263898 191414 264134
rect 190499 262444 190565 262445
rect 190499 262380 190500 262444
rect 190564 262380 190565 262444
rect 190499 262379 190565 262380
rect 189211 199748 189277 199749
rect 189211 199684 189212 199748
rect 189276 199684 189277 199748
rect 189211 199683 189277 199684
rect 188846 142430 189090 142490
rect 188846 142085 188906 142430
rect 189027 142220 189093 142221
rect 189027 142156 189028 142220
rect 189092 142156 189093 142220
rect 189027 142155 189093 142156
rect 188843 142084 188909 142085
rect 188843 142020 188844 142084
rect 188908 142020 188909 142084
rect 188843 142019 188909 142020
rect 189030 137325 189090 142155
rect 189027 137324 189093 137325
rect 189027 137260 189028 137324
rect 189092 137260 189093 137324
rect 189027 137259 189093 137260
rect 189214 79253 189274 199683
rect 189395 147524 189461 147525
rect 189395 147460 189396 147524
rect 189460 147460 189461 147524
rect 189395 147459 189461 147460
rect 189211 79252 189277 79253
rect 189211 79188 189212 79252
rect 189276 79188 189277 79252
rect 189211 79187 189277 79188
rect 189398 76533 189458 147459
rect 190502 144261 190562 262379
rect 190794 262000 191414 263898
rect 191971 263124 192037 263125
rect 191971 263060 191972 263124
rect 192036 263060 192037 263124
rect 191971 263059 192037 263060
rect 191787 262580 191853 262581
rect 191787 262516 191788 262580
rect 191852 262516 191853 262580
rect 191787 262515 191853 262516
rect 190794 192454 191414 198000
rect 190794 192218 190826 192454
rect 191062 192218 191146 192454
rect 191382 192218 191414 192454
rect 190794 192134 191414 192218
rect 190794 191898 190826 192134
rect 191062 191898 191146 192134
rect 191382 191898 191414 192134
rect 190794 156454 191414 191898
rect 190794 156218 190826 156454
rect 191062 156218 191146 156454
rect 191382 156218 191414 156454
rect 190794 156134 191414 156218
rect 190794 155898 190826 156134
rect 191062 155898 191146 156134
rect 191382 155898 191414 156134
rect 190499 144260 190565 144261
rect 190499 144196 190500 144260
rect 190564 144196 190565 144260
rect 190499 144195 190565 144196
rect 190499 143580 190565 143581
rect 190499 143516 190500 143580
rect 190564 143516 190565 143580
rect 190499 143515 190565 143516
rect 189579 141268 189645 141269
rect 189579 141204 189580 141268
rect 189644 141204 189645 141268
rect 189579 141203 189645 141204
rect 189395 76532 189461 76533
rect 189395 76468 189396 76532
rect 189460 76468 189461 76532
rect 189395 76467 189461 76468
rect 188291 68780 188357 68781
rect 188291 68716 188292 68780
rect 188356 68716 188357 68780
rect 188291 68715 188357 68716
rect 187923 66196 187989 66197
rect 187923 66132 187924 66196
rect 187988 66132 187989 66196
rect 187923 66131 187989 66132
rect 188107 66196 188173 66197
rect 188107 66132 188108 66196
rect 188172 66132 188173 66196
rect 188107 66131 188173 66132
rect 187926 65653 187986 66131
rect 187923 65652 187989 65653
rect 187923 65588 187924 65652
rect 187988 65588 187989 65652
rect 187923 65587 187989 65588
rect 188110 65109 188170 66131
rect 188107 65108 188173 65109
rect 188107 65044 188108 65108
rect 188172 65044 188173 65108
rect 188107 65043 188173 65044
rect 187739 61980 187805 61981
rect 187739 61916 187740 61980
rect 187804 61916 187805 61980
rect 187739 61915 187805 61916
rect 187003 44028 187069 44029
rect 187003 43964 187004 44028
rect 187068 43964 187069 44028
rect 187003 43963 187069 43964
rect 186294 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 186914 43954
rect 186294 43634 186914 43718
rect 186294 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 186914 43634
rect 187006 43621 187066 43963
rect 187003 43620 187069 43621
rect 187003 43556 187004 43620
rect 187068 43556 187069 43620
rect 187003 43555 187069 43556
rect 186294 7954 186914 43398
rect 189582 31789 189642 141203
rect 190502 79117 190562 143515
rect 190794 142000 191414 155898
rect 191603 148476 191669 148477
rect 191603 148412 191604 148476
rect 191668 148412 191669 148476
rect 191603 148411 191669 148412
rect 190867 140860 190933 140861
rect 190867 140796 190868 140860
rect 190932 140796 190933 140860
rect 190867 140795 190933 140796
rect 190870 80613 190930 140795
rect 191051 114476 191117 114477
rect 191051 114412 191052 114476
rect 191116 114412 191117 114476
rect 191051 114411 191117 114412
rect 190867 80612 190933 80613
rect 190867 80548 190868 80612
rect 190932 80548 190933 80612
rect 190867 80547 190933 80548
rect 191054 79389 191114 114411
rect 191051 79388 191117 79389
rect 191051 79324 191052 79388
rect 191116 79324 191117 79388
rect 191051 79323 191117 79324
rect 190499 79116 190565 79117
rect 190499 79052 190500 79116
rect 190564 79052 190565 79116
rect 190499 79051 190565 79052
rect 190794 48454 191414 78000
rect 191606 70277 191666 148411
rect 191790 144533 191850 262515
rect 191974 144669 192034 263059
rect 192155 147388 192221 147389
rect 192155 147324 192156 147388
rect 192220 147324 192221 147388
rect 192155 147323 192221 147324
rect 191971 144668 192037 144669
rect 191971 144604 191972 144668
rect 192036 144604 192037 144668
rect 191971 144603 192037 144604
rect 191787 144532 191853 144533
rect 191787 144468 191788 144532
rect 191852 144468 191853 144532
rect 191787 144467 191853 144468
rect 192158 76805 192218 147323
rect 192339 141268 192405 141269
rect 192339 141204 192340 141268
rect 192404 141204 192405 141268
rect 192339 141203 192405 141204
rect 192155 76804 192221 76805
rect 192155 76740 192156 76804
rect 192220 76740 192221 76804
rect 192155 76739 192221 76740
rect 191603 70276 191669 70277
rect 191603 70212 191604 70276
rect 191668 70212 191669 70276
rect 191603 70211 191669 70212
rect 190794 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 191414 48454
rect 190794 48134 191414 48218
rect 190794 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 191414 48134
rect 189579 31788 189645 31789
rect 189579 31724 189580 31788
rect 189644 31724 189645 31788
rect 189579 31723 189645 31724
rect 186294 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 186914 7954
rect 186294 7634 186914 7718
rect 186294 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 186914 7634
rect 186294 -1306 186914 7398
rect 186294 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 186914 -1306
rect 186294 -1626 186914 -1542
rect 186294 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 186914 -1626
rect 186294 -7654 186914 -1862
rect 190794 12454 191414 47898
rect 192342 45661 192402 141203
rect 193262 140725 193322 265235
rect 194547 265164 194613 265165
rect 194547 265100 194548 265164
rect 194612 265100 194613 265164
rect 194547 265099 194613 265100
rect 193443 262716 193509 262717
rect 193443 262652 193444 262716
rect 193508 262652 193509 262716
rect 193443 262651 193509 262652
rect 193446 141541 193506 262651
rect 193627 147660 193693 147661
rect 193627 147596 193628 147660
rect 193692 147596 193693 147660
rect 193627 147595 193693 147596
rect 193443 141540 193509 141541
rect 193443 141476 193444 141540
rect 193508 141476 193509 141540
rect 193443 141475 193509 141476
rect 193259 140724 193325 140725
rect 193259 140660 193260 140724
rect 193324 140660 193325 140724
rect 193259 140659 193325 140660
rect 193443 140724 193509 140725
rect 193443 140660 193444 140724
rect 193508 140660 193509 140724
rect 193443 140659 193509 140660
rect 193259 140588 193325 140589
rect 193259 140524 193260 140588
rect 193324 140524 193325 140588
rect 193259 140523 193325 140524
rect 193262 76397 193322 140523
rect 193446 76941 193506 140659
rect 193630 78573 193690 147595
rect 194550 144397 194610 265099
rect 194731 265028 194797 265029
rect 194731 264964 194732 265028
rect 194796 264964 194797 265028
rect 194731 264963 194797 264964
rect 194734 145893 194794 264963
rect 195294 232954 195914 268398
rect 195294 232718 195326 232954
rect 195562 232718 195646 232954
rect 195882 232718 195914 232954
rect 195294 232634 195914 232718
rect 195294 232398 195326 232634
rect 195562 232398 195646 232634
rect 195882 232398 195914 232634
rect 195294 196954 195914 232398
rect 199794 708678 200414 711590
rect 199794 708442 199826 708678
rect 200062 708442 200146 708678
rect 200382 708442 200414 708678
rect 199794 708358 200414 708442
rect 199794 708122 199826 708358
rect 200062 708122 200146 708358
rect 200382 708122 200414 708358
rect 199794 669454 200414 708122
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 525454 200414 560898
rect 199794 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 200414 525454
rect 199794 525134 200414 525218
rect 199794 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 200414 525134
rect 199794 489454 200414 524898
rect 199794 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 200414 489454
rect 199794 489134 200414 489218
rect 199794 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 200414 489134
rect 199794 453454 200414 488898
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 199794 417454 200414 452898
rect 199794 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 200414 417454
rect 199794 417134 200414 417218
rect 199794 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 200414 417134
rect 199794 381454 200414 416898
rect 199794 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 200414 381454
rect 199794 381134 200414 381218
rect 199794 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 200414 381134
rect 199794 345454 200414 380898
rect 199794 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 200414 345454
rect 199794 345134 200414 345218
rect 199794 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 200414 345134
rect 199794 309454 200414 344898
rect 199794 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 200414 309454
rect 199794 309134 200414 309218
rect 199794 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 200414 309134
rect 199794 273454 200414 308898
rect 199794 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 200414 273454
rect 199794 273134 200414 273218
rect 199794 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 200414 273134
rect 199794 237454 200414 272898
rect 199794 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 200414 237454
rect 199794 237134 200414 237218
rect 199794 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 200414 237134
rect 199794 201454 200414 236898
rect 199794 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 200414 201454
rect 199794 201134 200414 201218
rect 199794 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 200414 201134
rect 196387 198252 196453 198253
rect 196387 198188 196388 198252
rect 196452 198188 196453 198252
rect 196387 198187 196453 198188
rect 195294 196718 195326 196954
rect 195562 196718 195646 196954
rect 195882 196718 195914 196954
rect 195294 196634 195914 196718
rect 195294 196398 195326 196634
rect 195562 196398 195646 196634
rect 195882 196398 195914 196634
rect 195294 160954 195914 196398
rect 196203 192812 196269 192813
rect 196203 192748 196204 192812
rect 196268 192748 196269 192812
rect 196203 192747 196269 192748
rect 196019 192540 196085 192541
rect 196019 192476 196020 192540
rect 196084 192476 196085 192540
rect 196019 192475 196085 192476
rect 195294 160718 195326 160954
rect 195562 160718 195646 160954
rect 195882 160718 195914 160954
rect 195294 160634 195914 160718
rect 195294 160398 195326 160634
rect 195562 160398 195646 160634
rect 195882 160398 195914 160634
rect 194731 145892 194797 145893
rect 194731 145828 194732 145892
rect 194796 145828 194797 145892
rect 194731 145827 194797 145828
rect 194547 144396 194613 144397
rect 194547 144332 194548 144396
rect 194612 144332 194613 144396
rect 194547 144331 194613 144332
rect 195099 139500 195165 139501
rect 195099 139436 195100 139500
rect 195164 139436 195165 139500
rect 195099 139435 195165 139436
rect 193627 78572 193693 78573
rect 193627 78508 193628 78572
rect 193692 78508 193693 78572
rect 193627 78507 193693 78508
rect 193443 76940 193509 76941
rect 193443 76876 193444 76940
rect 193508 76876 193509 76940
rect 193443 76875 193509 76876
rect 193259 76396 193325 76397
rect 193259 76332 193260 76396
rect 193324 76332 193325 76396
rect 193259 76331 193325 76332
rect 195102 70413 195162 139435
rect 195294 124954 195914 160398
rect 195294 124718 195326 124954
rect 195562 124718 195646 124954
rect 195882 124718 195914 124954
rect 195294 124634 195914 124718
rect 195294 124398 195326 124634
rect 195562 124398 195646 124634
rect 195882 124398 195914 124634
rect 195294 88954 195914 124398
rect 195294 88718 195326 88954
rect 195562 88718 195646 88954
rect 195882 88718 195914 88954
rect 195294 88634 195914 88718
rect 195294 88398 195326 88634
rect 195562 88398 195646 88634
rect 195882 88398 195914 88634
rect 195099 70412 195165 70413
rect 195099 70348 195100 70412
rect 195164 70348 195165 70412
rect 195099 70347 195165 70348
rect 195294 52954 195914 88398
rect 195294 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 195914 52954
rect 195294 52634 195914 52718
rect 195294 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 195914 52634
rect 192339 45660 192405 45661
rect 192339 45596 192340 45660
rect 192404 45596 192405 45660
rect 192339 45595 192405 45596
rect 190794 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 191414 12454
rect 190794 12134 191414 12218
rect 190794 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 191414 12134
rect 190794 -2266 191414 11898
rect 190794 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 191414 -2266
rect 190794 -2586 191414 -2502
rect 190794 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 191414 -2586
rect 190794 -7654 191414 -2822
rect 195294 16954 195914 52398
rect 196022 48245 196082 192475
rect 196206 54501 196266 192747
rect 196390 75445 196450 198187
rect 198779 198116 198845 198117
rect 198779 198052 198780 198116
rect 198844 198052 198845 198116
rect 198779 198051 198845 198052
rect 197859 185604 197925 185605
rect 197859 185540 197860 185604
rect 197924 185540 197925 185604
rect 197859 185539 197925 185540
rect 197675 185332 197741 185333
rect 197675 185268 197676 185332
rect 197740 185268 197741 185332
rect 197675 185267 197741 185268
rect 197307 185196 197373 185197
rect 197307 185132 197308 185196
rect 197372 185132 197373 185196
rect 197307 185131 197373 185132
rect 196571 147796 196637 147797
rect 196571 147732 196572 147796
rect 196636 147732 196637 147796
rect 196571 147731 196637 147732
rect 196387 75444 196453 75445
rect 196387 75380 196388 75444
rect 196452 75380 196453 75444
rect 196387 75379 196453 75380
rect 196574 62933 196634 147731
rect 197310 64565 197370 185131
rect 197491 174588 197557 174589
rect 197491 174524 197492 174588
rect 197556 174524 197557 174588
rect 197491 174523 197557 174524
rect 197494 65109 197554 174523
rect 197678 80069 197738 185267
rect 197675 80068 197741 80069
rect 197675 80004 197676 80068
rect 197740 80004 197741 80068
rect 197675 80003 197741 80004
rect 197862 79933 197922 185539
rect 197859 79932 197925 79933
rect 197859 79868 197860 79932
rect 197924 79868 197925 79932
rect 197859 79867 197925 79868
rect 197491 65108 197557 65109
rect 197491 65044 197492 65108
rect 197556 65044 197557 65108
rect 197491 65043 197557 65044
rect 197307 64564 197373 64565
rect 197307 64500 197308 64564
rect 197372 64500 197373 64564
rect 197307 64499 197373 64500
rect 196571 62932 196637 62933
rect 196571 62868 196572 62932
rect 196636 62868 196637 62932
rect 196571 62867 196637 62868
rect 196203 54500 196269 54501
rect 196203 54436 196204 54500
rect 196268 54436 196269 54500
rect 196203 54435 196269 54436
rect 198782 49469 198842 198051
rect 199794 165454 200414 200898
rect 204294 709638 204914 711590
rect 204294 709402 204326 709638
rect 204562 709402 204646 709638
rect 204882 709402 204914 709638
rect 204294 709318 204914 709402
rect 204294 709082 204326 709318
rect 204562 709082 204646 709318
rect 204882 709082 204914 709318
rect 204294 673954 204914 709082
rect 204294 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 204914 673954
rect 204294 673634 204914 673718
rect 204294 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 204914 673634
rect 204294 637954 204914 673398
rect 204294 637718 204326 637954
rect 204562 637718 204646 637954
rect 204882 637718 204914 637954
rect 204294 637634 204914 637718
rect 204294 637398 204326 637634
rect 204562 637398 204646 637634
rect 204882 637398 204914 637634
rect 204294 601954 204914 637398
rect 204294 601718 204326 601954
rect 204562 601718 204646 601954
rect 204882 601718 204914 601954
rect 204294 601634 204914 601718
rect 204294 601398 204326 601634
rect 204562 601398 204646 601634
rect 204882 601398 204914 601634
rect 204294 565954 204914 601398
rect 204294 565718 204326 565954
rect 204562 565718 204646 565954
rect 204882 565718 204914 565954
rect 204294 565634 204914 565718
rect 204294 565398 204326 565634
rect 204562 565398 204646 565634
rect 204882 565398 204914 565634
rect 204294 529954 204914 565398
rect 204294 529718 204326 529954
rect 204562 529718 204646 529954
rect 204882 529718 204914 529954
rect 204294 529634 204914 529718
rect 204294 529398 204326 529634
rect 204562 529398 204646 529634
rect 204882 529398 204914 529634
rect 204294 493954 204914 529398
rect 204294 493718 204326 493954
rect 204562 493718 204646 493954
rect 204882 493718 204914 493954
rect 204294 493634 204914 493718
rect 204294 493398 204326 493634
rect 204562 493398 204646 493634
rect 204882 493398 204914 493634
rect 204294 457954 204914 493398
rect 204294 457718 204326 457954
rect 204562 457718 204646 457954
rect 204882 457718 204914 457954
rect 204294 457634 204914 457718
rect 204294 457398 204326 457634
rect 204562 457398 204646 457634
rect 204882 457398 204914 457634
rect 204294 421954 204914 457398
rect 204294 421718 204326 421954
rect 204562 421718 204646 421954
rect 204882 421718 204914 421954
rect 204294 421634 204914 421718
rect 204294 421398 204326 421634
rect 204562 421398 204646 421634
rect 204882 421398 204914 421634
rect 204294 385954 204914 421398
rect 204294 385718 204326 385954
rect 204562 385718 204646 385954
rect 204882 385718 204914 385954
rect 204294 385634 204914 385718
rect 204294 385398 204326 385634
rect 204562 385398 204646 385634
rect 204882 385398 204914 385634
rect 204294 349954 204914 385398
rect 204294 349718 204326 349954
rect 204562 349718 204646 349954
rect 204882 349718 204914 349954
rect 204294 349634 204914 349718
rect 204294 349398 204326 349634
rect 204562 349398 204646 349634
rect 204882 349398 204914 349634
rect 204294 313954 204914 349398
rect 204294 313718 204326 313954
rect 204562 313718 204646 313954
rect 204882 313718 204914 313954
rect 204294 313634 204914 313718
rect 204294 313398 204326 313634
rect 204562 313398 204646 313634
rect 204882 313398 204914 313634
rect 204294 277954 204914 313398
rect 204294 277718 204326 277954
rect 204562 277718 204646 277954
rect 204882 277718 204914 277954
rect 204294 277634 204914 277718
rect 204294 277398 204326 277634
rect 204562 277398 204646 277634
rect 204882 277398 204914 277634
rect 204294 241954 204914 277398
rect 204294 241718 204326 241954
rect 204562 241718 204646 241954
rect 204882 241718 204914 241954
rect 204294 241634 204914 241718
rect 204294 241398 204326 241634
rect 204562 241398 204646 241634
rect 204882 241398 204914 241634
rect 204294 205954 204914 241398
rect 204294 205718 204326 205954
rect 204562 205718 204646 205954
rect 204882 205718 204914 205954
rect 204294 205634 204914 205718
rect 204294 205398 204326 205634
rect 204562 205398 204646 205634
rect 204882 205398 204914 205634
rect 200987 199884 201053 199885
rect 200987 199820 200988 199884
rect 201052 199820 201053 199884
rect 200987 199819 201053 199820
rect 200619 185740 200685 185741
rect 200619 185676 200620 185740
rect 200684 185676 200685 185740
rect 200619 185675 200685 185676
rect 199794 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 200414 165454
rect 199794 165134 200414 165218
rect 199794 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 200414 165134
rect 199331 147796 199397 147797
rect 199331 147732 199332 147796
rect 199396 147732 199397 147796
rect 199331 147731 199397 147732
rect 198963 147252 199029 147253
rect 198963 147188 198964 147252
rect 199028 147188 199029 147252
rect 198963 147187 199029 147188
rect 198966 74221 199026 147187
rect 198963 74220 199029 74221
rect 198963 74156 198964 74220
rect 199028 74156 199029 74220
rect 198963 74155 199029 74156
rect 199334 64890 199394 147731
rect 198966 64830 199394 64890
rect 199794 129454 200414 164898
rect 199794 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 200414 129454
rect 199794 129134 200414 129218
rect 199794 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 200414 129134
rect 199794 93454 200414 128898
rect 199794 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 200414 93454
rect 199794 93134 200414 93218
rect 199794 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 200414 93134
rect 198966 60349 199026 64830
rect 198963 60348 199029 60349
rect 198963 60284 198964 60348
rect 199028 60284 199029 60348
rect 198963 60283 199029 60284
rect 198966 59941 199026 60283
rect 198963 59940 199029 59941
rect 198963 59876 198964 59940
rect 199028 59876 199029 59940
rect 198963 59875 199029 59876
rect 199794 57454 200414 92898
rect 200622 66877 200682 185675
rect 200803 185468 200869 185469
rect 200803 185404 200804 185468
rect 200868 185404 200869 185468
rect 200803 185403 200869 185404
rect 200806 69597 200866 185403
rect 200803 69596 200869 69597
rect 200803 69532 200804 69596
rect 200868 69532 200869 69596
rect 200803 69531 200869 69532
rect 200990 68917 201050 199819
rect 201723 198796 201789 198797
rect 201723 198732 201724 198796
rect 201788 198732 201789 198796
rect 201723 198731 201789 198732
rect 201539 173500 201605 173501
rect 201539 173436 201540 173500
rect 201604 173436 201605 173500
rect 201539 173435 201605 173436
rect 200987 68916 201053 68917
rect 200987 68852 200988 68916
rect 201052 68852 201053 68916
rect 200987 68851 201053 68852
rect 200619 66876 200685 66877
rect 200619 66812 200620 66876
rect 200684 66812 200685 66876
rect 200619 66811 200685 66812
rect 201542 57629 201602 173435
rect 201726 64701 201786 198731
rect 203011 193900 203077 193901
rect 203011 193836 203012 193900
rect 203076 193836 203077 193900
rect 203011 193835 203077 193836
rect 201907 186556 201973 186557
rect 201907 186492 201908 186556
rect 201972 186492 201973 186556
rect 201907 186491 201973 186492
rect 201723 64700 201789 64701
rect 201723 64636 201724 64700
rect 201788 64636 201789 64700
rect 201723 64635 201789 64636
rect 201726 64157 201786 64635
rect 201723 64156 201789 64157
rect 201723 64092 201724 64156
rect 201788 64092 201789 64156
rect 201723 64091 201789 64092
rect 201910 62797 201970 186491
rect 203014 151830 203074 193835
rect 202830 151770 203074 151830
rect 204294 169954 204914 205398
rect 204294 169718 204326 169954
rect 204562 169718 204646 169954
rect 204882 169718 204914 169954
rect 204294 169634 204914 169718
rect 204294 169398 204326 169634
rect 204562 169398 204646 169634
rect 204882 169398 204914 169634
rect 202830 74550 202890 151770
rect 203011 150108 203077 150109
rect 203011 150044 203012 150108
rect 203076 150044 203077 150108
rect 203011 150043 203077 150044
rect 203014 75581 203074 150043
rect 203195 149972 203261 149973
rect 203195 149908 203196 149972
rect 203260 149908 203261 149972
rect 203195 149907 203261 149908
rect 203198 78981 203258 149907
rect 204294 133954 204914 169398
rect 204294 133718 204326 133954
rect 204562 133718 204646 133954
rect 204882 133718 204914 133954
rect 204294 133634 204914 133718
rect 204294 133398 204326 133634
rect 204562 133398 204646 133634
rect 204882 133398 204914 133634
rect 204294 97954 204914 133398
rect 204294 97718 204326 97954
rect 204562 97718 204646 97954
rect 204882 97718 204914 97954
rect 204294 97634 204914 97718
rect 204294 97398 204326 97634
rect 204562 97398 204646 97634
rect 204882 97398 204914 97634
rect 203195 78980 203261 78981
rect 203195 78916 203196 78980
rect 203260 78916 203261 78980
rect 203195 78915 203261 78916
rect 203011 75580 203077 75581
rect 203011 75516 203012 75580
rect 203076 75516 203077 75580
rect 203011 75515 203077 75516
rect 202830 74490 203074 74550
rect 201907 62796 201973 62797
rect 201907 62732 201908 62796
rect 201972 62732 201973 62796
rect 201907 62731 201973 62732
rect 201539 57628 201605 57629
rect 201539 57564 201540 57628
rect 201604 57564 201605 57628
rect 201539 57563 201605 57564
rect 202827 57628 202893 57629
rect 202827 57564 202828 57628
rect 202892 57564 202893 57628
rect 202827 57563 202893 57564
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 202830 57221 202890 57563
rect 199794 57134 200414 57218
rect 202827 57220 202893 57221
rect 202827 57156 202828 57220
rect 202892 57156 202893 57220
rect 202827 57155 202893 57156
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 198779 49468 198845 49469
rect 198779 49404 198780 49468
rect 198844 49404 198845 49468
rect 198779 49403 198845 49404
rect 198782 49061 198842 49403
rect 198779 49060 198845 49061
rect 198779 48996 198780 49060
rect 198844 48996 198845 49060
rect 198779 48995 198845 48996
rect 196019 48244 196085 48245
rect 196019 48180 196020 48244
rect 196084 48180 196085 48244
rect 196019 48179 196085 48180
rect 196022 47701 196082 48179
rect 196019 47700 196085 47701
rect 196019 47636 196020 47700
rect 196084 47636 196085 47700
rect 196019 47635 196085 47636
rect 195294 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 195914 16954
rect 195294 16634 195914 16718
rect 195294 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 195914 16634
rect 195294 -3226 195914 16398
rect 195294 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 195914 -3226
rect 195294 -3546 195914 -3462
rect 195294 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 195914 -3546
rect 195294 -7654 195914 -3782
rect 199794 21454 200414 56898
rect 203014 52325 203074 74490
rect 204294 61954 204914 97398
rect 204294 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 204914 61954
rect 204294 61634 204914 61718
rect 204294 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 204914 61634
rect 203011 52324 203077 52325
rect 203011 52260 203012 52324
rect 203076 52260 203077 52324
rect 203011 52259 203077 52260
rect 204115 52324 204181 52325
rect 204115 52260 204116 52324
rect 204180 52260 204181 52324
rect 204115 52259 204181 52260
rect 204118 51917 204178 52259
rect 204115 51916 204181 51917
rect 204115 51852 204116 51916
rect 204180 51852 204181 51916
rect 204115 51851 204181 51852
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -4186 200414 20898
rect 199794 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 200414 -4186
rect 199794 -4506 200414 -4422
rect 199794 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 200414 -4506
rect 199794 -7654 200414 -4742
rect 204294 25954 204914 61398
rect 204294 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 204914 25954
rect 204294 25634 204914 25718
rect 204294 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 204914 25634
rect 204294 -5146 204914 25398
rect 204294 -5382 204326 -5146
rect 204562 -5382 204646 -5146
rect 204882 -5382 204914 -5146
rect 204294 -5466 204914 -5382
rect 204294 -5702 204326 -5466
rect 204562 -5702 204646 -5466
rect 204882 -5702 204914 -5466
rect 204294 -7654 204914 -5702
rect 208794 710598 209414 711590
rect 208794 710362 208826 710598
rect 209062 710362 209146 710598
rect 209382 710362 209414 710598
rect 208794 710278 209414 710362
rect 208794 710042 208826 710278
rect 209062 710042 209146 710278
rect 209382 710042 209414 710278
rect 208794 678454 209414 710042
rect 208794 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 209414 678454
rect 208794 678134 209414 678218
rect 208794 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 209414 678134
rect 208794 642454 209414 677898
rect 208794 642218 208826 642454
rect 209062 642218 209146 642454
rect 209382 642218 209414 642454
rect 208794 642134 209414 642218
rect 208794 641898 208826 642134
rect 209062 641898 209146 642134
rect 209382 641898 209414 642134
rect 208794 606454 209414 641898
rect 208794 606218 208826 606454
rect 209062 606218 209146 606454
rect 209382 606218 209414 606454
rect 208794 606134 209414 606218
rect 208794 605898 208826 606134
rect 209062 605898 209146 606134
rect 209382 605898 209414 606134
rect 208794 570454 209414 605898
rect 208794 570218 208826 570454
rect 209062 570218 209146 570454
rect 209382 570218 209414 570454
rect 208794 570134 209414 570218
rect 208794 569898 208826 570134
rect 209062 569898 209146 570134
rect 209382 569898 209414 570134
rect 208794 534454 209414 569898
rect 208794 534218 208826 534454
rect 209062 534218 209146 534454
rect 209382 534218 209414 534454
rect 208794 534134 209414 534218
rect 208794 533898 208826 534134
rect 209062 533898 209146 534134
rect 209382 533898 209414 534134
rect 208794 498454 209414 533898
rect 208794 498218 208826 498454
rect 209062 498218 209146 498454
rect 209382 498218 209414 498454
rect 208794 498134 209414 498218
rect 208794 497898 208826 498134
rect 209062 497898 209146 498134
rect 209382 497898 209414 498134
rect 208794 462454 209414 497898
rect 208794 462218 208826 462454
rect 209062 462218 209146 462454
rect 209382 462218 209414 462454
rect 208794 462134 209414 462218
rect 208794 461898 208826 462134
rect 209062 461898 209146 462134
rect 209382 461898 209414 462134
rect 208794 426454 209414 461898
rect 208794 426218 208826 426454
rect 209062 426218 209146 426454
rect 209382 426218 209414 426454
rect 208794 426134 209414 426218
rect 208794 425898 208826 426134
rect 209062 425898 209146 426134
rect 209382 425898 209414 426134
rect 208794 390454 209414 425898
rect 208794 390218 208826 390454
rect 209062 390218 209146 390454
rect 209382 390218 209414 390454
rect 208794 390134 209414 390218
rect 208794 389898 208826 390134
rect 209062 389898 209146 390134
rect 209382 389898 209414 390134
rect 208794 354454 209414 389898
rect 208794 354218 208826 354454
rect 209062 354218 209146 354454
rect 209382 354218 209414 354454
rect 208794 354134 209414 354218
rect 208794 353898 208826 354134
rect 209062 353898 209146 354134
rect 209382 353898 209414 354134
rect 208794 318454 209414 353898
rect 208794 318218 208826 318454
rect 209062 318218 209146 318454
rect 209382 318218 209414 318454
rect 208794 318134 209414 318218
rect 208794 317898 208826 318134
rect 209062 317898 209146 318134
rect 209382 317898 209414 318134
rect 208794 282454 209414 317898
rect 208794 282218 208826 282454
rect 209062 282218 209146 282454
rect 209382 282218 209414 282454
rect 208794 282134 209414 282218
rect 208794 281898 208826 282134
rect 209062 281898 209146 282134
rect 209382 281898 209414 282134
rect 208794 246454 209414 281898
rect 208794 246218 208826 246454
rect 209062 246218 209146 246454
rect 209382 246218 209414 246454
rect 208794 246134 209414 246218
rect 208794 245898 208826 246134
rect 209062 245898 209146 246134
rect 209382 245898 209414 246134
rect 208794 210454 209414 245898
rect 208794 210218 208826 210454
rect 209062 210218 209146 210454
rect 209382 210218 209414 210454
rect 208794 210134 209414 210218
rect 208794 209898 208826 210134
rect 209062 209898 209146 210134
rect 209382 209898 209414 210134
rect 208794 174454 209414 209898
rect 208794 174218 208826 174454
rect 209062 174218 209146 174454
rect 209382 174218 209414 174454
rect 208794 174134 209414 174218
rect 208794 173898 208826 174134
rect 209062 173898 209146 174134
rect 209382 173898 209414 174134
rect 208794 138454 209414 173898
rect 208794 138218 208826 138454
rect 209062 138218 209146 138454
rect 209382 138218 209414 138454
rect 208794 138134 209414 138218
rect 208794 137898 208826 138134
rect 209062 137898 209146 138134
rect 209382 137898 209414 138134
rect 208794 102454 209414 137898
rect 208794 102218 208826 102454
rect 209062 102218 209146 102454
rect 209382 102218 209414 102454
rect 208794 102134 209414 102218
rect 208794 101898 208826 102134
rect 209062 101898 209146 102134
rect 209382 101898 209414 102134
rect 208794 66454 209414 101898
rect 208794 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 209414 66454
rect 208794 66134 209414 66218
rect 208794 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 209414 66134
rect 208794 30454 209414 65898
rect 208794 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 209414 30454
rect 208794 30134 209414 30218
rect 208794 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 209414 30134
rect 208794 -6106 209414 29898
rect 208794 -6342 208826 -6106
rect 209062 -6342 209146 -6106
rect 209382 -6342 209414 -6106
rect 208794 -6426 209414 -6342
rect 208794 -6662 208826 -6426
rect 209062 -6662 209146 -6426
rect 209382 -6662 209414 -6426
rect 208794 -7654 209414 -6662
rect 213294 711558 213914 711590
rect 213294 711322 213326 711558
rect 213562 711322 213646 711558
rect 213882 711322 213914 711558
rect 213294 711238 213914 711322
rect 213294 711002 213326 711238
rect 213562 711002 213646 711238
rect 213882 711002 213914 711238
rect 213294 682954 213914 711002
rect 213294 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 213914 682954
rect 213294 682634 213914 682718
rect 213294 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 213914 682634
rect 213294 646954 213914 682398
rect 213294 646718 213326 646954
rect 213562 646718 213646 646954
rect 213882 646718 213914 646954
rect 213294 646634 213914 646718
rect 213294 646398 213326 646634
rect 213562 646398 213646 646634
rect 213882 646398 213914 646634
rect 213294 610954 213914 646398
rect 213294 610718 213326 610954
rect 213562 610718 213646 610954
rect 213882 610718 213914 610954
rect 213294 610634 213914 610718
rect 213294 610398 213326 610634
rect 213562 610398 213646 610634
rect 213882 610398 213914 610634
rect 213294 574954 213914 610398
rect 213294 574718 213326 574954
rect 213562 574718 213646 574954
rect 213882 574718 213914 574954
rect 213294 574634 213914 574718
rect 213294 574398 213326 574634
rect 213562 574398 213646 574634
rect 213882 574398 213914 574634
rect 213294 538954 213914 574398
rect 213294 538718 213326 538954
rect 213562 538718 213646 538954
rect 213882 538718 213914 538954
rect 213294 538634 213914 538718
rect 213294 538398 213326 538634
rect 213562 538398 213646 538634
rect 213882 538398 213914 538634
rect 213294 502954 213914 538398
rect 213294 502718 213326 502954
rect 213562 502718 213646 502954
rect 213882 502718 213914 502954
rect 213294 502634 213914 502718
rect 213294 502398 213326 502634
rect 213562 502398 213646 502634
rect 213882 502398 213914 502634
rect 213294 466954 213914 502398
rect 213294 466718 213326 466954
rect 213562 466718 213646 466954
rect 213882 466718 213914 466954
rect 213294 466634 213914 466718
rect 213294 466398 213326 466634
rect 213562 466398 213646 466634
rect 213882 466398 213914 466634
rect 213294 430954 213914 466398
rect 213294 430718 213326 430954
rect 213562 430718 213646 430954
rect 213882 430718 213914 430954
rect 213294 430634 213914 430718
rect 213294 430398 213326 430634
rect 213562 430398 213646 430634
rect 213882 430398 213914 430634
rect 213294 394954 213914 430398
rect 213294 394718 213326 394954
rect 213562 394718 213646 394954
rect 213882 394718 213914 394954
rect 213294 394634 213914 394718
rect 213294 394398 213326 394634
rect 213562 394398 213646 394634
rect 213882 394398 213914 394634
rect 213294 358954 213914 394398
rect 213294 358718 213326 358954
rect 213562 358718 213646 358954
rect 213882 358718 213914 358954
rect 213294 358634 213914 358718
rect 213294 358398 213326 358634
rect 213562 358398 213646 358634
rect 213882 358398 213914 358634
rect 213294 322954 213914 358398
rect 213294 322718 213326 322954
rect 213562 322718 213646 322954
rect 213882 322718 213914 322954
rect 213294 322634 213914 322718
rect 213294 322398 213326 322634
rect 213562 322398 213646 322634
rect 213882 322398 213914 322634
rect 213294 286954 213914 322398
rect 213294 286718 213326 286954
rect 213562 286718 213646 286954
rect 213882 286718 213914 286954
rect 213294 286634 213914 286718
rect 213294 286398 213326 286634
rect 213562 286398 213646 286634
rect 213882 286398 213914 286634
rect 213294 250954 213914 286398
rect 213294 250718 213326 250954
rect 213562 250718 213646 250954
rect 213882 250718 213914 250954
rect 213294 250634 213914 250718
rect 213294 250398 213326 250634
rect 213562 250398 213646 250634
rect 213882 250398 213914 250634
rect 213294 214954 213914 250398
rect 213294 214718 213326 214954
rect 213562 214718 213646 214954
rect 213882 214718 213914 214954
rect 213294 214634 213914 214718
rect 213294 214398 213326 214634
rect 213562 214398 213646 214634
rect 213882 214398 213914 214634
rect 213294 178954 213914 214398
rect 213294 178718 213326 178954
rect 213562 178718 213646 178954
rect 213882 178718 213914 178954
rect 213294 178634 213914 178718
rect 213294 178398 213326 178634
rect 213562 178398 213646 178634
rect 213882 178398 213914 178634
rect 213294 142954 213914 178398
rect 213294 142718 213326 142954
rect 213562 142718 213646 142954
rect 213882 142718 213914 142954
rect 213294 142634 213914 142718
rect 213294 142398 213326 142634
rect 213562 142398 213646 142634
rect 213882 142398 213914 142634
rect 213294 106954 213914 142398
rect 213294 106718 213326 106954
rect 213562 106718 213646 106954
rect 213882 106718 213914 106954
rect 213294 106634 213914 106718
rect 213294 106398 213326 106634
rect 213562 106398 213646 106634
rect 213882 106398 213914 106634
rect 213294 70954 213914 106398
rect 213294 70718 213326 70954
rect 213562 70718 213646 70954
rect 213882 70718 213914 70954
rect 213294 70634 213914 70718
rect 213294 70398 213326 70634
rect 213562 70398 213646 70634
rect 213882 70398 213914 70634
rect 213294 34954 213914 70398
rect 213294 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 213914 34954
rect 213294 34634 213914 34718
rect 213294 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 213914 34634
rect 213294 -7066 213914 34398
rect 213294 -7302 213326 -7066
rect 213562 -7302 213646 -7066
rect 213882 -7302 213914 -7066
rect 213294 -7386 213914 -7302
rect 213294 -7622 213326 -7386
rect 213562 -7622 213646 -7386
rect 213882 -7622 213914 -7386
rect 213294 -7654 213914 -7622
rect 217794 704838 218414 711590
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 543454 218414 578898
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 507454 218414 542898
rect 217794 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 218414 507454
rect 217794 507134 218414 507218
rect 217794 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 218414 507134
rect 217794 471454 218414 506898
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 435454 218414 470898
rect 217794 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 218414 435454
rect 217794 435134 218414 435218
rect 217794 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 218414 435134
rect 217794 399454 218414 434898
rect 217794 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 218414 399454
rect 217794 399134 218414 399218
rect 217794 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 218414 399134
rect 217794 363454 218414 398898
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 327454 218414 362898
rect 217794 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 218414 327454
rect 217794 327134 218414 327218
rect 217794 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 218414 327134
rect 217794 291454 218414 326898
rect 217794 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 218414 291454
rect 217794 291134 218414 291218
rect 217794 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 218414 291134
rect 217794 255454 218414 290898
rect 217794 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 218414 255454
rect 217794 255134 218414 255218
rect 217794 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 218414 255134
rect 217794 219454 218414 254898
rect 217794 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 218414 219454
rect 217794 219134 218414 219218
rect 217794 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 218414 219134
rect 217794 183454 218414 218898
rect 217794 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 218414 183454
rect 217794 183134 218414 183218
rect 217794 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 218414 183134
rect 217794 147454 218414 182898
rect 217794 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 218414 147454
rect 217794 147134 218414 147218
rect 217794 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 218414 147134
rect 217794 111454 218414 146898
rect 217794 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 218414 111454
rect 217794 111134 218414 111218
rect 217794 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 218414 111134
rect 217794 75454 218414 110898
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -7654 218414 -902
rect 222294 705798 222914 711590
rect 222294 705562 222326 705798
rect 222562 705562 222646 705798
rect 222882 705562 222914 705798
rect 222294 705478 222914 705562
rect 222294 705242 222326 705478
rect 222562 705242 222646 705478
rect 222882 705242 222914 705478
rect 222294 691954 222914 705242
rect 222294 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 222914 691954
rect 222294 691634 222914 691718
rect 222294 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 222914 691634
rect 222294 655954 222914 691398
rect 222294 655718 222326 655954
rect 222562 655718 222646 655954
rect 222882 655718 222914 655954
rect 222294 655634 222914 655718
rect 222294 655398 222326 655634
rect 222562 655398 222646 655634
rect 222882 655398 222914 655634
rect 222294 619954 222914 655398
rect 222294 619718 222326 619954
rect 222562 619718 222646 619954
rect 222882 619718 222914 619954
rect 222294 619634 222914 619718
rect 222294 619398 222326 619634
rect 222562 619398 222646 619634
rect 222882 619398 222914 619634
rect 222294 583954 222914 619398
rect 222294 583718 222326 583954
rect 222562 583718 222646 583954
rect 222882 583718 222914 583954
rect 222294 583634 222914 583718
rect 222294 583398 222326 583634
rect 222562 583398 222646 583634
rect 222882 583398 222914 583634
rect 222294 547954 222914 583398
rect 222294 547718 222326 547954
rect 222562 547718 222646 547954
rect 222882 547718 222914 547954
rect 222294 547634 222914 547718
rect 222294 547398 222326 547634
rect 222562 547398 222646 547634
rect 222882 547398 222914 547634
rect 222294 511954 222914 547398
rect 222294 511718 222326 511954
rect 222562 511718 222646 511954
rect 222882 511718 222914 511954
rect 222294 511634 222914 511718
rect 222294 511398 222326 511634
rect 222562 511398 222646 511634
rect 222882 511398 222914 511634
rect 222294 475954 222914 511398
rect 222294 475718 222326 475954
rect 222562 475718 222646 475954
rect 222882 475718 222914 475954
rect 222294 475634 222914 475718
rect 222294 475398 222326 475634
rect 222562 475398 222646 475634
rect 222882 475398 222914 475634
rect 222294 439954 222914 475398
rect 222294 439718 222326 439954
rect 222562 439718 222646 439954
rect 222882 439718 222914 439954
rect 222294 439634 222914 439718
rect 222294 439398 222326 439634
rect 222562 439398 222646 439634
rect 222882 439398 222914 439634
rect 222294 403954 222914 439398
rect 222294 403718 222326 403954
rect 222562 403718 222646 403954
rect 222882 403718 222914 403954
rect 222294 403634 222914 403718
rect 222294 403398 222326 403634
rect 222562 403398 222646 403634
rect 222882 403398 222914 403634
rect 222294 367954 222914 403398
rect 222294 367718 222326 367954
rect 222562 367718 222646 367954
rect 222882 367718 222914 367954
rect 222294 367634 222914 367718
rect 222294 367398 222326 367634
rect 222562 367398 222646 367634
rect 222882 367398 222914 367634
rect 222294 331954 222914 367398
rect 222294 331718 222326 331954
rect 222562 331718 222646 331954
rect 222882 331718 222914 331954
rect 222294 331634 222914 331718
rect 222294 331398 222326 331634
rect 222562 331398 222646 331634
rect 222882 331398 222914 331634
rect 222294 295954 222914 331398
rect 222294 295718 222326 295954
rect 222562 295718 222646 295954
rect 222882 295718 222914 295954
rect 222294 295634 222914 295718
rect 222294 295398 222326 295634
rect 222562 295398 222646 295634
rect 222882 295398 222914 295634
rect 222294 259954 222914 295398
rect 222294 259718 222326 259954
rect 222562 259718 222646 259954
rect 222882 259718 222914 259954
rect 222294 259634 222914 259718
rect 222294 259398 222326 259634
rect 222562 259398 222646 259634
rect 222882 259398 222914 259634
rect 222294 223954 222914 259398
rect 222294 223718 222326 223954
rect 222562 223718 222646 223954
rect 222882 223718 222914 223954
rect 222294 223634 222914 223718
rect 222294 223398 222326 223634
rect 222562 223398 222646 223634
rect 222882 223398 222914 223634
rect 222294 187954 222914 223398
rect 222294 187718 222326 187954
rect 222562 187718 222646 187954
rect 222882 187718 222914 187954
rect 222294 187634 222914 187718
rect 222294 187398 222326 187634
rect 222562 187398 222646 187634
rect 222882 187398 222914 187634
rect 222294 151954 222914 187398
rect 222294 151718 222326 151954
rect 222562 151718 222646 151954
rect 222882 151718 222914 151954
rect 222294 151634 222914 151718
rect 222294 151398 222326 151634
rect 222562 151398 222646 151634
rect 222882 151398 222914 151634
rect 222294 115954 222914 151398
rect 222294 115718 222326 115954
rect 222562 115718 222646 115954
rect 222882 115718 222914 115954
rect 222294 115634 222914 115718
rect 222294 115398 222326 115634
rect 222562 115398 222646 115634
rect 222882 115398 222914 115634
rect 222294 79954 222914 115398
rect 222294 79718 222326 79954
rect 222562 79718 222646 79954
rect 222882 79718 222914 79954
rect 222294 79634 222914 79718
rect 222294 79398 222326 79634
rect 222562 79398 222646 79634
rect 222882 79398 222914 79634
rect 222294 43954 222914 79398
rect 222294 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 222914 43954
rect 222294 43634 222914 43718
rect 222294 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 222914 43634
rect 222294 7954 222914 43398
rect 222294 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 222914 7954
rect 222294 7634 222914 7718
rect 222294 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 222914 7634
rect 222294 -1306 222914 7398
rect 222294 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 222914 -1306
rect 222294 -1626 222914 -1542
rect 222294 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 222914 -1626
rect 222294 -7654 222914 -1862
rect 226794 706758 227414 711590
rect 226794 706522 226826 706758
rect 227062 706522 227146 706758
rect 227382 706522 227414 706758
rect 226794 706438 227414 706522
rect 226794 706202 226826 706438
rect 227062 706202 227146 706438
rect 227382 706202 227414 706438
rect 226794 696454 227414 706202
rect 226794 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 227414 696454
rect 226794 696134 227414 696218
rect 226794 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 227414 696134
rect 226794 660454 227414 695898
rect 226794 660218 226826 660454
rect 227062 660218 227146 660454
rect 227382 660218 227414 660454
rect 226794 660134 227414 660218
rect 226794 659898 226826 660134
rect 227062 659898 227146 660134
rect 227382 659898 227414 660134
rect 226794 624454 227414 659898
rect 226794 624218 226826 624454
rect 227062 624218 227146 624454
rect 227382 624218 227414 624454
rect 226794 624134 227414 624218
rect 226794 623898 226826 624134
rect 227062 623898 227146 624134
rect 227382 623898 227414 624134
rect 226794 588454 227414 623898
rect 226794 588218 226826 588454
rect 227062 588218 227146 588454
rect 227382 588218 227414 588454
rect 226794 588134 227414 588218
rect 226794 587898 226826 588134
rect 227062 587898 227146 588134
rect 227382 587898 227414 588134
rect 226794 552454 227414 587898
rect 226794 552218 226826 552454
rect 227062 552218 227146 552454
rect 227382 552218 227414 552454
rect 226794 552134 227414 552218
rect 226794 551898 226826 552134
rect 227062 551898 227146 552134
rect 227382 551898 227414 552134
rect 226794 516454 227414 551898
rect 226794 516218 226826 516454
rect 227062 516218 227146 516454
rect 227382 516218 227414 516454
rect 226794 516134 227414 516218
rect 226794 515898 226826 516134
rect 227062 515898 227146 516134
rect 227382 515898 227414 516134
rect 226794 480454 227414 515898
rect 226794 480218 226826 480454
rect 227062 480218 227146 480454
rect 227382 480218 227414 480454
rect 226794 480134 227414 480218
rect 226794 479898 226826 480134
rect 227062 479898 227146 480134
rect 227382 479898 227414 480134
rect 226794 444454 227414 479898
rect 226794 444218 226826 444454
rect 227062 444218 227146 444454
rect 227382 444218 227414 444454
rect 226794 444134 227414 444218
rect 226794 443898 226826 444134
rect 227062 443898 227146 444134
rect 227382 443898 227414 444134
rect 226794 408454 227414 443898
rect 226794 408218 226826 408454
rect 227062 408218 227146 408454
rect 227382 408218 227414 408454
rect 226794 408134 227414 408218
rect 226794 407898 226826 408134
rect 227062 407898 227146 408134
rect 227382 407898 227414 408134
rect 226794 372454 227414 407898
rect 226794 372218 226826 372454
rect 227062 372218 227146 372454
rect 227382 372218 227414 372454
rect 226794 372134 227414 372218
rect 226794 371898 226826 372134
rect 227062 371898 227146 372134
rect 227382 371898 227414 372134
rect 226794 336454 227414 371898
rect 226794 336218 226826 336454
rect 227062 336218 227146 336454
rect 227382 336218 227414 336454
rect 226794 336134 227414 336218
rect 226794 335898 226826 336134
rect 227062 335898 227146 336134
rect 227382 335898 227414 336134
rect 226794 300454 227414 335898
rect 226794 300218 226826 300454
rect 227062 300218 227146 300454
rect 227382 300218 227414 300454
rect 226794 300134 227414 300218
rect 226794 299898 226826 300134
rect 227062 299898 227146 300134
rect 227382 299898 227414 300134
rect 226794 264454 227414 299898
rect 226794 264218 226826 264454
rect 227062 264218 227146 264454
rect 227382 264218 227414 264454
rect 226794 264134 227414 264218
rect 226794 263898 226826 264134
rect 227062 263898 227146 264134
rect 227382 263898 227414 264134
rect 226794 228454 227414 263898
rect 226794 228218 226826 228454
rect 227062 228218 227146 228454
rect 227382 228218 227414 228454
rect 226794 228134 227414 228218
rect 226794 227898 226826 228134
rect 227062 227898 227146 228134
rect 227382 227898 227414 228134
rect 226794 192454 227414 227898
rect 226794 192218 226826 192454
rect 227062 192218 227146 192454
rect 227382 192218 227414 192454
rect 226794 192134 227414 192218
rect 226794 191898 226826 192134
rect 227062 191898 227146 192134
rect 227382 191898 227414 192134
rect 226794 156454 227414 191898
rect 226794 156218 226826 156454
rect 227062 156218 227146 156454
rect 227382 156218 227414 156454
rect 226794 156134 227414 156218
rect 226794 155898 226826 156134
rect 227062 155898 227146 156134
rect 227382 155898 227414 156134
rect 226794 120454 227414 155898
rect 226794 120218 226826 120454
rect 227062 120218 227146 120454
rect 227382 120218 227414 120454
rect 226794 120134 227414 120218
rect 226794 119898 226826 120134
rect 227062 119898 227146 120134
rect 227382 119898 227414 120134
rect 226794 84454 227414 119898
rect 226794 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 227414 84454
rect 226794 84134 227414 84218
rect 226794 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 227414 84134
rect 226794 48454 227414 83898
rect 226794 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 227414 48454
rect 226794 48134 227414 48218
rect 226794 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 227414 48134
rect 226794 12454 227414 47898
rect 226794 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 227414 12454
rect 226794 12134 227414 12218
rect 226794 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 227414 12134
rect 226794 -2266 227414 11898
rect 226794 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 227414 -2266
rect 226794 -2586 227414 -2502
rect 226794 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 227414 -2586
rect 226794 -7654 227414 -2822
rect 231294 707718 231914 711590
rect 231294 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 231914 707718
rect 231294 707398 231914 707482
rect 231294 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 231914 707398
rect 231294 700954 231914 707162
rect 231294 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 231914 700954
rect 231294 700634 231914 700718
rect 231294 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 231914 700634
rect 231294 664954 231914 700398
rect 231294 664718 231326 664954
rect 231562 664718 231646 664954
rect 231882 664718 231914 664954
rect 231294 664634 231914 664718
rect 231294 664398 231326 664634
rect 231562 664398 231646 664634
rect 231882 664398 231914 664634
rect 231294 628954 231914 664398
rect 231294 628718 231326 628954
rect 231562 628718 231646 628954
rect 231882 628718 231914 628954
rect 231294 628634 231914 628718
rect 231294 628398 231326 628634
rect 231562 628398 231646 628634
rect 231882 628398 231914 628634
rect 231294 592954 231914 628398
rect 231294 592718 231326 592954
rect 231562 592718 231646 592954
rect 231882 592718 231914 592954
rect 231294 592634 231914 592718
rect 231294 592398 231326 592634
rect 231562 592398 231646 592634
rect 231882 592398 231914 592634
rect 231294 556954 231914 592398
rect 231294 556718 231326 556954
rect 231562 556718 231646 556954
rect 231882 556718 231914 556954
rect 231294 556634 231914 556718
rect 231294 556398 231326 556634
rect 231562 556398 231646 556634
rect 231882 556398 231914 556634
rect 231294 520954 231914 556398
rect 231294 520718 231326 520954
rect 231562 520718 231646 520954
rect 231882 520718 231914 520954
rect 231294 520634 231914 520718
rect 231294 520398 231326 520634
rect 231562 520398 231646 520634
rect 231882 520398 231914 520634
rect 231294 484954 231914 520398
rect 231294 484718 231326 484954
rect 231562 484718 231646 484954
rect 231882 484718 231914 484954
rect 231294 484634 231914 484718
rect 231294 484398 231326 484634
rect 231562 484398 231646 484634
rect 231882 484398 231914 484634
rect 231294 448954 231914 484398
rect 231294 448718 231326 448954
rect 231562 448718 231646 448954
rect 231882 448718 231914 448954
rect 231294 448634 231914 448718
rect 231294 448398 231326 448634
rect 231562 448398 231646 448634
rect 231882 448398 231914 448634
rect 231294 412954 231914 448398
rect 231294 412718 231326 412954
rect 231562 412718 231646 412954
rect 231882 412718 231914 412954
rect 231294 412634 231914 412718
rect 231294 412398 231326 412634
rect 231562 412398 231646 412634
rect 231882 412398 231914 412634
rect 231294 376954 231914 412398
rect 231294 376718 231326 376954
rect 231562 376718 231646 376954
rect 231882 376718 231914 376954
rect 231294 376634 231914 376718
rect 231294 376398 231326 376634
rect 231562 376398 231646 376634
rect 231882 376398 231914 376634
rect 231294 340954 231914 376398
rect 231294 340718 231326 340954
rect 231562 340718 231646 340954
rect 231882 340718 231914 340954
rect 231294 340634 231914 340718
rect 231294 340398 231326 340634
rect 231562 340398 231646 340634
rect 231882 340398 231914 340634
rect 231294 304954 231914 340398
rect 231294 304718 231326 304954
rect 231562 304718 231646 304954
rect 231882 304718 231914 304954
rect 231294 304634 231914 304718
rect 231294 304398 231326 304634
rect 231562 304398 231646 304634
rect 231882 304398 231914 304634
rect 231294 268954 231914 304398
rect 231294 268718 231326 268954
rect 231562 268718 231646 268954
rect 231882 268718 231914 268954
rect 231294 268634 231914 268718
rect 231294 268398 231326 268634
rect 231562 268398 231646 268634
rect 231882 268398 231914 268634
rect 231294 232954 231914 268398
rect 231294 232718 231326 232954
rect 231562 232718 231646 232954
rect 231882 232718 231914 232954
rect 231294 232634 231914 232718
rect 231294 232398 231326 232634
rect 231562 232398 231646 232634
rect 231882 232398 231914 232634
rect 231294 196954 231914 232398
rect 231294 196718 231326 196954
rect 231562 196718 231646 196954
rect 231882 196718 231914 196954
rect 231294 196634 231914 196718
rect 231294 196398 231326 196634
rect 231562 196398 231646 196634
rect 231882 196398 231914 196634
rect 231294 160954 231914 196398
rect 231294 160718 231326 160954
rect 231562 160718 231646 160954
rect 231882 160718 231914 160954
rect 231294 160634 231914 160718
rect 231294 160398 231326 160634
rect 231562 160398 231646 160634
rect 231882 160398 231914 160634
rect 231294 124954 231914 160398
rect 231294 124718 231326 124954
rect 231562 124718 231646 124954
rect 231882 124718 231914 124954
rect 231294 124634 231914 124718
rect 231294 124398 231326 124634
rect 231562 124398 231646 124634
rect 231882 124398 231914 124634
rect 231294 88954 231914 124398
rect 231294 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 231914 88954
rect 231294 88634 231914 88718
rect 231294 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 231914 88634
rect 231294 52954 231914 88398
rect 231294 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 231914 52954
rect 231294 52634 231914 52718
rect 231294 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 231914 52634
rect 231294 16954 231914 52398
rect 231294 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 231914 16954
rect 231294 16634 231914 16718
rect 231294 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 231914 16634
rect 231294 -3226 231914 16398
rect 231294 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 231914 -3226
rect 231294 -3546 231914 -3462
rect 231294 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 231914 -3546
rect 231294 -7654 231914 -3782
rect 235794 708678 236414 711590
rect 235794 708442 235826 708678
rect 236062 708442 236146 708678
rect 236382 708442 236414 708678
rect 235794 708358 236414 708442
rect 235794 708122 235826 708358
rect 236062 708122 236146 708358
rect 236382 708122 236414 708358
rect 235794 669454 236414 708122
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 561454 236414 596898
rect 235794 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 236414 561454
rect 235794 561134 236414 561218
rect 235794 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 236414 561134
rect 235794 525454 236414 560898
rect 235794 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 236414 525454
rect 235794 525134 236414 525218
rect 235794 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 236414 525134
rect 235794 489454 236414 524898
rect 235794 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 236414 489454
rect 235794 489134 236414 489218
rect 235794 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 236414 489134
rect 235794 453454 236414 488898
rect 235794 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 236414 453454
rect 235794 453134 236414 453218
rect 235794 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 236414 453134
rect 235794 417454 236414 452898
rect 235794 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 236414 417454
rect 235794 417134 236414 417218
rect 235794 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 236414 417134
rect 235794 381454 236414 416898
rect 235794 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 236414 381454
rect 235794 381134 236414 381218
rect 235794 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 236414 381134
rect 235794 345454 236414 380898
rect 235794 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 236414 345454
rect 235794 345134 236414 345218
rect 235794 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 236414 345134
rect 235794 309454 236414 344898
rect 235794 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 236414 309454
rect 235794 309134 236414 309218
rect 235794 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 236414 309134
rect 235794 273454 236414 308898
rect 235794 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 236414 273454
rect 235794 273134 236414 273218
rect 235794 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 236414 273134
rect 235794 237454 236414 272898
rect 235794 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 236414 237454
rect 235794 237134 236414 237218
rect 235794 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 236414 237134
rect 235794 201454 236414 236898
rect 235794 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 236414 201454
rect 235794 201134 236414 201218
rect 235794 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 236414 201134
rect 235794 165454 236414 200898
rect 235794 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 236414 165454
rect 235794 165134 236414 165218
rect 235794 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 236414 165134
rect 235794 129454 236414 164898
rect 235794 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 236414 129454
rect 235794 129134 236414 129218
rect 235794 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 236414 129134
rect 235794 93454 236414 128898
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 235794 57454 236414 92898
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -4186 236414 20898
rect 235794 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 236414 -4186
rect 235794 -4506 236414 -4422
rect 235794 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 236414 -4506
rect 235794 -7654 236414 -4742
rect 240294 709638 240914 711590
rect 240294 709402 240326 709638
rect 240562 709402 240646 709638
rect 240882 709402 240914 709638
rect 240294 709318 240914 709402
rect 240294 709082 240326 709318
rect 240562 709082 240646 709318
rect 240882 709082 240914 709318
rect 240294 673954 240914 709082
rect 240294 673718 240326 673954
rect 240562 673718 240646 673954
rect 240882 673718 240914 673954
rect 240294 673634 240914 673718
rect 240294 673398 240326 673634
rect 240562 673398 240646 673634
rect 240882 673398 240914 673634
rect 240294 637954 240914 673398
rect 240294 637718 240326 637954
rect 240562 637718 240646 637954
rect 240882 637718 240914 637954
rect 240294 637634 240914 637718
rect 240294 637398 240326 637634
rect 240562 637398 240646 637634
rect 240882 637398 240914 637634
rect 240294 601954 240914 637398
rect 240294 601718 240326 601954
rect 240562 601718 240646 601954
rect 240882 601718 240914 601954
rect 240294 601634 240914 601718
rect 240294 601398 240326 601634
rect 240562 601398 240646 601634
rect 240882 601398 240914 601634
rect 240294 565954 240914 601398
rect 240294 565718 240326 565954
rect 240562 565718 240646 565954
rect 240882 565718 240914 565954
rect 240294 565634 240914 565718
rect 240294 565398 240326 565634
rect 240562 565398 240646 565634
rect 240882 565398 240914 565634
rect 240294 529954 240914 565398
rect 240294 529718 240326 529954
rect 240562 529718 240646 529954
rect 240882 529718 240914 529954
rect 240294 529634 240914 529718
rect 240294 529398 240326 529634
rect 240562 529398 240646 529634
rect 240882 529398 240914 529634
rect 240294 493954 240914 529398
rect 240294 493718 240326 493954
rect 240562 493718 240646 493954
rect 240882 493718 240914 493954
rect 240294 493634 240914 493718
rect 240294 493398 240326 493634
rect 240562 493398 240646 493634
rect 240882 493398 240914 493634
rect 240294 457954 240914 493398
rect 240294 457718 240326 457954
rect 240562 457718 240646 457954
rect 240882 457718 240914 457954
rect 240294 457634 240914 457718
rect 240294 457398 240326 457634
rect 240562 457398 240646 457634
rect 240882 457398 240914 457634
rect 240294 421954 240914 457398
rect 240294 421718 240326 421954
rect 240562 421718 240646 421954
rect 240882 421718 240914 421954
rect 240294 421634 240914 421718
rect 240294 421398 240326 421634
rect 240562 421398 240646 421634
rect 240882 421398 240914 421634
rect 240294 385954 240914 421398
rect 240294 385718 240326 385954
rect 240562 385718 240646 385954
rect 240882 385718 240914 385954
rect 240294 385634 240914 385718
rect 240294 385398 240326 385634
rect 240562 385398 240646 385634
rect 240882 385398 240914 385634
rect 240294 349954 240914 385398
rect 240294 349718 240326 349954
rect 240562 349718 240646 349954
rect 240882 349718 240914 349954
rect 240294 349634 240914 349718
rect 240294 349398 240326 349634
rect 240562 349398 240646 349634
rect 240882 349398 240914 349634
rect 240294 313954 240914 349398
rect 240294 313718 240326 313954
rect 240562 313718 240646 313954
rect 240882 313718 240914 313954
rect 240294 313634 240914 313718
rect 240294 313398 240326 313634
rect 240562 313398 240646 313634
rect 240882 313398 240914 313634
rect 240294 277954 240914 313398
rect 240294 277718 240326 277954
rect 240562 277718 240646 277954
rect 240882 277718 240914 277954
rect 240294 277634 240914 277718
rect 240294 277398 240326 277634
rect 240562 277398 240646 277634
rect 240882 277398 240914 277634
rect 240294 241954 240914 277398
rect 240294 241718 240326 241954
rect 240562 241718 240646 241954
rect 240882 241718 240914 241954
rect 240294 241634 240914 241718
rect 240294 241398 240326 241634
rect 240562 241398 240646 241634
rect 240882 241398 240914 241634
rect 240294 205954 240914 241398
rect 240294 205718 240326 205954
rect 240562 205718 240646 205954
rect 240882 205718 240914 205954
rect 240294 205634 240914 205718
rect 240294 205398 240326 205634
rect 240562 205398 240646 205634
rect 240882 205398 240914 205634
rect 240294 169954 240914 205398
rect 240294 169718 240326 169954
rect 240562 169718 240646 169954
rect 240882 169718 240914 169954
rect 240294 169634 240914 169718
rect 240294 169398 240326 169634
rect 240562 169398 240646 169634
rect 240882 169398 240914 169634
rect 240294 133954 240914 169398
rect 240294 133718 240326 133954
rect 240562 133718 240646 133954
rect 240882 133718 240914 133954
rect 240294 133634 240914 133718
rect 240294 133398 240326 133634
rect 240562 133398 240646 133634
rect 240882 133398 240914 133634
rect 240294 97954 240914 133398
rect 240294 97718 240326 97954
rect 240562 97718 240646 97954
rect 240882 97718 240914 97954
rect 240294 97634 240914 97718
rect 240294 97398 240326 97634
rect 240562 97398 240646 97634
rect 240882 97398 240914 97634
rect 240294 61954 240914 97398
rect 240294 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 240914 61954
rect 240294 61634 240914 61718
rect 240294 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 240914 61634
rect 240294 25954 240914 61398
rect 240294 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 240914 25954
rect 240294 25634 240914 25718
rect 240294 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 240914 25634
rect 240294 -5146 240914 25398
rect 240294 -5382 240326 -5146
rect 240562 -5382 240646 -5146
rect 240882 -5382 240914 -5146
rect 240294 -5466 240914 -5382
rect 240294 -5702 240326 -5466
rect 240562 -5702 240646 -5466
rect 240882 -5702 240914 -5466
rect 240294 -7654 240914 -5702
rect 244794 710598 245414 711590
rect 244794 710362 244826 710598
rect 245062 710362 245146 710598
rect 245382 710362 245414 710598
rect 244794 710278 245414 710362
rect 244794 710042 244826 710278
rect 245062 710042 245146 710278
rect 245382 710042 245414 710278
rect 244794 678454 245414 710042
rect 244794 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 245414 678454
rect 244794 678134 245414 678218
rect 244794 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 245414 678134
rect 244794 642454 245414 677898
rect 244794 642218 244826 642454
rect 245062 642218 245146 642454
rect 245382 642218 245414 642454
rect 244794 642134 245414 642218
rect 244794 641898 244826 642134
rect 245062 641898 245146 642134
rect 245382 641898 245414 642134
rect 244794 606454 245414 641898
rect 244794 606218 244826 606454
rect 245062 606218 245146 606454
rect 245382 606218 245414 606454
rect 244794 606134 245414 606218
rect 244794 605898 244826 606134
rect 245062 605898 245146 606134
rect 245382 605898 245414 606134
rect 244794 570454 245414 605898
rect 244794 570218 244826 570454
rect 245062 570218 245146 570454
rect 245382 570218 245414 570454
rect 244794 570134 245414 570218
rect 244794 569898 244826 570134
rect 245062 569898 245146 570134
rect 245382 569898 245414 570134
rect 244794 534454 245414 569898
rect 244794 534218 244826 534454
rect 245062 534218 245146 534454
rect 245382 534218 245414 534454
rect 244794 534134 245414 534218
rect 244794 533898 244826 534134
rect 245062 533898 245146 534134
rect 245382 533898 245414 534134
rect 244794 498454 245414 533898
rect 244794 498218 244826 498454
rect 245062 498218 245146 498454
rect 245382 498218 245414 498454
rect 244794 498134 245414 498218
rect 244794 497898 244826 498134
rect 245062 497898 245146 498134
rect 245382 497898 245414 498134
rect 244794 462454 245414 497898
rect 244794 462218 244826 462454
rect 245062 462218 245146 462454
rect 245382 462218 245414 462454
rect 244794 462134 245414 462218
rect 244794 461898 244826 462134
rect 245062 461898 245146 462134
rect 245382 461898 245414 462134
rect 244794 426454 245414 461898
rect 244794 426218 244826 426454
rect 245062 426218 245146 426454
rect 245382 426218 245414 426454
rect 244794 426134 245414 426218
rect 244794 425898 244826 426134
rect 245062 425898 245146 426134
rect 245382 425898 245414 426134
rect 244794 390454 245414 425898
rect 244794 390218 244826 390454
rect 245062 390218 245146 390454
rect 245382 390218 245414 390454
rect 244794 390134 245414 390218
rect 244794 389898 244826 390134
rect 245062 389898 245146 390134
rect 245382 389898 245414 390134
rect 244794 354454 245414 389898
rect 244794 354218 244826 354454
rect 245062 354218 245146 354454
rect 245382 354218 245414 354454
rect 244794 354134 245414 354218
rect 244794 353898 244826 354134
rect 245062 353898 245146 354134
rect 245382 353898 245414 354134
rect 244794 318454 245414 353898
rect 244794 318218 244826 318454
rect 245062 318218 245146 318454
rect 245382 318218 245414 318454
rect 244794 318134 245414 318218
rect 244794 317898 244826 318134
rect 245062 317898 245146 318134
rect 245382 317898 245414 318134
rect 244794 282454 245414 317898
rect 244794 282218 244826 282454
rect 245062 282218 245146 282454
rect 245382 282218 245414 282454
rect 244794 282134 245414 282218
rect 244794 281898 244826 282134
rect 245062 281898 245146 282134
rect 245382 281898 245414 282134
rect 244794 246454 245414 281898
rect 244794 246218 244826 246454
rect 245062 246218 245146 246454
rect 245382 246218 245414 246454
rect 244794 246134 245414 246218
rect 244794 245898 244826 246134
rect 245062 245898 245146 246134
rect 245382 245898 245414 246134
rect 244794 210454 245414 245898
rect 244794 210218 244826 210454
rect 245062 210218 245146 210454
rect 245382 210218 245414 210454
rect 244794 210134 245414 210218
rect 244794 209898 244826 210134
rect 245062 209898 245146 210134
rect 245382 209898 245414 210134
rect 244794 174454 245414 209898
rect 244794 174218 244826 174454
rect 245062 174218 245146 174454
rect 245382 174218 245414 174454
rect 244794 174134 245414 174218
rect 244794 173898 244826 174134
rect 245062 173898 245146 174134
rect 245382 173898 245414 174134
rect 244794 138454 245414 173898
rect 244794 138218 244826 138454
rect 245062 138218 245146 138454
rect 245382 138218 245414 138454
rect 244794 138134 245414 138218
rect 244794 137898 244826 138134
rect 245062 137898 245146 138134
rect 245382 137898 245414 138134
rect 244794 102454 245414 137898
rect 244794 102218 244826 102454
rect 245062 102218 245146 102454
rect 245382 102218 245414 102454
rect 244794 102134 245414 102218
rect 244794 101898 244826 102134
rect 245062 101898 245146 102134
rect 245382 101898 245414 102134
rect 244794 66454 245414 101898
rect 244794 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 245414 66454
rect 244794 66134 245414 66218
rect 244794 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 245414 66134
rect 244794 30454 245414 65898
rect 244794 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 245414 30454
rect 244794 30134 245414 30218
rect 244794 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 245414 30134
rect 244794 -6106 245414 29898
rect 244794 -6342 244826 -6106
rect 245062 -6342 245146 -6106
rect 245382 -6342 245414 -6106
rect 244794 -6426 245414 -6342
rect 244794 -6662 244826 -6426
rect 245062 -6662 245146 -6426
rect 245382 -6662 245414 -6426
rect 244794 -7654 245414 -6662
rect 249294 711558 249914 711590
rect 249294 711322 249326 711558
rect 249562 711322 249646 711558
rect 249882 711322 249914 711558
rect 249294 711238 249914 711322
rect 249294 711002 249326 711238
rect 249562 711002 249646 711238
rect 249882 711002 249914 711238
rect 249294 682954 249914 711002
rect 249294 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 249914 682954
rect 249294 682634 249914 682718
rect 249294 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 249914 682634
rect 249294 646954 249914 682398
rect 249294 646718 249326 646954
rect 249562 646718 249646 646954
rect 249882 646718 249914 646954
rect 249294 646634 249914 646718
rect 249294 646398 249326 646634
rect 249562 646398 249646 646634
rect 249882 646398 249914 646634
rect 249294 610954 249914 646398
rect 249294 610718 249326 610954
rect 249562 610718 249646 610954
rect 249882 610718 249914 610954
rect 249294 610634 249914 610718
rect 249294 610398 249326 610634
rect 249562 610398 249646 610634
rect 249882 610398 249914 610634
rect 249294 574954 249914 610398
rect 249294 574718 249326 574954
rect 249562 574718 249646 574954
rect 249882 574718 249914 574954
rect 249294 574634 249914 574718
rect 249294 574398 249326 574634
rect 249562 574398 249646 574634
rect 249882 574398 249914 574634
rect 249294 538954 249914 574398
rect 249294 538718 249326 538954
rect 249562 538718 249646 538954
rect 249882 538718 249914 538954
rect 249294 538634 249914 538718
rect 249294 538398 249326 538634
rect 249562 538398 249646 538634
rect 249882 538398 249914 538634
rect 249294 502954 249914 538398
rect 249294 502718 249326 502954
rect 249562 502718 249646 502954
rect 249882 502718 249914 502954
rect 249294 502634 249914 502718
rect 249294 502398 249326 502634
rect 249562 502398 249646 502634
rect 249882 502398 249914 502634
rect 249294 466954 249914 502398
rect 249294 466718 249326 466954
rect 249562 466718 249646 466954
rect 249882 466718 249914 466954
rect 249294 466634 249914 466718
rect 249294 466398 249326 466634
rect 249562 466398 249646 466634
rect 249882 466398 249914 466634
rect 249294 430954 249914 466398
rect 249294 430718 249326 430954
rect 249562 430718 249646 430954
rect 249882 430718 249914 430954
rect 249294 430634 249914 430718
rect 249294 430398 249326 430634
rect 249562 430398 249646 430634
rect 249882 430398 249914 430634
rect 249294 394954 249914 430398
rect 249294 394718 249326 394954
rect 249562 394718 249646 394954
rect 249882 394718 249914 394954
rect 249294 394634 249914 394718
rect 249294 394398 249326 394634
rect 249562 394398 249646 394634
rect 249882 394398 249914 394634
rect 249294 358954 249914 394398
rect 249294 358718 249326 358954
rect 249562 358718 249646 358954
rect 249882 358718 249914 358954
rect 249294 358634 249914 358718
rect 249294 358398 249326 358634
rect 249562 358398 249646 358634
rect 249882 358398 249914 358634
rect 249294 322954 249914 358398
rect 249294 322718 249326 322954
rect 249562 322718 249646 322954
rect 249882 322718 249914 322954
rect 249294 322634 249914 322718
rect 249294 322398 249326 322634
rect 249562 322398 249646 322634
rect 249882 322398 249914 322634
rect 249294 286954 249914 322398
rect 249294 286718 249326 286954
rect 249562 286718 249646 286954
rect 249882 286718 249914 286954
rect 249294 286634 249914 286718
rect 249294 286398 249326 286634
rect 249562 286398 249646 286634
rect 249882 286398 249914 286634
rect 249294 250954 249914 286398
rect 249294 250718 249326 250954
rect 249562 250718 249646 250954
rect 249882 250718 249914 250954
rect 249294 250634 249914 250718
rect 249294 250398 249326 250634
rect 249562 250398 249646 250634
rect 249882 250398 249914 250634
rect 249294 214954 249914 250398
rect 249294 214718 249326 214954
rect 249562 214718 249646 214954
rect 249882 214718 249914 214954
rect 249294 214634 249914 214718
rect 249294 214398 249326 214634
rect 249562 214398 249646 214634
rect 249882 214398 249914 214634
rect 249294 178954 249914 214398
rect 249294 178718 249326 178954
rect 249562 178718 249646 178954
rect 249882 178718 249914 178954
rect 249294 178634 249914 178718
rect 249294 178398 249326 178634
rect 249562 178398 249646 178634
rect 249882 178398 249914 178634
rect 249294 142954 249914 178398
rect 249294 142718 249326 142954
rect 249562 142718 249646 142954
rect 249882 142718 249914 142954
rect 249294 142634 249914 142718
rect 249294 142398 249326 142634
rect 249562 142398 249646 142634
rect 249882 142398 249914 142634
rect 249294 106954 249914 142398
rect 249294 106718 249326 106954
rect 249562 106718 249646 106954
rect 249882 106718 249914 106954
rect 249294 106634 249914 106718
rect 249294 106398 249326 106634
rect 249562 106398 249646 106634
rect 249882 106398 249914 106634
rect 249294 70954 249914 106398
rect 249294 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 249914 70954
rect 249294 70634 249914 70718
rect 249294 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 249914 70634
rect 249294 34954 249914 70398
rect 249294 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 249914 34954
rect 249294 34634 249914 34718
rect 249294 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 249914 34634
rect 249294 -7066 249914 34398
rect 249294 -7302 249326 -7066
rect 249562 -7302 249646 -7066
rect 249882 -7302 249914 -7066
rect 249294 -7386 249914 -7302
rect 249294 -7622 249326 -7386
rect 249562 -7622 249646 -7386
rect 249882 -7622 249914 -7386
rect 249294 -7654 249914 -7622
rect 253794 704838 254414 711590
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 543454 254414 578898
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 507454 254414 542898
rect 253794 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 254414 507454
rect 253794 507134 254414 507218
rect 253794 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 254414 507134
rect 253794 471454 254414 506898
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 253794 435454 254414 470898
rect 253794 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 254414 435454
rect 253794 435134 254414 435218
rect 253794 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 254414 435134
rect 253794 399454 254414 434898
rect 253794 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 254414 399454
rect 253794 399134 254414 399218
rect 253794 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 254414 399134
rect 253794 363454 254414 398898
rect 253794 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 254414 363454
rect 253794 363134 254414 363218
rect 253794 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 254414 363134
rect 253794 327454 254414 362898
rect 253794 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 254414 327454
rect 253794 327134 254414 327218
rect 253794 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 254414 327134
rect 253794 291454 254414 326898
rect 253794 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 254414 291454
rect 253794 291134 254414 291218
rect 253794 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 254414 291134
rect 253794 255454 254414 290898
rect 253794 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 254414 255454
rect 253794 255134 254414 255218
rect 253794 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 254414 255134
rect 253794 219454 254414 254898
rect 253794 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 254414 219454
rect 253794 219134 254414 219218
rect 253794 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 254414 219134
rect 253794 183454 254414 218898
rect 253794 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 254414 183454
rect 253794 183134 254414 183218
rect 253794 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 254414 183134
rect 253794 147454 254414 182898
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 253794 111454 254414 146898
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 253794 75454 254414 110898
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -7654 254414 -902
rect 258294 705798 258914 711590
rect 258294 705562 258326 705798
rect 258562 705562 258646 705798
rect 258882 705562 258914 705798
rect 258294 705478 258914 705562
rect 258294 705242 258326 705478
rect 258562 705242 258646 705478
rect 258882 705242 258914 705478
rect 258294 691954 258914 705242
rect 258294 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 258914 691954
rect 258294 691634 258914 691718
rect 258294 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 258914 691634
rect 258294 655954 258914 691398
rect 258294 655718 258326 655954
rect 258562 655718 258646 655954
rect 258882 655718 258914 655954
rect 258294 655634 258914 655718
rect 258294 655398 258326 655634
rect 258562 655398 258646 655634
rect 258882 655398 258914 655634
rect 258294 619954 258914 655398
rect 258294 619718 258326 619954
rect 258562 619718 258646 619954
rect 258882 619718 258914 619954
rect 258294 619634 258914 619718
rect 258294 619398 258326 619634
rect 258562 619398 258646 619634
rect 258882 619398 258914 619634
rect 258294 583954 258914 619398
rect 258294 583718 258326 583954
rect 258562 583718 258646 583954
rect 258882 583718 258914 583954
rect 258294 583634 258914 583718
rect 258294 583398 258326 583634
rect 258562 583398 258646 583634
rect 258882 583398 258914 583634
rect 258294 547954 258914 583398
rect 258294 547718 258326 547954
rect 258562 547718 258646 547954
rect 258882 547718 258914 547954
rect 258294 547634 258914 547718
rect 258294 547398 258326 547634
rect 258562 547398 258646 547634
rect 258882 547398 258914 547634
rect 258294 511954 258914 547398
rect 258294 511718 258326 511954
rect 258562 511718 258646 511954
rect 258882 511718 258914 511954
rect 258294 511634 258914 511718
rect 258294 511398 258326 511634
rect 258562 511398 258646 511634
rect 258882 511398 258914 511634
rect 258294 475954 258914 511398
rect 258294 475718 258326 475954
rect 258562 475718 258646 475954
rect 258882 475718 258914 475954
rect 258294 475634 258914 475718
rect 258294 475398 258326 475634
rect 258562 475398 258646 475634
rect 258882 475398 258914 475634
rect 258294 439954 258914 475398
rect 258294 439718 258326 439954
rect 258562 439718 258646 439954
rect 258882 439718 258914 439954
rect 258294 439634 258914 439718
rect 258294 439398 258326 439634
rect 258562 439398 258646 439634
rect 258882 439398 258914 439634
rect 258294 403954 258914 439398
rect 258294 403718 258326 403954
rect 258562 403718 258646 403954
rect 258882 403718 258914 403954
rect 258294 403634 258914 403718
rect 258294 403398 258326 403634
rect 258562 403398 258646 403634
rect 258882 403398 258914 403634
rect 258294 367954 258914 403398
rect 258294 367718 258326 367954
rect 258562 367718 258646 367954
rect 258882 367718 258914 367954
rect 258294 367634 258914 367718
rect 258294 367398 258326 367634
rect 258562 367398 258646 367634
rect 258882 367398 258914 367634
rect 258294 331954 258914 367398
rect 258294 331718 258326 331954
rect 258562 331718 258646 331954
rect 258882 331718 258914 331954
rect 258294 331634 258914 331718
rect 258294 331398 258326 331634
rect 258562 331398 258646 331634
rect 258882 331398 258914 331634
rect 258294 295954 258914 331398
rect 258294 295718 258326 295954
rect 258562 295718 258646 295954
rect 258882 295718 258914 295954
rect 258294 295634 258914 295718
rect 258294 295398 258326 295634
rect 258562 295398 258646 295634
rect 258882 295398 258914 295634
rect 258294 259954 258914 295398
rect 258294 259718 258326 259954
rect 258562 259718 258646 259954
rect 258882 259718 258914 259954
rect 258294 259634 258914 259718
rect 258294 259398 258326 259634
rect 258562 259398 258646 259634
rect 258882 259398 258914 259634
rect 258294 223954 258914 259398
rect 258294 223718 258326 223954
rect 258562 223718 258646 223954
rect 258882 223718 258914 223954
rect 258294 223634 258914 223718
rect 258294 223398 258326 223634
rect 258562 223398 258646 223634
rect 258882 223398 258914 223634
rect 258294 187954 258914 223398
rect 258294 187718 258326 187954
rect 258562 187718 258646 187954
rect 258882 187718 258914 187954
rect 258294 187634 258914 187718
rect 258294 187398 258326 187634
rect 258562 187398 258646 187634
rect 258882 187398 258914 187634
rect 258294 151954 258914 187398
rect 258294 151718 258326 151954
rect 258562 151718 258646 151954
rect 258882 151718 258914 151954
rect 258294 151634 258914 151718
rect 258294 151398 258326 151634
rect 258562 151398 258646 151634
rect 258882 151398 258914 151634
rect 258294 115954 258914 151398
rect 258294 115718 258326 115954
rect 258562 115718 258646 115954
rect 258882 115718 258914 115954
rect 258294 115634 258914 115718
rect 258294 115398 258326 115634
rect 258562 115398 258646 115634
rect 258882 115398 258914 115634
rect 258294 79954 258914 115398
rect 258294 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 258914 79954
rect 258294 79634 258914 79718
rect 258294 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 258914 79634
rect 258294 43954 258914 79398
rect 258294 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 258914 43954
rect 258294 43634 258914 43718
rect 258294 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 258914 43634
rect 258294 7954 258914 43398
rect 258294 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 258914 7954
rect 258294 7634 258914 7718
rect 258294 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 258914 7634
rect 258294 -1306 258914 7398
rect 258294 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 258914 -1306
rect 258294 -1626 258914 -1542
rect 258294 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 258914 -1626
rect 258294 -7654 258914 -1862
rect 262794 706758 263414 711590
rect 262794 706522 262826 706758
rect 263062 706522 263146 706758
rect 263382 706522 263414 706758
rect 262794 706438 263414 706522
rect 262794 706202 262826 706438
rect 263062 706202 263146 706438
rect 263382 706202 263414 706438
rect 262794 696454 263414 706202
rect 262794 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 263414 696454
rect 262794 696134 263414 696218
rect 262794 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 263414 696134
rect 262794 660454 263414 695898
rect 262794 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 263414 660454
rect 262794 660134 263414 660218
rect 262794 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 263414 660134
rect 262794 624454 263414 659898
rect 262794 624218 262826 624454
rect 263062 624218 263146 624454
rect 263382 624218 263414 624454
rect 262794 624134 263414 624218
rect 262794 623898 262826 624134
rect 263062 623898 263146 624134
rect 263382 623898 263414 624134
rect 262794 588454 263414 623898
rect 262794 588218 262826 588454
rect 263062 588218 263146 588454
rect 263382 588218 263414 588454
rect 262794 588134 263414 588218
rect 262794 587898 262826 588134
rect 263062 587898 263146 588134
rect 263382 587898 263414 588134
rect 262794 552454 263414 587898
rect 262794 552218 262826 552454
rect 263062 552218 263146 552454
rect 263382 552218 263414 552454
rect 262794 552134 263414 552218
rect 262794 551898 262826 552134
rect 263062 551898 263146 552134
rect 263382 551898 263414 552134
rect 262794 516454 263414 551898
rect 262794 516218 262826 516454
rect 263062 516218 263146 516454
rect 263382 516218 263414 516454
rect 262794 516134 263414 516218
rect 262794 515898 262826 516134
rect 263062 515898 263146 516134
rect 263382 515898 263414 516134
rect 262794 480454 263414 515898
rect 262794 480218 262826 480454
rect 263062 480218 263146 480454
rect 263382 480218 263414 480454
rect 262794 480134 263414 480218
rect 262794 479898 262826 480134
rect 263062 479898 263146 480134
rect 263382 479898 263414 480134
rect 262794 444454 263414 479898
rect 262794 444218 262826 444454
rect 263062 444218 263146 444454
rect 263382 444218 263414 444454
rect 262794 444134 263414 444218
rect 262794 443898 262826 444134
rect 263062 443898 263146 444134
rect 263382 443898 263414 444134
rect 262794 408454 263414 443898
rect 262794 408218 262826 408454
rect 263062 408218 263146 408454
rect 263382 408218 263414 408454
rect 262794 408134 263414 408218
rect 262794 407898 262826 408134
rect 263062 407898 263146 408134
rect 263382 407898 263414 408134
rect 262794 372454 263414 407898
rect 262794 372218 262826 372454
rect 263062 372218 263146 372454
rect 263382 372218 263414 372454
rect 262794 372134 263414 372218
rect 262794 371898 262826 372134
rect 263062 371898 263146 372134
rect 263382 371898 263414 372134
rect 262794 336454 263414 371898
rect 262794 336218 262826 336454
rect 263062 336218 263146 336454
rect 263382 336218 263414 336454
rect 262794 336134 263414 336218
rect 262794 335898 262826 336134
rect 263062 335898 263146 336134
rect 263382 335898 263414 336134
rect 262794 300454 263414 335898
rect 262794 300218 262826 300454
rect 263062 300218 263146 300454
rect 263382 300218 263414 300454
rect 262794 300134 263414 300218
rect 262794 299898 262826 300134
rect 263062 299898 263146 300134
rect 263382 299898 263414 300134
rect 262794 264454 263414 299898
rect 262794 264218 262826 264454
rect 263062 264218 263146 264454
rect 263382 264218 263414 264454
rect 262794 264134 263414 264218
rect 262794 263898 262826 264134
rect 263062 263898 263146 264134
rect 263382 263898 263414 264134
rect 262794 228454 263414 263898
rect 262794 228218 262826 228454
rect 263062 228218 263146 228454
rect 263382 228218 263414 228454
rect 262794 228134 263414 228218
rect 262794 227898 262826 228134
rect 263062 227898 263146 228134
rect 263382 227898 263414 228134
rect 262794 192454 263414 227898
rect 262794 192218 262826 192454
rect 263062 192218 263146 192454
rect 263382 192218 263414 192454
rect 262794 192134 263414 192218
rect 262794 191898 262826 192134
rect 263062 191898 263146 192134
rect 263382 191898 263414 192134
rect 262794 156454 263414 191898
rect 262794 156218 262826 156454
rect 263062 156218 263146 156454
rect 263382 156218 263414 156454
rect 262794 156134 263414 156218
rect 262794 155898 262826 156134
rect 263062 155898 263146 156134
rect 263382 155898 263414 156134
rect 262794 120454 263414 155898
rect 262794 120218 262826 120454
rect 263062 120218 263146 120454
rect 263382 120218 263414 120454
rect 262794 120134 263414 120218
rect 262794 119898 262826 120134
rect 263062 119898 263146 120134
rect 263382 119898 263414 120134
rect 262794 84454 263414 119898
rect 262794 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 263414 84454
rect 262794 84134 263414 84218
rect 262794 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 263414 84134
rect 262794 48454 263414 83898
rect 262794 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 263414 48454
rect 262794 48134 263414 48218
rect 262794 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 263414 48134
rect 262794 12454 263414 47898
rect 262794 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 263414 12454
rect 262794 12134 263414 12218
rect 262794 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 263414 12134
rect 262794 -2266 263414 11898
rect 262794 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 263414 -2266
rect 262794 -2586 263414 -2502
rect 262794 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 263414 -2586
rect 262794 -7654 263414 -2822
rect 267294 707718 267914 711590
rect 267294 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 267914 707718
rect 267294 707398 267914 707482
rect 267294 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 267914 707398
rect 267294 700954 267914 707162
rect 267294 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 267914 700954
rect 267294 700634 267914 700718
rect 267294 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 267914 700634
rect 267294 664954 267914 700398
rect 267294 664718 267326 664954
rect 267562 664718 267646 664954
rect 267882 664718 267914 664954
rect 267294 664634 267914 664718
rect 267294 664398 267326 664634
rect 267562 664398 267646 664634
rect 267882 664398 267914 664634
rect 267294 628954 267914 664398
rect 267294 628718 267326 628954
rect 267562 628718 267646 628954
rect 267882 628718 267914 628954
rect 267294 628634 267914 628718
rect 267294 628398 267326 628634
rect 267562 628398 267646 628634
rect 267882 628398 267914 628634
rect 267294 592954 267914 628398
rect 267294 592718 267326 592954
rect 267562 592718 267646 592954
rect 267882 592718 267914 592954
rect 267294 592634 267914 592718
rect 267294 592398 267326 592634
rect 267562 592398 267646 592634
rect 267882 592398 267914 592634
rect 267294 556954 267914 592398
rect 267294 556718 267326 556954
rect 267562 556718 267646 556954
rect 267882 556718 267914 556954
rect 267294 556634 267914 556718
rect 267294 556398 267326 556634
rect 267562 556398 267646 556634
rect 267882 556398 267914 556634
rect 267294 520954 267914 556398
rect 267294 520718 267326 520954
rect 267562 520718 267646 520954
rect 267882 520718 267914 520954
rect 267294 520634 267914 520718
rect 267294 520398 267326 520634
rect 267562 520398 267646 520634
rect 267882 520398 267914 520634
rect 267294 484954 267914 520398
rect 267294 484718 267326 484954
rect 267562 484718 267646 484954
rect 267882 484718 267914 484954
rect 267294 484634 267914 484718
rect 267294 484398 267326 484634
rect 267562 484398 267646 484634
rect 267882 484398 267914 484634
rect 267294 448954 267914 484398
rect 267294 448718 267326 448954
rect 267562 448718 267646 448954
rect 267882 448718 267914 448954
rect 267294 448634 267914 448718
rect 267294 448398 267326 448634
rect 267562 448398 267646 448634
rect 267882 448398 267914 448634
rect 267294 412954 267914 448398
rect 267294 412718 267326 412954
rect 267562 412718 267646 412954
rect 267882 412718 267914 412954
rect 267294 412634 267914 412718
rect 267294 412398 267326 412634
rect 267562 412398 267646 412634
rect 267882 412398 267914 412634
rect 267294 376954 267914 412398
rect 267294 376718 267326 376954
rect 267562 376718 267646 376954
rect 267882 376718 267914 376954
rect 267294 376634 267914 376718
rect 267294 376398 267326 376634
rect 267562 376398 267646 376634
rect 267882 376398 267914 376634
rect 267294 340954 267914 376398
rect 267294 340718 267326 340954
rect 267562 340718 267646 340954
rect 267882 340718 267914 340954
rect 267294 340634 267914 340718
rect 267294 340398 267326 340634
rect 267562 340398 267646 340634
rect 267882 340398 267914 340634
rect 267294 304954 267914 340398
rect 267294 304718 267326 304954
rect 267562 304718 267646 304954
rect 267882 304718 267914 304954
rect 267294 304634 267914 304718
rect 267294 304398 267326 304634
rect 267562 304398 267646 304634
rect 267882 304398 267914 304634
rect 267294 268954 267914 304398
rect 267294 268718 267326 268954
rect 267562 268718 267646 268954
rect 267882 268718 267914 268954
rect 267294 268634 267914 268718
rect 267294 268398 267326 268634
rect 267562 268398 267646 268634
rect 267882 268398 267914 268634
rect 267294 232954 267914 268398
rect 267294 232718 267326 232954
rect 267562 232718 267646 232954
rect 267882 232718 267914 232954
rect 267294 232634 267914 232718
rect 267294 232398 267326 232634
rect 267562 232398 267646 232634
rect 267882 232398 267914 232634
rect 267294 196954 267914 232398
rect 267294 196718 267326 196954
rect 267562 196718 267646 196954
rect 267882 196718 267914 196954
rect 267294 196634 267914 196718
rect 267294 196398 267326 196634
rect 267562 196398 267646 196634
rect 267882 196398 267914 196634
rect 267294 160954 267914 196398
rect 267294 160718 267326 160954
rect 267562 160718 267646 160954
rect 267882 160718 267914 160954
rect 267294 160634 267914 160718
rect 267294 160398 267326 160634
rect 267562 160398 267646 160634
rect 267882 160398 267914 160634
rect 267294 124954 267914 160398
rect 267294 124718 267326 124954
rect 267562 124718 267646 124954
rect 267882 124718 267914 124954
rect 267294 124634 267914 124718
rect 267294 124398 267326 124634
rect 267562 124398 267646 124634
rect 267882 124398 267914 124634
rect 267294 88954 267914 124398
rect 267294 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 267914 88954
rect 267294 88634 267914 88718
rect 267294 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 267914 88634
rect 267294 52954 267914 88398
rect 267294 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 267914 52954
rect 267294 52634 267914 52718
rect 267294 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 267914 52634
rect 267294 16954 267914 52398
rect 267294 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 267914 16954
rect 267294 16634 267914 16718
rect 267294 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 267914 16634
rect 267294 -3226 267914 16398
rect 267294 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 267914 -3226
rect 267294 -3546 267914 -3462
rect 267294 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 267914 -3546
rect 267294 -7654 267914 -3782
rect 271794 708678 272414 711590
rect 271794 708442 271826 708678
rect 272062 708442 272146 708678
rect 272382 708442 272414 708678
rect 271794 708358 272414 708442
rect 271794 708122 271826 708358
rect 272062 708122 272146 708358
rect 272382 708122 272414 708358
rect 271794 669454 272414 708122
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 561454 272414 596898
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 525454 272414 560898
rect 271794 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 272414 525454
rect 271794 525134 272414 525218
rect 271794 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 272414 525134
rect 271794 489454 272414 524898
rect 271794 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 272414 489454
rect 271794 489134 272414 489218
rect 271794 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 272414 489134
rect 271794 453454 272414 488898
rect 271794 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 272414 453454
rect 271794 453134 272414 453218
rect 271794 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 272414 453134
rect 271794 417454 272414 452898
rect 271794 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 272414 417454
rect 271794 417134 272414 417218
rect 271794 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 272414 417134
rect 271794 381454 272414 416898
rect 271794 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 272414 381454
rect 271794 381134 272414 381218
rect 271794 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 272414 381134
rect 271794 345454 272414 380898
rect 271794 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 272414 345454
rect 271794 345134 272414 345218
rect 271794 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 272414 345134
rect 271794 309454 272414 344898
rect 271794 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 272414 309454
rect 271794 309134 272414 309218
rect 271794 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 272414 309134
rect 271794 273454 272414 308898
rect 271794 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 272414 273454
rect 271794 273134 272414 273218
rect 271794 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 272414 273134
rect 271794 237454 272414 272898
rect 271794 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 272414 237454
rect 271794 237134 272414 237218
rect 271794 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 272414 237134
rect 271794 201454 272414 236898
rect 271794 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 272414 201454
rect 271794 201134 272414 201218
rect 271794 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 272414 201134
rect 271794 165454 272414 200898
rect 271794 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 272414 165454
rect 271794 165134 272414 165218
rect 271794 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 272414 165134
rect 271794 129454 272414 164898
rect 271794 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 272414 129454
rect 271794 129134 272414 129218
rect 271794 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 272414 129134
rect 271794 93454 272414 128898
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271794 57454 272414 92898
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -4186 272414 20898
rect 271794 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 272414 -4186
rect 271794 -4506 272414 -4422
rect 271794 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 272414 -4506
rect 271794 -7654 272414 -4742
rect 276294 709638 276914 711590
rect 276294 709402 276326 709638
rect 276562 709402 276646 709638
rect 276882 709402 276914 709638
rect 276294 709318 276914 709402
rect 276294 709082 276326 709318
rect 276562 709082 276646 709318
rect 276882 709082 276914 709318
rect 276294 673954 276914 709082
rect 276294 673718 276326 673954
rect 276562 673718 276646 673954
rect 276882 673718 276914 673954
rect 276294 673634 276914 673718
rect 276294 673398 276326 673634
rect 276562 673398 276646 673634
rect 276882 673398 276914 673634
rect 276294 637954 276914 673398
rect 276294 637718 276326 637954
rect 276562 637718 276646 637954
rect 276882 637718 276914 637954
rect 276294 637634 276914 637718
rect 276294 637398 276326 637634
rect 276562 637398 276646 637634
rect 276882 637398 276914 637634
rect 276294 601954 276914 637398
rect 276294 601718 276326 601954
rect 276562 601718 276646 601954
rect 276882 601718 276914 601954
rect 276294 601634 276914 601718
rect 276294 601398 276326 601634
rect 276562 601398 276646 601634
rect 276882 601398 276914 601634
rect 276294 565954 276914 601398
rect 276294 565718 276326 565954
rect 276562 565718 276646 565954
rect 276882 565718 276914 565954
rect 276294 565634 276914 565718
rect 276294 565398 276326 565634
rect 276562 565398 276646 565634
rect 276882 565398 276914 565634
rect 276294 529954 276914 565398
rect 276294 529718 276326 529954
rect 276562 529718 276646 529954
rect 276882 529718 276914 529954
rect 276294 529634 276914 529718
rect 276294 529398 276326 529634
rect 276562 529398 276646 529634
rect 276882 529398 276914 529634
rect 276294 493954 276914 529398
rect 276294 493718 276326 493954
rect 276562 493718 276646 493954
rect 276882 493718 276914 493954
rect 276294 493634 276914 493718
rect 276294 493398 276326 493634
rect 276562 493398 276646 493634
rect 276882 493398 276914 493634
rect 276294 457954 276914 493398
rect 276294 457718 276326 457954
rect 276562 457718 276646 457954
rect 276882 457718 276914 457954
rect 276294 457634 276914 457718
rect 276294 457398 276326 457634
rect 276562 457398 276646 457634
rect 276882 457398 276914 457634
rect 276294 421954 276914 457398
rect 276294 421718 276326 421954
rect 276562 421718 276646 421954
rect 276882 421718 276914 421954
rect 276294 421634 276914 421718
rect 276294 421398 276326 421634
rect 276562 421398 276646 421634
rect 276882 421398 276914 421634
rect 276294 385954 276914 421398
rect 276294 385718 276326 385954
rect 276562 385718 276646 385954
rect 276882 385718 276914 385954
rect 276294 385634 276914 385718
rect 276294 385398 276326 385634
rect 276562 385398 276646 385634
rect 276882 385398 276914 385634
rect 276294 349954 276914 385398
rect 276294 349718 276326 349954
rect 276562 349718 276646 349954
rect 276882 349718 276914 349954
rect 276294 349634 276914 349718
rect 276294 349398 276326 349634
rect 276562 349398 276646 349634
rect 276882 349398 276914 349634
rect 276294 313954 276914 349398
rect 276294 313718 276326 313954
rect 276562 313718 276646 313954
rect 276882 313718 276914 313954
rect 276294 313634 276914 313718
rect 276294 313398 276326 313634
rect 276562 313398 276646 313634
rect 276882 313398 276914 313634
rect 276294 277954 276914 313398
rect 276294 277718 276326 277954
rect 276562 277718 276646 277954
rect 276882 277718 276914 277954
rect 276294 277634 276914 277718
rect 276294 277398 276326 277634
rect 276562 277398 276646 277634
rect 276882 277398 276914 277634
rect 276294 241954 276914 277398
rect 276294 241718 276326 241954
rect 276562 241718 276646 241954
rect 276882 241718 276914 241954
rect 276294 241634 276914 241718
rect 276294 241398 276326 241634
rect 276562 241398 276646 241634
rect 276882 241398 276914 241634
rect 276294 205954 276914 241398
rect 276294 205718 276326 205954
rect 276562 205718 276646 205954
rect 276882 205718 276914 205954
rect 276294 205634 276914 205718
rect 276294 205398 276326 205634
rect 276562 205398 276646 205634
rect 276882 205398 276914 205634
rect 276294 169954 276914 205398
rect 276294 169718 276326 169954
rect 276562 169718 276646 169954
rect 276882 169718 276914 169954
rect 276294 169634 276914 169718
rect 276294 169398 276326 169634
rect 276562 169398 276646 169634
rect 276882 169398 276914 169634
rect 276294 133954 276914 169398
rect 276294 133718 276326 133954
rect 276562 133718 276646 133954
rect 276882 133718 276914 133954
rect 276294 133634 276914 133718
rect 276294 133398 276326 133634
rect 276562 133398 276646 133634
rect 276882 133398 276914 133634
rect 276294 97954 276914 133398
rect 276294 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 276914 97954
rect 276294 97634 276914 97718
rect 276294 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 276914 97634
rect 276294 61954 276914 97398
rect 276294 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 276914 61954
rect 276294 61634 276914 61718
rect 276294 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 276914 61634
rect 276294 25954 276914 61398
rect 276294 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 276914 25954
rect 276294 25634 276914 25718
rect 276294 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 276914 25634
rect 276294 -5146 276914 25398
rect 276294 -5382 276326 -5146
rect 276562 -5382 276646 -5146
rect 276882 -5382 276914 -5146
rect 276294 -5466 276914 -5382
rect 276294 -5702 276326 -5466
rect 276562 -5702 276646 -5466
rect 276882 -5702 276914 -5466
rect 276294 -7654 276914 -5702
rect 280794 710598 281414 711590
rect 280794 710362 280826 710598
rect 281062 710362 281146 710598
rect 281382 710362 281414 710598
rect 280794 710278 281414 710362
rect 280794 710042 280826 710278
rect 281062 710042 281146 710278
rect 281382 710042 281414 710278
rect 280794 678454 281414 710042
rect 280794 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 281414 678454
rect 280794 678134 281414 678218
rect 280794 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 281414 678134
rect 280794 642454 281414 677898
rect 280794 642218 280826 642454
rect 281062 642218 281146 642454
rect 281382 642218 281414 642454
rect 280794 642134 281414 642218
rect 280794 641898 280826 642134
rect 281062 641898 281146 642134
rect 281382 641898 281414 642134
rect 280794 606454 281414 641898
rect 280794 606218 280826 606454
rect 281062 606218 281146 606454
rect 281382 606218 281414 606454
rect 280794 606134 281414 606218
rect 280794 605898 280826 606134
rect 281062 605898 281146 606134
rect 281382 605898 281414 606134
rect 280794 570454 281414 605898
rect 280794 570218 280826 570454
rect 281062 570218 281146 570454
rect 281382 570218 281414 570454
rect 280794 570134 281414 570218
rect 280794 569898 280826 570134
rect 281062 569898 281146 570134
rect 281382 569898 281414 570134
rect 280794 534454 281414 569898
rect 280794 534218 280826 534454
rect 281062 534218 281146 534454
rect 281382 534218 281414 534454
rect 280794 534134 281414 534218
rect 280794 533898 280826 534134
rect 281062 533898 281146 534134
rect 281382 533898 281414 534134
rect 280794 498454 281414 533898
rect 280794 498218 280826 498454
rect 281062 498218 281146 498454
rect 281382 498218 281414 498454
rect 280794 498134 281414 498218
rect 280794 497898 280826 498134
rect 281062 497898 281146 498134
rect 281382 497898 281414 498134
rect 280794 462454 281414 497898
rect 280794 462218 280826 462454
rect 281062 462218 281146 462454
rect 281382 462218 281414 462454
rect 280794 462134 281414 462218
rect 280794 461898 280826 462134
rect 281062 461898 281146 462134
rect 281382 461898 281414 462134
rect 280794 426454 281414 461898
rect 280794 426218 280826 426454
rect 281062 426218 281146 426454
rect 281382 426218 281414 426454
rect 280794 426134 281414 426218
rect 280794 425898 280826 426134
rect 281062 425898 281146 426134
rect 281382 425898 281414 426134
rect 280794 390454 281414 425898
rect 280794 390218 280826 390454
rect 281062 390218 281146 390454
rect 281382 390218 281414 390454
rect 280794 390134 281414 390218
rect 280794 389898 280826 390134
rect 281062 389898 281146 390134
rect 281382 389898 281414 390134
rect 280794 354454 281414 389898
rect 280794 354218 280826 354454
rect 281062 354218 281146 354454
rect 281382 354218 281414 354454
rect 280794 354134 281414 354218
rect 280794 353898 280826 354134
rect 281062 353898 281146 354134
rect 281382 353898 281414 354134
rect 280794 318454 281414 353898
rect 280794 318218 280826 318454
rect 281062 318218 281146 318454
rect 281382 318218 281414 318454
rect 280794 318134 281414 318218
rect 280794 317898 280826 318134
rect 281062 317898 281146 318134
rect 281382 317898 281414 318134
rect 280794 282454 281414 317898
rect 280794 282218 280826 282454
rect 281062 282218 281146 282454
rect 281382 282218 281414 282454
rect 280794 282134 281414 282218
rect 280794 281898 280826 282134
rect 281062 281898 281146 282134
rect 281382 281898 281414 282134
rect 280794 246454 281414 281898
rect 280794 246218 280826 246454
rect 281062 246218 281146 246454
rect 281382 246218 281414 246454
rect 280794 246134 281414 246218
rect 280794 245898 280826 246134
rect 281062 245898 281146 246134
rect 281382 245898 281414 246134
rect 280794 210454 281414 245898
rect 280794 210218 280826 210454
rect 281062 210218 281146 210454
rect 281382 210218 281414 210454
rect 280794 210134 281414 210218
rect 280794 209898 280826 210134
rect 281062 209898 281146 210134
rect 281382 209898 281414 210134
rect 280794 174454 281414 209898
rect 280794 174218 280826 174454
rect 281062 174218 281146 174454
rect 281382 174218 281414 174454
rect 280794 174134 281414 174218
rect 280794 173898 280826 174134
rect 281062 173898 281146 174134
rect 281382 173898 281414 174134
rect 280794 138454 281414 173898
rect 280794 138218 280826 138454
rect 281062 138218 281146 138454
rect 281382 138218 281414 138454
rect 280794 138134 281414 138218
rect 280794 137898 280826 138134
rect 281062 137898 281146 138134
rect 281382 137898 281414 138134
rect 280794 102454 281414 137898
rect 280794 102218 280826 102454
rect 281062 102218 281146 102454
rect 281382 102218 281414 102454
rect 280794 102134 281414 102218
rect 280794 101898 280826 102134
rect 281062 101898 281146 102134
rect 281382 101898 281414 102134
rect 280794 66454 281414 101898
rect 280794 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 281414 66454
rect 280794 66134 281414 66218
rect 280794 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 281414 66134
rect 280794 30454 281414 65898
rect 280794 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 281414 30454
rect 280794 30134 281414 30218
rect 280794 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 281414 30134
rect 280794 -6106 281414 29898
rect 280794 -6342 280826 -6106
rect 281062 -6342 281146 -6106
rect 281382 -6342 281414 -6106
rect 280794 -6426 281414 -6342
rect 280794 -6662 280826 -6426
rect 281062 -6662 281146 -6426
rect 281382 -6662 281414 -6426
rect 280794 -7654 281414 -6662
rect 285294 711558 285914 711590
rect 285294 711322 285326 711558
rect 285562 711322 285646 711558
rect 285882 711322 285914 711558
rect 285294 711238 285914 711322
rect 285294 711002 285326 711238
rect 285562 711002 285646 711238
rect 285882 711002 285914 711238
rect 285294 682954 285914 711002
rect 285294 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 285914 682954
rect 285294 682634 285914 682718
rect 285294 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 285914 682634
rect 285294 646954 285914 682398
rect 285294 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 285914 646954
rect 285294 646634 285914 646718
rect 285294 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 285914 646634
rect 285294 610954 285914 646398
rect 285294 610718 285326 610954
rect 285562 610718 285646 610954
rect 285882 610718 285914 610954
rect 285294 610634 285914 610718
rect 285294 610398 285326 610634
rect 285562 610398 285646 610634
rect 285882 610398 285914 610634
rect 285294 574954 285914 610398
rect 285294 574718 285326 574954
rect 285562 574718 285646 574954
rect 285882 574718 285914 574954
rect 285294 574634 285914 574718
rect 285294 574398 285326 574634
rect 285562 574398 285646 574634
rect 285882 574398 285914 574634
rect 285294 538954 285914 574398
rect 285294 538718 285326 538954
rect 285562 538718 285646 538954
rect 285882 538718 285914 538954
rect 285294 538634 285914 538718
rect 285294 538398 285326 538634
rect 285562 538398 285646 538634
rect 285882 538398 285914 538634
rect 285294 502954 285914 538398
rect 285294 502718 285326 502954
rect 285562 502718 285646 502954
rect 285882 502718 285914 502954
rect 285294 502634 285914 502718
rect 285294 502398 285326 502634
rect 285562 502398 285646 502634
rect 285882 502398 285914 502634
rect 285294 466954 285914 502398
rect 285294 466718 285326 466954
rect 285562 466718 285646 466954
rect 285882 466718 285914 466954
rect 285294 466634 285914 466718
rect 285294 466398 285326 466634
rect 285562 466398 285646 466634
rect 285882 466398 285914 466634
rect 285294 430954 285914 466398
rect 285294 430718 285326 430954
rect 285562 430718 285646 430954
rect 285882 430718 285914 430954
rect 285294 430634 285914 430718
rect 285294 430398 285326 430634
rect 285562 430398 285646 430634
rect 285882 430398 285914 430634
rect 285294 394954 285914 430398
rect 285294 394718 285326 394954
rect 285562 394718 285646 394954
rect 285882 394718 285914 394954
rect 285294 394634 285914 394718
rect 285294 394398 285326 394634
rect 285562 394398 285646 394634
rect 285882 394398 285914 394634
rect 285294 358954 285914 394398
rect 285294 358718 285326 358954
rect 285562 358718 285646 358954
rect 285882 358718 285914 358954
rect 285294 358634 285914 358718
rect 285294 358398 285326 358634
rect 285562 358398 285646 358634
rect 285882 358398 285914 358634
rect 285294 322954 285914 358398
rect 285294 322718 285326 322954
rect 285562 322718 285646 322954
rect 285882 322718 285914 322954
rect 285294 322634 285914 322718
rect 285294 322398 285326 322634
rect 285562 322398 285646 322634
rect 285882 322398 285914 322634
rect 285294 286954 285914 322398
rect 285294 286718 285326 286954
rect 285562 286718 285646 286954
rect 285882 286718 285914 286954
rect 285294 286634 285914 286718
rect 285294 286398 285326 286634
rect 285562 286398 285646 286634
rect 285882 286398 285914 286634
rect 285294 250954 285914 286398
rect 285294 250718 285326 250954
rect 285562 250718 285646 250954
rect 285882 250718 285914 250954
rect 285294 250634 285914 250718
rect 285294 250398 285326 250634
rect 285562 250398 285646 250634
rect 285882 250398 285914 250634
rect 285294 214954 285914 250398
rect 285294 214718 285326 214954
rect 285562 214718 285646 214954
rect 285882 214718 285914 214954
rect 285294 214634 285914 214718
rect 285294 214398 285326 214634
rect 285562 214398 285646 214634
rect 285882 214398 285914 214634
rect 285294 178954 285914 214398
rect 285294 178718 285326 178954
rect 285562 178718 285646 178954
rect 285882 178718 285914 178954
rect 285294 178634 285914 178718
rect 285294 178398 285326 178634
rect 285562 178398 285646 178634
rect 285882 178398 285914 178634
rect 285294 142954 285914 178398
rect 285294 142718 285326 142954
rect 285562 142718 285646 142954
rect 285882 142718 285914 142954
rect 285294 142634 285914 142718
rect 285294 142398 285326 142634
rect 285562 142398 285646 142634
rect 285882 142398 285914 142634
rect 285294 106954 285914 142398
rect 285294 106718 285326 106954
rect 285562 106718 285646 106954
rect 285882 106718 285914 106954
rect 285294 106634 285914 106718
rect 285294 106398 285326 106634
rect 285562 106398 285646 106634
rect 285882 106398 285914 106634
rect 285294 70954 285914 106398
rect 285294 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 285914 70954
rect 285294 70634 285914 70718
rect 285294 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 285914 70634
rect 285294 34954 285914 70398
rect 285294 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 285914 34954
rect 285294 34634 285914 34718
rect 285294 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 285914 34634
rect 285294 -7066 285914 34398
rect 285294 -7302 285326 -7066
rect 285562 -7302 285646 -7066
rect 285882 -7302 285914 -7066
rect 285294 -7386 285914 -7302
rect 285294 -7622 285326 -7386
rect 285562 -7622 285646 -7386
rect 285882 -7622 285914 -7386
rect 285294 -7654 285914 -7622
rect 289794 704838 290414 711590
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 289794 471454 290414 506898
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 435454 290414 470898
rect 289794 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 290414 435454
rect 289794 435134 290414 435218
rect 289794 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 290414 435134
rect 289794 399454 290414 434898
rect 289794 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 290414 399454
rect 289794 399134 290414 399218
rect 289794 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 290414 399134
rect 289794 363454 290414 398898
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 289794 327454 290414 362898
rect 289794 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 290414 327454
rect 289794 327134 290414 327218
rect 289794 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 290414 327134
rect 289794 291454 290414 326898
rect 289794 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 290414 291454
rect 289794 291134 290414 291218
rect 289794 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 290414 291134
rect 289794 255454 290414 290898
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 289794 219454 290414 254898
rect 289794 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 290414 219454
rect 289794 219134 290414 219218
rect 289794 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 290414 219134
rect 289794 183454 290414 218898
rect 289794 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 290414 183454
rect 289794 183134 290414 183218
rect 289794 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 290414 183134
rect 289794 147454 290414 182898
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 111454 290414 146898
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 289794 75454 290414 110898
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -7654 290414 -902
rect 294294 705798 294914 711590
rect 294294 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 294914 705798
rect 294294 705478 294914 705562
rect 294294 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 294914 705478
rect 294294 691954 294914 705242
rect 294294 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 294914 691954
rect 294294 691634 294914 691718
rect 294294 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 294914 691634
rect 294294 655954 294914 691398
rect 294294 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 294914 655954
rect 294294 655634 294914 655718
rect 294294 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 294914 655634
rect 294294 619954 294914 655398
rect 294294 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 294914 619954
rect 294294 619634 294914 619718
rect 294294 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 294914 619634
rect 294294 583954 294914 619398
rect 294294 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 294914 583954
rect 294294 583634 294914 583718
rect 294294 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 294914 583634
rect 294294 547954 294914 583398
rect 294294 547718 294326 547954
rect 294562 547718 294646 547954
rect 294882 547718 294914 547954
rect 294294 547634 294914 547718
rect 294294 547398 294326 547634
rect 294562 547398 294646 547634
rect 294882 547398 294914 547634
rect 294294 511954 294914 547398
rect 294294 511718 294326 511954
rect 294562 511718 294646 511954
rect 294882 511718 294914 511954
rect 294294 511634 294914 511718
rect 294294 511398 294326 511634
rect 294562 511398 294646 511634
rect 294882 511398 294914 511634
rect 294294 475954 294914 511398
rect 294294 475718 294326 475954
rect 294562 475718 294646 475954
rect 294882 475718 294914 475954
rect 294294 475634 294914 475718
rect 294294 475398 294326 475634
rect 294562 475398 294646 475634
rect 294882 475398 294914 475634
rect 294294 439954 294914 475398
rect 294294 439718 294326 439954
rect 294562 439718 294646 439954
rect 294882 439718 294914 439954
rect 294294 439634 294914 439718
rect 294294 439398 294326 439634
rect 294562 439398 294646 439634
rect 294882 439398 294914 439634
rect 294294 403954 294914 439398
rect 294294 403718 294326 403954
rect 294562 403718 294646 403954
rect 294882 403718 294914 403954
rect 294294 403634 294914 403718
rect 294294 403398 294326 403634
rect 294562 403398 294646 403634
rect 294882 403398 294914 403634
rect 294294 367954 294914 403398
rect 294294 367718 294326 367954
rect 294562 367718 294646 367954
rect 294882 367718 294914 367954
rect 294294 367634 294914 367718
rect 294294 367398 294326 367634
rect 294562 367398 294646 367634
rect 294882 367398 294914 367634
rect 294294 331954 294914 367398
rect 294294 331718 294326 331954
rect 294562 331718 294646 331954
rect 294882 331718 294914 331954
rect 294294 331634 294914 331718
rect 294294 331398 294326 331634
rect 294562 331398 294646 331634
rect 294882 331398 294914 331634
rect 294294 295954 294914 331398
rect 294294 295718 294326 295954
rect 294562 295718 294646 295954
rect 294882 295718 294914 295954
rect 294294 295634 294914 295718
rect 294294 295398 294326 295634
rect 294562 295398 294646 295634
rect 294882 295398 294914 295634
rect 294294 259954 294914 295398
rect 294294 259718 294326 259954
rect 294562 259718 294646 259954
rect 294882 259718 294914 259954
rect 294294 259634 294914 259718
rect 294294 259398 294326 259634
rect 294562 259398 294646 259634
rect 294882 259398 294914 259634
rect 294294 223954 294914 259398
rect 294294 223718 294326 223954
rect 294562 223718 294646 223954
rect 294882 223718 294914 223954
rect 294294 223634 294914 223718
rect 294294 223398 294326 223634
rect 294562 223398 294646 223634
rect 294882 223398 294914 223634
rect 294294 187954 294914 223398
rect 294294 187718 294326 187954
rect 294562 187718 294646 187954
rect 294882 187718 294914 187954
rect 294294 187634 294914 187718
rect 294294 187398 294326 187634
rect 294562 187398 294646 187634
rect 294882 187398 294914 187634
rect 294294 151954 294914 187398
rect 294294 151718 294326 151954
rect 294562 151718 294646 151954
rect 294882 151718 294914 151954
rect 294294 151634 294914 151718
rect 294294 151398 294326 151634
rect 294562 151398 294646 151634
rect 294882 151398 294914 151634
rect 294294 115954 294914 151398
rect 294294 115718 294326 115954
rect 294562 115718 294646 115954
rect 294882 115718 294914 115954
rect 294294 115634 294914 115718
rect 294294 115398 294326 115634
rect 294562 115398 294646 115634
rect 294882 115398 294914 115634
rect 294294 79954 294914 115398
rect 294294 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 294914 79954
rect 294294 79634 294914 79718
rect 294294 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 294914 79634
rect 294294 43954 294914 79398
rect 294294 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 294914 43954
rect 294294 43634 294914 43718
rect 294294 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 294914 43634
rect 294294 7954 294914 43398
rect 294294 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 294914 7954
rect 294294 7634 294914 7718
rect 294294 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 294914 7634
rect 294294 -1306 294914 7398
rect 294294 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 294914 -1306
rect 294294 -1626 294914 -1542
rect 294294 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 294914 -1626
rect 294294 -7654 294914 -1862
rect 298794 706758 299414 711590
rect 298794 706522 298826 706758
rect 299062 706522 299146 706758
rect 299382 706522 299414 706758
rect 298794 706438 299414 706522
rect 298794 706202 298826 706438
rect 299062 706202 299146 706438
rect 299382 706202 299414 706438
rect 298794 696454 299414 706202
rect 298794 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 299414 696454
rect 298794 696134 299414 696218
rect 298794 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 299414 696134
rect 298794 660454 299414 695898
rect 298794 660218 298826 660454
rect 299062 660218 299146 660454
rect 299382 660218 299414 660454
rect 298794 660134 299414 660218
rect 298794 659898 298826 660134
rect 299062 659898 299146 660134
rect 299382 659898 299414 660134
rect 298794 624454 299414 659898
rect 298794 624218 298826 624454
rect 299062 624218 299146 624454
rect 299382 624218 299414 624454
rect 298794 624134 299414 624218
rect 298794 623898 298826 624134
rect 299062 623898 299146 624134
rect 299382 623898 299414 624134
rect 298794 588454 299414 623898
rect 298794 588218 298826 588454
rect 299062 588218 299146 588454
rect 299382 588218 299414 588454
rect 298794 588134 299414 588218
rect 298794 587898 298826 588134
rect 299062 587898 299146 588134
rect 299382 587898 299414 588134
rect 298794 552454 299414 587898
rect 298794 552218 298826 552454
rect 299062 552218 299146 552454
rect 299382 552218 299414 552454
rect 298794 552134 299414 552218
rect 298794 551898 298826 552134
rect 299062 551898 299146 552134
rect 299382 551898 299414 552134
rect 298794 516454 299414 551898
rect 298794 516218 298826 516454
rect 299062 516218 299146 516454
rect 299382 516218 299414 516454
rect 298794 516134 299414 516218
rect 298794 515898 298826 516134
rect 299062 515898 299146 516134
rect 299382 515898 299414 516134
rect 298794 480454 299414 515898
rect 298794 480218 298826 480454
rect 299062 480218 299146 480454
rect 299382 480218 299414 480454
rect 298794 480134 299414 480218
rect 298794 479898 298826 480134
rect 299062 479898 299146 480134
rect 299382 479898 299414 480134
rect 298794 444454 299414 479898
rect 298794 444218 298826 444454
rect 299062 444218 299146 444454
rect 299382 444218 299414 444454
rect 298794 444134 299414 444218
rect 298794 443898 298826 444134
rect 299062 443898 299146 444134
rect 299382 443898 299414 444134
rect 298794 408454 299414 443898
rect 298794 408218 298826 408454
rect 299062 408218 299146 408454
rect 299382 408218 299414 408454
rect 298794 408134 299414 408218
rect 298794 407898 298826 408134
rect 299062 407898 299146 408134
rect 299382 407898 299414 408134
rect 298794 372454 299414 407898
rect 298794 372218 298826 372454
rect 299062 372218 299146 372454
rect 299382 372218 299414 372454
rect 298794 372134 299414 372218
rect 298794 371898 298826 372134
rect 299062 371898 299146 372134
rect 299382 371898 299414 372134
rect 298794 336454 299414 371898
rect 298794 336218 298826 336454
rect 299062 336218 299146 336454
rect 299382 336218 299414 336454
rect 298794 336134 299414 336218
rect 298794 335898 298826 336134
rect 299062 335898 299146 336134
rect 299382 335898 299414 336134
rect 298794 300454 299414 335898
rect 298794 300218 298826 300454
rect 299062 300218 299146 300454
rect 299382 300218 299414 300454
rect 298794 300134 299414 300218
rect 298794 299898 298826 300134
rect 299062 299898 299146 300134
rect 299382 299898 299414 300134
rect 298794 264454 299414 299898
rect 298794 264218 298826 264454
rect 299062 264218 299146 264454
rect 299382 264218 299414 264454
rect 298794 264134 299414 264218
rect 298794 263898 298826 264134
rect 299062 263898 299146 264134
rect 299382 263898 299414 264134
rect 298794 228454 299414 263898
rect 298794 228218 298826 228454
rect 299062 228218 299146 228454
rect 299382 228218 299414 228454
rect 298794 228134 299414 228218
rect 298794 227898 298826 228134
rect 299062 227898 299146 228134
rect 299382 227898 299414 228134
rect 298794 192454 299414 227898
rect 298794 192218 298826 192454
rect 299062 192218 299146 192454
rect 299382 192218 299414 192454
rect 298794 192134 299414 192218
rect 298794 191898 298826 192134
rect 299062 191898 299146 192134
rect 299382 191898 299414 192134
rect 298794 156454 299414 191898
rect 298794 156218 298826 156454
rect 299062 156218 299146 156454
rect 299382 156218 299414 156454
rect 298794 156134 299414 156218
rect 298794 155898 298826 156134
rect 299062 155898 299146 156134
rect 299382 155898 299414 156134
rect 298794 120454 299414 155898
rect 298794 120218 298826 120454
rect 299062 120218 299146 120454
rect 299382 120218 299414 120454
rect 298794 120134 299414 120218
rect 298794 119898 298826 120134
rect 299062 119898 299146 120134
rect 299382 119898 299414 120134
rect 298794 84454 299414 119898
rect 298794 84218 298826 84454
rect 299062 84218 299146 84454
rect 299382 84218 299414 84454
rect 298794 84134 299414 84218
rect 298794 83898 298826 84134
rect 299062 83898 299146 84134
rect 299382 83898 299414 84134
rect 298794 48454 299414 83898
rect 298794 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 299414 48454
rect 298794 48134 299414 48218
rect 298794 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 299414 48134
rect 298794 12454 299414 47898
rect 298794 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 299414 12454
rect 298794 12134 299414 12218
rect 298794 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 299414 12134
rect 298794 -2266 299414 11898
rect 298794 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 299414 -2266
rect 298794 -2586 299414 -2502
rect 298794 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 299414 -2586
rect 298794 -7654 299414 -2822
rect 303294 707718 303914 711590
rect 303294 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 303914 707718
rect 303294 707398 303914 707482
rect 303294 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 303914 707398
rect 303294 700954 303914 707162
rect 303294 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 303914 700954
rect 303294 700634 303914 700718
rect 303294 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 303914 700634
rect 303294 664954 303914 700398
rect 303294 664718 303326 664954
rect 303562 664718 303646 664954
rect 303882 664718 303914 664954
rect 303294 664634 303914 664718
rect 303294 664398 303326 664634
rect 303562 664398 303646 664634
rect 303882 664398 303914 664634
rect 303294 628954 303914 664398
rect 303294 628718 303326 628954
rect 303562 628718 303646 628954
rect 303882 628718 303914 628954
rect 303294 628634 303914 628718
rect 303294 628398 303326 628634
rect 303562 628398 303646 628634
rect 303882 628398 303914 628634
rect 303294 592954 303914 628398
rect 303294 592718 303326 592954
rect 303562 592718 303646 592954
rect 303882 592718 303914 592954
rect 303294 592634 303914 592718
rect 303294 592398 303326 592634
rect 303562 592398 303646 592634
rect 303882 592398 303914 592634
rect 303294 556954 303914 592398
rect 303294 556718 303326 556954
rect 303562 556718 303646 556954
rect 303882 556718 303914 556954
rect 303294 556634 303914 556718
rect 303294 556398 303326 556634
rect 303562 556398 303646 556634
rect 303882 556398 303914 556634
rect 303294 520954 303914 556398
rect 303294 520718 303326 520954
rect 303562 520718 303646 520954
rect 303882 520718 303914 520954
rect 303294 520634 303914 520718
rect 303294 520398 303326 520634
rect 303562 520398 303646 520634
rect 303882 520398 303914 520634
rect 303294 484954 303914 520398
rect 303294 484718 303326 484954
rect 303562 484718 303646 484954
rect 303882 484718 303914 484954
rect 303294 484634 303914 484718
rect 303294 484398 303326 484634
rect 303562 484398 303646 484634
rect 303882 484398 303914 484634
rect 303294 448954 303914 484398
rect 303294 448718 303326 448954
rect 303562 448718 303646 448954
rect 303882 448718 303914 448954
rect 303294 448634 303914 448718
rect 303294 448398 303326 448634
rect 303562 448398 303646 448634
rect 303882 448398 303914 448634
rect 303294 412954 303914 448398
rect 303294 412718 303326 412954
rect 303562 412718 303646 412954
rect 303882 412718 303914 412954
rect 303294 412634 303914 412718
rect 303294 412398 303326 412634
rect 303562 412398 303646 412634
rect 303882 412398 303914 412634
rect 303294 376954 303914 412398
rect 303294 376718 303326 376954
rect 303562 376718 303646 376954
rect 303882 376718 303914 376954
rect 303294 376634 303914 376718
rect 303294 376398 303326 376634
rect 303562 376398 303646 376634
rect 303882 376398 303914 376634
rect 303294 340954 303914 376398
rect 303294 340718 303326 340954
rect 303562 340718 303646 340954
rect 303882 340718 303914 340954
rect 303294 340634 303914 340718
rect 303294 340398 303326 340634
rect 303562 340398 303646 340634
rect 303882 340398 303914 340634
rect 303294 304954 303914 340398
rect 303294 304718 303326 304954
rect 303562 304718 303646 304954
rect 303882 304718 303914 304954
rect 303294 304634 303914 304718
rect 303294 304398 303326 304634
rect 303562 304398 303646 304634
rect 303882 304398 303914 304634
rect 303294 268954 303914 304398
rect 303294 268718 303326 268954
rect 303562 268718 303646 268954
rect 303882 268718 303914 268954
rect 303294 268634 303914 268718
rect 303294 268398 303326 268634
rect 303562 268398 303646 268634
rect 303882 268398 303914 268634
rect 303294 232954 303914 268398
rect 303294 232718 303326 232954
rect 303562 232718 303646 232954
rect 303882 232718 303914 232954
rect 303294 232634 303914 232718
rect 303294 232398 303326 232634
rect 303562 232398 303646 232634
rect 303882 232398 303914 232634
rect 303294 196954 303914 232398
rect 303294 196718 303326 196954
rect 303562 196718 303646 196954
rect 303882 196718 303914 196954
rect 303294 196634 303914 196718
rect 303294 196398 303326 196634
rect 303562 196398 303646 196634
rect 303882 196398 303914 196634
rect 303294 160954 303914 196398
rect 303294 160718 303326 160954
rect 303562 160718 303646 160954
rect 303882 160718 303914 160954
rect 303294 160634 303914 160718
rect 303294 160398 303326 160634
rect 303562 160398 303646 160634
rect 303882 160398 303914 160634
rect 303294 124954 303914 160398
rect 303294 124718 303326 124954
rect 303562 124718 303646 124954
rect 303882 124718 303914 124954
rect 303294 124634 303914 124718
rect 303294 124398 303326 124634
rect 303562 124398 303646 124634
rect 303882 124398 303914 124634
rect 303294 88954 303914 124398
rect 303294 88718 303326 88954
rect 303562 88718 303646 88954
rect 303882 88718 303914 88954
rect 303294 88634 303914 88718
rect 303294 88398 303326 88634
rect 303562 88398 303646 88634
rect 303882 88398 303914 88634
rect 303294 52954 303914 88398
rect 303294 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 303914 52954
rect 303294 52634 303914 52718
rect 303294 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 303914 52634
rect 303294 16954 303914 52398
rect 303294 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 303914 16954
rect 303294 16634 303914 16718
rect 303294 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 303914 16634
rect 303294 -3226 303914 16398
rect 303294 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 303914 -3226
rect 303294 -3546 303914 -3462
rect 303294 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 303914 -3546
rect 303294 -7654 303914 -3782
rect 307794 708678 308414 711590
rect 307794 708442 307826 708678
rect 308062 708442 308146 708678
rect 308382 708442 308414 708678
rect 307794 708358 308414 708442
rect 307794 708122 307826 708358
rect 308062 708122 308146 708358
rect 308382 708122 308414 708358
rect 307794 669454 308414 708122
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 525454 308414 560898
rect 307794 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 308414 525454
rect 307794 525134 308414 525218
rect 307794 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 308414 525134
rect 307794 489454 308414 524898
rect 307794 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 308414 489454
rect 307794 489134 308414 489218
rect 307794 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 308414 489134
rect 307794 453454 308414 488898
rect 307794 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 308414 453454
rect 307794 453134 308414 453218
rect 307794 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 308414 453134
rect 307794 417454 308414 452898
rect 307794 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 308414 417454
rect 307794 417134 308414 417218
rect 307794 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 308414 417134
rect 307794 381454 308414 416898
rect 307794 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 308414 381454
rect 307794 381134 308414 381218
rect 307794 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 308414 381134
rect 307794 345454 308414 380898
rect 307794 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 308414 345454
rect 307794 345134 308414 345218
rect 307794 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 308414 345134
rect 307794 309454 308414 344898
rect 307794 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 308414 309454
rect 307794 309134 308414 309218
rect 307794 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 308414 309134
rect 307794 273454 308414 308898
rect 307794 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 308414 273454
rect 307794 273134 308414 273218
rect 307794 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 308414 273134
rect 307794 237454 308414 272898
rect 307794 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 308414 237454
rect 307794 237134 308414 237218
rect 307794 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 308414 237134
rect 307794 201454 308414 236898
rect 307794 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 308414 201454
rect 307794 201134 308414 201218
rect 307794 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 308414 201134
rect 307794 165454 308414 200898
rect 307794 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 308414 165454
rect 307794 165134 308414 165218
rect 307794 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 308414 165134
rect 307794 129454 308414 164898
rect 307794 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 308414 129454
rect 307794 129134 308414 129218
rect 307794 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 308414 129134
rect 307794 93454 308414 128898
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -4186 308414 20898
rect 307794 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 308414 -4186
rect 307794 -4506 308414 -4422
rect 307794 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 308414 -4506
rect 307794 -7654 308414 -4742
rect 312294 709638 312914 711590
rect 312294 709402 312326 709638
rect 312562 709402 312646 709638
rect 312882 709402 312914 709638
rect 312294 709318 312914 709402
rect 312294 709082 312326 709318
rect 312562 709082 312646 709318
rect 312882 709082 312914 709318
rect 312294 673954 312914 709082
rect 312294 673718 312326 673954
rect 312562 673718 312646 673954
rect 312882 673718 312914 673954
rect 312294 673634 312914 673718
rect 312294 673398 312326 673634
rect 312562 673398 312646 673634
rect 312882 673398 312914 673634
rect 312294 637954 312914 673398
rect 312294 637718 312326 637954
rect 312562 637718 312646 637954
rect 312882 637718 312914 637954
rect 312294 637634 312914 637718
rect 312294 637398 312326 637634
rect 312562 637398 312646 637634
rect 312882 637398 312914 637634
rect 312294 601954 312914 637398
rect 312294 601718 312326 601954
rect 312562 601718 312646 601954
rect 312882 601718 312914 601954
rect 312294 601634 312914 601718
rect 312294 601398 312326 601634
rect 312562 601398 312646 601634
rect 312882 601398 312914 601634
rect 312294 565954 312914 601398
rect 312294 565718 312326 565954
rect 312562 565718 312646 565954
rect 312882 565718 312914 565954
rect 312294 565634 312914 565718
rect 312294 565398 312326 565634
rect 312562 565398 312646 565634
rect 312882 565398 312914 565634
rect 312294 529954 312914 565398
rect 312294 529718 312326 529954
rect 312562 529718 312646 529954
rect 312882 529718 312914 529954
rect 312294 529634 312914 529718
rect 312294 529398 312326 529634
rect 312562 529398 312646 529634
rect 312882 529398 312914 529634
rect 312294 493954 312914 529398
rect 312294 493718 312326 493954
rect 312562 493718 312646 493954
rect 312882 493718 312914 493954
rect 312294 493634 312914 493718
rect 312294 493398 312326 493634
rect 312562 493398 312646 493634
rect 312882 493398 312914 493634
rect 312294 457954 312914 493398
rect 312294 457718 312326 457954
rect 312562 457718 312646 457954
rect 312882 457718 312914 457954
rect 312294 457634 312914 457718
rect 312294 457398 312326 457634
rect 312562 457398 312646 457634
rect 312882 457398 312914 457634
rect 312294 421954 312914 457398
rect 312294 421718 312326 421954
rect 312562 421718 312646 421954
rect 312882 421718 312914 421954
rect 312294 421634 312914 421718
rect 312294 421398 312326 421634
rect 312562 421398 312646 421634
rect 312882 421398 312914 421634
rect 312294 385954 312914 421398
rect 312294 385718 312326 385954
rect 312562 385718 312646 385954
rect 312882 385718 312914 385954
rect 312294 385634 312914 385718
rect 312294 385398 312326 385634
rect 312562 385398 312646 385634
rect 312882 385398 312914 385634
rect 312294 349954 312914 385398
rect 312294 349718 312326 349954
rect 312562 349718 312646 349954
rect 312882 349718 312914 349954
rect 312294 349634 312914 349718
rect 312294 349398 312326 349634
rect 312562 349398 312646 349634
rect 312882 349398 312914 349634
rect 312294 313954 312914 349398
rect 312294 313718 312326 313954
rect 312562 313718 312646 313954
rect 312882 313718 312914 313954
rect 312294 313634 312914 313718
rect 312294 313398 312326 313634
rect 312562 313398 312646 313634
rect 312882 313398 312914 313634
rect 312294 277954 312914 313398
rect 312294 277718 312326 277954
rect 312562 277718 312646 277954
rect 312882 277718 312914 277954
rect 312294 277634 312914 277718
rect 312294 277398 312326 277634
rect 312562 277398 312646 277634
rect 312882 277398 312914 277634
rect 312294 241954 312914 277398
rect 312294 241718 312326 241954
rect 312562 241718 312646 241954
rect 312882 241718 312914 241954
rect 312294 241634 312914 241718
rect 312294 241398 312326 241634
rect 312562 241398 312646 241634
rect 312882 241398 312914 241634
rect 312294 205954 312914 241398
rect 312294 205718 312326 205954
rect 312562 205718 312646 205954
rect 312882 205718 312914 205954
rect 312294 205634 312914 205718
rect 312294 205398 312326 205634
rect 312562 205398 312646 205634
rect 312882 205398 312914 205634
rect 312294 169954 312914 205398
rect 312294 169718 312326 169954
rect 312562 169718 312646 169954
rect 312882 169718 312914 169954
rect 312294 169634 312914 169718
rect 312294 169398 312326 169634
rect 312562 169398 312646 169634
rect 312882 169398 312914 169634
rect 312294 133954 312914 169398
rect 312294 133718 312326 133954
rect 312562 133718 312646 133954
rect 312882 133718 312914 133954
rect 312294 133634 312914 133718
rect 312294 133398 312326 133634
rect 312562 133398 312646 133634
rect 312882 133398 312914 133634
rect 312294 97954 312914 133398
rect 312294 97718 312326 97954
rect 312562 97718 312646 97954
rect 312882 97718 312914 97954
rect 312294 97634 312914 97718
rect 312294 97398 312326 97634
rect 312562 97398 312646 97634
rect 312882 97398 312914 97634
rect 312294 61954 312914 97398
rect 312294 61718 312326 61954
rect 312562 61718 312646 61954
rect 312882 61718 312914 61954
rect 312294 61634 312914 61718
rect 312294 61398 312326 61634
rect 312562 61398 312646 61634
rect 312882 61398 312914 61634
rect 312294 25954 312914 61398
rect 312294 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 312914 25954
rect 312294 25634 312914 25718
rect 312294 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 312914 25634
rect 312294 -5146 312914 25398
rect 312294 -5382 312326 -5146
rect 312562 -5382 312646 -5146
rect 312882 -5382 312914 -5146
rect 312294 -5466 312914 -5382
rect 312294 -5702 312326 -5466
rect 312562 -5702 312646 -5466
rect 312882 -5702 312914 -5466
rect 312294 -7654 312914 -5702
rect 316794 710598 317414 711590
rect 316794 710362 316826 710598
rect 317062 710362 317146 710598
rect 317382 710362 317414 710598
rect 316794 710278 317414 710362
rect 316794 710042 316826 710278
rect 317062 710042 317146 710278
rect 317382 710042 317414 710278
rect 316794 678454 317414 710042
rect 316794 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 317414 678454
rect 316794 678134 317414 678218
rect 316794 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 317414 678134
rect 316794 642454 317414 677898
rect 316794 642218 316826 642454
rect 317062 642218 317146 642454
rect 317382 642218 317414 642454
rect 316794 642134 317414 642218
rect 316794 641898 316826 642134
rect 317062 641898 317146 642134
rect 317382 641898 317414 642134
rect 316794 606454 317414 641898
rect 316794 606218 316826 606454
rect 317062 606218 317146 606454
rect 317382 606218 317414 606454
rect 316794 606134 317414 606218
rect 316794 605898 316826 606134
rect 317062 605898 317146 606134
rect 317382 605898 317414 606134
rect 316794 570454 317414 605898
rect 316794 570218 316826 570454
rect 317062 570218 317146 570454
rect 317382 570218 317414 570454
rect 316794 570134 317414 570218
rect 316794 569898 316826 570134
rect 317062 569898 317146 570134
rect 317382 569898 317414 570134
rect 316794 534454 317414 569898
rect 316794 534218 316826 534454
rect 317062 534218 317146 534454
rect 317382 534218 317414 534454
rect 316794 534134 317414 534218
rect 316794 533898 316826 534134
rect 317062 533898 317146 534134
rect 317382 533898 317414 534134
rect 316794 498454 317414 533898
rect 316794 498218 316826 498454
rect 317062 498218 317146 498454
rect 317382 498218 317414 498454
rect 316794 498134 317414 498218
rect 316794 497898 316826 498134
rect 317062 497898 317146 498134
rect 317382 497898 317414 498134
rect 316794 462454 317414 497898
rect 316794 462218 316826 462454
rect 317062 462218 317146 462454
rect 317382 462218 317414 462454
rect 316794 462134 317414 462218
rect 316794 461898 316826 462134
rect 317062 461898 317146 462134
rect 317382 461898 317414 462134
rect 316794 426454 317414 461898
rect 316794 426218 316826 426454
rect 317062 426218 317146 426454
rect 317382 426218 317414 426454
rect 316794 426134 317414 426218
rect 316794 425898 316826 426134
rect 317062 425898 317146 426134
rect 317382 425898 317414 426134
rect 316794 390454 317414 425898
rect 316794 390218 316826 390454
rect 317062 390218 317146 390454
rect 317382 390218 317414 390454
rect 316794 390134 317414 390218
rect 316794 389898 316826 390134
rect 317062 389898 317146 390134
rect 317382 389898 317414 390134
rect 316794 354454 317414 389898
rect 316794 354218 316826 354454
rect 317062 354218 317146 354454
rect 317382 354218 317414 354454
rect 316794 354134 317414 354218
rect 316794 353898 316826 354134
rect 317062 353898 317146 354134
rect 317382 353898 317414 354134
rect 316794 318454 317414 353898
rect 316794 318218 316826 318454
rect 317062 318218 317146 318454
rect 317382 318218 317414 318454
rect 316794 318134 317414 318218
rect 316794 317898 316826 318134
rect 317062 317898 317146 318134
rect 317382 317898 317414 318134
rect 316794 282454 317414 317898
rect 316794 282218 316826 282454
rect 317062 282218 317146 282454
rect 317382 282218 317414 282454
rect 316794 282134 317414 282218
rect 316794 281898 316826 282134
rect 317062 281898 317146 282134
rect 317382 281898 317414 282134
rect 316794 246454 317414 281898
rect 316794 246218 316826 246454
rect 317062 246218 317146 246454
rect 317382 246218 317414 246454
rect 316794 246134 317414 246218
rect 316794 245898 316826 246134
rect 317062 245898 317146 246134
rect 317382 245898 317414 246134
rect 316794 210454 317414 245898
rect 316794 210218 316826 210454
rect 317062 210218 317146 210454
rect 317382 210218 317414 210454
rect 316794 210134 317414 210218
rect 316794 209898 316826 210134
rect 317062 209898 317146 210134
rect 317382 209898 317414 210134
rect 316794 174454 317414 209898
rect 316794 174218 316826 174454
rect 317062 174218 317146 174454
rect 317382 174218 317414 174454
rect 316794 174134 317414 174218
rect 316794 173898 316826 174134
rect 317062 173898 317146 174134
rect 317382 173898 317414 174134
rect 316794 138454 317414 173898
rect 316794 138218 316826 138454
rect 317062 138218 317146 138454
rect 317382 138218 317414 138454
rect 316794 138134 317414 138218
rect 316794 137898 316826 138134
rect 317062 137898 317146 138134
rect 317382 137898 317414 138134
rect 316794 102454 317414 137898
rect 316794 102218 316826 102454
rect 317062 102218 317146 102454
rect 317382 102218 317414 102454
rect 316794 102134 317414 102218
rect 316794 101898 316826 102134
rect 317062 101898 317146 102134
rect 317382 101898 317414 102134
rect 316794 66454 317414 101898
rect 316794 66218 316826 66454
rect 317062 66218 317146 66454
rect 317382 66218 317414 66454
rect 316794 66134 317414 66218
rect 316794 65898 316826 66134
rect 317062 65898 317146 66134
rect 317382 65898 317414 66134
rect 316794 30454 317414 65898
rect 316794 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 317414 30454
rect 316794 30134 317414 30218
rect 316794 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 317414 30134
rect 316794 -6106 317414 29898
rect 316794 -6342 316826 -6106
rect 317062 -6342 317146 -6106
rect 317382 -6342 317414 -6106
rect 316794 -6426 317414 -6342
rect 316794 -6662 316826 -6426
rect 317062 -6662 317146 -6426
rect 317382 -6662 317414 -6426
rect 316794 -7654 317414 -6662
rect 321294 711558 321914 711590
rect 321294 711322 321326 711558
rect 321562 711322 321646 711558
rect 321882 711322 321914 711558
rect 321294 711238 321914 711322
rect 321294 711002 321326 711238
rect 321562 711002 321646 711238
rect 321882 711002 321914 711238
rect 321294 682954 321914 711002
rect 321294 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 321914 682954
rect 321294 682634 321914 682718
rect 321294 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 321914 682634
rect 321294 646954 321914 682398
rect 321294 646718 321326 646954
rect 321562 646718 321646 646954
rect 321882 646718 321914 646954
rect 321294 646634 321914 646718
rect 321294 646398 321326 646634
rect 321562 646398 321646 646634
rect 321882 646398 321914 646634
rect 321294 610954 321914 646398
rect 321294 610718 321326 610954
rect 321562 610718 321646 610954
rect 321882 610718 321914 610954
rect 321294 610634 321914 610718
rect 321294 610398 321326 610634
rect 321562 610398 321646 610634
rect 321882 610398 321914 610634
rect 321294 574954 321914 610398
rect 321294 574718 321326 574954
rect 321562 574718 321646 574954
rect 321882 574718 321914 574954
rect 321294 574634 321914 574718
rect 321294 574398 321326 574634
rect 321562 574398 321646 574634
rect 321882 574398 321914 574634
rect 321294 538954 321914 574398
rect 321294 538718 321326 538954
rect 321562 538718 321646 538954
rect 321882 538718 321914 538954
rect 321294 538634 321914 538718
rect 321294 538398 321326 538634
rect 321562 538398 321646 538634
rect 321882 538398 321914 538634
rect 321294 502954 321914 538398
rect 321294 502718 321326 502954
rect 321562 502718 321646 502954
rect 321882 502718 321914 502954
rect 321294 502634 321914 502718
rect 321294 502398 321326 502634
rect 321562 502398 321646 502634
rect 321882 502398 321914 502634
rect 321294 466954 321914 502398
rect 321294 466718 321326 466954
rect 321562 466718 321646 466954
rect 321882 466718 321914 466954
rect 321294 466634 321914 466718
rect 321294 466398 321326 466634
rect 321562 466398 321646 466634
rect 321882 466398 321914 466634
rect 321294 430954 321914 466398
rect 321294 430718 321326 430954
rect 321562 430718 321646 430954
rect 321882 430718 321914 430954
rect 321294 430634 321914 430718
rect 321294 430398 321326 430634
rect 321562 430398 321646 430634
rect 321882 430398 321914 430634
rect 321294 394954 321914 430398
rect 321294 394718 321326 394954
rect 321562 394718 321646 394954
rect 321882 394718 321914 394954
rect 321294 394634 321914 394718
rect 321294 394398 321326 394634
rect 321562 394398 321646 394634
rect 321882 394398 321914 394634
rect 321294 358954 321914 394398
rect 321294 358718 321326 358954
rect 321562 358718 321646 358954
rect 321882 358718 321914 358954
rect 321294 358634 321914 358718
rect 321294 358398 321326 358634
rect 321562 358398 321646 358634
rect 321882 358398 321914 358634
rect 321294 322954 321914 358398
rect 321294 322718 321326 322954
rect 321562 322718 321646 322954
rect 321882 322718 321914 322954
rect 321294 322634 321914 322718
rect 321294 322398 321326 322634
rect 321562 322398 321646 322634
rect 321882 322398 321914 322634
rect 321294 286954 321914 322398
rect 321294 286718 321326 286954
rect 321562 286718 321646 286954
rect 321882 286718 321914 286954
rect 321294 286634 321914 286718
rect 321294 286398 321326 286634
rect 321562 286398 321646 286634
rect 321882 286398 321914 286634
rect 321294 250954 321914 286398
rect 321294 250718 321326 250954
rect 321562 250718 321646 250954
rect 321882 250718 321914 250954
rect 321294 250634 321914 250718
rect 321294 250398 321326 250634
rect 321562 250398 321646 250634
rect 321882 250398 321914 250634
rect 321294 214954 321914 250398
rect 321294 214718 321326 214954
rect 321562 214718 321646 214954
rect 321882 214718 321914 214954
rect 321294 214634 321914 214718
rect 321294 214398 321326 214634
rect 321562 214398 321646 214634
rect 321882 214398 321914 214634
rect 321294 178954 321914 214398
rect 321294 178718 321326 178954
rect 321562 178718 321646 178954
rect 321882 178718 321914 178954
rect 321294 178634 321914 178718
rect 321294 178398 321326 178634
rect 321562 178398 321646 178634
rect 321882 178398 321914 178634
rect 321294 142954 321914 178398
rect 321294 142718 321326 142954
rect 321562 142718 321646 142954
rect 321882 142718 321914 142954
rect 321294 142634 321914 142718
rect 321294 142398 321326 142634
rect 321562 142398 321646 142634
rect 321882 142398 321914 142634
rect 321294 106954 321914 142398
rect 321294 106718 321326 106954
rect 321562 106718 321646 106954
rect 321882 106718 321914 106954
rect 321294 106634 321914 106718
rect 321294 106398 321326 106634
rect 321562 106398 321646 106634
rect 321882 106398 321914 106634
rect 321294 70954 321914 106398
rect 321294 70718 321326 70954
rect 321562 70718 321646 70954
rect 321882 70718 321914 70954
rect 321294 70634 321914 70718
rect 321294 70398 321326 70634
rect 321562 70398 321646 70634
rect 321882 70398 321914 70634
rect 321294 34954 321914 70398
rect 321294 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 321914 34954
rect 321294 34634 321914 34718
rect 321294 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 321914 34634
rect 321294 -7066 321914 34398
rect 321294 -7302 321326 -7066
rect 321562 -7302 321646 -7066
rect 321882 -7302 321914 -7066
rect 321294 -7386 321914 -7302
rect 321294 -7622 321326 -7386
rect 321562 -7622 321646 -7386
rect 321882 -7622 321914 -7386
rect 321294 -7654 321914 -7622
rect 325794 704838 326414 711590
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 507454 326414 542898
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 325794 435454 326414 470898
rect 325794 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 326414 435454
rect 325794 435134 326414 435218
rect 325794 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 326414 435134
rect 325794 399454 326414 434898
rect 325794 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 326414 399454
rect 325794 399134 326414 399218
rect 325794 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 326414 399134
rect 325794 363454 326414 398898
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 325794 327454 326414 362898
rect 325794 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 326414 327454
rect 325794 327134 326414 327218
rect 325794 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 326414 327134
rect 325794 291454 326414 326898
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 325794 219454 326414 254898
rect 325794 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 326414 219454
rect 325794 219134 326414 219218
rect 325794 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 326414 219134
rect 325794 183454 326414 218898
rect 325794 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 326414 183454
rect 325794 183134 326414 183218
rect 325794 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 326414 183134
rect 325794 147454 326414 182898
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 111454 326414 146898
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -7654 326414 -902
rect 330294 705798 330914 711590
rect 330294 705562 330326 705798
rect 330562 705562 330646 705798
rect 330882 705562 330914 705798
rect 330294 705478 330914 705562
rect 330294 705242 330326 705478
rect 330562 705242 330646 705478
rect 330882 705242 330914 705478
rect 330294 691954 330914 705242
rect 330294 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 330914 691954
rect 330294 691634 330914 691718
rect 330294 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 330914 691634
rect 330294 655954 330914 691398
rect 330294 655718 330326 655954
rect 330562 655718 330646 655954
rect 330882 655718 330914 655954
rect 330294 655634 330914 655718
rect 330294 655398 330326 655634
rect 330562 655398 330646 655634
rect 330882 655398 330914 655634
rect 330294 619954 330914 655398
rect 330294 619718 330326 619954
rect 330562 619718 330646 619954
rect 330882 619718 330914 619954
rect 330294 619634 330914 619718
rect 330294 619398 330326 619634
rect 330562 619398 330646 619634
rect 330882 619398 330914 619634
rect 330294 583954 330914 619398
rect 330294 583718 330326 583954
rect 330562 583718 330646 583954
rect 330882 583718 330914 583954
rect 330294 583634 330914 583718
rect 330294 583398 330326 583634
rect 330562 583398 330646 583634
rect 330882 583398 330914 583634
rect 330294 547954 330914 583398
rect 330294 547718 330326 547954
rect 330562 547718 330646 547954
rect 330882 547718 330914 547954
rect 330294 547634 330914 547718
rect 330294 547398 330326 547634
rect 330562 547398 330646 547634
rect 330882 547398 330914 547634
rect 330294 511954 330914 547398
rect 330294 511718 330326 511954
rect 330562 511718 330646 511954
rect 330882 511718 330914 511954
rect 330294 511634 330914 511718
rect 330294 511398 330326 511634
rect 330562 511398 330646 511634
rect 330882 511398 330914 511634
rect 330294 475954 330914 511398
rect 330294 475718 330326 475954
rect 330562 475718 330646 475954
rect 330882 475718 330914 475954
rect 330294 475634 330914 475718
rect 330294 475398 330326 475634
rect 330562 475398 330646 475634
rect 330882 475398 330914 475634
rect 330294 439954 330914 475398
rect 330294 439718 330326 439954
rect 330562 439718 330646 439954
rect 330882 439718 330914 439954
rect 330294 439634 330914 439718
rect 330294 439398 330326 439634
rect 330562 439398 330646 439634
rect 330882 439398 330914 439634
rect 330294 403954 330914 439398
rect 330294 403718 330326 403954
rect 330562 403718 330646 403954
rect 330882 403718 330914 403954
rect 330294 403634 330914 403718
rect 330294 403398 330326 403634
rect 330562 403398 330646 403634
rect 330882 403398 330914 403634
rect 330294 367954 330914 403398
rect 330294 367718 330326 367954
rect 330562 367718 330646 367954
rect 330882 367718 330914 367954
rect 330294 367634 330914 367718
rect 330294 367398 330326 367634
rect 330562 367398 330646 367634
rect 330882 367398 330914 367634
rect 330294 331954 330914 367398
rect 330294 331718 330326 331954
rect 330562 331718 330646 331954
rect 330882 331718 330914 331954
rect 330294 331634 330914 331718
rect 330294 331398 330326 331634
rect 330562 331398 330646 331634
rect 330882 331398 330914 331634
rect 330294 295954 330914 331398
rect 330294 295718 330326 295954
rect 330562 295718 330646 295954
rect 330882 295718 330914 295954
rect 330294 295634 330914 295718
rect 330294 295398 330326 295634
rect 330562 295398 330646 295634
rect 330882 295398 330914 295634
rect 330294 259954 330914 295398
rect 330294 259718 330326 259954
rect 330562 259718 330646 259954
rect 330882 259718 330914 259954
rect 330294 259634 330914 259718
rect 330294 259398 330326 259634
rect 330562 259398 330646 259634
rect 330882 259398 330914 259634
rect 330294 223954 330914 259398
rect 330294 223718 330326 223954
rect 330562 223718 330646 223954
rect 330882 223718 330914 223954
rect 330294 223634 330914 223718
rect 330294 223398 330326 223634
rect 330562 223398 330646 223634
rect 330882 223398 330914 223634
rect 330294 187954 330914 223398
rect 330294 187718 330326 187954
rect 330562 187718 330646 187954
rect 330882 187718 330914 187954
rect 330294 187634 330914 187718
rect 330294 187398 330326 187634
rect 330562 187398 330646 187634
rect 330882 187398 330914 187634
rect 330294 151954 330914 187398
rect 330294 151718 330326 151954
rect 330562 151718 330646 151954
rect 330882 151718 330914 151954
rect 330294 151634 330914 151718
rect 330294 151398 330326 151634
rect 330562 151398 330646 151634
rect 330882 151398 330914 151634
rect 330294 115954 330914 151398
rect 330294 115718 330326 115954
rect 330562 115718 330646 115954
rect 330882 115718 330914 115954
rect 330294 115634 330914 115718
rect 330294 115398 330326 115634
rect 330562 115398 330646 115634
rect 330882 115398 330914 115634
rect 330294 79954 330914 115398
rect 330294 79718 330326 79954
rect 330562 79718 330646 79954
rect 330882 79718 330914 79954
rect 330294 79634 330914 79718
rect 330294 79398 330326 79634
rect 330562 79398 330646 79634
rect 330882 79398 330914 79634
rect 330294 43954 330914 79398
rect 330294 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 330914 43954
rect 330294 43634 330914 43718
rect 330294 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 330914 43634
rect 330294 7954 330914 43398
rect 330294 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 330914 7954
rect 330294 7634 330914 7718
rect 330294 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 330914 7634
rect 330294 -1306 330914 7398
rect 330294 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 330914 -1306
rect 330294 -1626 330914 -1542
rect 330294 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 330914 -1626
rect 330294 -7654 330914 -1862
rect 334794 706758 335414 711590
rect 334794 706522 334826 706758
rect 335062 706522 335146 706758
rect 335382 706522 335414 706758
rect 334794 706438 335414 706522
rect 334794 706202 334826 706438
rect 335062 706202 335146 706438
rect 335382 706202 335414 706438
rect 334794 696454 335414 706202
rect 334794 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 335414 696454
rect 334794 696134 335414 696218
rect 334794 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 335414 696134
rect 334794 660454 335414 695898
rect 334794 660218 334826 660454
rect 335062 660218 335146 660454
rect 335382 660218 335414 660454
rect 334794 660134 335414 660218
rect 334794 659898 334826 660134
rect 335062 659898 335146 660134
rect 335382 659898 335414 660134
rect 334794 624454 335414 659898
rect 334794 624218 334826 624454
rect 335062 624218 335146 624454
rect 335382 624218 335414 624454
rect 334794 624134 335414 624218
rect 334794 623898 334826 624134
rect 335062 623898 335146 624134
rect 335382 623898 335414 624134
rect 334794 588454 335414 623898
rect 334794 588218 334826 588454
rect 335062 588218 335146 588454
rect 335382 588218 335414 588454
rect 334794 588134 335414 588218
rect 334794 587898 334826 588134
rect 335062 587898 335146 588134
rect 335382 587898 335414 588134
rect 334794 552454 335414 587898
rect 334794 552218 334826 552454
rect 335062 552218 335146 552454
rect 335382 552218 335414 552454
rect 334794 552134 335414 552218
rect 334794 551898 334826 552134
rect 335062 551898 335146 552134
rect 335382 551898 335414 552134
rect 334794 516454 335414 551898
rect 334794 516218 334826 516454
rect 335062 516218 335146 516454
rect 335382 516218 335414 516454
rect 334794 516134 335414 516218
rect 334794 515898 334826 516134
rect 335062 515898 335146 516134
rect 335382 515898 335414 516134
rect 334794 480454 335414 515898
rect 334794 480218 334826 480454
rect 335062 480218 335146 480454
rect 335382 480218 335414 480454
rect 334794 480134 335414 480218
rect 334794 479898 334826 480134
rect 335062 479898 335146 480134
rect 335382 479898 335414 480134
rect 334794 444454 335414 479898
rect 334794 444218 334826 444454
rect 335062 444218 335146 444454
rect 335382 444218 335414 444454
rect 334794 444134 335414 444218
rect 334794 443898 334826 444134
rect 335062 443898 335146 444134
rect 335382 443898 335414 444134
rect 334794 408454 335414 443898
rect 334794 408218 334826 408454
rect 335062 408218 335146 408454
rect 335382 408218 335414 408454
rect 334794 408134 335414 408218
rect 334794 407898 334826 408134
rect 335062 407898 335146 408134
rect 335382 407898 335414 408134
rect 334794 372454 335414 407898
rect 334794 372218 334826 372454
rect 335062 372218 335146 372454
rect 335382 372218 335414 372454
rect 334794 372134 335414 372218
rect 334794 371898 334826 372134
rect 335062 371898 335146 372134
rect 335382 371898 335414 372134
rect 334794 336454 335414 371898
rect 334794 336218 334826 336454
rect 335062 336218 335146 336454
rect 335382 336218 335414 336454
rect 334794 336134 335414 336218
rect 334794 335898 334826 336134
rect 335062 335898 335146 336134
rect 335382 335898 335414 336134
rect 334794 300454 335414 335898
rect 334794 300218 334826 300454
rect 335062 300218 335146 300454
rect 335382 300218 335414 300454
rect 334794 300134 335414 300218
rect 334794 299898 334826 300134
rect 335062 299898 335146 300134
rect 335382 299898 335414 300134
rect 334794 264454 335414 299898
rect 334794 264218 334826 264454
rect 335062 264218 335146 264454
rect 335382 264218 335414 264454
rect 334794 264134 335414 264218
rect 334794 263898 334826 264134
rect 335062 263898 335146 264134
rect 335382 263898 335414 264134
rect 334794 228454 335414 263898
rect 334794 228218 334826 228454
rect 335062 228218 335146 228454
rect 335382 228218 335414 228454
rect 334794 228134 335414 228218
rect 334794 227898 334826 228134
rect 335062 227898 335146 228134
rect 335382 227898 335414 228134
rect 334794 192454 335414 227898
rect 334794 192218 334826 192454
rect 335062 192218 335146 192454
rect 335382 192218 335414 192454
rect 334794 192134 335414 192218
rect 334794 191898 334826 192134
rect 335062 191898 335146 192134
rect 335382 191898 335414 192134
rect 334794 156454 335414 191898
rect 334794 156218 334826 156454
rect 335062 156218 335146 156454
rect 335382 156218 335414 156454
rect 334794 156134 335414 156218
rect 334794 155898 334826 156134
rect 335062 155898 335146 156134
rect 335382 155898 335414 156134
rect 334794 120454 335414 155898
rect 334794 120218 334826 120454
rect 335062 120218 335146 120454
rect 335382 120218 335414 120454
rect 334794 120134 335414 120218
rect 334794 119898 334826 120134
rect 335062 119898 335146 120134
rect 335382 119898 335414 120134
rect 334794 84454 335414 119898
rect 334794 84218 334826 84454
rect 335062 84218 335146 84454
rect 335382 84218 335414 84454
rect 334794 84134 335414 84218
rect 334794 83898 334826 84134
rect 335062 83898 335146 84134
rect 335382 83898 335414 84134
rect 334794 48454 335414 83898
rect 334794 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 335414 48454
rect 334794 48134 335414 48218
rect 334794 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 335414 48134
rect 334794 12454 335414 47898
rect 334794 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 335414 12454
rect 334794 12134 335414 12218
rect 334794 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 335414 12134
rect 334794 -2266 335414 11898
rect 334794 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 335414 -2266
rect 334794 -2586 335414 -2502
rect 334794 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 335414 -2586
rect 334794 -7654 335414 -2822
rect 339294 707718 339914 711590
rect 339294 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 339914 707718
rect 339294 707398 339914 707482
rect 339294 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 339914 707398
rect 339294 700954 339914 707162
rect 339294 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 339914 700954
rect 339294 700634 339914 700718
rect 339294 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 339914 700634
rect 339294 664954 339914 700398
rect 339294 664718 339326 664954
rect 339562 664718 339646 664954
rect 339882 664718 339914 664954
rect 339294 664634 339914 664718
rect 339294 664398 339326 664634
rect 339562 664398 339646 664634
rect 339882 664398 339914 664634
rect 339294 628954 339914 664398
rect 339294 628718 339326 628954
rect 339562 628718 339646 628954
rect 339882 628718 339914 628954
rect 339294 628634 339914 628718
rect 339294 628398 339326 628634
rect 339562 628398 339646 628634
rect 339882 628398 339914 628634
rect 339294 592954 339914 628398
rect 339294 592718 339326 592954
rect 339562 592718 339646 592954
rect 339882 592718 339914 592954
rect 339294 592634 339914 592718
rect 339294 592398 339326 592634
rect 339562 592398 339646 592634
rect 339882 592398 339914 592634
rect 339294 556954 339914 592398
rect 339294 556718 339326 556954
rect 339562 556718 339646 556954
rect 339882 556718 339914 556954
rect 339294 556634 339914 556718
rect 339294 556398 339326 556634
rect 339562 556398 339646 556634
rect 339882 556398 339914 556634
rect 339294 520954 339914 556398
rect 339294 520718 339326 520954
rect 339562 520718 339646 520954
rect 339882 520718 339914 520954
rect 339294 520634 339914 520718
rect 339294 520398 339326 520634
rect 339562 520398 339646 520634
rect 339882 520398 339914 520634
rect 339294 484954 339914 520398
rect 339294 484718 339326 484954
rect 339562 484718 339646 484954
rect 339882 484718 339914 484954
rect 339294 484634 339914 484718
rect 339294 484398 339326 484634
rect 339562 484398 339646 484634
rect 339882 484398 339914 484634
rect 339294 448954 339914 484398
rect 339294 448718 339326 448954
rect 339562 448718 339646 448954
rect 339882 448718 339914 448954
rect 339294 448634 339914 448718
rect 339294 448398 339326 448634
rect 339562 448398 339646 448634
rect 339882 448398 339914 448634
rect 339294 412954 339914 448398
rect 339294 412718 339326 412954
rect 339562 412718 339646 412954
rect 339882 412718 339914 412954
rect 339294 412634 339914 412718
rect 339294 412398 339326 412634
rect 339562 412398 339646 412634
rect 339882 412398 339914 412634
rect 339294 376954 339914 412398
rect 339294 376718 339326 376954
rect 339562 376718 339646 376954
rect 339882 376718 339914 376954
rect 339294 376634 339914 376718
rect 339294 376398 339326 376634
rect 339562 376398 339646 376634
rect 339882 376398 339914 376634
rect 339294 340954 339914 376398
rect 339294 340718 339326 340954
rect 339562 340718 339646 340954
rect 339882 340718 339914 340954
rect 339294 340634 339914 340718
rect 339294 340398 339326 340634
rect 339562 340398 339646 340634
rect 339882 340398 339914 340634
rect 339294 304954 339914 340398
rect 339294 304718 339326 304954
rect 339562 304718 339646 304954
rect 339882 304718 339914 304954
rect 339294 304634 339914 304718
rect 339294 304398 339326 304634
rect 339562 304398 339646 304634
rect 339882 304398 339914 304634
rect 339294 268954 339914 304398
rect 339294 268718 339326 268954
rect 339562 268718 339646 268954
rect 339882 268718 339914 268954
rect 339294 268634 339914 268718
rect 339294 268398 339326 268634
rect 339562 268398 339646 268634
rect 339882 268398 339914 268634
rect 339294 232954 339914 268398
rect 339294 232718 339326 232954
rect 339562 232718 339646 232954
rect 339882 232718 339914 232954
rect 339294 232634 339914 232718
rect 339294 232398 339326 232634
rect 339562 232398 339646 232634
rect 339882 232398 339914 232634
rect 339294 196954 339914 232398
rect 339294 196718 339326 196954
rect 339562 196718 339646 196954
rect 339882 196718 339914 196954
rect 339294 196634 339914 196718
rect 339294 196398 339326 196634
rect 339562 196398 339646 196634
rect 339882 196398 339914 196634
rect 339294 160954 339914 196398
rect 339294 160718 339326 160954
rect 339562 160718 339646 160954
rect 339882 160718 339914 160954
rect 339294 160634 339914 160718
rect 339294 160398 339326 160634
rect 339562 160398 339646 160634
rect 339882 160398 339914 160634
rect 339294 124954 339914 160398
rect 339294 124718 339326 124954
rect 339562 124718 339646 124954
rect 339882 124718 339914 124954
rect 339294 124634 339914 124718
rect 339294 124398 339326 124634
rect 339562 124398 339646 124634
rect 339882 124398 339914 124634
rect 339294 88954 339914 124398
rect 339294 88718 339326 88954
rect 339562 88718 339646 88954
rect 339882 88718 339914 88954
rect 339294 88634 339914 88718
rect 339294 88398 339326 88634
rect 339562 88398 339646 88634
rect 339882 88398 339914 88634
rect 339294 52954 339914 88398
rect 339294 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 339914 52954
rect 339294 52634 339914 52718
rect 339294 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 339914 52634
rect 339294 16954 339914 52398
rect 339294 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 339914 16954
rect 339294 16634 339914 16718
rect 339294 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 339914 16634
rect 339294 -3226 339914 16398
rect 339294 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 339914 -3226
rect 339294 -3546 339914 -3462
rect 339294 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 339914 -3546
rect 339294 -7654 339914 -3782
rect 343794 708678 344414 711590
rect 343794 708442 343826 708678
rect 344062 708442 344146 708678
rect 344382 708442 344414 708678
rect 343794 708358 344414 708442
rect 343794 708122 343826 708358
rect 344062 708122 344146 708358
rect 344382 708122 344414 708358
rect 343794 669454 344414 708122
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561454 344414 596898
rect 343794 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 344414 561454
rect 343794 561134 344414 561218
rect 343794 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 344414 561134
rect 343794 525454 344414 560898
rect 343794 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 344414 525454
rect 343794 525134 344414 525218
rect 343794 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 344414 525134
rect 343794 489454 344414 524898
rect 343794 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 344414 489454
rect 343794 489134 344414 489218
rect 343794 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 344414 489134
rect 343794 453454 344414 488898
rect 343794 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 344414 453454
rect 343794 453134 344414 453218
rect 343794 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 344414 453134
rect 343794 417454 344414 452898
rect 343794 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 344414 417454
rect 343794 417134 344414 417218
rect 343794 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 344414 417134
rect 343794 381454 344414 416898
rect 343794 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 344414 381454
rect 343794 381134 344414 381218
rect 343794 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 344414 381134
rect 343794 345454 344414 380898
rect 343794 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 344414 345454
rect 343794 345134 344414 345218
rect 343794 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 344414 345134
rect 343794 309454 344414 344898
rect 343794 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 344414 309454
rect 343794 309134 344414 309218
rect 343794 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 344414 309134
rect 343794 273454 344414 308898
rect 343794 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 344414 273454
rect 343794 273134 344414 273218
rect 343794 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 344414 273134
rect 343794 237454 344414 272898
rect 343794 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 344414 237454
rect 343794 237134 344414 237218
rect 343794 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 344414 237134
rect 343794 201454 344414 236898
rect 343794 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 344414 201454
rect 343794 201134 344414 201218
rect 343794 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 344414 201134
rect 343794 165454 344414 200898
rect 343794 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 344414 165454
rect 343794 165134 344414 165218
rect 343794 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 344414 165134
rect 343794 129454 344414 164898
rect 343794 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 344414 129454
rect 343794 129134 344414 129218
rect 343794 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 344414 129134
rect 343794 93454 344414 128898
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -4186 344414 20898
rect 343794 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 344414 -4186
rect 343794 -4506 344414 -4422
rect 343794 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 344414 -4506
rect 343794 -7654 344414 -4742
rect 348294 709638 348914 711590
rect 348294 709402 348326 709638
rect 348562 709402 348646 709638
rect 348882 709402 348914 709638
rect 348294 709318 348914 709402
rect 348294 709082 348326 709318
rect 348562 709082 348646 709318
rect 348882 709082 348914 709318
rect 348294 673954 348914 709082
rect 348294 673718 348326 673954
rect 348562 673718 348646 673954
rect 348882 673718 348914 673954
rect 348294 673634 348914 673718
rect 348294 673398 348326 673634
rect 348562 673398 348646 673634
rect 348882 673398 348914 673634
rect 348294 637954 348914 673398
rect 348294 637718 348326 637954
rect 348562 637718 348646 637954
rect 348882 637718 348914 637954
rect 348294 637634 348914 637718
rect 348294 637398 348326 637634
rect 348562 637398 348646 637634
rect 348882 637398 348914 637634
rect 348294 601954 348914 637398
rect 348294 601718 348326 601954
rect 348562 601718 348646 601954
rect 348882 601718 348914 601954
rect 348294 601634 348914 601718
rect 348294 601398 348326 601634
rect 348562 601398 348646 601634
rect 348882 601398 348914 601634
rect 348294 565954 348914 601398
rect 348294 565718 348326 565954
rect 348562 565718 348646 565954
rect 348882 565718 348914 565954
rect 348294 565634 348914 565718
rect 348294 565398 348326 565634
rect 348562 565398 348646 565634
rect 348882 565398 348914 565634
rect 348294 529954 348914 565398
rect 348294 529718 348326 529954
rect 348562 529718 348646 529954
rect 348882 529718 348914 529954
rect 348294 529634 348914 529718
rect 348294 529398 348326 529634
rect 348562 529398 348646 529634
rect 348882 529398 348914 529634
rect 348294 493954 348914 529398
rect 348294 493718 348326 493954
rect 348562 493718 348646 493954
rect 348882 493718 348914 493954
rect 348294 493634 348914 493718
rect 348294 493398 348326 493634
rect 348562 493398 348646 493634
rect 348882 493398 348914 493634
rect 348294 457954 348914 493398
rect 348294 457718 348326 457954
rect 348562 457718 348646 457954
rect 348882 457718 348914 457954
rect 348294 457634 348914 457718
rect 348294 457398 348326 457634
rect 348562 457398 348646 457634
rect 348882 457398 348914 457634
rect 348294 421954 348914 457398
rect 348294 421718 348326 421954
rect 348562 421718 348646 421954
rect 348882 421718 348914 421954
rect 348294 421634 348914 421718
rect 348294 421398 348326 421634
rect 348562 421398 348646 421634
rect 348882 421398 348914 421634
rect 348294 385954 348914 421398
rect 348294 385718 348326 385954
rect 348562 385718 348646 385954
rect 348882 385718 348914 385954
rect 348294 385634 348914 385718
rect 348294 385398 348326 385634
rect 348562 385398 348646 385634
rect 348882 385398 348914 385634
rect 348294 349954 348914 385398
rect 348294 349718 348326 349954
rect 348562 349718 348646 349954
rect 348882 349718 348914 349954
rect 348294 349634 348914 349718
rect 348294 349398 348326 349634
rect 348562 349398 348646 349634
rect 348882 349398 348914 349634
rect 348294 313954 348914 349398
rect 348294 313718 348326 313954
rect 348562 313718 348646 313954
rect 348882 313718 348914 313954
rect 348294 313634 348914 313718
rect 348294 313398 348326 313634
rect 348562 313398 348646 313634
rect 348882 313398 348914 313634
rect 348294 277954 348914 313398
rect 348294 277718 348326 277954
rect 348562 277718 348646 277954
rect 348882 277718 348914 277954
rect 348294 277634 348914 277718
rect 348294 277398 348326 277634
rect 348562 277398 348646 277634
rect 348882 277398 348914 277634
rect 348294 241954 348914 277398
rect 348294 241718 348326 241954
rect 348562 241718 348646 241954
rect 348882 241718 348914 241954
rect 348294 241634 348914 241718
rect 348294 241398 348326 241634
rect 348562 241398 348646 241634
rect 348882 241398 348914 241634
rect 348294 205954 348914 241398
rect 348294 205718 348326 205954
rect 348562 205718 348646 205954
rect 348882 205718 348914 205954
rect 348294 205634 348914 205718
rect 348294 205398 348326 205634
rect 348562 205398 348646 205634
rect 348882 205398 348914 205634
rect 348294 169954 348914 205398
rect 348294 169718 348326 169954
rect 348562 169718 348646 169954
rect 348882 169718 348914 169954
rect 348294 169634 348914 169718
rect 348294 169398 348326 169634
rect 348562 169398 348646 169634
rect 348882 169398 348914 169634
rect 348294 133954 348914 169398
rect 348294 133718 348326 133954
rect 348562 133718 348646 133954
rect 348882 133718 348914 133954
rect 348294 133634 348914 133718
rect 348294 133398 348326 133634
rect 348562 133398 348646 133634
rect 348882 133398 348914 133634
rect 348294 97954 348914 133398
rect 348294 97718 348326 97954
rect 348562 97718 348646 97954
rect 348882 97718 348914 97954
rect 348294 97634 348914 97718
rect 348294 97398 348326 97634
rect 348562 97398 348646 97634
rect 348882 97398 348914 97634
rect 348294 61954 348914 97398
rect 348294 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 348914 61954
rect 348294 61634 348914 61718
rect 348294 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 348914 61634
rect 348294 25954 348914 61398
rect 348294 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 348914 25954
rect 348294 25634 348914 25718
rect 348294 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 348914 25634
rect 348294 -5146 348914 25398
rect 348294 -5382 348326 -5146
rect 348562 -5382 348646 -5146
rect 348882 -5382 348914 -5146
rect 348294 -5466 348914 -5382
rect 348294 -5702 348326 -5466
rect 348562 -5702 348646 -5466
rect 348882 -5702 348914 -5466
rect 348294 -7654 348914 -5702
rect 352794 710598 353414 711590
rect 352794 710362 352826 710598
rect 353062 710362 353146 710598
rect 353382 710362 353414 710598
rect 352794 710278 353414 710362
rect 352794 710042 352826 710278
rect 353062 710042 353146 710278
rect 353382 710042 353414 710278
rect 352794 678454 353414 710042
rect 352794 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 353414 678454
rect 352794 678134 353414 678218
rect 352794 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 353414 678134
rect 352794 642454 353414 677898
rect 352794 642218 352826 642454
rect 353062 642218 353146 642454
rect 353382 642218 353414 642454
rect 352794 642134 353414 642218
rect 352794 641898 352826 642134
rect 353062 641898 353146 642134
rect 353382 641898 353414 642134
rect 352794 606454 353414 641898
rect 352794 606218 352826 606454
rect 353062 606218 353146 606454
rect 353382 606218 353414 606454
rect 352794 606134 353414 606218
rect 352794 605898 352826 606134
rect 353062 605898 353146 606134
rect 353382 605898 353414 606134
rect 352794 570454 353414 605898
rect 352794 570218 352826 570454
rect 353062 570218 353146 570454
rect 353382 570218 353414 570454
rect 352794 570134 353414 570218
rect 352794 569898 352826 570134
rect 353062 569898 353146 570134
rect 353382 569898 353414 570134
rect 352794 534454 353414 569898
rect 352794 534218 352826 534454
rect 353062 534218 353146 534454
rect 353382 534218 353414 534454
rect 352794 534134 353414 534218
rect 352794 533898 352826 534134
rect 353062 533898 353146 534134
rect 353382 533898 353414 534134
rect 352794 498454 353414 533898
rect 352794 498218 352826 498454
rect 353062 498218 353146 498454
rect 353382 498218 353414 498454
rect 352794 498134 353414 498218
rect 352794 497898 352826 498134
rect 353062 497898 353146 498134
rect 353382 497898 353414 498134
rect 352794 462454 353414 497898
rect 352794 462218 352826 462454
rect 353062 462218 353146 462454
rect 353382 462218 353414 462454
rect 352794 462134 353414 462218
rect 352794 461898 352826 462134
rect 353062 461898 353146 462134
rect 353382 461898 353414 462134
rect 352794 426454 353414 461898
rect 352794 426218 352826 426454
rect 353062 426218 353146 426454
rect 353382 426218 353414 426454
rect 352794 426134 353414 426218
rect 352794 425898 352826 426134
rect 353062 425898 353146 426134
rect 353382 425898 353414 426134
rect 352794 390454 353414 425898
rect 352794 390218 352826 390454
rect 353062 390218 353146 390454
rect 353382 390218 353414 390454
rect 352794 390134 353414 390218
rect 352794 389898 352826 390134
rect 353062 389898 353146 390134
rect 353382 389898 353414 390134
rect 352794 354454 353414 389898
rect 352794 354218 352826 354454
rect 353062 354218 353146 354454
rect 353382 354218 353414 354454
rect 352794 354134 353414 354218
rect 352794 353898 352826 354134
rect 353062 353898 353146 354134
rect 353382 353898 353414 354134
rect 352794 318454 353414 353898
rect 352794 318218 352826 318454
rect 353062 318218 353146 318454
rect 353382 318218 353414 318454
rect 352794 318134 353414 318218
rect 352794 317898 352826 318134
rect 353062 317898 353146 318134
rect 353382 317898 353414 318134
rect 352794 282454 353414 317898
rect 352794 282218 352826 282454
rect 353062 282218 353146 282454
rect 353382 282218 353414 282454
rect 352794 282134 353414 282218
rect 352794 281898 352826 282134
rect 353062 281898 353146 282134
rect 353382 281898 353414 282134
rect 352794 246454 353414 281898
rect 352794 246218 352826 246454
rect 353062 246218 353146 246454
rect 353382 246218 353414 246454
rect 352794 246134 353414 246218
rect 352794 245898 352826 246134
rect 353062 245898 353146 246134
rect 353382 245898 353414 246134
rect 352794 210454 353414 245898
rect 352794 210218 352826 210454
rect 353062 210218 353146 210454
rect 353382 210218 353414 210454
rect 352794 210134 353414 210218
rect 352794 209898 352826 210134
rect 353062 209898 353146 210134
rect 353382 209898 353414 210134
rect 352794 174454 353414 209898
rect 352794 174218 352826 174454
rect 353062 174218 353146 174454
rect 353382 174218 353414 174454
rect 352794 174134 353414 174218
rect 352794 173898 352826 174134
rect 353062 173898 353146 174134
rect 353382 173898 353414 174134
rect 352794 138454 353414 173898
rect 352794 138218 352826 138454
rect 353062 138218 353146 138454
rect 353382 138218 353414 138454
rect 352794 138134 353414 138218
rect 352794 137898 352826 138134
rect 353062 137898 353146 138134
rect 353382 137898 353414 138134
rect 352794 102454 353414 137898
rect 352794 102218 352826 102454
rect 353062 102218 353146 102454
rect 353382 102218 353414 102454
rect 352794 102134 353414 102218
rect 352794 101898 352826 102134
rect 353062 101898 353146 102134
rect 353382 101898 353414 102134
rect 352794 66454 353414 101898
rect 352794 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 353414 66454
rect 352794 66134 353414 66218
rect 352794 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 353414 66134
rect 352794 30454 353414 65898
rect 352794 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 353414 30454
rect 352794 30134 353414 30218
rect 352794 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 353414 30134
rect 352794 -6106 353414 29898
rect 352794 -6342 352826 -6106
rect 353062 -6342 353146 -6106
rect 353382 -6342 353414 -6106
rect 352794 -6426 353414 -6342
rect 352794 -6662 352826 -6426
rect 353062 -6662 353146 -6426
rect 353382 -6662 353414 -6426
rect 352794 -7654 353414 -6662
rect 357294 711558 357914 711590
rect 357294 711322 357326 711558
rect 357562 711322 357646 711558
rect 357882 711322 357914 711558
rect 357294 711238 357914 711322
rect 357294 711002 357326 711238
rect 357562 711002 357646 711238
rect 357882 711002 357914 711238
rect 357294 682954 357914 711002
rect 357294 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 357914 682954
rect 357294 682634 357914 682718
rect 357294 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 357914 682634
rect 357294 646954 357914 682398
rect 357294 646718 357326 646954
rect 357562 646718 357646 646954
rect 357882 646718 357914 646954
rect 357294 646634 357914 646718
rect 357294 646398 357326 646634
rect 357562 646398 357646 646634
rect 357882 646398 357914 646634
rect 357294 610954 357914 646398
rect 357294 610718 357326 610954
rect 357562 610718 357646 610954
rect 357882 610718 357914 610954
rect 357294 610634 357914 610718
rect 357294 610398 357326 610634
rect 357562 610398 357646 610634
rect 357882 610398 357914 610634
rect 357294 574954 357914 610398
rect 357294 574718 357326 574954
rect 357562 574718 357646 574954
rect 357882 574718 357914 574954
rect 357294 574634 357914 574718
rect 357294 574398 357326 574634
rect 357562 574398 357646 574634
rect 357882 574398 357914 574634
rect 357294 538954 357914 574398
rect 357294 538718 357326 538954
rect 357562 538718 357646 538954
rect 357882 538718 357914 538954
rect 357294 538634 357914 538718
rect 357294 538398 357326 538634
rect 357562 538398 357646 538634
rect 357882 538398 357914 538634
rect 357294 502954 357914 538398
rect 357294 502718 357326 502954
rect 357562 502718 357646 502954
rect 357882 502718 357914 502954
rect 357294 502634 357914 502718
rect 357294 502398 357326 502634
rect 357562 502398 357646 502634
rect 357882 502398 357914 502634
rect 357294 466954 357914 502398
rect 357294 466718 357326 466954
rect 357562 466718 357646 466954
rect 357882 466718 357914 466954
rect 357294 466634 357914 466718
rect 357294 466398 357326 466634
rect 357562 466398 357646 466634
rect 357882 466398 357914 466634
rect 357294 430954 357914 466398
rect 357294 430718 357326 430954
rect 357562 430718 357646 430954
rect 357882 430718 357914 430954
rect 357294 430634 357914 430718
rect 357294 430398 357326 430634
rect 357562 430398 357646 430634
rect 357882 430398 357914 430634
rect 357294 394954 357914 430398
rect 357294 394718 357326 394954
rect 357562 394718 357646 394954
rect 357882 394718 357914 394954
rect 357294 394634 357914 394718
rect 357294 394398 357326 394634
rect 357562 394398 357646 394634
rect 357882 394398 357914 394634
rect 357294 358954 357914 394398
rect 357294 358718 357326 358954
rect 357562 358718 357646 358954
rect 357882 358718 357914 358954
rect 357294 358634 357914 358718
rect 357294 358398 357326 358634
rect 357562 358398 357646 358634
rect 357882 358398 357914 358634
rect 357294 322954 357914 358398
rect 357294 322718 357326 322954
rect 357562 322718 357646 322954
rect 357882 322718 357914 322954
rect 357294 322634 357914 322718
rect 357294 322398 357326 322634
rect 357562 322398 357646 322634
rect 357882 322398 357914 322634
rect 357294 286954 357914 322398
rect 357294 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 357914 286954
rect 357294 286634 357914 286718
rect 357294 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 357914 286634
rect 357294 250954 357914 286398
rect 357294 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 357914 250954
rect 357294 250634 357914 250718
rect 357294 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 357914 250634
rect 357294 214954 357914 250398
rect 357294 214718 357326 214954
rect 357562 214718 357646 214954
rect 357882 214718 357914 214954
rect 357294 214634 357914 214718
rect 357294 214398 357326 214634
rect 357562 214398 357646 214634
rect 357882 214398 357914 214634
rect 357294 178954 357914 214398
rect 357294 178718 357326 178954
rect 357562 178718 357646 178954
rect 357882 178718 357914 178954
rect 357294 178634 357914 178718
rect 357294 178398 357326 178634
rect 357562 178398 357646 178634
rect 357882 178398 357914 178634
rect 357294 142954 357914 178398
rect 357294 142718 357326 142954
rect 357562 142718 357646 142954
rect 357882 142718 357914 142954
rect 357294 142634 357914 142718
rect 357294 142398 357326 142634
rect 357562 142398 357646 142634
rect 357882 142398 357914 142634
rect 357294 106954 357914 142398
rect 357294 106718 357326 106954
rect 357562 106718 357646 106954
rect 357882 106718 357914 106954
rect 357294 106634 357914 106718
rect 357294 106398 357326 106634
rect 357562 106398 357646 106634
rect 357882 106398 357914 106634
rect 357294 70954 357914 106398
rect 357294 70718 357326 70954
rect 357562 70718 357646 70954
rect 357882 70718 357914 70954
rect 357294 70634 357914 70718
rect 357294 70398 357326 70634
rect 357562 70398 357646 70634
rect 357882 70398 357914 70634
rect 357294 34954 357914 70398
rect 357294 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 357914 34954
rect 357294 34634 357914 34718
rect 357294 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 357914 34634
rect 357294 -7066 357914 34398
rect 357294 -7302 357326 -7066
rect 357562 -7302 357646 -7066
rect 357882 -7302 357914 -7066
rect 357294 -7386 357914 -7302
rect 357294 -7622 357326 -7386
rect 357562 -7622 357646 -7386
rect 357882 -7622 357914 -7386
rect 357294 -7654 357914 -7622
rect 361794 704838 362414 711590
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 361794 363454 362414 398898
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -7654 362414 -902
rect 366294 705798 366914 711590
rect 366294 705562 366326 705798
rect 366562 705562 366646 705798
rect 366882 705562 366914 705798
rect 366294 705478 366914 705562
rect 366294 705242 366326 705478
rect 366562 705242 366646 705478
rect 366882 705242 366914 705478
rect 366294 691954 366914 705242
rect 366294 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 366914 691954
rect 366294 691634 366914 691718
rect 366294 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 366914 691634
rect 366294 655954 366914 691398
rect 366294 655718 366326 655954
rect 366562 655718 366646 655954
rect 366882 655718 366914 655954
rect 366294 655634 366914 655718
rect 366294 655398 366326 655634
rect 366562 655398 366646 655634
rect 366882 655398 366914 655634
rect 366294 619954 366914 655398
rect 366294 619718 366326 619954
rect 366562 619718 366646 619954
rect 366882 619718 366914 619954
rect 366294 619634 366914 619718
rect 366294 619398 366326 619634
rect 366562 619398 366646 619634
rect 366882 619398 366914 619634
rect 366294 583954 366914 619398
rect 366294 583718 366326 583954
rect 366562 583718 366646 583954
rect 366882 583718 366914 583954
rect 366294 583634 366914 583718
rect 366294 583398 366326 583634
rect 366562 583398 366646 583634
rect 366882 583398 366914 583634
rect 366294 547954 366914 583398
rect 366294 547718 366326 547954
rect 366562 547718 366646 547954
rect 366882 547718 366914 547954
rect 366294 547634 366914 547718
rect 366294 547398 366326 547634
rect 366562 547398 366646 547634
rect 366882 547398 366914 547634
rect 366294 511954 366914 547398
rect 366294 511718 366326 511954
rect 366562 511718 366646 511954
rect 366882 511718 366914 511954
rect 366294 511634 366914 511718
rect 366294 511398 366326 511634
rect 366562 511398 366646 511634
rect 366882 511398 366914 511634
rect 366294 475954 366914 511398
rect 366294 475718 366326 475954
rect 366562 475718 366646 475954
rect 366882 475718 366914 475954
rect 366294 475634 366914 475718
rect 366294 475398 366326 475634
rect 366562 475398 366646 475634
rect 366882 475398 366914 475634
rect 366294 439954 366914 475398
rect 366294 439718 366326 439954
rect 366562 439718 366646 439954
rect 366882 439718 366914 439954
rect 366294 439634 366914 439718
rect 366294 439398 366326 439634
rect 366562 439398 366646 439634
rect 366882 439398 366914 439634
rect 366294 403954 366914 439398
rect 366294 403718 366326 403954
rect 366562 403718 366646 403954
rect 366882 403718 366914 403954
rect 366294 403634 366914 403718
rect 366294 403398 366326 403634
rect 366562 403398 366646 403634
rect 366882 403398 366914 403634
rect 366294 367954 366914 403398
rect 366294 367718 366326 367954
rect 366562 367718 366646 367954
rect 366882 367718 366914 367954
rect 366294 367634 366914 367718
rect 366294 367398 366326 367634
rect 366562 367398 366646 367634
rect 366882 367398 366914 367634
rect 366294 331954 366914 367398
rect 366294 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 366914 331954
rect 366294 331634 366914 331718
rect 366294 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 366914 331634
rect 366294 295954 366914 331398
rect 366294 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 366914 295954
rect 366294 295634 366914 295718
rect 366294 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 366914 295634
rect 366294 259954 366914 295398
rect 366294 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 366914 259954
rect 366294 259634 366914 259718
rect 366294 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 366914 259634
rect 366294 223954 366914 259398
rect 366294 223718 366326 223954
rect 366562 223718 366646 223954
rect 366882 223718 366914 223954
rect 366294 223634 366914 223718
rect 366294 223398 366326 223634
rect 366562 223398 366646 223634
rect 366882 223398 366914 223634
rect 366294 187954 366914 223398
rect 366294 187718 366326 187954
rect 366562 187718 366646 187954
rect 366882 187718 366914 187954
rect 366294 187634 366914 187718
rect 366294 187398 366326 187634
rect 366562 187398 366646 187634
rect 366882 187398 366914 187634
rect 366294 151954 366914 187398
rect 366294 151718 366326 151954
rect 366562 151718 366646 151954
rect 366882 151718 366914 151954
rect 366294 151634 366914 151718
rect 366294 151398 366326 151634
rect 366562 151398 366646 151634
rect 366882 151398 366914 151634
rect 366294 115954 366914 151398
rect 366294 115718 366326 115954
rect 366562 115718 366646 115954
rect 366882 115718 366914 115954
rect 366294 115634 366914 115718
rect 366294 115398 366326 115634
rect 366562 115398 366646 115634
rect 366882 115398 366914 115634
rect 366294 79954 366914 115398
rect 366294 79718 366326 79954
rect 366562 79718 366646 79954
rect 366882 79718 366914 79954
rect 366294 79634 366914 79718
rect 366294 79398 366326 79634
rect 366562 79398 366646 79634
rect 366882 79398 366914 79634
rect 366294 43954 366914 79398
rect 366294 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 366914 43954
rect 366294 43634 366914 43718
rect 366294 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 366914 43634
rect 366294 7954 366914 43398
rect 366294 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 366914 7954
rect 366294 7634 366914 7718
rect 366294 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 366914 7634
rect 366294 -1306 366914 7398
rect 366294 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 366914 -1306
rect 366294 -1626 366914 -1542
rect 366294 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 366914 -1626
rect 366294 -7654 366914 -1862
rect 370794 706758 371414 711590
rect 370794 706522 370826 706758
rect 371062 706522 371146 706758
rect 371382 706522 371414 706758
rect 370794 706438 371414 706522
rect 370794 706202 370826 706438
rect 371062 706202 371146 706438
rect 371382 706202 371414 706438
rect 370794 696454 371414 706202
rect 370794 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 371414 696454
rect 370794 696134 371414 696218
rect 370794 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 371414 696134
rect 370794 660454 371414 695898
rect 370794 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 371414 660454
rect 370794 660134 371414 660218
rect 370794 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 371414 660134
rect 370794 624454 371414 659898
rect 370794 624218 370826 624454
rect 371062 624218 371146 624454
rect 371382 624218 371414 624454
rect 370794 624134 371414 624218
rect 370794 623898 370826 624134
rect 371062 623898 371146 624134
rect 371382 623898 371414 624134
rect 370794 588454 371414 623898
rect 370794 588218 370826 588454
rect 371062 588218 371146 588454
rect 371382 588218 371414 588454
rect 370794 588134 371414 588218
rect 370794 587898 370826 588134
rect 371062 587898 371146 588134
rect 371382 587898 371414 588134
rect 370794 552454 371414 587898
rect 370794 552218 370826 552454
rect 371062 552218 371146 552454
rect 371382 552218 371414 552454
rect 370794 552134 371414 552218
rect 370794 551898 370826 552134
rect 371062 551898 371146 552134
rect 371382 551898 371414 552134
rect 370794 516454 371414 551898
rect 370794 516218 370826 516454
rect 371062 516218 371146 516454
rect 371382 516218 371414 516454
rect 370794 516134 371414 516218
rect 370794 515898 370826 516134
rect 371062 515898 371146 516134
rect 371382 515898 371414 516134
rect 370794 480454 371414 515898
rect 370794 480218 370826 480454
rect 371062 480218 371146 480454
rect 371382 480218 371414 480454
rect 370794 480134 371414 480218
rect 370794 479898 370826 480134
rect 371062 479898 371146 480134
rect 371382 479898 371414 480134
rect 370794 444454 371414 479898
rect 370794 444218 370826 444454
rect 371062 444218 371146 444454
rect 371382 444218 371414 444454
rect 370794 444134 371414 444218
rect 370794 443898 370826 444134
rect 371062 443898 371146 444134
rect 371382 443898 371414 444134
rect 370794 408454 371414 443898
rect 370794 408218 370826 408454
rect 371062 408218 371146 408454
rect 371382 408218 371414 408454
rect 370794 408134 371414 408218
rect 370794 407898 370826 408134
rect 371062 407898 371146 408134
rect 371382 407898 371414 408134
rect 370794 372454 371414 407898
rect 370794 372218 370826 372454
rect 371062 372218 371146 372454
rect 371382 372218 371414 372454
rect 370794 372134 371414 372218
rect 370794 371898 370826 372134
rect 371062 371898 371146 372134
rect 371382 371898 371414 372134
rect 370794 336454 371414 371898
rect 370794 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 371414 336454
rect 370794 336134 371414 336218
rect 370794 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 371414 336134
rect 370794 300454 371414 335898
rect 370794 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 371414 300454
rect 370794 300134 371414 300218
rect 370794 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 371414 300134
rect 370794 264454 371414 299898
rect 370794 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 371414 264454
rect 370794 264134 371414 264218
rect 370794 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 371414 264134
rect 370794 228454 371414 263898
rect 370794 228218 370826 228454
rect 371062 228218 371146 228454
rect 371382 228218 371414 228454
rect 370794 228134 371414 228218
rect 370794 227898 370826 228134
rect 371062 227898 371146 228134
rect 371382 227898 371414 228134
rect 370794 192454 371414 227898
rect 370794 192218 370826 192454
rect 371062 192218 371146 192454
rect 371382 192218 371414 192454
rect 370794 192134 371414 192218
rect 370794 191898 370826 192134
rect 371062 191898 371146 192134
rect 371382 191898 371414 192134
rect 370794 156454 371414 191898
rect 370794 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 371414 156454
rect 370794 156134 371414 156218
rect 370794 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 371414 156134
rect 370794 120454 371414 155898
rect 370794 120218 370826 120454
rect 371062 120218 371146 120454
rect 371382 120218 371414 120454
rect 370794 120134 371414 120218
rect 370794 119898 370826 120134
rect 371062 119898 371146 120134
rect 371382 119898 371414 120134
rect 370794 84454 371414 119898
rect 370794 84218 370826 84454
rect 371062 84218 371146 84454
rect 371382 84218 371414 84454
rect 370794 84134 371414 84218
rect 370794 83898 370826 84134
rect 371062 83898 371146 84134
rect 371382 83898 371414 84134
rect 370794 48454 371414 83898
rect 370794 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 371414 48454
rect 370794 48134 371414 48218
rect 370794 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 371414 48134
rect 370794 12454 371414 47898
rect 370794 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 371414 12454
rect 370794 12134 371414 12218
rect 370794 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 371414 12134
rect 370794 -2266 371414 11898
rect 370794 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 371414 -2266
rect 370794 -2586 371414 -2502
rect 370794 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 371414 -2586
rect 370794 -7654 371414 -2822
rect 375294 707718 375914 711590
rect 375294 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 375914 707718
rect 375294 707398 375914 707482
rect 375294 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 375914 707398
rect 375294 700954 375914 707162
rect 375294 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 375914 700954
rect 375294 700634 375914 700718
rect 375294 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 375914 700634
rect 375294 664954 375914 700398
rect 375294 664718 375326 664954
rect 375562 664718 375646 664954
rect 375882 664718 375914 664954
rect 375294 664634 375914 664718
rect 375294 664398 375326 664634
rect 375562 664398 375646 664634
rect 375882 664398 375914 664634
rect 375294 628954 375914 664398
rect 375294 628718 375326 628954
rect 375562 628718 375646 628954
rect 375882 628718 375914 628954
rect 375294 628634 375914 628718
rect 375294 628398 375326 628634
rect 375562 628398 375646 628634
rect 375882 628398 375914 628634
rect 375294 592954 375914 628398
rect 375294 592718 375326 592954
rect 375562 592718 375646 592954
rect 375882 592718 375914 592954
rect 375294 592634 375914 592718
rect 375294 592398 375326 592634
rect 375562 592398 375646 592634
rect 375882 592398 375914 592634
rect 375294 556954 375914 592398
rect 375294 556718 375326 556954
rect 375562 556718 375646 556954
rect 375882 556718 375914 556954
rect 375294 556634 375914 556718
rect 375294 556398 375326 556634
rect 375562 556398 375646 556634
rect 375882 556398 375914 556634
rect 375294 520954 375914 556398
rect 375294 520718 375326 520954
rect 375562 520718 375646 520954
rect 375882 520718 375914 520954
rect 375294 520634 375914 520718
rect 375294 520398 375326 520634
rect 375562 520398 375646 520634
rect 375882 520398 375914 520634
rect 375294 484954 375914 520398
rect 375294 484718 375326 484954
rect 375562 484718 375646 484954
rect 375882 484718 375914 484954
rect 375294 484634 375914 484718
rect 375294 484398 375326 484634
rect 375562 484398 375646 484634
rect 375882 484398 375914 484634
rect 375294 448954 375914 484398
rect 375294 448718 375326 448954
rect 375562 448718 375646 448954
rect 375882 448718 375914 448954
rect 375294 448634 375914 448718
rect 375294 448398 375326 448634
rect 375562 448398 375646 448634
rect 375882 448398 375914 448634
rect 375294 412954 375914 448398
rect 375294 412718 375326 412954
rect 375562 412718 375646 412954
rect 375882 412718 375914 412954
rect 375294 412634 375914 412718
rect 375294 412398 375326 412634
rect 375562 412398 375646 412634
rect 375882 412398 375914 412634
rect 375294 376954 375914 412398
rect 375294 376718 375326 376954
rect 375562 376718 375646 376954
rect 375882 376718 375914 376954
rect 375294 376634 375914 376718
rect 375294 376398 375326 376634
rect 375562 376398 375646 376634
rect 375882 376398 375914 376634
rect 375294 340954 375914 376398
rect 375294 340718 375326 340954
rect 375562 340718 375646 340954
rect 375882 340718 375914 340954
rect 375294 340634 375914 340718
rect 375294 340398 375326 340634
rect 375562 340398 375646 340634
rect 375882 340398 375914 340634
rect 375294 304954 375914 340398
rect 375294 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 375914 304954
rect 375294 304634 375914 304718
rect 375294 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 375914 304634
rect 375294 268954 375914 304398
rect 375294 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 375914 268954
rect 375294 268634 375914 268718
rect 375294 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 375914 268634
rect 375294 232954 375914 268398
rect 375294 232718 375326 232954
rect 375562 232718 375646 232954
rect 375882 232718 375914 232954
rect 375294 232634 375914 232718
rect 375294 232398 375326 232634
rect 375562 232398 375646 232634
rect 375882 232398 375914 232634
rect 375294 196954 375914 232398
rect 375294 196718 375326 196954
rect 375562 196718 375646 196954
rect 375882 196718 375914 196954
rect 375294 196634 375914 196718
rect 375294 196398 375326 196634
rect 375562 196398 375646 196634
rect 375882 196398 375914 196634
rect 375294 160954 375914 196398
rect 375294 160718 375326 160954
rect 375562 160718 375646 160954
rect 375882 160718 375914 160954
rect 375294 160634 375914 160718
rect 375294 160398 375326 160634
rect 375562 160398 375646 160634
rect 375882 160398 375914 160634
rect 375294 124954 375914 160398
rect 375294 124718 375326 124954
rect 375562 124718 375646 124954
rect 375882 124718 375914 124954
rect 375294 124634 375914 124718
rect 375294 124398 375326 124634
rect 375562 124398 375646 124634
rect 375882 124398 375914 124634
rect 375294 88954 375914 124398
rect 375294 88718 375326 88954
rect 375562 88718 375646 88954
rect 375882 88718 375914 88954
rect 375294 88634 375914 88718
rect 375294 88398 375326 88634
rect 375562 88398 375646 88634
rect 375882 88398 375914 88634
rect 375294 52954 375914 88398
rect 375294 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 375914 52954
rect 375294 52634 375914 52718
rect 375294 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 375914 52634
rect 375294 16954 375914 52398
rect 375294 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 375914 16954
rect 375294 16634 375914 16718
rect 375294 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 375914 16634
rect 375294 -3226 375914 16398
rect 375294 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 375914 -3226
rect 375294 -3546 375914 -3462
rect 375294 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 375914 -3546
rect 375294 -7654 375914 -3782
rect 379794 708678 380414 711590
rect 379794 708442 379826 708678
rect 380062 708442 380146 708678
rect 380382 708442 380414 708678
rect 379794 708358 380414 708442
rect 379794 708122 379826 708358
rect 380062 708122 380146 708358
rect 380382 708122 380414 708358
rect 379794 669454 380414 708122
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 453454 380414 488898
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 379794 417454 380414 452898
rect 379794 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 380414 417454
rect 379794 417134 380414 417218
rect 379794 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 380414 417134
rect 379794 381454 380414 416898
rect 379794 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 380414 381454
rect 379794 381134 380414 381218
rect 379794 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 380414 381134
rect 379794 345454 380414 380898
rect 379794 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 380414 345454
rect 379794 345134 380414 345218
rect 379794 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 380414 345134
rect 379794 309454 380414 344898
rect 379794 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 380414 309454
rect 379794 309134 380414 309218
rect 379794 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 380414 309134
rect 379794 273454 380414 308898
rect 379794 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 380414 273454
rect 379794 273134 380414 273218
rect 379794 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 380414 273134
rect 379794 237454 380414 272898
rect 379794 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 380414 237454
rect 379794 237134 380414 237218
rect 379794 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 380414 237134
rect 379794 201454 380414 236898
rect 379794 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 380414 201454
rect 379794 201134 380414 201218
rect 379794 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 380414 201134
rect 379794 165454 380414 200898
rect 379794 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 380414 165454
rect 379794 165134 380414 165218
rect 379794 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 380414 165134
rect 379794 129454 380414 164898
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -4186 380414 20898
rect 379794 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 380414 -4186
rect 379794 -4506 380414 -4422
rect 379794 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 380414 -4506
rect 379794 -7654 380414 -4742
rect 384294 709638 384914 711590
rect 384294 709402 384326 709638
rect 384562 709402 384646 709638
rect 384882 709402 384914 709638
rect 384294 709318 384914 709402
rect 384294 709082 384326 709318
rect 384562 709082 384646 709318
rect 384882 709082 384914 709318
rect 384294 673954 384914 709082
rect 384294 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 384914 673954
rect 384294 673634 384914 673718
rect 384294 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 384914 673634
rect 384294 637954 384914 673398
rect 384294 637718 384326 637954
rect 384562 637718 384646 637954
rect 384882 637718 384914 637954
rect 384294 637634 384914 637718
rect 384294 637398 384326 637634
rect 384562 637398 384646 637634
rect 384882 637398 384914 637634
rect 384294 601954 384914 637398
rect 384294 601718 384326 601954
rect 384562 601718 384646 601954
rect 384882 601718 384914 601954
rect 384294 601634 384914 601718
rect 384294 601398 384326 601634
rect 384562 601398 384646 601634
rect 384882 601398 384914 601634
rect 384294 565954 384914 601398
rect 384294 565718 384326 565954
rect 384562 565718 384646 565954
rect 384882 565718 384914 565954
rect 384294 565634 384914 565718
rect 384294 565398 384326 565634
rect 384562 565398 384646 565634
rect 384882 565398 384914 565634
rect 384294 529954 384914 565398
rect 384294 529718 384326 529954
rect 384562 529718 384646 529954
rect 384882 529718 384914 529954
rect 384294 529634 384914 529718
rect 384294 529398 384326 529634
rect 384562 529398 384646 529634
rect 384882 529398 384914 529634
rect 384294 493954 384914 529398
rect 384294 493718 384326 493954
rect 384562 493718 384646 493954
rect 384882 493718 384914 493954
rect 384294 493634 384914 493718
rect 384294 493398 384326 493634
rect 384562 493398 384646 493634
rect 384882 493398 384914 493634
rect 384294 457954 384914 493398
rect 384294 457718 384326 457954
rect 384562 457718 384646 457954
rect 384882 457718 384914 457954
rect 384294 457634 384914 457718
rect 384294 457398 384326 457634
rect 384562 457398 384646 457634
rect 384882 457398 384914 457634
rect 384294 421954 384914 457398
rect 384294 421718 384326 421954
rect 384562 421718 384646 421954
rect 384882 421718 384914 421954
rect 384294 421634 384914 421718
rect 384294 421398 384326 421634
rect 384562 421398 384646 421634
rect 384882 421398 384914 421634
rect 384294 385954 384914 421398
rect 384294 385718 384326 385954
rect 384562 385718 384646 385954
rect 384882 385718 384914 385954
rect 384294 385634 384914 385718
rect 384294 385398 384326 385634
rect 384562 385398 384646 385634
rect 384882 385398 384914 385634
rect 384294 349954 384914 385398
rect 384294 349718 384326 349954
rect 384562 349718 384646 349954
rect 384882 349718 384914 349954
rect 384294 349634 384914 349718
rect 384294 349398 384326 349634
rect 384562 349398 384646 349634
rect 384882 349398 384914 349634
rect 384294 313954 384914 349398
rect 384294 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 384914 313954
rect 384294 313634 384914 313718
rect 384294 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 384914 313634
rect 384294 277954 384914 313398
rect 384294 277718 384326 277954
rect 384562 277718 384646 277954
rect 384882 277718 384914 277954
rect 384294 277634 384914 277718
rect 384294 277398 384326 277634
rect 384562 277398 384646 277634
rect 384882 277398 384914 277634
rect 384294 241954 384914 277398
rect 384294 241718 384326 241954
rect 384562 241718 384646 241954
rect 384882 241718 384914 241954
rect 384294 241634 384914 241718
rect 384294 241398 384326 241634
rect 384562 241398 384646 241634
rect 384882 241398 384914 241634
rect 384294 205954 384914 241398
rect 384294 205718 384326 205954
rect 384562 205718 384646 205954
rect 384882 205718 384914 205954
rect 384294 205634 384914 205718
rect 384294 205398 384326 205634
rect 384562 205398 384646 205634
rect 384882 205398 384914 205634
rect 384294 169954 384914 205398
rect 384294 169718 384326 169954
rect 384562 169718 384646 169954
rect 384882 169718 384914 169954
rect 384294 169634 384914 169718
rect 384294 169398 384326 169634
rect 384562 169398 384646 169634
rect 384882 169398 384914 169634
rect 384294 133954 384914 169398
rect 384294 133718 384326 133954
rect 384562 133718 384646 133954
rect 384882 133718 384914 133954
rect 384294 133634 384914 133718
rect 384294 133398 384326 133634
rect 384562 133398 384646 133634
rect 384882 133398 384914 133634
rect 384294 97954 384914 133398
rect 384294 97718 384326 97954
rect 384562 97718 384646 97954
rect 384882 97718 384914 97954
rect 384294 97634 384914 97718
rect 384294 97398 384326 97634
rect 384562 97398 384646 97634
rect 384882 97398 384914 97634
rect 384294 61954 384914 97398
rect 384294 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 384914 61954
rect 384294 61634 384914 61718
rect 384294 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 384914 61634
rect 384294 25954 384914 61398
rect 384294 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 384914 25954
rect 384294 25634 384914 25718
rect 384294 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 384914 25634
rect 384294 -5146 384914 25398
rect 384294 -5382 384326 -5146
rect 384562 -5382 384646 -5146
rect 384882 -5382 384914 -5146
rect 384294 -5466 384914 -5382
rect 384294 -5702 384326 -5466
rect 384562 -5702 384646 -5466
rect 384882 -5702 384914 -5466
rect 384294 -7654 384914 -5702
rect 388794 710598 389414 711590
rect 388794 710362 388826 710598
rect 389062 710362 389146 710598
rect 389382 710362 389414 710598
rect 388794 710278 389414 710362
rect 388794 710042 388826 710278
rect 389062 710042 389146 710278
rect 389382 710042 389414 710278
rect 388794 678454 389414 710042
rect 388794 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 389414 678454
rect 388794 678134 389414 678218
rect 388794 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 389414 678134
rect 388794 642454 389414 677898
rect 388794 642218 388826 642454
rect 389062 642218 389146 642454
rect 389382 642218 389414 642454
rect 388794 642134 389414 642218
rect 388794 641898 388826 642134
rect 389062 641898 389146 642134
rect 389382 641898 389414 642134
rect 388794 606454 389414 641898
rect 388794 606218 388826 606454
rect 389062 606218 389146 606454
rect 389382 606218 389414 606454
rect 388794 606134 389414 606218
rect 388794 605898 388826 606134
rect 389062 605898 389146 606134
rect 389382 605898 389414 606134
rect 388794 570454 389414 605898
rect 388794 570218 388826 570454
rect 389062 570218 389146 570454
rect 389382 570218 389414 570454
rect 388794 570134 389414 570218
rect 388794 569898 388826 570134
rect 389062 569898 389146 570134
rect 389382 569898 389414 570134
rect 388794 534454 389414 569898
rect 388794 534218 388826 534454
rect 389062 534218 389146 534454
rect 389382 534218 389414 534454
rect 388794 534134 389414 534218
rect 388794 533898 388826 534134
rect 389062 533898 389146 534134
rect 389382 533898 389414 534134
rect 388794 498454 389414 533898
rect 388794 498218 388826 498454
rect 389062 498218 389146 498454
rect 389382 498218 389414 498454
rect 388794 498134 389414 498218
rect 388794 497898 388826 498134
rect 389062 497898 389146 498134
rect 389382 497898 389414 498134
rect 388794 462454 389414 497898
rect 388794 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 389414 462454
rect 388794 462134 389414 462218
rect 388794 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 389414 462134
rect 388794 426454 389414 461898
rect 388794 426218 388826 426454
rect 389062 426218 389146 426454
rect 389382 426218 389414 426454
rect 388794 426134 389414 426218
rect 388794 425898 388826 426134
rect 389062 425898 389146 426134
rect 389382 425898 389414 426134
rect 388794 390454 389414 425898
rect 388794 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 389414 390454
rect 388794 390134 389414 390218
rect 388794 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 389414 390134
rect 388794 354454 389414 389898
rect 388794 354218 388826 354454
rect 389062 354218 389146 354454
rect 389382 354218 389414 354454
rect 388794 354134 389414 354218
rect 388794 353898 388826 354134
rect 389062 353898 389146 354134
rect 389382 353898 389414 354134
rect 388794 318454 389414 353898
rect 388794 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 389414 318454
rect 388794 318134 389414 318218
rect 388794 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 389414 318134
rect 388794 282454 389414 317898
rect 388794 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 389414 282454
rect 388794 282134 389414 282218
rect 388794 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 389414 282134
rect 388794 246454 389414 281898
rect 388794 246218 388826 246454
rect 389062 246218 389146 246454
rect 389382 246218 389414 246454
rect 388794 246134 389414 246218
rect 388794 245898 388826 246134
rect 389062 245898 389146 246134
rect 389382 245898 389414 246134
rect 388794 210454 389414 245898
rect 388794 210218 388826 210454
rect 389062 210218 389146 210454
rect 389382 210218 389414 210454
rect 388794 210134 389414 210218
rect 388794 209898 388826 210134
rect 389062 209898 389146 210134
rect 389382 209898 389414 210134
rect 388794 174454 389414 209898
rect 388794 174218 388826 174454
rect 389062 174218 389146 174454
rect 389382 174218 389414 174454
rect 388794 174134 389414 174218
rect 388794 173898 388826 174134
rect 389062 173898 389146 174134
rect 389382 173898 389414 174134
rect 388794 138454 389414 173898
rect 388794 138218 388826 138454
rect 389062 138218 389146 138454
rect 389382 138218 389414 138454
rect 388794 138134 389414 138218
rect 388794 137898 388826 138134
rect 389062 137898 389146 138134
rect 389382 137898 389414 138134
rect 388794 102454 389414 137898
rect 388794 102218 388826 102454
rect 389062 102218 389146 102454
rect 389382 102218 389414 102454
rect 388794 102134 389414 102218
rect 388794 101898 388826 102134
rect 389062 101898 389146 102134
rect 389382 101898 389414 102134
rect 388794 66454 389414 101898
rect 388794 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 389414 66454
rect 388794 66134 389414 66218
rect 388794 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 389414 66134
rect 388794 30454 389414 65898
rect 388794 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 389414 30454
rect 388794 30134 389414 30218
rect 388794 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 389414 30134
rect 388794 -6106 389414 29898
rect 388794 -6342 388826 -6106
rect 389062 -6342 389146 -6106
rect 389382 -6342 389414 -6106
rect 388794 -6426 389414 -6342
rect 388794 -6662 388826 -6426
rect 389062 -6662 389146 -6426
rect 389382 -6662 389414 -6426
rect 388794 -7654 389414 -6662
rect 393294 711558 393914 711590
rect 393294 711322 393326 711558
rect 393562 711322 393646 711558
rect 393882 711322 393914 711558
rect 393294 711238 393914 711322
rect 393294 711002 393326 711238
rect 393562 711002 393646 711238
rect 393882 711002 393914 711238
rect 393294 682954 393914 711002
rect 393294 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 393914 682954
rect 393294 682634 393914 682718
rect 393294 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 393914 682634
rect 393294 646954 393914 682398
rect 393294 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 393914 646954
rect 393294 646634 393914 646718
rect 393294 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 393914 646634
rect 393294 610954 393914 646398
rect 393294 610718 393326 610954
rect 393562 610718 393646 610954
rect 393882 610718 393914 610954
rect 393294 610634 393914 610718
rect 393294 610398 393326 610634
rect 393562 610398 393646 610634
rect 393882 610398 393914 610634
rect 393294 574954 393914 610398
rect 393294 574718 393326 574954
rect 393562 574718 393646 574954
rect 393882 574718 393914 574954
rect 393294 574634 393914 574718
rect 393294 574398 393326 574634
rect 393562 574398 393646 574634
rect 393882 574398 393914 574634
rect 393294 538954 393914 574398
rect 393294 538718 393326 538954
rect 393562 538718 393646 538954
rect 393882 538718 393914 538954
rect 393294 538634 393914 538718
rect 393294 538398 393326 538634
rect 393562 538398 393646 538634
rect 393882 538398 393914 538634
rect 393294 502954 393914 538398
rect 393294 502718 393326 502954
rect 393562 502718 393646 502954
rect 393882 502718 393914 502954
rect 393294 502634 393914 502718
rect 393294 502398 393326 502634
rect 393562 502398 393646 502634
rect 393882 502398 393914 502634
rect 393294 466954 393914 502398
rect 393294 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 393914 466954
rect 393294 466634 393914 466718
rect 393294 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 393914 466634
rect 393294 430954 393914 466398
rect 393294 430718 393326 430954
rect 393562 430718 393646 430954
rect 393882 430718 393914 430954
rect 393294 430634 393914 430718
rect 393294 430398 393326 430634
rect 393562 430398 393646 430634
rect 393882 430398 393914 430634
rect 393294 394954 393914 430398
rect 393294 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 393914 394954
rect 393294 394634 393914 394718
rect 393294 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 393914 394634
rect 393294 358954 393914 394398
rect 393294 358718 393326 358954
rect 393562 358718 393646 358954
rect 393882 358718 393914 358954
rect 393294 358634 393914 358718
rect 393294 358398 393326 358634
rect 393562 358398 393646 358634
rect 393882 358398 393914 358634
rect 393294 322954 393914 358398
rect 393294 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 393914 322954
rect 393294 322634 393914 322718
rect 393294 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 393914 322634
rect 393294 286954 393914 322398
rect 393294 286718 393326 286954
rect 393562 286718 393646 286954
rect 393882 286718 393914 286954
rect 393294 286634 393914 286718
rect 393294 286398 393326 286634
rect 393562 286398 393646 286634
rect 393882 286398 393914 286634
rect 393294 250954 393914 286398
rect 393294 250718 393326 250954
rect 393562 250718 393646 250954
rect 393882 250718 393914 250954
rect 393294 250634 393914 250718
rect 393294 250398 393326 250634
rect 393562 250398 393646 250634
rect 393882 250398 393914 250634
rect 393294 214954 393914 250398
rect 393294 214718 393326 214954
rect 393562 214718 393646 214954
rect 393882 214718 393914 214954
rect 393294 214634 393914 214718
rect 393294 214398 393326 214634
rect 393562 214398 393646 214634
rect 393882 214398 393914 214634
rect 393294 178954 393914 214398
rect 393294 178718 393326 178954
rect 393562 178718 393646 178954
rect 393882 178718 393914 178954
rect 393294 178634 393914 178718
rect 393294 178398 393326 178634
rect 393562 178398 393646 178634
rect 393882 178398 393914 178634
rect 393294 142954 393914 178398
rect 393294 142718 393326 142954
rect 393562 142718 393646 142954
rect 393882 142718 393914 142954
rect 393294 142634 393914 142718
rect 393294 142398 393326 142634
rect 393562 142398 393646 142634
rect 393882 142398 393914 142634
rect 393294 106954 393914 142398
rect 393294 106718 393326 106954
rect 393562 106718 393646 106954
rect 393882 106718 393914 106954
rect 393294 106634 393914 106718
rect 393294 106398 393326 106634
rect 393562 106398 393646 106634
rect 393882 106398 393914 106634
rect 393294 70954 393914 106398
rect 393294 70718 393326 70954
rect 393562 70718 393646 70954
rect 393882 70718 393914 70954
rect 393294 70634 393914 70718
rect 393294 70398 393326 70634
rect 393562 70398 393646 70634
rect 393882 70398 393914 70634
rect 393294 34954 393914 70398
rect 393294 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 393914 34954
rect 393294 34634 393914 34718
rect 393294 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 393914 34634
rect 393294 -7066 393914 34398
rect 393294 -7302 393326 -7066
rect 393562 -7302 393646 -7066
rect 393882 -7302 393914 -7066
rect 393294 -7386 393914 -7302
rect 393294 -7622 393326 -7386
rect 393562 -7622 393646 -7386
rect 393882 -7622 393914 -7386
rect 393294 -7654 393914 -7622
rect 397794 704838 398414 711590
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -7654 398414 -902
rect 402294 705798 402914 711590
rect 402294 705562 402326 705798
rect 402562 705562 402646 705798
rect 402882 705562 402914 705798
rect 402294 705478 402914 705562
rect 402294 705242 402326 705478
rect 402562 705242 402646 705478
rect 402882 705242 402914 705478
rect 402294 691954 402914 705242
rect 402294 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 402914 691954
rect 402294 691634 402914 691718
rect 402294 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 402914 691634
rect 402294 655954 402914 691398
rect 402294 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 402914 655954
rect 402294 655634 402914 655718
rect 402294 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 402914 655634
rect 402294 619954 402914 655398
rect 402294 619718 402326 619954
rect 402562 619718 402646 619954
rect 402882 619718 402914 619954
rect 402294 619634 402914 619718
rect 402294 619398 402326 619634
rect 402562 619398 402646 619634
rect 402882 619398 402914 619634
rect 402294 583954 402914 619398
rect 402294 583718 402326 583954
rect 402562 583718 402646 583954
rect 402882 583718 402914 583954
rect 402294 583634 402914 583718
rect 402294 583398 402326 583634
rect 402562 583398 402646 583634
rect 402882 583398 402914 583634
rect 402294 547954 402914 583398
rect 402294 547718 402326 547954
rect 402562 547718 402646 547954
rect 402882 547718 402914 547954
rect 402294 547634 402914 547718
rect 402294 547398 402326 547634
rect 402562 547398 402646 547634
rect 402882 547398 402914 547634
rect 402294 511954 402914 547398
rect 402294 511718 402326 511954
rect 402562 511718 402646 511954
rect 402882 511718 402914 511954
rect 402294 511634 402914 511718
rect 402294 511398 402326 511634
rect 402562 511398 402646 511634
rect 402882 511398 402914 511634
rect 402294 475954 402914 511398
rect 402294 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 402914 475954
rect 402294 475634 402914 475718
rect 402294 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 402914 475634
rect 402294 439954 402914 475398
rect 402294 439718 402326 439954
rect 402562 439718 402646 439954
rect 402882 439718 402914 439954
rect 402294 439634 402914 439718
rect 402294 439398 402326 439634
rect 402562 439398 402646 439634
rect 402882 439398 402914 439634
rect 402294 403954 402914 439398
rect 402294 403718 402326 403954
rect 402562 403718 402646 403954
rect 402882 403718 402914 403954
rect 402294 403634 402914 403718
rect 402294 403398 402326 403634
rect 402562 403398 402646 403634
rect 402882 403398 402914 403634
rect 402294 367954 402914 403398
rect 402294 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 402914 367954
rect 402294 367634 402914 367718
rect 402294 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 402914 367634
rect 402294 331954 402914 367398
rect 402294 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 402914 331954
rect 402294 331634 402914 331718
rect 402294 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 402914 331634
rect 402294 295954 402914 331398
rect 402294 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 402914 295954
rect 402294 295634 402914 295718
rect 402294 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 402914 295634
rect 402294 259954 402914 295398
rect 402294 259718 402326 259954
rect 402562 259718 402646 259954
rect 402882 259718 402914 259954
rect 402294 259634 402914 259718
rect 402294 259398 402326 259634
rect 402562 259398 402646 259634
rect 402882 259398 402914 259634
rect 402294 223954 402914 259398
rect 402294 223718 402326 223954
rect 402562 223718 402646 223954
rect 402882 223718 402914 223954
rect 402294 223634 402914 223718
rect 402294 223398 402326 223634
rect 402562 223398 402646 223634
rect 402882 223398 402914 223634
rect 402294 187954 402914 223398
rect 402294 187718 402326 187954
rect 402562 187718 402646 187954
rect 402882 187718 402914 187954
rect 402294 187634 402914 187718
rect 402294 187398 402326 187634
rect 402562 187398 402646 187634
rect 402882 187398 402914 187634
rect 402294 151954 402914 187398
rect 402294 151718 402326 151954
rect 402562 151718 402646 151954
rect 402882 151718 402914 151954
rect 402294 151634 402914 151718
rect 402294 151398 402326 151634
rect 402562 151398 402646 151634
rect 402882 151398 402914 151634
rect 402294 115954 402914 151398
rect 402294 115718 402326 115954
rect 402562 115718 402646 115954
rect 402882 115718 402914 115954
rect 402294 115634 402914 115718
rect 402294 115398 402326 115634
rect 402562 115398 402646 115634
rect 402882 115398 402914 115634
rect 402294 79954 402914 115398
rect 402294 79718 402326 79954
rect 402562 79718 402646 79954
rect 402882 79718 402914 79954
rect 402294 79634 402914 79718
rect 402294 79398 402326 79634
rect 402562 79398 402646 79634
rect 402882 79398 402914 79634
rect 402294 43954 402914 79398
rect 402294 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 402914 43954
rect 402294 43634 402914 43718
rect 402294 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 402914 43634
rect 402294 7954 402914 43398
rect 402294 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 402914 7954
rect 402294 7634 402914 7718
rect 402294 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 402914 7634
rect 402294 -1306 402914 7398
rect 402294 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 402914 -1306
rect 402294 -1626 402914 -1542
rect 402294 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 402914 -1626
rect 402294 -7654 402914 -1862
rect 406794 706758 407414 711590
rect 406794 706522 406826 706758
rect 407062 706522 407146 706758
rect 407382 706522 407414 706758
rect 406794 706438 407414 706522
rect 406794 706202 406826 706438
rect 407062 706202 407146 706438
rect 407382 706202 407414 706438
rect 406794 696454 407414 706202
rect 406794 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 407414 696454
rect 406794 696134 407414 696218
rect 406794 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 407414 696134
rect 406794 660454 407414 695898
rect 406794 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 407414 660454
rect 406794 660134 407414 660218
rect 406794 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 407414 660134
rect 406794 624454 407414 659898
rect 406794 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 407414 624454
rect 406794 624134 407414 624218
rect 406794 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 407414 624134
rect 406794 588454 407414 623898
rect 406794 588218 406826 588454
rect 407062 588218 407146 588454
rect 407382 588218 407414 588454
rect 406794 588134 407414 588218
rect 406794 587898 406826 588134
rect 407062 587898 407146 588134
rect 407382 587898 407414 588134
rect 406794 552454 407414 587898
rect 406794 552218 406826 552454
rect 407062 552218 407146 552454
rect 407382 552218 407414 552454
rect 406794 552134 407414 552218
rect 406794 551898 406826 552134
rect 407062 551898 407146 552134
rect 407382 551898 407414 552134
rect 406794 516454 407414 551898
rect 406794 516218 406826 516454
rect 407062 516218 407146 516454
rect 407382 516218 407414 516454
rect 406794 516134 407414 516218
rect 406794 515898 406826 516134
rect 407062 515898 407146 516134
rect 407382 515898 407414 516134
rect 406794 480454 407414 515898
rect 406794 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 407414 480454
rect 406794 480134 407414 480218
rect 406794 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 407414 480134
rect 406794 444454 407414 479898
rect 406794 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 407414 444454
rect 406794 444134 407414 444218
rect 406794 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 407414 444134
rect 406794 408454 407414 443898
rect 406794 408218 406826 408454
rect 407062 408218 407146 408454
rect 407382 408218 407414 408454
rect 406794 408134 407414 408218
rect 406794 407898 406826 408134
rect 407062 407898 407146 408134
rect 407382 407898 407414 408134
rect 406794 372454 407414 407898
rect 406794 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 407414 372454
rect 406794 372134 407414 372218
rect 406794 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 407414 372134
rect 406794 336454 407414 371898
rect 406794 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 407414 336454
rect 406794 336134 407414 336218
rect 406794 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 407414 336134
rect 406794 300454 407414 335898
rect 406794 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 407414 300454
rect 406794 300134 407414 300218
rect 406794 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 407414 300134
rect 406794 264454 407414 299898
rect 406794 264218 406826 264454
rect 407062 264218 407146 264454
rect 407382 264218 407414 264454
rect 406794 264134 407414 264218
rect 406794 263898 406826 264134
rect 407062 263898 407146 264134
rect 407382 263898 407414 264134
rect 406794 228454 407414 263898
rect 406794 228218 406826 228454
rect 407062 228218 407146 228454
rect 407382 228218 407414 228454
rect 406794 228134 407414 228218
rect 406794 227898 406826 228134
rect 407062 227898 407146 228134
rect 407382 227898 407414 228134
rect 406794 192454 407414 227898
rect 406794 192218 406826 192454
rect 407062 192218 407146 192454
rect 407382 192218 407414 192454
rect 406794 192134 407414 192218
rect 406794 191898 406826 192134
rect 407062 191898 407146 192134
rect 407382 191898 407414 192134
rect 406794 156454 407414 191898
rect 406794 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 407414 156454
rect 406794 156134 407414 156218
rect 406794 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 407414 156134
rect 406794 120454 407414 155898
rect 406794 120218 406826 120454
rect 407062 120218 407146 120454
rect 407382 120218 407414 120454
rect 406794 120134 407414 120218
rect 406794 119898 406826 120134
rect 407062 119898 407146 120134
rect 407382 119898 407414 120134
rect 406794 84454 407414 119898
rect 406794 84218 406826 84454
rect 407062 84218 407146 84454
rect 407382 84218 407414 84454
rect 406794 84134 407414 84218
rect 406794 83898 406826 84134
rect 407062 83898 407146 84134
rect 407382 83898 407414 84134
rect 406794 48454 407414 83898
rect 406794 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 407414 48454
rect 406794 48134 407414 48218
rect 406794 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 407414 48134
rect 406794 12454 407414 47898
rect 406794 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 407414 12454
rect 406794 12134 407414 12218
rect 406794 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 407414 12134
rect 406794 -2266 407414 11898
rect 406794 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 407414 -2266
rect 406794 -2586 407414 -2502
rect 406794 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 407414 -2586
rect 406794 -7654 407414 -2822
rect 411294 707718 411914 711590
rect 411294 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 411914 707718
rect 411294 707398 411914 707482
rect 411294 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 411914 707398
rect 411294 700954 411914 707162
rect 411294 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 411914 700954
rect 411294 700634 411914 700718
rect 411294 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 411914 700634
rect 411294 664954 411914 700398
rect 411294 664718 411326 664954
rect 411562 664718 411646 664954
rect 411882 664718 411914 664954
rect 411294 664634 411914 664718
rect 411294 664398 411326 664634
rect 411562 664398 411646 664634
rect 411882 664398 411914 664634
rect 411294 628954 411914 664398
rect 411294 628718 411326 628954
rect 411562 628718 411646 628954
rect 411882 628718 411914 628954
rect 411294 628634 411914 628718
rect 411294 628398 411326 628634
rect 411562 628398 411646 628634
rect 411882 628398 411914 628634
rect 411294 592954 411914 628398
rect 411294 592718 411326 592954
rect 411562 592718 411646 592954
rect 411882 592718 411914 592954
rect 411294 592634 411914 592718
rect 411294 592398 411326 592634
rect 411562 592398 411646 592634
rect 411882 592398 411914 592634
rect 411294 556954 411914 592398
rect 411294 556718 411326 556954
rect 411562 556718 411646 556954
rect 411882 556718 411914 556954
rect 411294 556634 411914 556718
rect 411294 556398 411326 556634
rect 411562 556398 411646 556634
rect 411882 556398 411914 556634
rect 411294 520954 411914 556398
rect 411294 520718 411326 520954
rect 411562 520718 411646 520954
rect 411882 520718 411914 520954
rect 411294 520634 411914 520718
rect 411294 520398 411326 520634
rect 411562 520398 411646 520634
rect 411882 520398 411914 520634
rect 411294 484954 411914 520398
rect 411294 484718 411326 484954
rect 411562 484718 411646 484954
rect 411882 484718 411914 484954
rect 411294 484634 411914 484718
rect 411294 484398 411326 484634
rect 411562 484398 411646 484634
rect 411882 484398 411914 484634
rect 411294 448954 411914 484398
rect 411294 448718 411326 448954
rect 411562 448718 411646 448954
rect 411882 448718 411914 448954
rect 411294 448634 411914 448718
rect 411294 448398 411326 448634
rect 411562 448398 411646 448634
rect 411882 448398 411914 448634
rect 411294 412954 411914 448398
rect 411294 412718 411326 412954
rect 411562 412718 411646 412954
rect 411882 412718 411914 412954
rect 411294 412634 411914 412718
rect 411294 412398 411326 412634
rect 411562 412398 411646 412634
rect 411882 412398 411914 412634
rect 411294 376954 411914 412398
rect 411294 376718 411326 376954
rect 411562 376718 411646 376954
rect 411882 376718 411914 376954
rect 411294 376634 411914 376718
rect 411294 376398 411326 376634
rect 411562 376398 411646 376634
rect 411882 376398 411914 376634
rect 411294 340954 411914 376398
rect 411294 340718 411326 340954
rect 411562 340718 411646 340954
rect 411882 340718 411914 340954
rect 411294 340634 411914 340718
rect 411294 340398 411326 340634
rect 411562 340398 411646 340634
rect 411882 340398 411914 340634
rect 411294 304954 411914 340398
rect 411294 304718 411326 304954
rect 411562 304718 411646 304954
rect 411882 304718 411914 304954
rect 411294 304634 411914 304718
rect 411294 304398 411326 304634
rect 411562 304398 411646 304634
rect 411882 304398 411914 304634
rect 411294 268954 411914 304398
rect 411294 268718 411326 268954
rect 411562 268718 411646 268954
rect 411882 268718 411914 268954
rect 411294 268634 411914 268718
rect 411294 268398 411326 268634
rect 411562 268398 411646 268634
rect 411882 268398 411914 268634
rect 411294 232954 411914 268398
rect 411294 232718 411326 232954
rect 411562 232718 411646 232954
rect 411882 232718 411914 232954
rect 411294 232634 411914 232718
rect 411294 232398 411326 232634
rect 411562 232398 411646 232634
rect 411882 232398 411914 232634
rect 411294 196954 411914 232398
rect 411294 196718 411326 196954
rect 411562 196718 411646 196954
rect 411882 196718 411914 196954
rect 411294 196634 411914 196718
rect 411294 196398 411326 196634
rect 411562 196398 411646 196634
rect 411882 196398 411914 196634
rect 411294 160954 411914 196398
rect 411294 160718 411326 160954
rect 411562 160718 411646 160954
rect 411882 160718 411914 160954
rect 411294 160634 411914 160718
rect 411294 160398 411326 160634
rect 411562 160398 411646 160634
rect 411882 160398 411914 160634
rect 411294 124954 411914 160398
rect 411294 124718 411326 124954
rect 411562 124718 411646 124954
rect 411882 124718 411914 124954
rect 411294 124634 411914 124718
rect 411294 124398 411326 124634
rect 411562 124398 411646 124634
rect 411882 124398 411914 124634
rect 411294 88954 411914 124398
rect 411294 88718 411326 88954
rect 411562 88718 411646 88954
rect 411882 88718 411914 88954
rect 411294 88634 411914 88718
rect 411294 88398 411326 88634
rect 411562 88398 411646 88634
rect 411882 88398 411914 88634
rect 411294 52954 411914 88398
rect 411294 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 411914 52954
rect 411294 52634 411914 52718
rect 411294 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 411914 52634
rect 411294 16954 411914 52398
rect 411294 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 411914 16954
rect 411294 16634 411914 16718
rect 411294 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 411914 16634
rect 411294 -3226 411914 16398
rect 411294 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 411914 -3226
rect 411294 -3546 411914 -3462
rect 411294 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 411914 -3546
rect 411294 -7654 411914 -3782
rect 415794 708678 416414 711590
rect 415794 708442 415826 708678
rect 416062 708442 416146 708678
rect 416382 708442 416414 708678
rect 415794 708358 416414 708442
rect 415794 708122 415826 708358
rect 416062 708122 416146 708358
rect 416382 708122 416414 708358
rect 415794 669454 416414 708122
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 525454 416414 560898
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 453454 416414 488898
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 417454 416414 452898
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 381454 416414 416898
rect 415794 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 416414 381454
rect 415794 381134 416414 381218
rect 415794 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 416414 381134
rect 415794 345454 416414 380898
rect 415794 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 416414 345454
rect 415794 345134 416414 345218
rect 415794 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 416414 345134
rect 415794 309454 416414 344898
rect 415794 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 416414 309454
rect 415794 309134 416414 309218
rect 415794 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 416414 309134
rect 415794 273454 416414 308898
rect 415794 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 416414 273454
rect 415794 273134 416414 273218
rect 415794 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 416414 273134
rect 415794 237454 416414 272898
rect 415794 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 416414 237454
rect 415794 237134 416414 237218
rect 415794 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 416414 237134
rect 415794 201454 416414 236898
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 415794 165454 416414 200898
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 415794 129454 416414 164898
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 415794 93454 416414 128898
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -4186 416414 20898
rect 415794 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 416414 -4186
rect 415794 -4506 416414 -4422
rect 415794 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 416414 -4506
rect 415794 -7654 416414 -4742
rect 420294 709638 420914 711590
rect 420294 709402 420326 709638
rect 420562 709402 420646 709638
rect 420882 709402 420914 709638
rect 420294 709318 420914 709402
rect 420294 709082 420326 709318
rect 420562 709082 420646 709318
rect 420882 709082 420914 709318
rect 420294 673954 420914 709082
rect 420294 673718 420326 673954
rect 420562 673718 420646 673954
rect 420882 673718 420914 673954
rect 420294 673634 420914 673718
rect 420294 673398 420326 673634
rect 420562 673398 420646 673634
rect 420882 673398 420914 673634
rect 420294 637954 420914 673398
rect 420294 637718 420326 637954
rect 420562 637718 420646 637954
rect 420882 637718 420914 637954
rect 420294 637634 420914 637718
rect 420294 637398 420326 637634
rect 420562 637398 420646 637634
rect 420882 637398 420914 637634
rect 420294 601954 420914 637398
rect 420294 601718 420326 601954
rect 420562 601718 420646 601954
rect 420882 601718 420914 601954
rect 420294 601634 420914 601718
rect 420294 601398 420326 601634
rect 420562 601398 420646 601634
rect 420882 601398 420914 601634
rect 420294 565954 420914 601398
rect 420294 565718 420326 565954
rect 420562 565718 420646 565954
rect 420882 565718 420914 565954
rect 420294 565634 420914 565718
rect 420294 565398 420326 565634
rect 420562 565398 420646 565634
rect 420882 565398 420914 565634
rect 420294 529954 420914 565398
rect 420294 529718 420326 529954
rect 420562 529718 420646 529954
rect 420882 529718 420914 529954
rect 420294 529634 420914 529718
rect 420294 529398 420326 529634
rect 420562 529398 420646 529634
rect 420882 529398 420914 529634
rect 420294 493954 420914 529398
rect 420294 493718 420326 493954
rect 420562 493718 420646 493954
rect 420882 493718 420914 493954
rect 420294 493634 420914 493718
rect 420294 493398 420326 493634
rect 420562 493398 420646 493634
rect 420882 493398 420914 493634
rect 420294 457954 420914 493398
rect 420294 457718 420326 457954
rect 420562 457718 420646 457954
rect 420882 457718 420914 457954
rect 420294 457634 420914 457718
rect 420294 457398 420326 457634
rect 420562 457398 420646 457634
rect 420882 457398 420914 457634
rect 420294 421954 420914 457398
rect 420294 421718 420326 421954
rect 420562 421718 420646 421954
rect 420882 421718 420914 421954
rect 420294 421634 420914 421718
rect 420294 421398 420326 421634
rect 420562 421398 420646 421634
rect 420882 421398 420914 421634
rect 420294 385954 420914 421398
rect 420294 385718 420326 385954
rect 420562 385718 420646 385954
rect 420882 385718 420914 385954
rect 420294 385634 420914 385718
rect 420294 385398 420326 385634
rect 420562 385398 420646 385634
rect 420882 385398 420914 385634
rect 420294 349954 420914 385398
rect 420294 349718 420326 349954
rect 420562 349718 420646 349954
rect 420882 349718 420914 349954
rect 420294 349634 420914 349718
rect 420294 349398 420326 349634
rect 420562 349398 420646 349634
rect 420882 349398 420914 349634
rect 420294 313954 420914 349398
rect 420294 313718 420326 313954
rect 420562 313718 420646 313954
rect 420882 313718 420914 313954
rect 420294 313634 420914 313718
rect 420294 313398 420326 313634
rect 420562 313398 420646 313634
rect 420882 313398 420914 313634
rect 420294 277954 420914 313398
rect 420294 277718 420326 277954
rect 420562 277718 420646 277954
rect 420882 277718 420914 277954
rect 420294 277634 420914 277718
rect 420294 277398 420326 277634
rect 420562 277398 420646 277634
rect 420882 277398 420914 277634
rect 420294 241954 420914 277398
rect 420294 241718 420326 241954
rect 420562 241718 420646 241954
rect 420882 241718 420914 241954
rect 420294 241634 420914 241718
rect 420294 241398 420326 241634
rect 420562 241398 420646 241634
rect 420882 241398 420914 241634
rect 420294 205954 420914 241398
rect 420294 205718 420326 205954
rect 420562 205718 420646 205954
rect 420882 205718 420914 205954
rect 420294 205634 420914 205718
rect 420294 205398 420326 205634
rect 420562 205398 420646 205634
rect 420882 205398 420914 205634
rect 420294 169954 420914 205398
rect 420294 169718 420326 169954
rect 420562 169718 420646 169954
rect 420882 169718 420914 169954
rect 420294 169634 420914 169718
rect 420294 169398 420326 169634
rect 420562 169398 420646 169634
rect 420882 169398 420914 169634
rect 420294 133954 420914 169398
rect 420294 133718 420326 133954
rect 420562 133718 420646 133954
rect 420882 133718 420914 133954
rect 420294 133634 420914 133718
rect 420294 133398 420326 133634
rect 420562 133398 420646 133634
rect 420882 133398 420914 133634
rect 420294 97954 420914 133398
rect 420294 97718 420326 97954
rect 420562 97718 420646 97954
rect 420882 97718 420914 97954
rect 420294 97634 420914 97718
rect 420294 97398 420326 97634
rect 420562 97398 420646 97634
rect 420882 97398 420914 97634
rect 420294 61954 420914 97398
rect 420294 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 420914 61954
rect 420294 61634 420914 61718
rect 420294 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 420914 61634
rect 420294 25954 420914 61398
rect 420294 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 420914 25954
rect 420294 25634 420914 25718
rect 420294 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 420914 25634
rect 420294 -5146 420914 25398
rect 420294 -5382 420326 -5146
rect 420562 -5382 420646 -5146
rect 420882 -5382 420914 -5146
rect 420294 -5466 420914 -5382
rect 420294 -5702 420326 -5466
rect 420562 -5702 420646 -5466
rect 420882 -5702 420914 -5466
rect 420294 -7654 420914 -5702
rect 424794 710598 425414 711590
rect 424794 710362 424826 710598
rect 425062 710362 425146 710598
rect 425382 710362 425414 710598
rect 424794 710278 425414 710362
rect 424794 710042 424826 710278
rect 425062 710042 425146 710278
rect 425382 710042 425414 710278
rect 424794 678454 425414 710042
rect 424794 678218 424826 678454
rect 425062 678218 425146 678454
rect 425382 678218 425414 678454
rect 424794 678134 425414 678218
rect 424794 677898 424826 678134
rect 425062 677898 425146 678134
rect 425382 677898 425414 678134
rect 424794 642454 425414 677898
rect 424794 642218 424826 642454
rect 425062 642218 425146 642454
rect 425382 642218 425414 642454
rect 424794 642134 425414 642218
rect 424794 641898 424826 642134
rect 425062 641898 425146 642134
rect 425382 641898 425414 642134
rect 424794 606454 425414 641898
rect 424794 606218 424826 606454
rect 425062 606218 425146 606454
rect 425382 606218 425414 606454
rect 424794 606134 425414 606218
rect 424794 605898 424826 606134
rect 425062 605898 425146 606134
rect 425382 605898 425414 606134
rect 424794 570454 425414 605898
rect 424794 570218 424826 570454
rect 425062 570218 425146 570454
rect 425382 570218 425414 570454
rect 424794 570134 425414 570218
rect 424794 569898 424826 570134
rect 425062 569898 425146 570134
rect 425382 569898 425414 570134
rect 424794 534454 425414 569898
rect 424794 534218 424826 534454
rect 425062 534218 425146 534454
rect 425382 534218 425414 534454
rect 424794 534134 425414 534218
rect 424794 533898 424826 534134
rect 425062 533898 425146 534134
rect 425382 533898 425414 534134
rect 424794 498454 425414 533898
rect 424794 498218 424826 498454
rect 425062 498218 425146 498454
rect 425382 498218 425414 498454
rect 424794 498134 425414 498218
rect 424794 497898 424826 498134
rect 425062 497898 425146 498134
rect 425382 497898 425414 498134
rect 424794 462454 425414 497898
rect 424794 462218 424826 462454
rect 425062 462218 425146 462454
rect 425382 462218 425414 462454
rect 424794 462134 425414 462218
rect 424794 461898 424826 462134
rect 425062 461898 425146 462134
rect 425382 461898 425414 462134
rect 424794 426454 425414 461898
rect 424794 426218 424826 426454
rect 425062 426218 425146 426454
rect 425382 426218 425414 426454
rect 424794 426134 425414 426218
rect 424794 425898 424826 426134
rect 425062 425898 425146 426134
rect 425382 425898 425414 426134
rect 424794 390454 425414 425898
rect 424794 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 425414 390454
rect 424794 390134 425414 390218
rect 424794 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 425414 390134
rect 424794 354454 425414 389898
rect 424794 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 425414 354454
rect 424794 354134 425414 354218
rect 424794 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 425414 354134
rect 424794 318454 425414 353898
rect 424794 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 425414 318454
rect 424794 318134 425414 318218
rect 424794 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 425414 318134
rect 424794 282454 425414 317898
rect 424794 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 425414 282454
rect 424794 282134 425414 282218
rect 424794 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 425414 282134
rect 424794 246454 425414 281898
rect 424794 246218 424826 246454
rect 425062 246218 425146 246454
rect 425382 246218 425414 246454
rect 424794 246134 425414 246218
rect 424794 245898 424826 246134
rect 425062 245898 425146 246134
rect 425382 245898 425414 246134
rect 424794 210454 425414 245898
rect 424794 210218 424826 210454
rect 425062 210218 425146 210454
rect 425382 210218 425414 210454
rect 424794 210134 425414 210218
rect 424794 209898 424826 210134
rect 425062 209898 425146 210134
rect 425382 209898 425414 210134
rect 424794 174454 425414 209898
rect 424794 174218 424826 174454
rect 425062 174218 425146 174454
rect 425382 174218 425414 174454
rect 424794 174134 425414 174218
rect 424794 173898 424826 174134
rect 425062 173898 425146 174134
rect 425382 173898 425414 174134
rect 424794 138454 425414 173898
rect 424794 138218 424826 138454
rect 425062 138218 425146 138454
rect 425382 138218 425414 138454
rect 424794 138134 425414 138218
rect 424794 137898 424826 138134
rect 425062 137898 425146 138134
rect 425382 137898 425414 138134
rect 424794 102454 425414 137898
rect 424794 102218 424826 102454
rect 425062 102218 425146 102454
rect 425382 102218 425414 102454
rect 424794 102134 425414 102218
rect 424794 101898 424826 102134
rect 425062 101898 425146 102134
rect 425382 101898 425414 102134
rect 424794 66454 425414 101898
rect 424794 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 425414 66454
rect 424794 66134 425414 66218
rect 424794 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 425414 66134
rect 424794 30454 425414 65898
rect 424794 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 425414 30454
rect 424794 30134 425414 30218
rect 424794 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 425414 30134
rect 424794 -6106 425414 29898
rect 424794 -6342 424826 -6106
rect 425062 -6342 425146 -6106
rect 425382 -6342 425414 -6106
rect 424794 -6426 425414 -6342
rect 424794 -6662 424826 -6426
rect 425062 -6662 425146 -6426
rect 425382 -6662 425414 -6426
rect 424794 -7654 425414 -6662
rect 429294 711558 429914 711590
rect 429294 711322 429326 711558
rect 429562 711322 429646 711558
rect 429882 711322 429914 711558
rect 429294 711238 429914 711322
rect 429294 711002 429326 711238
rect 429562 711002 429646 711238
rect 429882 711002 429914 711238
rect 429294 682954 429914 711002
rect 429294 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 429914 682954
rect 429294 682634 429914 682718
rect 429294 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 429914 682634
rect 429294 646954 429914 682398
rect 429294 646718 429326 646954
rect 429562 646718 429646 646954
rect 429882 646718 429914 646954
rect 429294 646634 429914 646718
rect 429294 646398 429326 646634
rect 429562 646398 429646 646634
rect 429882 646398 429914 646634
rect 429294 610954 429914 646398
rect 429294 610718 429326 610954
rect 429562 610718 429646 610954
rect 429882 610718 429914 610954
rect 429294 610634 429914 610718
rect 429294 610398 429326 610634
rect 429562 610398 429646 610634
rect 429882 610398 429914 610634
rect 429294 574954 429914 610398
rect 429294 574718 429326 574954
rect 429562 574718 429646 574954
rect 429882 574718 429914 574954
rect 429294 574634 429914 574718
rect 429294 574398 429326 574634
rect 429562 574398 429646 574634
rect 429882 574398 429914 574634
rect 429294 538954 429914 574398
rect 429294 538718 429326 538954
rect 429562 538718 429646 538954
rect 429882 538718 429914 538954
rect 429294 538634 429914 538718
rect 429294 538398 429326 538634
rect 429562 538398 429646 538634
rect 429882 538398 429914 538634
rect 429294 502954 429914 538398
rect 429294 502718 429326 502954
rect 429562 502718 429646 502954
rect 429882 502718 429914 502954
rect 429294 502634 429914 502718
rect 429294 502398 429326 502634
rect 429562 502398 429646 502634
rect 429882 502398 429914 502634
rect 429294 466954 429914 502398
rect 429294 466718 429326 466954
rect 429562 466718 429646 466954
rect 429882 466718 429914 466954
rect 429294 466634 429914 466718
rect 429294 466398 429326 466634
rect 429562 466398 429646 466634
rect 429882 466398 429914 466634
rect 429294 430954 429914 466398
rect 429294 430718 429326 430954
rect 429562 430718 429646 430954
rect 429882 430718 429914 430954
rect 429294 430634 429914 430718
rect 429294 430398 429326 430634
rect 429562 430398 429646 430634
rect 429882 430398 429914 430634
rect 429294 394954 429914 430398
rect 429294 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 429914 394954
rect 429294 394634 429914 394718
rect 429294 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 429914 394634
rect 429294 358954 429914 394398
rect 429294 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 429914 358954
rect 429294 358634 429914 358718
rect 429294 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 429914 358634
rect 429294 322954 429914 358398
rect 429294 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 429914 322954
rect 429294 322634 429914 322718
rect 429294 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 429914 322634
rect 429294 286954 429914 322398
rect 429294 286718 429326 286954
rect 429562 286718 429646 286954
rect 429882 286718 429914 286954
rect 429294 286634 429914 286718
rect 429294 286398 429326 286634
rect 429562 286398 429646 286634
rect 429882 286398 429914 286634
rect 429294 250954 429914 286398
rect 429294 250718 429326 250954
rect 429562 250718 429646 250954
rect 429882 250718 429914 250954
rect 429294 250634 429914 250718
rect 429294 250398 429326 250634
rect 429562 250398 429646 250634
rect 429882 250398 429914 250634
rect 429294 214954 429914 250398
rect 429294 214718 429326 214954
rect 429562 214718 429646 214954
rect 429882 214718 429914 214954
rect 429294 214634 429914 214718
rect 429294 214398 429326 214634
rect 429562 214398 429646 214634
rect 429882 214398 429914 214634
rect 429294 178954 429914 214398
rect 429294 178718 429326 178954
rect 429562 178718 429646 178954
rect 429882 178718 429914 178954
rect 429294 178634 429914 178718
rect 429294 178398 429326 178634
rect 429562 178398 429646 178634
rect 429882 178398 429914 178634
rect 429294 142954 429914 178398
rect 429294 142718 429326 142954
rect 429562 142718 429646 142954
rect 429882 142718 429914 142954
rect 429294 142634 429914 142718
rect 429294 142398 429326 142634
rect 429562 142398 429646 142634
rect 429882 142398 429914 142634
rect 429294 106954 429914 142398
rect 429294 106718 429326 106954
rect 429562 106718 429646 106954
rect 429882 106718 429914 106954
rect 429294 106634 429914 106718
rect 429294 106398 429326 106634
rect 429562 106398 429646 106634
rect 429882 106398 429914 106634
rect 429294 70954 429914 106398
rect 429294 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 429914 70954
rect 429294 70634 429914 70718
rect 429294 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 429914 70634
rect 429294 34954 429914 70398
rect 429294 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 429914 34954
rect 429294 34634 429914 34718
rect 429294 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 429914 34634
rect 429294 -7066 429914 34398
rect 429294 -7302 429326 -7066
rect 429562 -7302 429646 -7066
rect 429882 -7302 429914 -7066
rect 429294 -7386 429914 -7302
rect 429294 -7622 429326 -7386
rect 429562 -7622 429646 -7386
rect 429882 -7622 429914 -7386
rect 429294 -7654 429914 -7622
rect 433794 704838 434414 711590
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 147454 434414 182898
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -7654 434414 -902
rect 438294 705798 438914 711590
rect 438294 705562 438326 705798
rect 438562 705562 438646 705798
rect 438882 705562 438914 705798
rect 438294 705478 438914 705562
rect 438294 705242 438326 705478
rect 438562 705242 438646 705478
rect 438882 705242 438914 705478
rect 438294 691954 438914 705242
rect 438294 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 438914 691954
rect 438294 691634 438914 691718
rect 438294 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 438914 691634
rect 438294 655954 438914 691398
rect 438294 655718 438326 655954
rect 438562 655718 438646 655954
rect 438882 655718 438914 655954
rect 438294 655634 438914 655718
rect 438294 655398 438326 655634
rect 438562 655398 438646 655634
rect 438882 655398 438914 655634
rect 438294 619954 438914 655398
rect 438294 619718 438326 619954
rect 438562 619718 438646 619954
rect 438882 619718 438914 619954
rect 438294 619634 438914 619718
rect 438294 619398 438326 619634
rect 438562 619398 438646 619634
rect 438882 619398 438914 619634
rect 438294 583954 438914 619398
rect 438294 583718 438326 583954
rect 438562 583718 438646 583954
rect 438882 583718 438914 583954
rect 438294 583634 438914 583718
rect 438294 583398 438326 583634
rect 438562 583398 438646 583634
rect 438882 583398 438914 583634
rect 438294 547954 438914 583398
rect 438294 547718 438326 547954
rect 438562 547718 438646 547954
rect 438882 547718 438914 547954
rect 438294 547634 438914 547718
rect 438294 547398 438326 547634
rect 438562 547398 438646 547634
rect 438882 547398 438914 547634
rect 438294 511954 438914 547398
rect 438294 511718 438326 511954
rect 438562 511718 438646 511954
rect 438882 511718 438914 511954
rect 438294 511634 438914 511718
rect 438294 511398 438326 511634
rect 438562 511398 438646 511634
rect 438882 511398 438914 511634
rect 438294 475954 438914 511398
rect 438294 475718 438326 475954
rect 438562 475718 438646 475954
rect 438882 475718 438914 475954
rect 438294 475634 438914 475718
rect 438294 475398 438326 475634
rect 438562 475398 438646 475634
rect 438882 475398 438914 475634
rect 438294 439954 438914 475398
rect 438294 439718 438326 439954
rect 438562 439718 438646 439954
rect 438882 439718 438914 439954
rect 438294 439634 438914 439718
rect 438294 439398 438326 439634
rect 438562 439398 438646 439634
rect 438882 439398 438914 439634
rect 438294 403954 438914 439398
rect 438294 403718 438326 403954
rect 438562 403718 438646 403954
rect 438882 403718 438914 403954
rect 438294 403634 438914 403718
rect 438294 403398 438326 403634
rect 438562 403398 438646 403634
rect 438882 403398 438914 403634
rect 438294 367954 438914 403398
rect 438294 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 438914 367954
rect 438294 367634 438914 367718
rect 438294 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 438914 367634
rect 438294 331954 438914 367398
rect 438294 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 438914 331954
rect 438294 331634 438914 331718
rect 438294 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 438914 331634
rect 438294 295954 438914 331398
rect 438294 295718 438326 295954
rect 438562 295718 438646 295954
rect 438882 295718 438914 295954
rect 438294 295634 438914 295718
rect 438294 295398 438326 295634
rect 438562 295398 438646 295634
rect 438882 295398 438914 295634
rect 438294 259954 438914 295398
rect 438294 259718 438326 259954
rect 438562 259718 438646 259954
rect 438882 259718 438914 259954
rect 438294 259634 438914 259718
rect 438294 259398 438326 259634
rect 438562 259398 438646 259634
rect 438882 259398 438914 259634
rect 438294 223954 438914 259398
rect 438294 223718 438326 223954
rect 438562 223718 438646 223954
rect 438882 223718 438914 223954
rect 438294 223634 438914 223718
rect 438294 223398 438326 223634
rect 438562 223398 438646 223634
rect 438882 223398 438914 223634
rect 438294 187954 438914 223398
rect 438294 187718 438326 187954
rect 438562 187718 438646 187954
rect 438882 187718 438914 187954
rect 438294 187634 438914 187718
rect 438294 187398 438326 187634
rect 438562 187398 438646 187634
rect 438882 187398 438914 187634
rect 438294 151954 438914 187398
rect 438294 151718 438326 151954
rect 438562 151718 438646 151954
rect 438882 151718 438914 151954
rect 438294 151634 438914 151718
rect 438294 151398 438326 151634
rect 438562 151398 438646 151634
rect 438882 151398 438914 151634
rect 438294 115954 438914 151398
rect 438294 115718 438326 115954
rect 438562 115718 438646 115954
rect 438882 115718 438914 115954
rect 438294 115634 438914 115718
rect 438294 115398 438326 115634
rect 438562 115398 438646 115634
rect 438882 115398 438914 115634
rect 438294 79954 438914 115398
rect 438294 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 438914 79954
rect 438294 79634 438914 79718
rect 438294 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 438914 79634
rect 438294 43954 438914 79398
rect 438294 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 438914 43954
rect 438294 43634 438914 43718
rect 438294 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 438914 43634
rect 438294 7954 438914 43398
rect 438294 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 438914 7954
rect 438294 7634 438914 7718
rect 438294 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 438914 7634
rect 438294 -1306 438914 7398
rect 438294 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 438914 -1306
rect 438294 -1626 438914 -1542
rect 438294 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 438914 -1626
rect 438294 -7654 438914 -1862
rect 442794 706758 443414 711590
rect 442794 706522 442826 706758
rect 443062 706522 443146 706758
rect 443382 706522 443414 706758
rect 442794 706438 443414 706522
rect 442794 706202 442826 706438
rect 443062 706202 443146 706438
rect 443382 706202 443414 706438
rect 442794 696454 443414 706202
rect 442794 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 443414 696454
rect 442794 696134 443414 696218
rect 442794 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 443414 696134
rect 442794 660454 443414 695898
rect 442794 660218 442826 660454
rect 443062 660218 443146 660454
rect 443382 660218 443414 660454
rect 442794 660134 443414 660218
rect 442794 659898 442826 660134
rect 443062 659898 443146 660134
rect 443382 659898 443414 660134
rect 442794 624454 443414 659898
rect 442794 624218 442826 624454
rect 443062 624218 443146 624454
rect 443382 624218 443414 624454
rect 442794 624134 443414 624218
rect 442794 623898 442826 624134
rect 443062 623898 443146 624134
rect 443382 623898 443414 624134
rect 442794 588454 443414 623898
rect 442794 588218 442826 588454
rect 443062 588218 443146 588454
rect 443382 588218 443414 588454
rect 442794 588134 443414 588218
rect 442794 587898 442826 588134
rect 443062 587898 443146 588134
rect 443382 587898 443414 588134
rect 442794 552454 443414 587898
rect 442794 552218 442826 552454
rect 443062 552218 443146 552454
rect 443382 552218 443414 552454
rect 442794 552134 443414 552218
rect 442794 551898 442826 552134
rect 443062 551898 443146 552134
rect 443382 551898 443414 552134
rect 442794 516454 443414 551898
rect 442794 516218 442826 516454
rect 443062 516218 443146 516454
rect 443382 516218 443414 516454
rect 442794 516134 443414 516218
rect 442794 515898 442826 516134
rect 443062 515898 443146 516134
rect 443382 515898 443414 516134
rect 442794 480454 443414 515898
rect 442794 480218 442826 480454
rect 443062 480218 443146 480454
rect 443382 480218 443414 480454
rect 442794 480134 443414 480218
rect 442794 479898 442826 480134
rect 443062 479898 443146 480134
rect 443382 479898 443414 480134
rect 442794 444454 443414 479898
rect 442794 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 443414 444454
rect 442794 444134 443414 444218
rect 442794 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 443414 444134
rect 442794 408454 443414 443898
rect 442794 408218 442826 408454
rect 443062 408218 443146 408454
rect 443382 408218 443414 408454
rect 442794 408134 443414 408218
rect 442794 407898 442826 408134
rect 443062 407898 443146 408134
rect 443382 407898 443414 408134
rect 442794 372454 443414 407898
rect 442794 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 443414 372454
rect 442794 372134 443414 372218
rect 442794 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 443414 372134
rect 442794 336454 443414 371898
rect 442794 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 443414 336454
rect 442794 336134 443414 336218
rect 442794 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 443414 336134
rect 442794 300454 443414 335898
rect 442794 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 443414 300454
rect 442794 300134 443414 300218
rect 442794 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 443414 300134
rect 442794 264454 443414 299898
rect 442794 264218 442826 264454
rect 443062 264218 443146 264454
rect 443382 264218 443414 264454
rect 442794 264134 443414 264218
rect 442794 263898 442826 264134
rect 443062 263898 443146 264134
rect 443382 263898 443414 264134
rect 442794 228454 443414 263898
rect 442794 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 443414 228454
rect 442794 228134 443414 228218
rect 442794 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 443414 228134
rect 442794 192454 443414 227898
rect 442794 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 443414 192454
rect 442794 192134 443414 192218
rect 442794 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 443414 192134
rect 442794 156454 443414 191898
rect 442794 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 443414 156454
rect 442794 156134 443414 156218
rect 442794 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 443414 156134
rect 442794 120454 443414 155898
rect 442794 120218 442826 120454
rect 443062 120218 443146 120454
rect 443382 120218 443414 120454
rect 442794 120134 443414 120218
rect 442794 119898 442826 120134
rect 443062 119898 443146 120134
rect 443382 119898 443414 120134
rect 442794 84454 443414 119898
rect 442794 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 443414 84454
rect 442794 84134 443414 84218
rect 442794 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 443414 84134
rect 442794 48454 443414 83898
rect 442794 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 443414 48454
rect 442794 48134 443414 48218
rect 442794 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 443414 48134
rect 442794 12454 443414 47898
rect 442794 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 443414 12454
rect 442794 12134 443414 12218
rect 442794 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 443414 12134
rect 442794 -2266 443414 11898
rect 442794 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 443414 -2266
rect 442794 -2586 443414 -2502
rect 442794 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 443414 -2586
rect 442794 -7654 443414 -2822
rect 447294 707718 447914 711590
rect 447294 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 447914 707718
rect 447294 707398 447914 707482
rect 447294 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 447914 707398
rect 447294 700954 447914 707162
rect 447294 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 447914 700954
rect 447294 700634 447914 700718
rect 447294 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 447914 700634
rect 447294 664954 447914 700398
rect 447294 664718 447326 664954
rect 447562 664718 447646 664954
rect 447882 664718 447914 664954
rect 447294 664634 447914 664718
rect 447294 664398 447326 664634
rect 447562 664398 447646 664634
rect 447882 664398 447914 664634
rect 447294 628954 447914 664398
rect 447294 628718 447326 628954
rect 447562 628718 447646 628954
rect 447882 628718 447914 628954
rect 447294 628634 447914 628718
rect 447294 628398 447326 628634
rect 447562 628398 447646 628634
rect 447882 628398 447914 628634
rect 447294 592954 447914 628398
rect 447294 592718 447326 592954
rect 447562 592718 447646 592954
rect 447882 592718 447914 592954
rect 447294 592634 447914 592718
rect 447294 592398 447326 592634
rect 447562 592398 447646 592634
rect 447882 592398 447914 592634
rect 447294 556954 447914 592398
rect 447294 556718 447326 556954
rect 447562 556718 447646 556954
rect 447882 556718 447914 556954
rect 447294 556634 447914 556718
rect 447294 556398 447326 556634
rect 447562 556398 447646 556634
rect 447882 556398 447914 556634
rect 447294 520954 447914 556398
rect 447294 520718 447326 520954
rect 447562 520718 447646 520954
rect 447882 520718 447914 520954
rect 447294 520634 447914 520718
rect 447294 520398 447326 520634
rect 447562 520398 447646 520634
rect 447882 520398 447914 520634
rect 447294 484954 447914 520398
rect 447294 484718 447326 484954
rect 447562 484718 447646 484954
rect 447882 484718 447914 484954
rect 447294 484634 447914 484718
rect 447294 484398 447326 484634
rect 447562 484398 447646 484634
rect 447882 484398 447914 484634
rect 447294 448954 447914 484398
rect 447294 448718 447326 448954
rect 447562 448718 447646 448954
rect 447882 448718 447914 448954
rect 447294 448634 447914 448718
rect 447294 448398 447326 448634
rect 447562 448398 447646 448634
rect 447882 448398 447914 448634
rect 447294 412954 447914 448398
rect 447294 412718 447326 412954
rect 447562 412718 447646 412954
rect 447882 412718 447914 412954
rect 447294 412634 447914 412718
rect 447294 412398 447326 412634
rect 447562 412398 447646 412634
rect 447882 412398 447914 412634
rect 447294 376954 447914 412398
rect 447294 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 447914 376954
rect 447294 376634 447914 376718
rect 447294 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 447914 376634
rect 447294 340954 447914 376398
rect 447294 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 447914 340954
rect 447294 340634 447914 340718
rect 447294 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 447914 340634
rect 447294 304954 447914 340398
rect 447294 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 447914 304954
rect 447294 304634 447914 304718
rect 447294 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 447914 304634
rect 447294 268954 447914 304398
rect 447294 268718 447326 268954
rect 447562 268718 447646 268954
rect 447882 268718 447914 268954
rect 447294 268634 447914 268718
rect 447294 268398 447326 268634
rect 447562 268398 447646 268634
rect 447882 268398 447914 268634
rect 447294 232954 447914 268398
rect 447294 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 447914 232954
rect 447294 232634 447914 232718
rect 447294 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 447914 232634
rect 447294 196954 447914 232398
rect 447294 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 447914 196954
rect 447294 196634 447914 196718
rect 447294 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 447914 196634
rect 447294 160954 447914 196398
rect 447294 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 447914 160954
rect 447294 160634 447914 160718
rect 447294 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 447914 160634
rect 447294 124954 447914 160398
rect 447294 124718 447326 124954
rect 447562 124718 447646 124954
rect 447882 124718 447914 124954
rect 447294 124634 447914 124718
rect 447294 124398 447326 124634
rect 447562 124398 447646 124634
rect 447882 124398 447914 124634
rect 447294 88954 447914 124398
rect 447294 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 447914 88954
rect 447294 88634 447914 88718
rect 447294 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 447914 88634
rect 447294 52954 447914 88398
rect 447294 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 447914 52954
rect 447294 52634 447914 52718
rect 447294 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 447914 52634
rect 447294 16954 447914 52398
rect 447294 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 447914 16954
rect 447294 16634 447914 16718
rect 447294 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 447914 16634
rect 447294 -3226 447914 16398
rect 447294 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 447914 -3226
rect 447294 -3546 447914 -3462
rect 447294 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 447914 -3546
rect 447294 -7654 447914 -3782
rect 451794 708678 452414 711590
rect 451794 708442 451826 708678
rect 452062 708442 452146 708678
rect 452382 708442 452414 708678
rect 451794 708358 452414 708442
rect 451794 708122 451826 708358
rect 452062 708122 452146 708358
rect 452382 708122 452414 708358
rect 451794 669454 452414 708122
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 451794 309454 452414 344898
rect 451794 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 452414 309454
rect 451794 309134 452414 309218
rect 451794 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 452414 309134
rect 451794 273454 452414 308898
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 129454 452414 164898
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -4186 452414 20898
rect 451794 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 452414 -4186
rect 451794 -4506 452414 -4422
rect 451794 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 452414 -4506
rect 451794 -7654 452414 -4742
rect 456294 709638 456914 711590
rect 456294 709402 456326 709638
rect 456562 709402 456646 709638
rect 456882 709402 456914 709638
rect 456294 709318 456914 709402
rect 456294 709082 456326 709318
rect 456562 709082 456646 709318
rect 456882 709082 456914 709318
rect 456294 673954 456914 709082
rect 456294 673718 456326 673954
rect 456562 673718 456646 673954
rect 456882 673718 456914 673954
rect 456294 673634 456914 673718
rect 456294 673398 456326 673634
rect 456562 673398 456646 673634
rect 456882 673398 456914 673634
rect 456294 637954 456914 673398
rect 456294 637718 456326 637954
rect 456562 637718 456646 637954
rect 456882 637718 456914 637954
rect 456294 637634 456914 637718
rect 456294 637398 456326 637634
rect 456562 637398 456646 637634
rect 456882 637398 456914 637634
rect 456294 601954 456914 637398
rect 456294 601718 456326 601954
rect 456562 601718 456646 601954
rect 456882 601718 456914 601954
rect 456294 601634 456914 601718
rect 456294 601398 456326 601634
rect 456562 601398 456646 601634
rect 456882 601398 456914 601634
rect 456294 565954 456914 601398
rect 456294 565718 456326 565954
rect 456562 565718 456646 565954
rect 456882 565718 456914 565954
rect 456294 565634 456914 565718
rect 456294 565398 456326 565634
rect 456562 565398 456646 565634
rect 456882 565398 456914 565634
rect 456294 529954 456914 565398
rect 456294 529718 456326 529954
rect 456562 529718 456646 529954
rect 456882 529718 456914 529954
rect 456294 529634 456914 529718
rect 456294 529398 456326 529634
rect 456562 529398 456646 529634
rect 456882 529398 456914 529634
rect 456294 493954 456914 529398
rect 456294 493718 456326 493954
rect 456562 493718 456646 493954
rect 456882 493718 456914 493954
rect 456294 493634 456914 493718
rect 456294 493398 456326 493634
rect 456562 493398 456646 493634
rect 456882 493398 456914 493634
rect 456294 457954 456914 493398
rect 456294 457718 456326 457954
rect 456562 457718 456646 457954
rect 456882 457718 456914 457954
rect 456294 457634 456914 457718
rect 456294 457398 456326 457634
rect 456562 457398 456646 457634
rect 456882 457398 456914 457634
rect 456294 421954 456914 457398
rect 456294 421718 456326 421954
rect 456562 421718 456646 421954
rect 456882 421718 456914 421954
rect 456294 421634 456914 421718
rect 456294 421398 456326 421634
rect 456562 421398 456646 421634
rect 456882 421398 456914 421634
rect 456294 385954 456914 421398
rect 456294 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 456914 385954
rect 456294 385634 456914 385718
rect 456294 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 456914 385634
rect 456294 349954 456914 385398
rect 456294 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 456914 349954
rect 456294 349634 456914 349718
rect 456294 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 456914 349634
rect 456294 313954 456914 349398
rect 456294 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 456914 313954
rect 456294 313634 456914 313718
rect 456294 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 456914 313634
rect 456294 277954 456914 313398
rect 456294 277718 456326 277954
rect 456562 277718 456646 277954
rect 456882 277718 456914 277954
rect 456294 277634 456914 277718
rect 456294 277398 456326 277634
rect 456562 277398 456646 277634
rect 456882 277398 456914 277634
rect 456294 241954 456914 277398
rect 456294 241718 456326 241954
rect 456562 241718 456646 241954
rect 456882 241718 456914 241954
rect 456294 241634 456914 241718
rect 456294 241398 456326 241634
rect 456562 241398 456646 241634
rect 456882 241398 456914 241634
rect 456294 205954 456914 241398
rect 456294 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 456914 205954
rect 456294 205634 456914 205718
rect 456294 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 456914 205634
rect 456294 169954 456914 205398
rect 456294 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 456914 169954
rect 456294 169634 456914 169718
rect 456294 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 456914 169634
rect 456294 133954 456914 169398
rect 456294 133718 456326 133954
rect 456562 133718 456646 133954
rect 456882 133718 456914 133954
rect 456294 133634 456914 133718
rect 456294 133398 456326 133634
rect 456562 133398 456646 133634
rect 456882 133398 456914 133634
rect 456294 97954 456914 133398
rect 456294 97718 456326 97954
rect 456562 97718 456646 97954
rect 456882 97718 456914 97954
rect 456294 97634 456914 97718
rect 456294 97398 456326 97634
rect 456562 97398 456646 97634
rect 456882 97398 456914 97634
rect 456294 61954 456914 97398
rect 456294 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 456914 61954
rect 456294 61634 456914 61718
rect 456294 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 456914 61634
rect 456294 25954 456914 61398
rect 456294 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 456914 25954
rect 456294 25634 456914 25718
rect 456294 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 456914 25634
rect 456294 -5146 456914 25398
rect 456294 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 456914 -5146
rect 456294 -5466 456914 -5382
rect 456294 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 456914 -5466
rect 456294 -7654 456914 -5702
rect 460794 710598 461414 711590
rect 460794 710362 460826 710598
rect 461062 710362 461146 710598
rect 461382 710362 461414 710598
rect 460794 710278 461414 710362
rect 460794 710042 460826 710278
rect 461062 710042 461146 710278
rect 461382 710042 461414 710278
rect 460794 678454 461414 710042
rect 460794 678218 460826 678454
rect 461062 678218 461146 678454
rect 461382 678218 461414 678454
rect 460794 678134 461414 678218
rect 460794 677898 460826 678134
rect 461062 677898 461146 678134
rect 461382 677898 461414 678134
rect 460794 642454 461414 677898
rect 460794 642218 460826 642454
rect 461062 642218 461146 642454
rect 461382 642218 461414 642454
rect 460794 642134 461414 642218
rect 460794 641898 460826 642134
rect 461062 641898 461146 642134
rect 461382 641898 461414 642134
rect 460794 606454 461414 641898
rect 460794 606218 460826 606454
rect 461062 606218 461146 606454
rect 461382 606218 461414 606454
rect 460794 606134 461414 606218
rect 460794 605898 460826 606134
rect 461062 605898 461146 606134
rect 461382 605898 461414 606134
rect 460794 570454 461414 605898
rect 460794 570218 460826 570454
rect 461062 570218 461146 570454
rect 461382 570218 461414 570454
rect 460794 570134 461414 570218
rect 460794 569898 460826 570134
rect 461062 569898 461146 570134
rect 461382 569898 461414 570134
rect 460794 534454 461414 569898
rect 460794 534218 460826 534454
rect 461062 534218 461146 534454
rect 461382 534218 461414 534454
rect 460794 534134 461414 534218
rect 460794 533898 460826 534134
rect 461062 533898 461146 534134
rect 461382 533898 461414 534134
rect 460794 498454 461414 533898
rect 460794 498218 460826 498454
rect 461062 498218 461146 498454
rect 461382 498218 461414 498454
rect 460794 498134 461414 498218
rect 460794 497898 460826 498134
rect 461062 497898 461146 498134
rect 461382 497898 461414 498134
rect 460794 462454 461414 497898
rect 460794 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 461414 462454
rect 460794 462134 461414 462218
rect 460794 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 461414 462134
rect 460794 426454 461414 461898
rect 460794 426218 460826 426454
rect 461062 426218 461146 426454
rect 461382 426218 461414 426454
rect 460794 426134 461414 426218
rect 460794 425898 460826 426134
rect 461062 425898 461146 426134
rect 461382 425898 461414 426134
rect 460794 390454 461414 425898
rect 460794 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 461414 390454
rect 460794 390134 461414 390218
rect 460794 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 461414 390134
rect 460794 354454 461414 389898
rect 460794 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 461414 354454
rect 460794 354134 461414 354218
rect 460794 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 461414 354134
rect 460794 318454 461414 353898
rect 460794 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 461414 318454
rect 460794 318134 461414 318218
rect 460794 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 461414 318134
rect 460794 282454 461414 317898
rect 460794 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 461414 282454
rect 460794 282134 461414 282218
rect 460794 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 461414 282134
rect 460794 246454 461414 281898
rect 460794 246218 460826 246454
rect 461062 246218 461146 246454
rect 461382 246218 461414 246454
rect 460794 246134 461414 246218
rect 460794 245898 460826 246134
rect 461062 245898 461146 246134
rect 461382 245898 461414 246134
rect 460794 210454 461414 245898
rect 460794 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 461414 210454
rect 460794 210134 461414 210218
rect 460794 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 461414 210134
rect 460794 174454 461414 209898
rect 460794 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 461414 174454
rect 460794 174134 461414 174218
rect 460794 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 461414 174134
rect 460794 138454 461414 173898
rect 460794 138218 460826 138454
rect 461062 138218 461146 138454
rect 461382 138218 461414 138454
rect 460794 138134 461414 138218
rect 460794 137898 460826 138134
rect 461062 137898 461146 138134
rect 461382 137898 461414 138134
rect 460794 102454 461414 137898
rect 460794 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 461414 102454
rect 460794 102134 461414 102218
rect 460794 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 461414 102134
rect 460794 66454 461414 101898
rect 460794 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 461414 66454
rect 460794 66134 461414 66218
rect 460794 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 461414 66134
rect 460794 30454 461414 65898
rect 460794 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 461414 30454
rect 460794 30134 461414 30218
rect 460794 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 461414 30134
rect 460794 -6106 461414 29898
rect 460794 -6342 460826 -6106
rect 461062 -6342 461146 -6106
rect 461382 -6342 461414 -6106
rect 460794 -6426 461414 -6342
rect 460794 -6662 460826 -6426
rect 461062 -6662 461146 -6426
rect 461382 -6662 461414 -6426
rect 460794 -7654 461414 -6662
rect 465294 711558 465914 711590
rect 465294 711322 465326 711558
rect 465562 711322 465646 711558
rect 465882 711322 465914 711558
rect 465294 711238 465914 711322
rect 465294 711002 465326 711238
rect 465562 711002 465646 711238
rect 465882 711002 465914 711238
rect 465294 682954 465914 711002
rect 465294 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 465914 682954
rect 465294 682634 465914 682718
rect 465294 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 465914 682634
rect 465294 646954 465914 682398
rect 465294 646718 465326 646954
rect 465562 646718 465646 646954
rect 465882 646718 465914 646954
rect 465294 646634 465914 646718
rect 465294 646398 465326 646634
rect 465562 646398 465646 646634
rect 465882 646398 465914 646634
rect 465294 610954 465914 646398
rect 465294 610718 465326 610954
rect 465562 610718 465646 610954
rect 465882 610718 465914 610954
rect 465294 610634 465914 610718
rect 465294 610398 465326 610634
rect 465562 610398 465646 610634
rect 465882 610398 465914 610634
rect 465294 574954 465914 610398
rect 465294 574718 465326 574954
rect 465562 574718 465646 574954
rect 465882 574718 465914 574954
rect 465294 574634 465914 574718
rect 465294 574398 465326 574634
rect 465562 574398 465646 574634
rect 465882 574398 465914 574634
rect 465294 538954 465914 574398
rect 465294 538718 465326 538954
rect 465562 538718 465646 538954
rect 465882 538718 465914 538954
rect 465294 538634 465914 538718
rect 465294 538398 465326 538634
rect 465562 538398 465646 538634
rect 465882 538398 465914 538634
rect 465294 502954 465914 538398
rect 465294 502718 465326 502954
rect 465562 502718 465646 502954
rect 465882 502718 465914 502954
rect 465294 502634 465914 502718
rect 465294 502398 465326 502634
rect 465562 502398 465646 502634
rect 465882 502398 465914 502634
rect 465294 466954 465914 502398
rect 465294 466718 465326 466954
rect 465562 466718 465646 466954
rect 465882 466718 465914 466954
rect 465294 466634 465914 466718
rect 465294 466398 465326 466634
rect 465562 466398 465646 466634
rect 465882 466398 465914 466634
rect 465294 430954 465914 466398
rect 465294 430718 465326 430954
rect 465562 430718 465646 430954
rect 465882 430718 465914 430954
rect 465294 430634 465914 430718
rect 465294 430398 465326 430634
rect 465562 430398 465646 430634
rect 465882 430398 465914 430634
rect 465294 394954 465914 430398
rect 465294 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 465914 394954
rect 465294 394634 465914 394718
rect 465294 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 465914 394634
rect 465294 358954 465914 394398
rect 465294 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 465914 358954
rect 465294 358634 465914 358718
rect 465294 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 465914 358634
rect 465294 322954 465914 358398
rect 465294 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 465914 322954
rect 465294 322634 465914 322718
rect 465294 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 465914 322634
rect 465294 286954 465914 322398
rect 465294 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 465914 286954
rect 465294 286634 465914 286718
rect 465294 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 465914 286634
rect 465294 250954 465914 286398
rect 465294 250718 465326 250954
rect 465562 250718 465646 250954
rect 465882 250718 465914 250954
rect 465294 250634 465914 250718
rect 465294 250398 465326 250634
rect 465562 250398 465646 250634
rect 465882 250398 465914 250634
rect 465294 214954 465914 250398
rect 465294 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 465914 214954
rect 465294 214634 465914 214718
rect 465294 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 465914 214634
rect 465294 178954 465914 214398
rect 465294 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 465914 178954
rect 465294 178634 465914 178718
rect 465294 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 465914 178634
rect 465294 142954 465914 178398
rect 465294 142718 465326 142954
rect 465562 142718 465646 142954
rect 465882 142718 465914 142954
rect 465294 142634 465914 142718
rect 465294 142398 465326 142634
rect 465562 142398 465646 142634
rect 465882 142398 465914 142634
rect 465294 106954 465914 142398
rect 465294 106718 465326 106954
rect 465562 106718 465646 106954
rect 465882 106718 465914 106954
rect 465294 106634 465914 106718
rect 465294 106398 465326 106634
rect 465562 106398 465646 106634
rect 465882 106398 465914 106634
rect 465294 70954 465914 106398
rect 465294 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 465914 70954
rect 465294 70634 465914 70718
rect 465294 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 465914 70634
rect 465294 34954 465914 70398
rect 465294 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 465914 34954
rect 465294 34634 465914 34718
rect 465294 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 465914 34634
rect 465294 -7066 465914 34398
rect 465294 -7302 465326 -7066
rect 465562 -7302 465646 -7066
rect 465882 -7302 465914 -7066
rect 465294 -7386 465914 -7302
rect 465294 -7622 465326 -7386
rect 465562 -7622 465646 -7386
rect 465882 -7622 465914 -7386
rect 465294 -7654 465914 -7622
rect 469794 704838 470414 711590
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -7654 470414 -902
rect 474294 705798 474914 711590
rect 474294 705562 474326 705798
rect 474562 705562 474646 705798
rect 474882 705562 474914 705798
rect 474294 705478 474914 705562
rect 474294 705242 474326 705478
rect 474562 705242 474646 705478
rect 474882 705242 474914 705478
rect 474294 691954 474914 705242
rect 474294 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 474914 691954
rect 474294 691634 474914 691718
rect 474294 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 474914 691634
rect 474294 655954 474914 691398
rect 474294 655718 474326 655954
rect 474562 655718 474646 655954
rect 474882 655718 474914 655954
rect 474294 655634 474914 655718
rect 474294 655398 474326 655634
rect 474562 655398 474646 655634
rect 474882 655398 474914 655634
rect 474294 619954 474914 655398
rect 474294 619718 474326 619954
rect 474562 619718 474646 619954
rect 474882 619718 474914 619954
rect 474294 619634 474914 619718
rect 474294 619398 474326 619634
rect 474562 619398 474646 619634
rect 474882 619398 474914 619634
rect 474294 583954 474914 619398
rect 474294 583718 474326 583954
rect 474562 583718 474646 583954
rect 474882 583718 474914 583954
rect 474294 583634 474914 583718
rect 474294 583398 474326 583634
rect 474562 583398 474646 583634
rect 474882 583398 474914 583634
rect 474294 547954 474914 583398
rect 474294 547718 474326 547954
rect 474562 547718 474646 547954
rect 474882 547718 474914 547954
rect 474294 547634 474914 547718
rect 474294 547398 474326 547634
rect 474562 547398 474646 547634
rect 474882 547398 474914 547634
rect 474294 511954 474914 547398
rect 474294 511718 474326 511954
rect 474562 511718 474646 511954
rect 474882 511718 474914 511954
rect 474294 511634 474914 511718
rect 474294 511398 474326 511634
rect 474562 511398 474646 511634
rect 474882 511398 474914 511634
rect 474294 475954 474914 511398
rect 474294 475718 474326 475954
rect 474562 475718 474646 475954
rect 474882 475718 474914 475954
rect 474294 475634 474914 475718
rect 474294 475398 474326 475634
rect 474562 475398 474646 475634
rect 474882 475398 474914 475634
rect 474294 439954 474914 475398
rect 474294 439718 474326 439954
rect 474562 439718 474646 439954
rect 474882 439718 474914 439954
rect 474294 439634 474914 439718
rect 474294 439398 474326 439634
rect 474562 439398 474646 439634
rect 474882 439398 474914 439634
rect 474294 403954 474914 439398
rect 474294 403718 474326 403954
rect 474562 403718 474646 403954
rect 474882 403718 474914 403954
rect 474294 403634 474914 403718
rect 474294 403398 474326 403634
rect 474562 403398 474646 403634
rect 474882 403398 474914 403634
rect 474294 367954 474914 403398
rect 474294 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 474914 367954
rect 474294 367634 474914 367718
rect 474294 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 474914 367634
rect 474294 331954 474914 367398
rect 474294 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 474914 331954
rect 474294 331634 474914 331718
rect 474294 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 474914 331634
rect 474294 295954 474914 331398
rect 474294 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 474914 295954
rect 474294 295634 474914 295718
rect 474294 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 474914 295634
rect 474294 259954 474914 295398
rect 474294 259718 474326 259954
rect 474562 259718 474646 259954
rect 474882 259718 474914 259954
rect 474294 259634 474914 259718
rect 474294 259398 474326 259634
rect 474562 259398 474646 259634
rect 474882 259398 474914 259634
rect 474294 223954 474914 259398
rect 474294 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 474914 223954
rect 474294 223634 474914 223718
rect 474294 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 474914 223634
rect 474294 187954 474914 223398
rect 474294 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 474914 187954
rect 474294 187634 474914 187718
rect 474294 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 474914 187634
rect 474294 151954 474914 187398
rect 474294 151718 474326 151954
rect 474562 151718 474646 151954
rect 474882 151718 474914 151954
rect 474294 151634 474914 151718
rect 474294 151398 474326 151634
rect 474562 151398 474646 151634
rect 474882 151398 474914 151634
rect 474294 115954 474914 151398
rect 474294 115718 474326 115954
rect 474562 115718 474646 115954
rect 474882 115718 474914 115954
rect 474294 115634 474914 115718
rect 474294 115398 474326 115634
rect 474562 115398 474646 115634
rect 474882 115398 474914 115634
rect 474294 79954 474914 115398
rect 474294 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 474914 79954
rect 474294 79634 474914 79718
rect 474294 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 474914 79634
rect 474294 43954 474914 79398
rect 474294 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 474914 43954
rect 474294 43634 474914 43718
rect 474294 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 474914 43634
rect 474294 7954 474914 43398
rect 474294 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 474914 7954
rect 474294 7634 474914 7718
rect 474294 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 474914 7634
rect 474294 -1306 474914 7398
rect 474294 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 474914 -1306
rect 474294 -1626 474914 -1542
rect 474294 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 474914 -1626
rect 474294 -7654 474914 -1862
rect 478794 706758 479414 711590
rect 478794 706522 478826 706758
rect 479062 706522 479146 706758
rect 479382 706522 479414 706758
rect 478794 706438 479414 706522
rect 478794 706202 478826 706438
rect 479062 706202 479146 706438
rect 479382 706202 479414 706438
rect 478794 696454 479414 706202
rect 478794 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 479414 696454
rect 478794 696134 479414 696218
rect 478794 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 479414 696134
rect 478794 660454 479414 695898
rect 478794 660218 478826 660454
rect 479062 660218 479146 660454
rect 479382 660218 479414 660454
rect 478794 660134 479414 660218
rect 478794 659898 478826 660134
rect 479062 659898 479146 660134
rect 479382 659898 479414 660134
rect 478794 624454 479414 659898
rect 478794 624218 478826 624454
rect 479062 624218 479146 624454
rect 479382 624218 479414 624454
rect 478794 624134 479414 624218
rect 478794 623898 478826 624134
rect 479062 623898 479146 624134
rect 479382 623898 479414 624134
rect 478794 588454 479414 623898
rect 478794 588218 478826 588454
rect 479062 588218 479146 588454
rect 479382 588218 479414 588454
rect 478794 588134 479414 588218
rect 478794 587898 478826 588134
rect 479062 587898 479146 588134
rect 479382 587898 479414 588134
rect 478794 552454 479414 587898
rect 478794 552218 478826 552454
rect 479062 552218 479146 552454
rect 479382 552218 479414 552454
rect 478794 552134 479414 552218
rect 478794 551898 478826 552134
rect 479062 551898 479146 552134
rect 479382 551898 479414 552134
rect 478794 516454 479414 551898
rect 478794 516218 478826 516454
rect 479062 516218 479146 516454
rect 479382 516218 479414 516454
rect 478794 516134 479414 516218
rect 478794 515898 478826 516134
rect 479062 515898 479146 516134
rect 479382 515898 479414 516134
rect 478794 480454 479414 515898
rect 478794 480218 478826 480454
rect 479062 480218 479146 480454
rect 479382 480218 479414 480454
rect 478794 480134 479414 480218
rect 478794 479898 478826 480134
rect 479062 479898 479146 480134
rect 479382 479898 479414 480134
rect 478794 444454 479414 479898
rect 478794 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 479414 444454
rect 478794 444134 479414 444218
rect 478794 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 479414 444134
rect 478794 408454 479414 443898
rect 478794 408218 478826 408454
rect 479062 408218 479146 408454
rect 479382 408218 479414 408454
rect 478794 408134 479414 408218
rect 478794 407898 478826 408134
rect 479062 407898 479146 408134
rect 479382 407898 479414 408134
rect 478794 372454 479414 407898
rect 478794 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 479414 372454
rect 478794 372134 479414 372218
rect 478794 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 479414 372134
rect 478794 336454 479414 371898
rect 478794 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 479414 336454
rect 478794 336134 479414 336218
rect 478794 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 479414 336134
rect 478794 300454 479414 335898
rect 478794 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 479414 300454
rect 478794 300134 479414 300218
rect 478794 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 479414 300134
rect 478794 264454 479414 299898
rect 478794 264218 478826 264454
rect 479062 264218 479146 264454
rect 479382 264218 479414 264454
rect 478794 264134 479414 264218
rect 478794 263898 478826 264134
rect 479062 263898 479146 264134
rect 479382 263898 479414 264134
rect 478794 228454 479414 263898
rect 478794 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 479414 228454
rect 478794 228134 479414 228218
rect 478794 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 479414 228134
rect 478794 192454 479414 227898
rect 478794 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 479414 192454
rect 478794 192134 479414 192218
rect 478794 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 479414 192134
rect 478794 156454 479414 191898
rect 478794 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 479414 156454
rect 478794 156134 479414 156218
rect 478794 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 479414 156134
rect 478794 120454 479414 155898
rect 478794 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 479414 120454
rect 478794 120134 479414 120218
rect 478794 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 479414 120134
rect 478794 84454 479414 119898
rect 478794 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 479414 84454
rect 478794 84134 479414 84218
rect 478794 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 479414 84134
rect 478794 48454 479414 83898
rect 478794 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 479414 48454
rect 478794 48134 479414 48218
rect 478794 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 479414 48134
rect 478794 12454 479414 47898
rect 478794 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 479414 12454
rect 478794 12134 479414 12218
rect 478794 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 479414 12134
rect 478794 -2266 479414 11898
rect 478794 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 479414 -2266
rect 478794 -2586 479414 -2502
rect 478794 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 479414 -2586
rect 478794 -7654 479414 -2822
rect 483294 707718 483914 711590
rect 483294 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 483914 707718
rect 483294 707398 483914 707482
rect 483294 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 483914 707398
rect 483294 700954 483914 707162
rect 483294 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 483914 700954
rect 483294 700634 483914 700718
rect 483294 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 483914 700634
rect 483294 664954 483914 700398
rect 483294 664718 483326 664954
rect 483562 664718 483646 664954
rect 483882 664718 483914 664954
rect 483294 664634 483914 664718
rect 483294 664398 483326 664634
rect 483562 664398 483646 664634
rect 483882 664398 483914 664634
rect 483294 628954 483914 664398
rect 483294 628718 483326 628954
rect 483562 628718 483646 628954
rect 483882 628718 483914 628954
rect 483294 628634 483914 628718
rect 483294 628398 483326 628634
rect 483562 628398 483646 628634
rect 483882 628398 483914 628634
rect 483294 592954 483914 628398
rect 483294 592718 483326 592954
rect 483562 592718 483646 592954
rect 483882 592718 483914 592954
rect 483294 592634 483914 592718
rect 483294 592398 483326 592634
rect 483562 592398 483646 592634
rect 483882 592398 483914 592634
rect 483294 556954 483914 592398
rect 483294 556718 483326 556954
rect 483562 556718 483646 556954
rect 483882 556718 483914 556954
rect 483294 556634 483914 556718
rect 483294 556398 483326 556634
rect 483562 556398 483646 556634
rect 483882 556398 483914 556634
rect 483294 520954 483914 556398
rect 483294 520718 483326 520954
rect 483562 520718 483646 520954
rect 483882 520718 483914 520954
rect 483294 520634 483914 520718
rect 483294 520398 483326 520634
rect 483562 520398 483646 520634
rect 483882 520398 483914 520634
rect 483294 484954 483914 520398
rect 483294 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 483914 484954
rect 483294 484634 483914 484718
rect 483294 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 483914 484634
rect 483294 448954 483914 484398
rect 483294 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 483914 448954
rect 483294 448634 483914 448718
rect 483294 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 483914 448634
rect 483294 412954 483914 448398
rect 483294 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 483914 412954
rect 483294 412634 483914 412718
rect 483294 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 483914 412634
rect 483294 376954 483914 412398
rect 483294 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 483914 376954
rect 483294 376634 483914 376718
rect 483294 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 483914 376634
rect 483294 340954 483914 376398
rect 483294 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 483914 340954
rect 483294 340634 483914 340718
rect 483294 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 483914 340634
rect 483294 304954 483914 340398
rect 483294 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 483914 304954
rect 483294 304634 483914 304718
rect 483294 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 483914 304634
rect 483294 268954 483914 304398
rect 483294 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 483914 268954
rect 483294 268634 483914 268718
rect 483294 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 483914 268634
rect 483294 232954 483914 268398
rect 483294 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 483914 232954
rect 483294 232634 483914 232718
rect 483294 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 483914 232634
rect 483294 196954 483914 232398
rect 483294 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 483914 196954
rect 483294 196634 483914 196718
rect 483294 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 483914 196634
rect 483294 160954 483914 196398
rect 483294 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 483914 160954
rect 483294 160634 483914 160718
rect 483294 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 483914 160634
rect 483294 124954 483914 160398
rect 483294 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 483914 124954
rect 483294 124634 483914 124718
rect 483294 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 483914 124634
rect 483294 88954 483914 124398
rect 483294 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 483914 88954
rect 483294 88634 483914 88718
rect 483294 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 483914 88634
rect 483294 52954 483914 88398
rect 483294 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 483914 52954
rect 483294 52634 483914 52718
rect 483294 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 483914 52634
rect 483294 16954 483914 52398
rect 483294 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 483914 16954
rect 483294 16634 483914 16718
rect 483294 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 483914 16634
rect 483294 -3226 483914 16398
rect 483294 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 483914 -3226
rect 483294 -3546 483914 -3462
rect 483294 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 483914 -3546
rect 483294 -7654 483914 -3782
rect 487794 708678 488414 711590
rect 487794 708442 487826 708678
rect 488062 708442 488146 708678
rect 488382 708442 488414 708678
rect 487794 708358 488414 708442
rect 487794 708122 487826 708358
rect 488062 708122 488146 708358
rect 488382 708122 488414 708358
rect 487794 669454 488414 708122
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -4186 488414 20898
rect 487794 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 488414 -4186
rect 487794 -4506 488414 -4422
rect 487794 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 488414 -4506
rect 487794 -7654 488414 -4742
rect 492294 709638 492914 711590
rect 492294 709402 492326 709638
rect 492562 709402 492646 709638
rect 492882 709402 492914 709638
rect 492294 709318 492914 709402
rect 492294 709082 492326 709318
rect 492562 709082 492646 709318
rect 492882 709082 492914 709318
rect 492294 673954 492914 709082
rect 492294 673718 492326 673954
rect 492562 673718 492646 673954
rect 492882 673718 492914 673954
rect 492294 673634 492914 673718
rect 492294 673398 492326 673634
rect 492562 673398 492646 673634
rect 492882 673398 492914 673634
rect 492294 637954 492914 673398
rect 492294 637718 492326 637954
rect 492562 637718 492646 637954
rect 492882 637718 492914 637954
rect 492294 637634 492914 637718
rect 492294 637398 492326 637634
rect 492562 637398 492646 637634
rect 492882 637398 492914 637634
rect 492294 601954 492914 637398
rect 492294 601718 492326 601954
rect 492562 601718 492646 601954
rect 492882 601718 492914 601954
rect 492294 601634 492914 601718
rect 492294 601398 492326 601634
rect 492562 601398 492646 601634
rect 492882 601398 492914 601634
rect 492294 565954 492914 601398
rect 492294 565718 492326 565954
rect 492562 565718 492646 565954
rect 492882 565718 492914 565954
rect 492294 565634 492914 565718
rect 492294 565398 492326 565634
rect 492562 565398 492646 565634
rect 492882 565398 492914 565634
rect 492294 529954 492914 565398
rect 492294 529718 492326 529954
rect 492562 529718 492646 529954
rect 492882 529718 492914 529954
rect 492294 529634 492914 529718
rect 492294 529398 492326 529634
rect 492562 529398 492646 529634
rect 492882 529398 492914 529634
rect 492294 493954 492914 529398
rect 492294 493718 492326 493954
rect 492562 493718 492646 493954
rect 492882 493718 492914 493954
rect 492294 493634 492914 493718
rect 492294 493398 492326 493634
rect 492562 493398 492646 493634
rect 492882 493398 492914 493634
rect 492294 457954 492914 493398
rect 492294 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 492914 457954
rect 492294 457634 492914 457718
rect 492294 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 492914 457634
rect 492294 421954 492914 457398
rect 492294 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 492914 421954
rect 492294 421634 492914 421718
rect 492294 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 492914 421634
rect 492294 385954 492914 421398
rect 492294 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 492914 385954
rect 492294 385634 492914 385718
rect 492294 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 492914 385634
rect 492294 349954 492914 385398
rect 492294 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 492914 349954
rect 492294 349634 492914 349718
rect 492294 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 492914 349634
rect 492294 313954 492914 349398
rect 492294 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 492914 313954
rect 492294 313634 492914 313718
rect 492294 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 492914 313634
rect 492294 277954 492914 313398
rect 492294 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 492914 277954
rect 492294 277634 492914 277718
rect 492294 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 492914 277634
rect 492294 241954 492914 277398
rect 492294 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 492914 241954
rect 492294 241634 492914 241718
rect 492294 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 492914 241634
rect 492294 205954 492914 241398
rect 492294 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 492914 205954
rect 492294 205634 492914 205718
rect 492294 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 492914 205634
rect 492294 169954 492914 205398
rect 492294 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 492914 169954
rect 492294 169634 492914 169718
rect 492294 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 492914 169634
rect 492294 133954 492914 169398
rect 492294 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 492914 133954
rect 492294 133634 492914 133718
rect 492294 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 492914 133634
rect 492294 97954 492914 133398
rect 492294 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 492914 97954
rect 492294 97634 492914 97718
rect 492294 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 492914 97634
rect 492294 61954 492914 97398
rect 492294 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 492914 61954
rect 492294 61634 492914 61718
rect 492294 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 492914 61634
rect 492294 25954 492914 61398
rect 492294 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 492914 25954
rect 492294 25634 492914 25718
rect 492294 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 492914 25634
rect 492294 -5146 492914 25398
rect 492294 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 492914 -5146
rect 492294 -5466 492914 -5382
rect 492294 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 492914 -5466
rect 492294 -7654 492914 -5702
rect 496794 710598 497414 711590
rect 496794 710362 496826 710598
rect 497062 710362 497146 710598
rect 497382 710362 497414 710598
rect 496794 710278 497414 710362
rect 496794 710042 496826 710278
rect 497062 710042 497146 710278
rect 497382 710042 497414 710278
rect 496794 678454 497414 710042
rect 496794 678218 496826 678454
rect 497062 678218 497146 678454
rect 497382 678218 497414 678454
rect 496794 678134 497414 678218
rect 496794 677898 496826 678134
rect 497062 677898 497146 678134
rect 497382 677898 497414 678134
rect 496794 642454 497414 677898
rect 496794 642218 496826 642454
rect 497062 642218 497146 642454
rect 497382 642218 497414 642454
rect 496794 642134 497414 642218
rect 496794 641898 496826 642134
rect 497062 641898 497146 642134
rect 497382 641898 497414 642134
rect 496794 606454 497414 641898
rect 496794 606218 496826 606454
rect 497062 606218 497146 606454
rect 497382 606218 497414 606454
rect 496794 606134 497414 606218
rect 496794 605898 496826 606134
rect 497062 605898 497146 606134
rect 497382 605898 497414 606134
rect 496794 570454 497414 605898
rect 496794 570218 496826 570454
rect 497062 570218 497146 570454
rect 497382 570218 497414 570454
rect 496794 570134 497414 570218
rect 496794 569898 496826 570134
rect 497062 569898 497146 570134
rect 497382 569898 497414 570134
rect 496794 534454 497414 569898
rect 496794 534218 496826 534454
rect 497062 534218 497146 534454
rect 497382 534218 497414 534454
rect 496794 534134 497414 534218
rect 496794 533898 496826 534134
rect 497062 533898 497146 534134
rect 497382 533898 497414 534134
rect 496794 498454 497414 533898
rect 496794 498218 496826 498454
rect 497062 498218 497146 498454
rect 497382 498218 497414 498454
rect 496794 498134 497414 498218
rect 496794 497898 496826 498134
rect 497062 497898 497146 498134
rect 497382 497898 497414 498134
rect 496794 462454 497414 497898
rect 496794 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 497414 462454
rect 496794 462134 497414 462218
rect 496794 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 497414 462134
rect 496794 426454 497414 461898
rect 496794 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 497414 426454
rect 496794 426134 497414 426218
rect 496794 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 497414 426134
rect 496794 390454 497414 425898
rect 496794 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 497414 390454
rect 496794 390134 497414 390218
rect 496794 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 497414 390134
rect 496794 354454 497414 389898
rect 496794 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 497414 354454
rect 496794 354134 497414 354218
rect 496794 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 497414 354134
rect 496794 318454 497414 353898
rect 496794 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 497414 318454
rect 496794 318134 497414 318218
rect 496794 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 497414 318134
rect 496794 282454 497414 317898
rect 496794 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 497414 282454
rect 496794 282134 497414 282218
rect 496794 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 497414 282134
rect 496794 246454 497414 281898
rect 496794 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 497414 246454
rect 496794 246134 497414 246218
rect 496794 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 497414 246134
rect 496794 210454 497414 245898
rect 496794 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 497414 210454
rect 496794 210134 497414 210218
rect 496794 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 497414 210134
rect 496794 174454 497414 209898
rect 496794 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 497414 174454
rect 496794 174134 497414 174218
rect 496794 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 497414 174134
rect 496794 138454 497414 173898
rect 496794 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 497414 138454
rect 496794 138134 497414 138218
rect 496794 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 497414 138134
rect 496794 102454 497414 137898
rect 496794 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 497414 102454
rect 496794 102134 497414 102218
rect 496794 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 497414 102134
rect 496794 66454 497414 101898
rect 496794 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 497414 66454
rect 496794 66134 497414 66218
rect 496794 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 497414 66134
rect 496794 30454 497414 65898
rect 496794 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 497414 30454
rect 496794 30134 497414 30218
rect 496794 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 497414 30134
rect 496794 -6106 497414 29898
rect 496794 -6342 496826 -6106
rect 497062 -6342 497146 -6106
rect 497382 -6342 497414 -6106
rect 496794 -6426 497414 -6342
rect 496794 -6662 496826 -6426
rect 497062 -6662 497146 -6426
rect 497382 -6662 497414 -6426
rect 496794 -7654 497414 -6662
rect 501294 711558 501914 711590
rect 501294 711322 501326 711558
rect 501562 711322 501646 711558
rect 501882 711322 501914 711558
rect 501294 711238 501914 711322
rect 501294 711002 501326 711238
rect 501562 711002 501646 711238
rect 501882 711002 501914 711238
rect 501294 682954 501914 711002
rect 501294 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 501914 682954
rect 501294 682634 501914 682718
rect 501294 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 501914 682634
rect 501294 646954 501914 682398
rect 501294 646718 501326 646954
rect 501562 646718 501646 646954
rect 501882 646718 501914 646954
rect 501294 646634 501914 646718
rect 501294 646398 501326 646634
rect 501562 646398 501646 646634
rect 501882 646398 501914 646634
rect 501294 610954 501914 646398
rect 501294 610718 501326 610954
rect 501562 610718 501646 610954
rect 501882 610718 501914 610954
rect 501294 610634 501914 610718
rect 501294 610398 501326 610634
rect 501562 610398 501646 610634
rect 501882 610398 501914 610634
rect 501294 574954 501914 610398
rect 501294 574718 501326 574954
rect 501562 574718 501646 574954
rect 501882 574718 501914 574954
rect 501294 574634 501914 574718
rect 501294 574398 501326 574634
rect 501562 574398 501646 574634
rect 501882 574398 501914 574634
rect 501294 538954 501914 574398
rect 501294 538718 501326 538954
rect 501562 538718 501646 538954
rect 501882 538718 501914 538954
rect 501294 538634 501914 538718
rect 501294 538398 501326 538634
rect 501562 538398 501646 538634
rect 501882 538398 501914 538634
rect 501294 502954 501914 538398
rect 501294 502718 501326 502954
rect 501562 502718 501646 502954
rect 501882 502718 501914 502954
rect 501294 502634 501914 502718
rect 501294 502398 501326 502634
rect 501562 502398 501646 502634
rect 501882 502398 501914 502634
rect 501294 466954 501914 502398
rect 501294 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 501914 466954
rect 501294 466634 501914 466718
rect 501294 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 501914 466634
rect 501294 430954 501914 466398
rect 501294 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 501914 430954
rect 501294 430634 501914 430718
rect 501294 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 501914 430634
rect 501294 394954 501914 430398
rect 501294 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 501914 394954
rect 501294 394634 501914 394718
rect 501294 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 501914 394634
rect 501294 358954 501914 394398
rect 501294 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 501914 358954
rect 501294 358634 501914 358718
rect 501294 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 501914 358634
rect 501294 322954 501914 358398
rect 501294 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 501914 322954
rect 501294 322634 501914 322718
rect 501294 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 501914 322634
rect 501294 286954 501914 322398
rect 501294 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 501914 286954
rect 501294 286634 501914 286718
rect 501294 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 501914 286634
rect 501294 250954 501914 286398
rect 501294 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 501914 250954
rect 501294 250634 501914 250718
rect 501294 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 501914 250634
rect 501294 214954 501914 250398
rect 501294 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 501914 214954
rect 501294 214634 501914 214718
rect 501294 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 501914 214634
rect 501294 178954 501914 214398
rect 501294 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 501914 178954
rect 501294 178634 501914 178718
rect 501294 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 501914 178634
rect 501294 142954 501914 178398
rect 501294 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 501914 142954
rect 501294 142634 501914 142718
rect 501294 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 501914 142634
rect 501294 106954 501914 142398
rect 501294 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 501914 106954
rect 501294 106634 501914 106718
rect 501294 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 501914 106634
rect 501294 70954 501914 106398
rect 501294 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 501914 70954
rect 501294 70634 501914 70718
rect 501294 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 501914 70634
rect 501294 34954 501914 70398
rect 501294 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 501914 34954
rect 501294 34634 501914 34718
rect 501294 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 501914 34634
rect 501294 -7066 501914 34398
rect 501294 -7302 501326 -7066
rect 501562 -7302 501646 -7066
rect 501882 -7302 501914 -7066
rect 501294 -7386 501914 -7302
rect 501294 -7622 501326 -7386
rect 501562 -7622 501646 -7386
rect 501882 -7622 501914 -7386
rect 501294 -7654 501914 -7622
rect 505794 704838 506414 711590
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -7654 506414 -902
rect 510294 705798 510914 711590
rect 510294 705562 510326 705798
rect 510562 705562 510646 705798
rect 510882 705562 510914 705798
rect 510294 705478 510914 705562
rect 510294 705242 510326 705478
rect 510562 705242 510646 705478
rect 510882 705242 510914 705478
rect 510294 691954 510914 705242
rect 510294 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 510914 691954
rect 510294 691634 510914 691718
rect 510294 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 510914 691634
rect 510294 655954 510914 691398
rect 510294 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 510914 655954
rect 510294 655634 510914 655718
rect 510294 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 510914 655634
rect 510294 619954 510914 655398
rect 510294 619718 510326 619954
rect 510562 619718 510646 619954
rect 510882 619718 510914 619954
rect 510294 619634 510914 619718
rect 510294 619398 510326 619634
rect 510562 619398 510646 619634
rect 510882 619398 510914 619634
rect 510294 583954 510914 619398
rect 510294 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 510914 583954
rect 510294 583634 510914 583718
rect 510294 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 510914 583634
rect 510294 547954 510914 583398
rect 510294 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 510914 547954
rect 510294 547634 510914 547718
rect 510294 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 510914 547634
rect 510294 511954 510914 547398
rect 510294 511718 510326 511954
rect 510562 511718 510646 511954
rect 510882 511718 510914 511954
rect 510294 511634 510914 511718
rect 510294 511398 510326 511634
rect 510562 511398 510646 511634
rect 510882 511398 510914 511634
rect 510294 475954 510914 511398
rect 510294 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 510914 475954
rect 510294 475634 510914 475718
rect 510294 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 510914 475634
rect 510294 439954 510914 475398
rect 510294 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 510914 439954
rect 510294 439634 510914 439718
rect 510294 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 510914 439634
rect 510294 403954 510914 439398
rect 510294 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 510914 403954
rect 510294 403634 510914 403718
rect 510294 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 510914 403634
rect 510294 367954 510914 403398
rect 510294 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 510914 367954
rect 510294 367634 510914 367718
rect 510294 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 510914 367634
rect 510294 331954 510914 367398
rect 510294 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 510914 331954
rect 510294 331634 510914 331718
rect 510294 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 510914 331634
rect 510294 295954 510914 331398
rect 510294 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 510914 295954
rect 510294 295634 510914 295718
rect 510294 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 510914 295634
rect 510294 259954 510914 295398
rect 510294 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 510914 259954
rect 510294 259634 510914 259718
rect 510294 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 510914 259634
rect 510294 223954 510914 259398
rect 510294 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 510914 223954
rect 510294 223634 510914 223718
rect 510294 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 510914 223634
rect 510294 187954 510914 223398
rect 510294 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 510914 187954
rect 510294 187634 510914 187718
rect 510294 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 510914 187634
rect 510294 151954 510914 187398
rect 510294 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 510914 151954
rect 510294 151634 510914 151718
rect 510294 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 510914 151634
rect 510294 115954 510914 151398
rect 510294 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 510914 115954
rect 510294 115634 510914 115718
rect 510294 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 510914 115634
rect 510294 79954 510914 115398
rect 510294 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 510914 79954
rect 510294 79634 510914 79718
rect 510294 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 510914 79634
rect 510294 43954 510914 79398
rect 510294 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 510914 43954
rect 510294 43634 510914 43718
rect 510294 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 510914 43634
rect 510294 7954 510914 43398
rect 510294 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 510914 7954
rect 510294 7634 510914 7718
rect 510294 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 510914 7634
rect 510294 -1306 510914 7398
rect 510294 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 510914 -1306
rect 510294 -1626 510914 -1542
rect 510294 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 510914 -1626
rect 510294 -7654 510914 -1862
rect 514794 706758 515414 711590
rect 514794 706522 514826 706758
rect 515062 706522 515146 706758
rect 515382 706522 515414 706758
rect 514794 706438 515414 706522
rect 514794 706202 514826 706438
rect 515062 706202 515146 706438
rect 515382 706202 515414 706438
rect 514794 696454 515414 706202
rect 514794 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 515414 696454
rect 514794 696134 515414 696218
rect 514794 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 515414 696134
rect 514794 660454 515414 695898
rect 514794 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 515414 660454
rect 514794 660134 515414 660218
rect 514794 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 515414 660134
rect 514794 624454 515414 659898
rect 514794 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 515414 624454
rect 514794 624134 515414 624218
rect 514794 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 515414 624134
rect 514794 588454 515414 623898
rect 514794 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 515414 588454
rect 514794 588134 515414 588218
rect 514794 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 515414 588134
rect 514794 552454 515414 587898
rect 514794 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 515414 552454
rect 514794 552134 515414 552218
rect 514794 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 515414 552134
rect 514794 516454 515414 551898
rect 514794 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 515414 516454
rect 514794 516134 515414 516218
rect 514794 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 515414 516134
rect 514794 480454 515414 515898
rect 514794 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 515414 480454
rect 514794 480134 515414 480218
rect 514794 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 515414 480134
rect 514794 444454 515414 479898
rect 514794 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 515414 444454
rect 514794 444134 515414 444218
rect 514794 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 515414 444134
rect 514794 408454 515414 443898
rect 514794 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 515414 408454
rect 514794 408134 515414 408218
rect 514794 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 515414 408134
rect 514794 372454 515414 407898
rect 514794 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 515414 372454
rect 514794 372134 515414 372218
rect 514794 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 515414 372134
rect 514794 336454 515414 371898
rect 514794 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 515414 336454
rect 514794 336134 515414 336218
rect 514794 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 515414 336134
rect 514794 300454 515414 335898
rect 514794 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 515414 300454
rect 514794 300134 515414 300218
rect 514794 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 515414 300134
rect 514794 264454 515414 299898
rect 514794 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 515414 264454
rect 514794 264134 515414 264218
rect 514794 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 515414 264134
rect 514794 228454 515414 263898
rect 514794 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 515414 228454
rect 514794 228134 515414 228218
rect 514794 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 515414 228134
rect 514794 192454 515414 227898
rect 514794 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 515414 192454
rect 514794 192134 515414 192218
rect 514794 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 515414 192134
rect 514794 156454 515414 191898
rect 514794 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 515414 156454
rect 514794 156134 515414 156218
rect 514794 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 515414 156134
rect 514794 120454 515414 155898
rect 514794 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 515414 120454
rect 514794 120134 515414 120218
rect 514794 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 515414 120134
rect 514794 84454 515414 119898
rect 514794 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 515414 84454
rect 514794 84134 515414 84218
rect 514794 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 515414 84134
rect 514794 48454 515414 83898
rect 514794 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 515414 48454
rect 514794 48134 515414 48218
rect 514794 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 515414 48134
rect 514794 12454 515414 47898
rect 514794 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 515414 12454
rect 514794 12134 515414 12218
rect 514794 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 515414 12134
rect 514794 -2266 515414 11898
rect 514794 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 515414 -2266
rect 514794 -2586 515414 -2502
rect 514794 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 515414 -2586
rect 514794 -7654 515414 -2822
rect 519294 707718 519914 711590
rect 519294 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 519914 707718
rect 519294 707398 519914 707482
rect 519294 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 519914 707398
rect 519294 700954 519914 707162
rect 519294 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 519914 700954
rect 519294 700634 519914 700718
rect 519294 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 519914 700634
rect 519294 664954 519914 700398
rect 519294 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 519914 664954
rect 519294 664634 519914 664718
rect 519294 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 519914 664634
rect 519294 628954 519914 664398
rect 519294 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 519914 628954
rect 519294 628634 519914 628718
rect 519294 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 519914 628634
rect 519294 592954 519914 628398
rect 519294 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 519914 592954
rect 519294 592634 519914 592718
rect 519294 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 519914 592634
rect 519294 556954 519914 592398
rect 519294 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 519914 556954
rect 519294 556634 519914 556718
rect 519294 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 519914 556634
rect 519294 520954 519914 556398
rect 519294 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 519914 520954
rect 519294 520634 519914 520718
rect 519294 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 519914 520634
rect 519294 484954 519914 520398
rect 519294 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 519914 484954
rect 519294 484634 519914 484718
rect 519294 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 519914 484634
rect 519294 448954 519914 484398
rect 519294 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 519914 448954
rect 519294 448634 519914 448718
rect 519294 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 519914 448634
rect 519294 412954 519914 448398
rect 519294 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 519914 412954
rect 519294 412634 519914 412718
rect 519294 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 519914 412634
rect 519294 376954 519914 412398
rect 519294 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 519914 376954
rect 519294 376634 519914 376718
rect 519294 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 519914 376634
rect 519294 340954 519914 376398
rect 519294 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 519914 340954
rect 519294 340634 519914 340718
rect 519294 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 519914 340634
rect 519294 304954 519914 340398
rect 519294 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 519914 304954
rect 519294 304634 519914 304718
rect 519294 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 519914 304634
rect 519294 268954 519914 304398
rect 519294 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 519914 268954
rect 519294 268634 519914 268718
rect 519294 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 519914 268634
rect 519294 232954 519914 268398
rect 519294 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 519914 232954
rect 519294 232634 519914 232718
rect 519294 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 519914 232634
rect 519294 196954 519914 232398
rect 519294 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 519914 196954
rect 519294 196634 519914 196718
rect 519294 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 519914 196634
rect 519294 160954 519914 196398
rect 519294 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 519914 160954
rect 519294 160634 519914 160718
rect 519294 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 519914 160634
rect 519294 124954 519914 160398
rect 519294 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 519914 124954
rect 519294 124634 519914 124718
rect 519294 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 519914 124634
rect 519294 88954 519914 124398
rect 519294 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 519914 88954
rect 519294 88634 519914 88718
rect 519294 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 519914 88634
rect 519294 52954 519914 88398
rect 519294 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 519914 52954
rect 519294 52634 519914 52718
rect 519294 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 519914 52634
rect 519294 16954 519914 52398
rect 519294 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 519914 16954
rect 519294 16634 519914 16718
rect 519294 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 519914 16634
rect 519294 -3226 519914 16398
rect 519294 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 519914 -3226
rect 519294 -3546 519914 -3462
rect 519294 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 519914 -3546
rect 519294 -7654 519914 -3782
rect 523794 708678 524414 711590
rect 523794 708442 523826 708678
rect 524062 708442 524146 708678
rect 524382 708442 524414 708678
rect 523794 708358 524414 708442
rect 523794 708122 523826 708358
rect 524062 708122 524146 708358
rect 524382 708122 524414 708358
rect 523794 669454 524414 708122
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -4186 524414 20898
rect 523794 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 524414 -4186
rect 523794 -4506 524414 -4422
rect 523794 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 524414 -4506
rect 523794 -7654 524414 -4742
rect 528294 709638 528914 711590
rect 528294 709402 528326 709638
rect 528562 709402 528646 709638
rect 528882 709402 528914 709638
rect 528294 709318 528914 709402
rect 528294 709082 528326 709318
rect 528562 709082 528646 709318
rect 528882 709082 528914 709318
rect 528294 673954 528914 709082
rect 528294 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 528914 673954
rect 528294 673634 528914 673718
rect 528294 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 528914 673634
rect 528294 637954 528914 673398
rect 528294 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 528914 637954
rect 528294 637634 528914 637718
rect 528294 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 528914 637634
rect 528294 601954 528914 637398
rect 528294 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 528914 601954
rect 528294 601634 528914 601718
rect 528294 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 528914 601634
rect 528294 565954 528914 601398
rect 528294 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 528914 565954
rect 528294 565634 528914 565718
rect 528294 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 528914 565634
rect 528294 529954 528914 565398
rect 528294 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 528914 529954
rect 528294 529634 528914 529718
rect 528294 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 528914 529634
rect 528294 493954 528914 529398
rect 528294 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 528914 493954
rect 528294 493634 528914 493718
rect 528294 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 528914 493634
rect 528294 457954 528914 493398
rect 528294 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 528914 457954
rect 528294 457634 528914 457718
rect 528294 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 528914 457634
rect 528294 421954 528914 457398
rect 528294 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 528914 421954
rect 528294 421634 528914 421718
rect 528294 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 528914 421634
rect 528294 385954 528914 421398
rect 528294 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 528914 385954
rect 528294 385634 528914 385718
rect 528294 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 528914 385634
rect 528294 349954 528914 385398
rect 528294 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 528914 349954
rect 528294 349634 528914 349718
rect 528294 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 528914 349634
rect 528294 313954 528914 349398
rect 528294 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 528914 313954
rect 528294 313634 528914 313718
rect 528294 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 528914 313634
rect 528294 277954 528914 313398
rect 528294 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 528914 277954
rect 528294 277634 528914 277718
rect 528294 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 528914 277634
rect 528294 241954 528914 277398
rect 528294 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 528914 241954
rect 528294 241634 528914 241718
rect 528294 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 528914 241634
rect 528294 205954 528914 241398
rect 528294 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 528914 205954
rect 528294 205634 528914 205718
rect 528294 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 528914 205634
rect 528294 169954 528914 205398
rect 528294 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 528914 169954
rect 528294 169634 528914 169718
rect 528294 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 528914 169634
rect 528294 133954 528914 169398
rect 528294 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 528914 133954
rect 528294 133634 528914 133718
rect 528294 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 528914 133634
rect 528294 97954 528914 133398
rect 528294 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 528914 97954
rect 528294 97634 528914 97718
rect 528294 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 528914 97634
rect 528294 61954 528914 97398
rect 528294 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 528914 61954
rect 528294 61634 528914 61718
rect 528294 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 528914 61634
rect 528294 25954 528914 61398
rect 528294 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 528914 25954
rect 528294 25634 528914 25718
rect 528294 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 528914 25634
rect 528294 -5146 528914 25398
rect 528294 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 528914 -5146
rect 528294 -5466 528914 -5382
rect 528294 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 528914 -5466
rect 528294 -7654 528914 -5702
rect 532794 710598 533414 711590
rect 532794 710362 532826 710598
rect 533062 710362 533146 710598
rect 533382 710362 533414 710598
rect 532794 710278 533414 710362
rect 532794 710042 532826 710278
rect 533062 710042 533146 710278
rect 533382 710042 533414 710278
rect 532794 678454 533414 710042
rect 532794 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 533414 678454
rect 532794 678134 533414 678218
rect 532794 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 533414 678134
rect 532794 642454 533414 677898
rect 532794 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 533414 642454
rect 532794 642134 533414 642218
rect 532794 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 533414 642134
rect 532794 606454 533414 641898
rect 532794 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 533414 606454
rect 532794 606134 533414 606218
rect 532794 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 533414 606134
rect 532794 570454 533414 605898
rect 532794 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 533414 570454
rect 532794 570134 533414 570218
rect 532794 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 533414 570134
rect 532794 534454 533414 569898
rect 532794 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 533414 534454
rect 532794 534134 533414 534218
rect 532794 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 533414 534134
rect 532794 498454 533414 533898
rect 532794 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 533414 498454
rect 532794 498134 533414 498218
rect 532794 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 533414 498134
rect 532794 462454 533414 497898
rect 532794 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 533414 462454
rect 532794 462134 533414 462218
rect 532794 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 533414 462134
rect 532794 426454 533414 461898
rect 532794 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 533414 426454
rect 532794 426134 533414 426218
rect 532794 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 533414 426134
rect 532794 390454 533414 425898
rect 532794 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 533414 390454
rect 532794 390134 533414 390218
rect 532794 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 533414 390134
rect 532794 354454 533414 389898
rect 532794 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 533414 354454
rect 532794 354134 533414 354218
rect 532794 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 533414 354134
rect 532794 318454 533414 353898
rect 532794 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 533414 318454
rect 532794 318134 533414 318218
rect 532794 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 533414 318134
rect 532794 282454 533414 317898
rect 532794 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 533414 282454
rect 532794 282134 533414 282218
rect 532794 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 533414 282134
rect 532794 246454 533414 281898
rect 532794 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 533414 246454
rect 532794 246134 533414 246218
rect 532794 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 533414 246134
rect 532794 210454 533414 245898
rect 532794 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 533414 210454
rect 532794 210134 533414 210218
rect 532794 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 533414 210134
rect 532794 174454 533414 209898
rect 532794 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 533414 174454
rect 532794 174134 533414 174218
rect 532794 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 533414 174134
rect 532794 138454 533414 173898
rect 532794 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 533414 138454
rect 532794 138134 533414 138218
rect 532794 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 533414 138134
rect 532794 102454 533414 137898
rect 532794 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 533414 102454
rect 532794 102134 533414 102218
rect 532794 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 533414 102134
rect 532794 66454 533414 101898
rect 532794 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 533414 66454
rect 532794 66134 533414 66218
rect 532794 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 533414 66134
rect 532794 30454 533414 65898
rect 532794 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 533414 30454
rect 532794 30134 533414 30218
rect 532794 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 533414 30134
rect 532794 -6106 533414 29898
rect 532794 -6342 532826 -6106
rect 533062 -6342 533146 -6106
rect 533382 -6342 533414 -6106
rect 532794 -6426 533414 -6342
rect 532794 -6662 532826 -6426
rect 533062 -6662 533146 -6426
rect 533382 -6662 533414 -6426
rect 532794 -7654 533414 -6662
rect 537294 711558 537914 711590
rect 537294 711322 537326 711558
rect 537562 711322 537646 711558
rect 537882 711322 537914 711558
rect 537294 711238 537914 711322
rect 537294 711002 537326 711238
rect 537562 711002 537646 711238
rect 537882 711002 537914 711238
rect 537294 682954 537914 711002
rect 537294 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 537914 682954
rect 537294 682634 537914 682718
rect 537294 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 537914 682634
rect 537294 646954 537914 682398
rect 537294 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 537914 646954
rect 537294 646634 537914 646718
rect 537294 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 537914 646634
rect 537294 610954 537914 646398
rect 537294 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 537914 610954
rect 537294 610634 537914 610718
rect 537294 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 537914 610634
rect 537294 574954 537914 610398
rect 537294 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 537914 574954
rect 537294 574634 537914 574718
rect 537294 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 537914 574634
rect 537294 538954 537914 574398
rect 537294 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 537914 538954
rect 537294 538634 537914 538718
rect 537294 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 537914 538634
rect 537294 502954 537914 538398
rect 537294 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 537914 502954
rect 537294 502634 537914 502718
rect 537294 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 537914 502634
rect 537294 466954 537914 502398
rect 537294 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 537914 466954
rect 537294 466634 537914 466718
rect 537294 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 537914 466634
rect 537294 430954 537914 466398
rect 537294 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 537914 430954
rect 537294 430634 537914 430718
rect 537294 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 537914 430634
rect 537294 394954 537914 430398
rect 537294 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 537914 394954
rect 537294 394634 537914 394718
rect 537294 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 537914 394634
rect 537294 358954 537914 394398
rect 537294 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 537914 358954
rect 537294 358634 537914 358718
rect 537294 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 537914 358634
rect 537294 322954 537914 358398
rect 537294 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 537914 322954
rect 537294 322634 537914 322718
rect 537294 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 537914 322634
rect 537294 286954 537914 322398
rect 537294 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 537914 286954
rect 537294 286634 537914 286718
rect 537294 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 537914 286634
rect 537294 250954 537914 286398
rect 537294 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 537914 250954
rect 537294 250634 537914 250718
rect 537294 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 537914 250634
rect 537294 214954 537914 250398
rect 537294 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 537914 214954
rect 537294 214634 537914 214718
rect 537294 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 537914 214634
rect 537294 178954 537914 214398
rect 537294 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 537914 178954
rect 537294 178634 537914 178718
rect 537294 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 537914 178634
rect 537294 142954 537914 178398
rect 537294 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 537914 142954
rect 537294 142634 537914 142718
rect 537294 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 537914 142634
rect 537294 106954 537914 142398
rect 537294 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 537914 106954
rect 537294 106634 537914 106718
rect 537294 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 537914 106634
rect 537294 70954 537914 106398
rect 537294 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 537914 70954
rect 537294 70634 537914 70718
rect 537294 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 537914 70634
rect 537294 34954 537914 70398
rect 537294 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 537914 34954
rect 537294 34634 537914 34718
rect 537294 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 537914 34634
rect 537294 -7066 537914 34398
rect 537294 -7302 537326 -7066
rect 537562 -7302 537646 -7066
rect 537882 -7302 537914 -7066
rect 537294 -7386 537914 -7302
rect 537294 -7622 537326 -7386
rect 537562 -7622 537646 -7386
rect 537882 -7622 537914 -7386
rect 537294 -7654 537914 -7622
rect 541794 704838 542414 711590
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -7654 542414 -902
rect 546294 705798 546914 711590
rect 546294 705562 546326 705798
rect 546562 705562 546646 705798
rect 546882 705562 546914 705798
rect 546294 705478 546914 705562
rect 546294 705242 546326 705478
rect 546562 705242 546646 705478
rect 546882 705242 546914 705478
rect 546294 691954 546914 705242
rect 546294 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 546914 691954
rect 546294 691634 546914 691718
rect 546294 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 546914 691634
rect 546294 655954 546914 691398
rect 546294 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 546914 655954
rect 546294 655634 546914 655718
rect 546294 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 546914 655634
rect 546294 619954 546914 655398
rect 546294 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 546914 619954
rect 546294 619634 546914 619718
rect 546294 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 546914 619634
rect 546294 583954 546914 619398
rect 546294 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 546914 583954
rect 546294 583634 546914 583718
rect 546294 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 546914 583634
rect 546294 547954 546914 583398
rect 546294 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 546914 547954
rect 546294 547634 546914 547718
rect 546294 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 546914 547634
rect 546294 511954 546914 547398
rect 546294 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 546914 511954
rect 546294 511634 546914 511718
rect 546294 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 546914 511634
rect 546294 475954 546914 511398
rect 546294 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 546914 475954
rect 546294 475634 546914 475718
rect 546294 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 546914 475634
rect 546294 439954 546914 475398
rect 546294 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 546914 439954
rect 546294 439634 546914 439718
rect 546294 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 546914 439634
rect 546294 403954 546914 439398
rect 546294 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 546914 403954
rect 546294 403634 546914 403718
rect 546294 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 546914 403634
rect 546294 367954 546914 403398
rect 546294 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 546914 367954
rect 546294 367634 546914 367718
rect 546294 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 546914 367634
rect 546294 331954 546914 367398
rect 546294 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 546914 331954
rect 546294 331634 546914 331718
rect 546294 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 546914 331634
rect 546294 295954 546914 331398
rect 546294 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 546914 295954
rect 546294 295634 546914 295718
rect 546294 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 546914 295634
rect 546294 259954 546914 295398
rect 546294 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 546914 259954
rect 546294 259634 546914 259718
rect 546294 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 546914 259634
rect 546294 223954 546914 259398
rect 546294 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 546914 223954
rect 546294 223634 546914 223718
rect 546294 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 546914 223634
rect 546294 187954 546914 223398
rect 546294 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 546914 187954
rect 546294 187634 546914 187718
rect 546294 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 546914 187634
rect 546294 151954 546914 187398
rect 546294 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 546914 151954
rect 546294 151634 546914 151718
rect 546294 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 546914 151634
rect 546294 115954 546914 151398
rect 546294 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 546914 115954
rect 546294 115634 546914 115718
rect 546294 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 546914 115634
rect 546294 79954 546914 115398
rect 546294 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 546914 79954
rect 546294 79634 546914 79718
rect 546294 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 546914 79634
rect 546294 43954 546914 79398
rect 546294 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 546914 43954
rect 546294 43634 546914 43718
rect 546294 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 546914 43634
rect 546294 7954 546914 43398
rect 546294 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 546914 7954
rect 546294 7634 546914 7718
rect 546294 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 546914 7634
rect 546294 -1306 546914 7398
rect 546294 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 546914 -1306
rect 546294 -1626 546914 -1542
rect 546294 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 546914 -1626
rect 546294 -7654 546914 -1862
rect 550794 706758 551414 711590
rect 550794 706522 550826 706758
rect 551062 706522 551146 706758
rect 551382 706522 551414 706758
rect 550794 706438 551414 706522
rect 550794 706202 550826 706438
rect 551062 706202 551146 706438
rect 551382 706202 551414 706438
rect 550794 696454 551414 706202
rect 550794 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 551414 696454
rect 550794 696134 551414 696218
rect 550794 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 551414 696134
rect 550794 660454 551414 695898
rect 550794 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 551414 660454
rect 550794 660134 551414 660218
rect 550794 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 551414 660134
rect 550794 624454 551414 659898
rect 550794 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 551414 624454
rect 550794 624134 551414 624218
rect 550794 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 551414 624134
rect 550794 588454 551414 623898
rect 550794 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 551414 588454
rect 550794 588134 551414 588218
rect 550794 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 551414 588134
rect 550794 552454 551414 587898
rect 550794 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 551414 552454
rect 550794 552134 551414 552218
rect 550794 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 551414 552134
rect 550794 516454 551414 551898
rect 550794 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 551414 516454
rect 550794 516134 551414 516218
rect 550794 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 551414 516134
rect 550794 480454 551414 515898
rect 550794 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 551414 480454
rect 550794 480134 551414 480218
rect 550794 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 551414 480134
rect 550794 444454 551414 479898
rect 550794 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 551414 444454
rect 550794 444134 551414 444218
rect 550794 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 551414 444134
rect 550794 408454 551414 443898
rect 550794 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 551414 408454
rect 550794 408134 551414 408218
rect 550794 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 551414 408134
rect 550794 372454 551414 407898
rect 550794 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 551414 372454
rect 550794 372134 551414 372218
rect 550794 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 551414 372134
rect 550794 336454 551414 371898
rect 550794 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 551414 336454
rect 550794 336134 551414 336218
rect 550794 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 551414 336134
rect 550794 300454 551414 335898
rect 550794 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 551414 300454
rect 550794 300134 551414 300218
rect 550794 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 551414 300134
rect 550794 264454 551414 299898
rect 550794 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 551414 264454
rect 550794 264134 551414 264218
rect 550794 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 551414 264134
rect 550794 228454 551414 263898
rect 550794 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 551414 228454
rect 550794 228134 551414 228218
rect 550794 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 551414 228134
rect 550794 192454 551414 227898
rect 550794 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 551414 192454
rect 550794 192134 551414 192218
rect 550794 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 551414 192134
rect 550794 156454 551414 191898
rect 550794 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 551414 156454
rect 550794 156134 551414 156218
rect 550794 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 551414 156134
rect 550794 120454 551414 155898
rect 550794 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 551414 120454
rect 550794 120134 551414 120218
rect 550794 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 551414 120134
rect 550794 84454 551414 119898
rect 550794 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 551414 84454
rect 550794 84134 551414 84218
rect 550794 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 551414 84134
rect 550794 48454 551414 83898
rect 550794 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 551414 48454
rect 550794 48134 551414 48218
rect 550794 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 551414 48134
rect 550794 12454 551414 47898
rect 550794 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 551414 12454
rect 550794 12134 551414 12218
rect 550794 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 551414 12134
rect 550794 -2266 551414 11898
rect 550794 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 551414 -2266
rect 550794 -2586 551414 -2502
rect 550794 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 551414 -2586
rect 550794 -7654 551414 -2822
rect 555294 707718 555914 711590
rect 555294 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 555914 707718
rect 555294 707398 555914 707482
rect 555294 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 555914 707398
rect 555294 700954 555914 707162
rect 555294 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 555914 700954
rect 555294 700634 555914 700718
rect 555294 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 555914 700634
rect 555294 664954 555914 700398
rect 555294 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 555914 664954
rect 555294 664634 555914 664718
rect 555294 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 555914 664634
rect 555294 628954 555914 664398
rect 555294 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 555914 628954
rect 555294 628634 555914 628718
rect 555294 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 555914 628634
rect 555294 592954 555914 628398
rect 555294 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 555914 592954
rect 555294 592634 555914 592718
rect 555294 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 555914 592634
rect 555294 556954 555914 592398
rect 555294 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 555914 556954
rect 555294 556634 555914 556718
rect 555294 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 555914 556634
rect 555294 520954 555914 556398
rect 555294 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 555914 520954
rect 555294 520634 555914 520718
rect 555294 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 555914 520634
rect 555294 484954 555914 520398
rect 555294 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 555914 484954
rect 555294 484634 555914 484718
rect 555294 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 555914 484634
rect 555294 448954 555914 484398
rect 555294 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 555914 448954
rect 555294 448634 555914 448718
rect 555294 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 555914 448634
rect 555294 412954 555914 448398
rect 555294 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 555914 412954
rect 555294 412634 555914 412718
rect 555294 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 555914 412634
rect 555294 376954 555914 412398
rect 555294 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 555914 376954
rect 555294 376634 555914 376718
rect 555294 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 555914 376634
rect 555294 340954 555914 376398
rect 555294 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 555914 340954
rect 555294 340634 555914 340718
rect 555294 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 555914 340634
rect 555294 304954 555914 340398
rect 555294 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 555914 304954
rect 555294 304634 555914 304718
rect 555294 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 555914 304634
rect 555294 268954 555914 304398
rect 555294 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 555914 268954
rect 555294 268634 555914 268718
rect 555294 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 555914 268634
rect 555294 232954 555914 268398
rect 555294 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 555914 232954
rect 555294 232634 555914 232718
rect 555294 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 555914 232634
rect 555294 196954 555914 232398
rect 555294 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 555914 196954
rect 555294 196634 555914 196718
rect 555294 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 555914 196634
rect 555294 160954 555914 196398
rect 555294 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 555914 160954
rect 555294 160634 555914 160718
rect 555294 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 555914 160634
rect 555294 124954 555914 160398
rect 555294 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 555914 124954
rect 555294 124634 555914 124718
rect 555294 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 555914 124634
rect 555294 88954 555914 124398
rect 555294 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 555914 88954
rect 555294 88634 555914 88718
rect 555294 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 555914 88634
rect 555294 52954 555914 88398
rect 555294 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 555914 52954
rect 555294 52634 555914 52718
rect 555294 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 555914 52634
rect 555294 16954 555914 52398
rect 555294 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 555914 16954
rect 555294 16634 555914 16718
rect 555294 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 555914 16634
rect 555294 -3226 555914 16398
rect 555294 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 555914 -3226
rect 555294 -3546 555914 -3462
rect 555294 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 555914 -3546
rect 555294 -7654 555914 -3782
rect 559794 708678 560414 711590
rect 559794 708442 559826 708678
rect 560062 708442 560146 708678
rect 560382 708442 560414 708678
rect 559794 708358 560414 708442
rect 559794 708122 559826 708358
rect 560062 708122 560146 708358
rect 560382 708122 560414 708358
rect 559794 669454 560414 708122
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -4186 560414 20898
rect 559794 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 560414 -4186
rect 559794 -4506 560414 -4422
rect 559794 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 560414 -4506
rect 559794 -7654 560414 -4742
rect 564294 709638 564914 711590
rect 564294 709402 564326 709638
rect 564562 709402 564646 709638
rect 564882 709402 564914 709638
rect 564294 709318 564914 709402
rect 564294 709082 564326 709318
rect 564562 709082 564646 709318
rect 564882 709082 564914 709318
rect 564294 673954 564914 709082
rect 564294 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 564914 673954
rect 564294 673634 564914 673718
rect 564294 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 564914 673634
rect 564294 637954 564914 673398
rect 564294 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 564914 637954
rect 564294 637634 564914 637718
rect 564294 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 564914 637634
rect 564294 601954 564914 637398
rect 564294 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 564914 601954
rect 564294 601634 564914 601718
rect 564294 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 564914 601634
rect 564294 565954 564914 601398
rect 564294 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 564914 565954
rect 564294 565634 564914 565718
rect 564294 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 564914 565634
rect 564294 529954 564914 565398
rect 564294 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 564914 529954
rect 564294 529634 564914 529718
rect 564294 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 564914 529634
rect 564294 493954 564914 529398
rect 564294 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 564914 493954
rect 564294 493634 564914 493718
rect 564294 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 564914 493634
rect 564294 457954 564914 493398
rect 564294 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 564914 457954
rect 564294 457634 564914 457718
rect 564294 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 564914 457634
rect 564294 421954 564914 457398
rect 564294 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 564914 421954
rect 564294 421634 564914 421718
rect 564294 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 564914 421634
rect 564294 385954 564914 421398
rect 564294 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 564914 385954
rect 564294 385634 564914 385718
rect 564294 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 564914 385634
rect 564294 349954 564914 385398
rect 564294 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 564914 349954
rect 564294 349634 564914 349718
rect 564294 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 564914 349634
rect 564294 313954 564914 349398
rect 564294 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 564914 313954
rect 564294 313634 564914 313718
rect 564294 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 564914 313634
rect 564294 277954 564914 313398
rect 564294 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 564914 277954
rect 564294 277634 564914 277718
rect 564294 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 564914 277634
rect 564294 241954 564914 277398
rect 564294 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 564914 241954
rect 564294 241634 564914 241718
rect 564294 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 564914 241634
rect 564294 205954 564914 241398
rect 564294 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 564914 205954
rect 564294 205634 564914 205718
rect 564294 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 564914 205634
rect 564294 169954 564914 205398
rect 564294 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 564914 169954
rect 564294 169634 564914 169718
rect 564294 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 564914 169634
rect 564294 133954 564914 169398
rect 564294 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 564914 133954
rect 564294 133634 564914 133718
rect 564294 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 564914 133634
rect 564294 97954 564914 133398
rect 564294 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 564914 97954
rect 564294 97634 564914 97718
rect 564294 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 564914 97634
rect 564294 61954 564914 97398
rect 564294 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 564914 61954
rect 564294 61634 564914 61718
rect 564294 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 564914 61634
rect 564294 25954 564914 61398
rect 564294 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 564914 25954
rect 564294 25634 564914 25718
rect 564294 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 564914 25634
rect 564294 -5146 564914 25398
rect 564294 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 564914 -5146
rect 564294 -5466 564914 -5382
rect 564294 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 564914 -5466
rect 564294 -7654 564914 -5702
rect 568794 710598 569414 711590
rect 568794 710362 568826 710598
rect 569062 710362 569146 710598
rect 569382 710362 569414 710598
rect 568794 710278 569414 710362
rect 568794 710042 568826 710278
rect 569062 710042 569146 710278
rect 569382 710042 569414 710278
rect 568794 678454 569414 710042
rect 568794 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 569414 678454
rect 568794 678134 569414 678218
rect 568794 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 569414 678134
rect 568794 642454 569414 677898
rect 568794 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 569414 642454
rect 568794 642134 569414 642218
rect 568794 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 569414 642134
rect 568794 606454 569414 641898
rect 568794 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 569414 606454
rect 568794 606134 569414 606218
rect 568794 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 569414 606134
rect 568794 570454 569414 605898
rect 568794 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 569414 570454
rect 568794 570134 569414 570218
rect 568794 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 569414 570134
rect 568794 534454 569414 569898
rect 568794 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 569414 534454
rect 568794 534134 569414 534218
rect 568794 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 569414 534134
rect 568794 498454 569414 533898
rect 568794 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 569414 498454
rect 568794 498134 569414 498218
rect 568794 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 569414 498134
rect 568794 462454 569414 497898
rect 568794 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 569414 462454
rect 568794 462134 569414 462218
rect 568794 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 569414 462134
rect 568794 426454 569414 461898
rect 568794 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 569414 426454
rect 568794 426134 569414 426218
rect 568794 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 569414 426134
rect 568794 390454 569414 425898
rect 568794 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 569414 390454
rect 568794 390134 569414 390218
rect 568794 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 569414 390134
rect 568794 354454 569414 389898
rect 568794 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 569414 354454
rect 568794 354134 569414 354218
rect 568794 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 569414 354134
rect 568794 318454 569414 353898
rect 568794 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 569414 318454
rect 568794 318134 569414 318218
rect 568794 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 569414 318134
rect 568794 282454 569414 317898
rect 568794 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 569414 282454
rect 568794 282134 569414 282218
rect 568794 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 569414 282134
rect 568794 246454 569414 281898
rect 568794 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 569414 246454
rect 568794 246134 569414 246218
rect 568794 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 569414 246134
rect 568794 210454 569414 245898
rect 568794 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 569414 210454
rect 568794 210134 569414 210218
rect 568794 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 569414 210134
rect 568794 174454 569414 209898
rect 568794 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 569414 174454
rect 568794 174134 569414 174218
rect 568794 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 569414 174134
rect 568794 138454 569414 173898
rect 568794 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 569414 138454
rect 568794 138134 569414 138218
rect 568794 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 569414 138134
rect 568794 102454 569414 137898
rect 568794 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 569414 102454
rect 568794 102134 569414 102218
rect 568794 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 569414 102134
rect 568794 66454 569414 101898
rect 568794 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 569414 66454
rect 568794 66134 569414 66218
rect 568794 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 569414 66134
rect 568794 30454 569414 65898
rect 568794 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 569414 30454
rect 568794 30134 569414 30218
rect 568794 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 569414 30134
rect 568794 -6106 569414 29898
rect 568794 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 569414 -6106
rect 568794 -6426 569414 -6342
rect 568794 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 569414 -6426
rect 568794 -7654 569414 -6662
rect 573294 711558 573914 711590
rect 573294 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 573914 711558
rect 573294 711238 573914 711322
rect 573294 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 573914 711238
rect 573294 682954 573914 711002
rect 573294 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 573914 682954
rect 573294 682634 573914 682718
rect 573294 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 573914 682634
rect 573294 646954 573914 682398
rect 573294 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 573914 646954
rect 573294 646634 573914 646718
rect 573294 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 573914 646634
rect 573294 610954 573914 646398
rect 573294 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 573914 610954
rect 573294 610634 573914 610718
rect 573294 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 573914 610634
rect 573294 574954 573914 610398
rect 573294 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 573914 574954
rect 573294 574634 573914 574718
rect 573294 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 573914 574634
rect 573294 538954 573914 574398
rect 573294 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 573914 538954
rect 573294 538634 573914 538718
rect 573294 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 573914 538634
rect 573294 502954 573914 538398
rect 573294 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 573914 502954
rect 573294 502634 573914 502718
rect 573294 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 573914 502634
rect 573294 466954 573914 502398
rect 573294 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 573914 466954
rect 573294 466634 573914 466718
rect 573294 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 573914 466634
rect 573294 430954 573914 466398
rect 573294 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 573914 430954
rect 573294 430634 573914 430718
rect 573294 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 573914 430634
rect 573294 394954 573914 430398
rect 573294 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 573914 394954
rect 573294 394634 573914 394718
rect 573294 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 573914 394634
rect 573294 358954 573914 394398
rect 573294 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 573914 358954
rect 573294 358634 573914 358718
rect 573294 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 573914 358634
rect 573294 322954 573914 358398
rect 573294 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 573914 322954
rect 573294 322634 573914 322718
rect 573294 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 573914 322634
rect 573294 286954 573914 322398
rect 573294 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 573914 286954
rect 573294 286634 573914 286718
rect 573294 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 573914 286634
rect 573294 250954 573914 286398
rect 573294 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 573914 250954
rect 573294 250634 573914 250718
rect 573294 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 573914 250634
rect 573294 214954 573914 250398
rect 573294 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 573914 214954
rect 573294 214634 573914 214718
rect 573294 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 573914 214634
rect 573294 178954 573914 214398
rect 573294 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 573914 178954
rect 573294 178634 573914 178718
rect 573294 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 573914 178634
rect 573294 142954 573914 178398
rect 573294 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 573914 142954
rect 573294 142634 573914 142718
rect 573294 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 573914 142634
rect 573294 106954 573914 142398
rect 573294 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 573914 106954
rect 573294 106634 573914 106718
rect 573294 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 573914 106634
rect 573294 70954 573914 106398
rect 573294 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 573914 70954
rect 573294 70634 573914 70718
rect 573294 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 573914 70634
rect 573294 34954 573914 70398
rect 573294 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 573914 34954
rect 573294 34634 573914 34718
rect 573294 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 573914 34634
rect 573294 -7066 573914 34398
rect 573294 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 573914 -7066
rect 573294 -7386 573914 -7302
rect 573294 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 573914 -7386
rect 573294 -7654 573914 -7622
rect 577794 704838 578414 711590
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -7654 578414 -902
rect 582294 705798 582914 711590
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 582294 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 582914 705798
rect 582294 705478 582914 705562
rect 582294 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 582914 705478
rect 582294 691954 582914 705242
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 582294 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 582914 691954
rect 582294 691634 582914 691718
rect 582294 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 582914 691634
rect 582294 655954 582914 691398
rect 582294 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 582914 655954
rect 582294 655634 582914 655718
rect 582294 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 582914 655634
rect 582294 619954 582914 655398
rect 582294 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 582914 619954
rect 582294 619634 582914 619718
rect 582294 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 582914 619634
rect 582294 583954 582914 619398
rect 582294 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 582914 583954
rect 582294 583634 582914 583718
rect 582294 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 582914 583634
rect 582294 547954 582914 583398
rect 582294 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 582914 547954
rect 582294 547634 582914 547718
rect 582294 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 582914 547634
rect 582294 511954 582914 547398
rect 582294 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 582914 511954
rect 582294 511634 582914 511718
rect 582294 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 582914 511634
rect 582294 475954 582914 511398
rect 582294 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 582914 475954
rect 582294 475634 582914 475718
rect 582294 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 582914 475634
rect 582294 439954 582914 475398
rect 582294 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 582914 439954
rect 582294 439634 582914 439718
rect 582294 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 582914 439634
rect 582294 403954 582914 439398
rect 582294 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 582914 403954
rect 582294 403634 582914 403718
rect 582294 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 582914 403634
rect 582294 367954 582914 403398
rect 582294 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 582914 367954
rect 582294 367634 582914 367718
rect 582294 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 582914 367634
rect 582294 331954 582914 367398
rect 582294 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 582914 331954
rect 582294 331634 582914 331718
rect 582294 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 582914 331634
rect 582294 295954 582914 331398
rect 582294 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 582914 295954
rect 582294 295634 582914 295718
rect 582294 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 582914 295634
rect 582294 259954 582914 295398
rect 582294 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 582914 259954
rect 582294 259634 582914 259718
rect 582294 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 582914 259634
rect 582294 223954 582914 259398
rect 582294 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 582914 223954
rect 582294 223634 582914 223718
rect 582294 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 582914 223634
rect 582294 187954 582914 223398
rect 582294 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 582914 187954
rect 582294 187634 582914 187718
rect 582294 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 582914 187634
rect 582294 151954 582914 187398
rect 582294 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 582914 151954
rect 582294 151634 582914 151718
rect 582294 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 582914 151634
rect 582294 115954 582914 151398
rect 582294 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 582914 115954
rect 582294 115634 582914 115718
rect 582294 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 582914 115634
rect 582294 79954 582914 115398
rect 582294 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 582914 79954
rect 582294 79634 582914 79718
rect 582294 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 582914 79634
rect 582294 43954 582914 79398
rect 582294 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 582914 43954
rect 582294 43634 582914 43718
rect 582294 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 582914 43634
rect 582294 7954 582914 43398
rect 582294 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 582914 7954
rect 582294 7634 582914 7718
rect 582294 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 582914 7634
rect 582294 -1306 582914 7398
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 691954 586890 705242
rect 586270 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 586890 691954
rect 586270 691634 586890 691718
rect 586270 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 586890 691634
rect 586270 655954 586890 691398
rect 586270 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 586890 655954
rect 586270 655634 586890 655718
rect 586270 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 586890 655634
rect 586270 619954 586890 655398
rect 586270 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 586890 619954
rect 586270 619634 586890 619718
rect 586270 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 586890 619634
rect 586270 583954 586890 619398
rect 586270 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 586890 583954
rect 586270 583634 586890 583718
rect 586270 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 586890 583634
rect 586270 547954 586890 583398
rect 586270 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 586890 547954
rect 586270 547634 586890 547718
rect 586270 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 586890 547634
rect 586270 511954 586890 547398
rect 586270 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 586890 511954
rect 586270 511634 586890 511718
rect 586270 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 586890 511634
rect 586270 475954 586890 511398
rect 586270 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 586890 475954
rect 586270 475634 586890 475718
rect 586270 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 586890 475634
rect 586270 439954 586890 475398
rect 586270 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 586890 439954
rect 586270 439634 586890 439718
rect 586270 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 586890 439634
rect 586270 403954 586890 439398
rect 586270 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 586890 403954
rect 586270 403634 586890 403718
rect 586270 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 586890 403634
rect 586270 367954 586890 403398
rect 586270 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 586890 367954
rect 586270 367634 586890 367718
rect 586270 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 586890 367634
rect 586270 331954 586890 367398
rect 586270 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 586890 331954
rect 586270 331634 586890 331718
rect 586270 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 586890 331634
rect 586270 295954 586890 331398
rect 586270 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 586890 295954
rect 586270 295634 586890 295718
rect 586270 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 586890 295634
rect 586270 259954 586890 295398
rect 586270 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 586890 259954
rect 586270 259634 586890 259718
rect 586270 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 586890 259634
rect 586270 223954 586890 259398
rect 586270 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 586890 223954
rect 586270 223634 586890 223718
rect 586270 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 586890 223634
rect 586270 187954 586890 223398
rect 586270 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 586890 187954
rect 586270 187634 586890 187718
rect 586270 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 586890 187634
rect 586270 151954 586890 187398
rect 586270 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 586890 151954
rect 586270 151634 586890 151718
rect 586270 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 586890 151634
rect 586270 115954 586890 151398
rect 586270 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 586890 115954
rect 586270 115634 586890 115718
rect 586270 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 586890 115634
rect 586270 79954 586890 115398
rect 586270 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 586890 79954
rect 586270 79634 586890 79718
rect 586270 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 586890 79634
rect 586270 43954 586890 79398
rect 586270 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 586890 43954
rect 586270 43634 586890 43718
rect 586270 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 586890 43634
rect 586270 7954 586890 43398
rect 586270 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 586890 7954
rect 586270 7634 586890 7718
rect 586270 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 586890 7634
rect 582294 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 582914 -1306
rect 582294 -1626 582914 -1542
rect 582294 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 582914 -1626
rect 582294 -7654 582914 -1862
rect 586270 -1306 586890 7398
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 696454 587850 706202
rect 587230 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 587850 696454
rect 587230 696134 587850 696218
rect 587230 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 587850 696134
rect 587230 660454 587850 695898
rect 587230 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 587850 660454
rect 587230 660134 587850 660218
rect 587230 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 587850 660134
rect 587230 624454 587850 659898
rect 587230 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 587850 624454
rect 587230 624134 587850 624218
rect 587230 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 587850 624134
rect 587230 588454 587850 623898
rect 587230 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 587850 588454
rect 587230 588134 587850 588218
rect 587230 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 587850 588134
rect 587230 552454 587850 587898
rect 587230 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 587850 552454
rect 587230 552134 587850 552218
rect 587230 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 587850 552134
rect 587230 516454 587850 551898
rect 587230 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 587850 516454
rect 587230 516134 587850 516218
rect 587230 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 587850 516134
rect 587230 480454 587850 515898
rect 587230 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 587850 480454
rect 587230 480134 587850 480218
rect 587230 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 587850 480134
rect 587230 444454 587850 479898
rect 587230 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 587850 444454
rect 587230 444134 587850 444218
rect 587230 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 587850 444134
rect 587230 408454 587850 443898
rect 587230 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 587850 408454
rect 587230 408134 587850 408218
rect 587230 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 587850 408134
rect 587230 372454 587850 407898
rect 587230 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 587850 372454
rect 587230 372134 587850 372218
rect 587230 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 587850 372134
rect 587230 336454 587850 371898
rect 587230 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 587850 336454
rect 587230 336134 587850 336218
rect 587230 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 587850 336134
rect 587230 300454 587850 335898
rect 587230 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 587850 300454
rect 587230 300134 587850 300218
rect 587230 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 587850 300134
rect 587230 264454 587850 299898
rect 587230 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 587850 264454
rect 587230 264134 587850 264218
rect 587230 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 587850 264134
rect 587230 228454 587850 263898
rect 587230 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 587850 228454
rect 587230 228134 587850 228218
rect 587230 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 587850 228134
rect 587230 192454 587850 227898
rect 587230 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 587850 192454
rect 587230 192134 587850 192218
rect 587230 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 587850 192134
rect 587230 156454 587850 191898
rect 587230 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 587850 156454
rect 587230 156134 587850 156218
rect 587230 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 587850 156134
rect 587230 120454 587850 155898
rect 587230 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 587850 120454
rect 587230 120134 587850 120218
rect 587230 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 587850 120134
rect 587230 84454 587850 119898
rect 587230 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 587850 84454
rect 587230 84134 587850 84218
rect 587230 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 587850 84134
rect 587230 48454 587850 83898
rect 587230 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 587850 48454
rect 587230 48134 587850 48218
rect 587230 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 587850 48134
rect 587230 12454 587850 47898
rect 587230 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 587850 12454
rect 587230 12134 587850 12218
rect 587230 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 587850 12134
rect 587230 -2266 587850 11898
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 700954 588810 707162
rect 588190 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 588810 700954
rect 588190 700634 588810 700718
rect 588190 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 588810 700634
rect 588190 664954 588810 700398
rect 588190 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 588810 664954
rect 588190 664634 588810 664718
rect 588190 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 588810 664634
rect 588190 628954 588810 664398
rect 588190 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 588810 628954
rect 588190 628634 588810 628718
rect 588190 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 588810 628634
rect 588190 592954 588810 628398
rect 588190 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 588810 592954
rect 588190 592634 588810 592718
rect 588190 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 588810 592634
rect 588190 556954 588810 592398
rect 588190 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 588810 556954
rect 588190 556634 588810 556718
rect 588190 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 588810 556634
rect 588190 520954 588810 556398
rect 588190 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 588810 520954
rect 588190 520634 588810 520718
rect 588190 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 588810 520634
rect 588190 484954 588810 520398
rect 588190 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 588810 484954
rect 588190 484634 588810 484718
rect 588190 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 588810 484634
rect 588190 448954 588810 484398
rect 588190 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 588810 448954
rect 588190 448634 588810 448718
rect 588190 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 588810 448634
rect 588190 412954 588810 448398
rect 588190 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 588810 412954
rect 588190 412634 588810 412718
rect 588190 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 588810 412634
rect 588190 376954 588810 412398
rect 588190 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 588810 376954
rect 588190 376634 588810 376718
rect 588190 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 588810 376634
rect 588190 340954 588810 376398
rect 588190 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 588810 340954
rect 588190 340634 588810 340718
rect 588190 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 588810 340634
rect 588190 304954 588810 340398
rect 588190 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 588810 304954
rect 588190 304634 588810 304718
rect 588190 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 588810 304634
rect 588190 268954 588810 304398
rect 588190 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 588810 268954
rect 588190 268634 588810 268718
rect 588190 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 588810 268634
rect 588190 232954 588810 268398
rect 588190 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 588810 232954
rect 588190 232634 588810 232718
rect 588190 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 588810 232634
rect 588190 196954 588810 232398
rect 588190 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 588810 196954
rect 588190 196634 588810 196718
rect 588190 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 588810 196634
rect 588190 160954 588810 196398
rect 588190 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 588810 160954
rect 588190 160634 588810 160718
rect 588190 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 588810 160634
rect 588190 124954 588810 160398
rect 588190 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 588810 124954
rect 588190 124634 588810 124718
rect 588190 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 588810 124634
rect 588190 88954 588810 124398
rect 588190 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 588810 88954
rect 588190 88634 588810 88718
rect 588190 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 588810 88634
rect 588190 52954 588810 88398
rect 588190 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 588810 52954
rect 588190 52634 588810 52718
rect 588190 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 588810 52634
rect 588190 16954 588810 52398
rect 588190 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 588810 16954
rect 588190 16634 588810 16718
rect 588190 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 588810 16634
rect 588190 -3226 588810 16398
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 669454 589770 708122
rect 589150 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 589770 669454
rect 589150 669134 589770 669218
rect 589150 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 589770 669134
rect 589150 633454 589770 668898
rect 589150 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 589770 633454
rect 589150 633134 589770 633218
rect 589150 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 589770 633134
rect 589150 597454 589770 632898
rect 589150 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 589770 597454
rect 589150 597134 589770 597218
rect 589150 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 589770 597134
rect 589150 561454 589770 596898
rect 589150 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 589770 561454
rect 589150 561134 589770 561218
rect 589150 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 589770 561134
rect 589150 525454 589770 560898
rect 589150 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 589770 525454
rect 589150 525134 589770 525218
rect 589150 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 589770 525134
rect 589150 489454 589770 524898
rect 589150 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 589770 489454
rect 589150 489134 589770 489218
rect 589150 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 589770 489134
rect 589150 453454 589770 488898
rect 589150 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 589770 453454
rect 589150 453134 589770 453218
rect 589150 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 589770 453134
rect 589150 417454 589770 452898
rect 589150 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 589770 417454
rect 589150 417134 589770 417218
rect 589150 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 589770 417134
rect 589150 381454 589770 416898
rect 589150 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 589770 381454
rect 589150 381134 589770 381218
rect 589150 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 589770 381134
rect 589150 345454 589770 380898
rect 589150 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 589770 345454
rect 589150 345134 589770 345218
rect 589150 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 589770 345134
rect 589150 309454 589770 344898
rect 589150 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 589770 309454
rect 589150 309134 589770 309218
rect 589150 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 589770 309134
rect 589150 273454 589770 308898
rect 589150 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 589770 273454
rect 589150 273134 589770 273218
rect 589150 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 589770 273134
rect 589150 237454 589770 272898
rect 589150 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 589770 237454
rect 589150 237134 589770 237218
rect 589150 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 589770 237134
rect 589150 201454 589770 236898
rect 589150 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 589770 201454
rect 589150 201134 589770 201218
rect 589150 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 589770 201134
rect 589150 165454 589770 200898
rect 589150 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 589770 165454
rect 589150 165134 589770 165218
rect 589150 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 589770 165134
rect 589150 129454 589770 164898
rect 589150 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 589770 129454
rect 589150 129134 589770 129218
rect 589150 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 589770 129134
rect 589150 93454 589770 128898
rect 589150 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 589770 93454
rect 589150 93134 589770 93218
rect 589150 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 589770 93134
rect 589150 57454 589770 92898
rect 589150 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 589770 57454
rect 589150 57134 589770 57218
rect 589150 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 589770 57134
rect 589150 21454 589770 56898
rect 589150 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 589770 21454
rect 589150 21134 589770 21218
rect 589150 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 589770 21134
rect 589150 -4186 589770 20898
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 673954 590730 709082
rect 590110 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 590730 673954
rect 590110 673634 590730 673718
rect 590110 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 590730 673634
rect 590110 637954 590730 673398
rect 590110 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 590730 637954
rect 590110 637634 590730 637718
rect 590110 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 590730 637634
rect 590110 601954 590730 637398
rect 590110 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 590730 601954
rect 590110 601634 590730 601718
rect 590110 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 590730 601634
rect 590110 565954 590730 601398
rect 590110 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 590730 565954
rect 590110 565634 590730 565718
rect 590110 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 590730 565634
rect 590110 529954 590730 565398
rect 590110 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 590730 529954
rect 590110 529634 590730 529718
rect 590110 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 590730 529634
rect 590110 493954 590730 529398
rect 590110 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 590730 493954
rect 590110 493634 590730 493718
rect 590110 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 590730 493634
rect 590110 457954 590730 493398
rect 590110 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 590730 457954
rect 590110 457634 590730 457718
rect 590110 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 590730 457634
rect 590110 421954 590730 457398
rect 590110 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 590730 421954
rect 590110 421634 590730 421718
rect 590110 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 590730 421634
rect 590110 385954 590730 421398
rect 590110 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 590730 385954
rect 590110 385634 590730 385718
rect 590110 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 590730 385634
rect 590110 349954 590730 385398
rect 590110 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 590730 349954
rect 590110 349634 590730 349718
rect 590110 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 590730 349634
rect 590110 313954 590730 349398
rect 590110 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 590730 313954
rect 590110 313634 590730 313718
rect 590110 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 590730 313634
rect 590110 277954 590730 313398
rect 590110 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 590730 277954
rect 590110 277634 590730 277718
rect 590110 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 590730 277634
rect 590110 241954 590730 277398
rect 590110 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 590730 241954
rect 590110 241634 590730 241718
rect 590110 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 590730 241634
rect 590110 205954 590730 241398
rect 590110 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 590730 205954
rect 590110 205634 590730 205718
rect 590110 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 590730 205634
rect 590110 169954 590730 205398
rect 590110 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 590730 169954
rect 590110 169634 590730 169718
rect 590110 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 590730 169634
rect 590110 133954 590730 169398
rect 590110 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 590730 133954
rect 590110 133634 590730 133718
rect 590110 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 590730 133634
rect 590110 97954 590730 133398
rect 590110 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 590730 97954
rect 590110 97634 590730 97718
rect 590110 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 590730 97634
rect 590110 61954 590730 97398
rect 590110 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 590730 61954
rect 590110 61634 590730 61718
rect 590110 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 590730 61634
rect 590110 25954 590730 61398
rect 590110 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 590730 25954
rect 590110 25634 590730 25718
rect 590110 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 590730 25634
rect 590110 -5146 590730 25398
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 678454 591690 710042
rect 591070 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 591690 678454
rect 591070 678134 591690 678218
rect 591070 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 591690 678134
rect 591070 642454 591690 677898
rect 591070 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 591690 642454
rect 591070 642134 591690 642218
rect 591070 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 591690 642134
rect 591070 606454 591690 641898
rect 591070 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 591690 606454
rect 591070 606134 591690 606218
rect 591070 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 591690 606134
rect 591070 570454 591690 605898
rect 591070 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 591690 570454
rect 591070 570134 591690 570218
rect 591070 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 591690 570134
rect 591070 534454 591690 569898
rect 591070 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 591690 534454
rect 591070 534134 591690 534218
rect 591070 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 591690 534134
rect 591070 498454 591690 533898
rect 591070 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 591690 498454
rect 591070 498134 591690 498218
rect 591070 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 591690 498134
rect 591070 462454 591690 497898
rect 591070 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 591690 462454
rect 591070 462134 591690 462218
rect 591070 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 591690 462134
rect 591070 426454 591690 461898
rect 591070 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 591690 426454
rect 591070 426134 591690 426218
rect 591070 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 591690 426134
rect 591070 390454 591690 425898
rect 591070 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 591690 390454
rect 591070 390134 591690 390218
rect 591070 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 591690 390134
rect 591070 354454 591690 389898
rect 591070 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 591690 354454
rect 591070 354134 591690 354218
rect 591070 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 591690 354134
rect 591070 318454 591690 353898
rect 591070 318218 591102 318454
rect 591338 318218 591422 318454
rect 591658 318218 591690 318454
rect 591070 318134 591690 318218
rect 591070 317898 591102 318134
rect 591338 317898 591422 318134
rect 591658 317898 591690 318134
rect 591070 282454 591690 317898
rect 591070 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 591690 282454
rect 591070 282134 591690 282218
rect 591070 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 591690 282134
rect 591070 246454 591690 281898
rect 591070 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 591690 246454
rect 591070 246134 591690 246218
rect 591070 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 591690 246134
rect 591070 210454 591690 245898
rect 591070 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 591690 210454
rect 591070 210134 591690 210218
rect 591070 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 591690 210134
rect 591070 174454 591690 209898
rect 591070 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 591690 174454
rect 591070 174134 591690 174218
rect 591070 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 591690 174134
rect 591070 138454 591690 173898
rect 591070 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 591690 138454
rect 591070 138134 591690 138218
rect 591070 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 591690 138134
rect 591070 102454 591690 137898
rect 591070 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 591690 102454
rect 591070 102134 591690 102218
rect 591070 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 591690 102134
rect 591070 66454 591690 101898
rect 591070 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 591690 66454
rect 591070 66134 591690 66218
rect 591070 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 591690 66134
rect 591070 30454 591690 65898
rect 591070 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 591690 30454
rect 591070 30134 591690 30218
rect 591070 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 591690 30134
rect 591070 -6106 591690 29898
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 682954 592650 711002
rect 592030 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect 592030 682634 592650 682718
rect 592030 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect 592030 646954 592650 682398
rect 592030 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect 592030 646634 592650 646718
rect 592030 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect 592030 610954 592650 646398
rect 592030 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect 592030 610634 592650 610718
rect 592030 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect 592030 574954 592650 610398
rect 592030 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect 592030 574634 592650 574718
rect 592030 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect 592030 538954 592650 574398
rect 592030 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect 592030 538634 592650 538718
rect 592030 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect 592030 502954 592650 538398
rect 592030 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect 592030 502634 592650 502718
rect 592030 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect 592030 466954 592650 502398
rect 592030 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect 592030 466634 592650 466718
rect 592030 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect 592030 430954 592650 466398
rect 592030 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect 592030 430634 592650 430718
rect 592030 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect 592030 394954 592650 430398
rect 592030 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect 592030 394634 592650 394718
rect 592030 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect 592030 358954 592650 394398
rect 592030 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect 592030 358634 592650 358718
rect 592030 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect 592030 322954 592650 358398
rect 592030 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect 592030 322634 592650 322718
rect 592030 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect 592030 286954 592650 322398
rect 592030 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect 592030 286634 592650 286718
rect 592030 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect 592030 250954 592650 286398
rect 592030 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect 592030 250634 592650 250718
rect 592030 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect 592030 214954 592650 250398
rect 592030 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect 592030 214634 592650 214718
rect 592030 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect 592030 178954 592650 214398
rect 592030 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect 592030 178634 592650 178718
rect 592030 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect 592030 142954 592650 178398
rect 592030 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect 592030 142634 592650 142718
rect 592030 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect 592030 106954 592650 142398
rect 592030 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect 592030 106634 592650 106718
rect 592030 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect 592030 70954 592650 106398
rect 592030 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect 592030 70634 592650 70718
rect 592030 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect 592030 34954 592650 70398
rect 592030 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect 592030 34634 592650 34718
rect 592030 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect 592030 -7066 592650 34398
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 682718 -8458 682954
rect -8374 682718 -8138 682954
rect -8694 682398 -8458 682634
rect -8374 682398 -8138 682634
rect -8694 646718 -8458 646954
rect -8374 646718 -8138 646954
rect -8694 646398 -8458 646634
rect -8374 646398 -8138 646634
rect -8694 610718 -8458 610954
rect -8374 610718 -8138 610954
rect -8694 610398 -8458 610634
rect -8374 610398 -8138 610634
rect -8694 574718 -8458 574954
rect -8374 574718 -8138 574954
rect -8694 574398 -8458 574634
rect -8374 574398 -8138 574634
rect -8694 538718 -8458 538954
rect -8374 538718 -8138 538954
rect -8694 538398 -8458 538634
rect -8374 538398 -8138 538634
rect -8694 502718 -8458 502954
rect -8374 502718 -8138 502954
rect -8694 502398 -8458 502634
rect -8374 502398 -8138 502634
rect -8694 466718 -8458 466954
rect -8374 466718 -8138 466954
rect -8694 466398 -8458 466634
rect -8374 466398 -8138 466634
rect -8694 430718 -8458 430954
rect -8374 430718 -8138 430954
rect -8694 430398 -8458 430634
rect -8374 430398 -8138 430634
rect -8694 394718 -8458 394954
rect -8374 394718 -8138 394954
rect -8694 394398 -8458 394634
rect -8374 394398 -8138 394634
rect -8694 358718 -8458 358954
rect -8374 358718 -8138 358954
rect -8694 358398 -8458 358634
rect -8374 358398 -8138 358634
rect -8694 322718 -8458 322954
rect -8374 322718 -8138 322954
rect -8694 322398 -8458 322634
rect -8374 322398 -8138 322634
rect -8694 286718 -8458 286954
rect -8374 286718 -8138 286954
rect -8694 286398 -8458 286634
rect -8374 286398 -8138 286634
rect -8694 250718 -8458 250954
rect -8374 250718 -8138 250954
rect -8694 250398 -8458 250634
rect -8374 250398 -8138 250634
rect -8694 214718 -8458 214954
rect -8374 214718 -8138 214954
rect -8694 214398 -8458 214634
rect -8374 214398 -8138 214634
rect -8694 178718 -8458 178954
rect -8374 178718 -8138 178954
rect -8694 178398 -8458 178634
rect -8374 178398 -8138 178634
rect -8694 142718 -8458 142954
rect -8374 142718 -8138 142954
rect -8694 142398 -8458 142634
rect -8374 142398 -8138 142634
rect -8694 106718 -8458 106954
rect -8374 106718 -8138 106954
rect -8694 106398 -8458 106634
rect -8374 106398 -8138 106634
rect -8694 70718 -8458 70954
rect -8374 70718 -8138 70954
rect -8694 70398 -8458 70634
rect -8374 70398 -8138 70634
rect -8694 34718 -8458 34954
rect -8374 34718 -8138 34954
rect -8694 34398 -8458 34634
rect -8374 34398 -8138 34634
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect -7734 678218 -7498 678454
rect -7414 678218 -7178 678454
rect -7734 677898 -7498 678134
rect -7414 677898 -7178 678134
rect -7734 642218 -7498 642454
rect -7414 642218 -7178 642454
rect -7734 641898 -7498 642134
rect -7414 641898 -7178 642134
rect -7734 606218 -7498 606454
rect -7414 606218 -7178 606454
rect -7734 605898 -7498 606134
rect -7414 605898 -7178 606134
rect -7734 570218 -7498 570454
rect -7414 570218 -7178 570454
rect -7734 569898 -7498 570134
rect -7414 569898 -7178 570134
rect -7734 534218 -7498 534454
rect -7414 534218 -7178 534454
rect -7734 533898 -7498 534134
rect -7414 533898 -7178 534134
rect -7734 498218 -7498 498454
rect -7414 498218 -7178 498454
rect -7734 497898 -7498 498134
rect -7414 497898 -7178 498134
rect -7734 462218 -7498 462454
rect -7414 462218 -7178 462454
rect -7734 461898 -7498 462134
rect -7414 461898 -7178 462134
rect -7734 426218 -7498 426454
rect -7414 426218 -7178 426454
rect -7734 425898 -7498 426134
rect -7414 425898 -7178 426134
rect -7734 390218 -7498 390454
rect -7414 390218 -7178 390454
rect -7734 389898 -7498 390134
rect -7414 389898 -7178 390134
rect -7734 354218 -7498 354454
rect -7414 354218 -7178 354454
rect -7734 353898 -7498 354134
rect -7414 353898 -7178 354134
rect -7734 318218 -7498 318454
rect -7414 318218 -7178 318454
rect -7734 317898 -7498 318134
rect -7414 317898 -7178 318134
rect -7734 282218 -7498 282454
rect -7414 282218 -7178 282454
rect -7734 281898 -7498 282134
rect -7414 281898 -7178 282134
rect -7734 246218 -7498 246454
rect -7414 246218 -7178 246454
rect -7734 245898 -7498 246134
rect -7414 245898 -7178 246134
rect -7734 210218 -7498 210454
rect -7414 210218 -7178 210454
rect -7734 209898 -7498 210134
rect -7414 209898 -7178 210134
rect -7734 174218 -7498 174454
rect -7414 174218 -7178 174454
rect -7734 173898 -7498 174134
rect -7414 173898 -7178 174134
rect -7734 138218 -7498 138454
rect -7414 138218 -7178 138454
rect -7734 137898 -7498 138134
rect -7414 137898 -7178 138134
rect -7734 102218 -7498 102454
rect -7414 102218 -7178 102454
rect -7734 101898 -7498 102134
rect -7414 101898 -7178 102134
rect -7734 66218 -7498 66454
rect -7414 66218 -7178 66454
rect -7734 65898 -7498 66134
rect -7414 65898 -7178 66134
rect -7734 30218 -7498 30454
rect -7414 30218 -7178 30454
rect -7734 29898 -7498 30134
rect -7414 29898 -7178 30134
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 673718 -6538 673954
rect -6454 673718 -6218 673954
rect -6774 673398 -6538 673634
rect -6454 673398 -6218 673634
rect -6774 637718 -6538 637954
rect -6454 637718 -6218 637954
rect -6774 637398 -6538 637634
rect -6454 637398 -6218 637634
rect -6774 601718 -6538 601954
rect -6454 601718 -6218 601954
rect -6774 601398 -6538 601634
rect -6454 601398 -6218 601634
rect -6774 565718 -6538 565954
rect -6454 565718 -6218 565954
rect -6774 565398 -6538 565634
rect -6454 565398 -6218 565634
rect -6774 529718 -6538 529954
rect -6454 529718 -6218 529954
rect -6774 529398 -6538 529634
rect -6454 529398 -6218 529634
rect -6774 493718 -6538 493954
rect -6454 493718 -6218 493954
rect -6774 493398 -6538 493634
rect -6454 493398 -6218 493634
rect -6774 457718 -6538 457954
rect -6454 457718 -6218 457954
rect -6774 457398 -6538 457634
rect -6454 457398 -6218 457634
rect -6774 421718 -6538 421954
rect -6454 421718 -6218 421954
rect -6774 421398 -6538 421634
rect -6454 421398 -6218 421634
rect -6774 385718 -6538 385954
rect -6454 385718 -6218 385954
rect -6774 385398 -6538 385634
rect -6454 385398 -6218 385634
rect -6774 349718 -6538 349954
rect -6454 349718 -6218 349954
rect -6774 349398 -6538 349634
rect -6454 349398 -6218 349634
rect -6774 313718 -6538 313954
rect -6454 313718 -6218 313954
rect -6774 313398 -6538 313634
rect -6454 313398 -6218 313634
rect -6774 277718 -6538 277954
rect -6454 277718 -6218 277954
rect -6774 277398 -6538 277634
rect -6454 277398 -6218 277634
rect -6774 241718 -6538 241954
rect -6454 241718 -6218 241954
rect -6774 241398 -6538 241634
rect -6454 241398 -6218 241634
rect -6774 205718 -6538 205954
rect -6454 205718 -6218 205954
rect -6774 205398 -6538 205634
rect -6454 205398 -6218 205634
rect -6774 169718 -6538 169954
rect -6454 169718 -6218 169954
rect -6774 169398 -6538 169634
rect -6454 169398 -6218 169634
rect -6774 133718 -6538 133954
rect -6454 133718 -6218 133954
rect -6774 133398 -6538 133634
rect -6454 133398 -6218 133634
rect -6774 97718 -6538 97954
rect -6454 97718 -6218 97954
rect -6774 97398 -6538 97634
rect -6454 97398 -6218 97634
rect -6774 61718 -6538 61954
rect -6454 61718 -6218 61954
rect -6774 61398 -6538 61634
rect -6454 61398 -6218 61634
rect -6774 25718 -6538 25954
rect -6454 25718 -6218 25954
rect -6774 25398 -6538 25634
rect -6454 25398 -6218 25634
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect -5814 669218 -5578 669454
rect -5494 669218 -5258 669454
rect -5814 668898 -5578 669134
rect -5494 668898 -5258 669134
rect -5814 633218 -5578 633454
rect -5494 633218 -5258 633454
rect -5814 632898 -5578 633134
rect -5494 632898 -5258 633134
rect -5814 597218 -5578 597454
rect -5494 597218 -5258 597454
rect -5814 596898 -5578 597134
rect -5494 596898 -5258 597134
rect -5814 561218 -5578 561454
rect -5494 561218 -5258 561454
rect -5814 560898 -5578 561134
rect -5494 560898 -5258 561134
rect -5814 525218 -5578 525454
rect -5494 525218 -5258 525454
rect -5814 524898 -5578 525134
rect -5494 524898 -5258 525134
rect -5814 489218 -5578 489454
rect -5494 489218 -5258 489454
rect -5814 488898 -5578 489134
rect -5494 488898 -5258 489134
rect -5814 453218 -5578 453454
rect -5494 453218 -5258 453454
rect -5814 452898 -5578 453134
rect -5494 452898 -5258 453134
rect -5814 417218 -5578 417454
rect -5494 417218 -5258 417454
rect -5814 416898 -5578 417134
rect -5494 416898 -5258 417134
rect -5814 381218 -5578 381454
rect -5494 381218 -5258 381454
rect -5814 380898 -5578 381134
rect -5494 380898 -5258 381134
rect -5814 345218 -5578 345454
rect -5494 345218 -5258 345454
rect -5814 344898 -5578 345134
rect -5494 344898 -5258 345134
rect -5814 309218 -5578 309454
rect -5494 309218 -5258 309454
rect -5814 308898 -5578 309134
rect -5494 308898 -5258 309134
rect -5814 273218 -5578 273454
rect -5494 273218 -5258 273454
rect -5814 272898 -5578 273134
rect -5494 272898 -5258 273134
rect -5814 237218 -5578 237454
rect -5494 237218 -5258 237454
rect -5814 236898 -5578 237134
rect -5494 236898 -5258 237134
rect -5814 201218 -5578 201454
rect -5494 201218 -5258 201454
rect -5814 200898 -5578 201134
rect -5494 200898 -5258 201134
rect -5814 165218 -5578 165454
rect -5494 165218 -5258 165454
rect -5814 164898 -5578 165134
rect -5494 164898 -5258 165134
rect -5814 129218 -5578 129454
rect -5494 129218 -5258 129454
rect -5814 128898 -5578 129134
rect -5494 128898 -5258 129134
rect -5814 93218 -5578 93454
rect -5494 93218 -5258 93454
rect -5814 92898 -5578 93134
rect -5494 92898 -5258 93134
rect -5814 57218 -5578 57454
rect -5494 57218 -5258 57454
rect -5814 56898 -5578 57134
rect -5494 56898 -5258 57134
rect -5814 21218 -5578 21454
rect -5494 21218 -5258 21454
rect -5814 20898 -5578 21134
rect -5494 20898 -5258 21134
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 700718 -4618 700954
rect -4534 700718 -4298 700954
rect -4854 700398 -4618 700634
rect -4534 700398 -4298 700634
rect -4854 664718 -4618 664954
rect -4534 664718 -4298 664954
rect -4854 664398 -4618 664634
rect -4534 664398 -4298 664634
rect -4854 628718 -4618 628954
rect -4534 628718 -4298 628954
rect -4854 628398 -4618 628634
rect -4534 628398 -4298 628634
rect -4854 592718 -4618 592954
rect -4534 592718 -4298 592954
rect -4854 592398 -4618 592634
rect -4534 592398 -4298 592634
rect -4854 556718 -4618 556954
rect -4534 556718 -4298 556954
rect -4854 556398 -4618 556634
rect -4534 556398 -4298 556634
rect -4854 520718 -4618 520954
rect -4534 520718 -4298 520954
rect -4854 520398 -4618 520634
rect -4534 520398 -4298 520634
rect -4854 484718 -4618 484954
rect -4534 484718 -4298 484954
rect -4854 484398 -4618 484634
rect -4534 484398 -4298 484634
rect -4854 448718 -4618 448954
rect -4534 448718 -4298 448954
rect -4854 448398 -4618 448634
rect -4534 448398 -4298 448634
rect -4854 412718 -4618 412954
rect -4534 412718 -4298 412954
rect -4854 412398 -4618 412634
rect -4534 412398 -4298 412634
rect -4854 376718 -4618 376954
rect -4534 376718 -4298 376954
rect -4854 376398 -4618 376634
rect -4534 376398 -4298 376634
rect -4854 340718 -4618 340954
rect -4534 340718 -4298 340954
rect -4854 340398 -4618 340634
rect -4534 340398 -4298 340634
rect -4854 304718 -4618 304954
rect -4534 304718 -4298 304954
rect -4854 304398 -4618 304634
rect -4534 304398 -4298 304634
rect -4854 268718 -4618 268954
rect -4534 268718 -4298 268954
rect -4854 268398 -4618 268634
rect -4534 268398 -4298 268634
rect -4854 232718 -4618 232954
rect -4534 232718 -4298 232954
rect -4854 232398 -4618 232634
rect -4534 232398 -4298 232634
rect -4854 196718 -4618 196954
rect -4534 196718 -4298 196954
rect -4854 196398 -4618 196634
rect -4534 196398 -4298 196634
rect -4854 160718 -4618 160954
rect -4534 160718 -4298 160954
rect -4854 160398 -4618 160634
rect -4534 160398 -4298 160634
rect -4854 124718 -4618 124954
rect -4534 124718 -4298 124954
rect -4854 124398 -4618 124634
rect -4534 124398 -4298 124634
rect -4854 88718 -4618 88954
rect -4534 88718 -4298 88954
rect -4854 88398 -4618 88634
rect -4534 88398 -4298 88634
rect -4854 52718 -4618 52954
rect -4534 52718 -4298 52954
rect -4854 52398 -4618 52634
rect -4534 52398 -4298 52634
rect -4854 16718 -4618 16954
rect -4534 16718 -4298 16954
rect -4854 16398 -4618 16634
rect -4534 16398 -4298 16634
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect -3894 696218 -3658 696454
rect -3574 696218 -3338 696454
rect -3894 695898 -3658 696134
rect -3574 695898 -3338 696134
rect -3894 660218 -3658 660454
rect -3574 660218 -3338 660454
rect -3894 659898 -3658 660134
rect -3574 659898 -3338 660134
rect -3894 624218 -3658 624454
rect -3574 624218 -3338 624454
rect -3894 623898 -3658 624134
rect -3574 623898 -3338 624134
rect -3894 588218 -3658 588454
rect -3574 588218 -3338 588454
rect -3894 587898 -3658 588134
rect -3574 587898 -3338 588134
rect -3894 552218 -3658 552454
rect -3574 552218 -3338 552454
rect -3894 551898 -3658 552134
rect -3574 551898 -3338 552134
rect -3894 516218 -3658 516454
rect -3574 516218 -3338 516454
rect -3894 515898 -3658 516134
rect -3574 515898 -3338 516134
rect -3894 480218 -3658 480454
rect -3574 480218 -3338 480454
rect -3894 479898 -3658 480134
rect -3574 479898 -3338 480134
rect -3894 444218 -3658 444454
rect -3574 444218 -3338 444454
rect -3894 443898 -3658 444134
rect -3574 443898 -3338 444134
rect -3894 408218 -3658 408454
rect -3574 408218 -3338 408454
rect -3894 407898 -3658 408134
rect -3574 407898 -3338 408134
rect -3894 372218 -3658 372454
rect -3574 372218 -3338 372454
rect -3894 371898 -3658 372134
rect -3574 371898 -3338 372134
rect -3894 336218 -3658 336454
rect -3574 336218 -3338 336454
rect -3894 335898 -3658 336134
rect -3574 335898 -3338 336134
rect -3894 300218 -3658 300454
rect -3574 300218 -3338 300454
rect -3894 299898 -3658 300134
rect -3574 299898 -3338 300134
rect -3894 264218 -3658 264454
rect -3574 264218 -3338 264454
rect -3894 263898 -3658 264134
rect -3574 263898 -3338 264134
rect -3894 228218 -3658 228454
rect -3574 228218 -3338 228454
rect -3894 227898 -3658 228134
rect -3574 227898 -3338 228134
rect -3894 192218 -3658 192454
rect -3574 192218 -3338 192454
rect -3894 191898 -3658 192134
rect -3574 191898 -3338 192134
rect -3894 156218 -3658 156454
rect -3574 156218 -3338 156454
rect -3894 155898 -3658 156134
rect -3574 155898 -3338 156134
rect -3894 120218 -3658 120454
rect -3574 120218 -3338 120454
rect -3894 119898 -3658 120134
rect -3574 119898 -3338 120134
rect -3894 84218 -3658 84454
rect -3574 84218 -3338 84454
rect -3894 83898 -3658 84134
rect -3574 83898 -3338 84134
rect -3894 48218 -3658 48454
rect -3574 48218 -3338 48454
rect -3894 47898 -3658 48134
rect -3574 47898 -3338 48134
rect -3894 12218 -3658 12454
rect -3574 12218 -3338 12454
rect -3894 11898 -3658 12134
rect -3574 11898 -3338 12134
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 691718 -2698 691954
rect -2614 691718 -2378 691954
rect -2934 691398 -2698 691634
rect -2614 691398 -2378 691634
rect -2934 655718 -2698 655954
rect -2614 655718 -2378 655954
rect -2934 655398 -2698 655634
rect -2614 655398 -2378 655634
rect -2934 619718 -2698 619954
rect -2614 619718 -2378 619954
rect -2934 619398 -2698 619634
rect -2614 619398 -2378 619634
rect -2934 583718 -2698 583954
rect -2614 583718 -2378 583954
rect -2934 583398 -2698 583634
rect -2614 583398 -2378 583634
rect -2934 547718 -2698 547954
rect -2614 547718 -2378 547954
rect -2934 547398 -2698 547634
rect -2614 547398 -2378 547634
rect -2934 511718 -2698 511954
rect -2614 511718 -2378 511954
rect -2934 511398 -2698 511634
rect -2614 511398 -2378 511634
rect -2934 475718 -2698 475954
rect -2614 475718 -2378 475954
rect -2934 475398 -2698 475634
rect -2614 475398 -2378 475634
rect -2934 439718 -2698 439954
rect -2614 439718 -2378 439954
rect -2934 439398 -2698 439634
rect -2614 439398 -2378 439634
rect -2934 403718 -2698 403954
rect -2614 403718 -2378 403954
rect -2934 403398 -2698 403634
rect -2614 403398 -2378 403634
rect -2934 367718 -2698 367954
rect -2614 367718 -2378 367954
rect -2934 367398 -2698 367634
rect -2614 367398 -2378 367634
rect -2934 331718 -2698 331954
rect -2614 331718 -2378 331954
rect -2934 331398 -2698 331634
rect -2614 331398 -2378 331634
rect -2934 295718 -2698 295954
rect -2614 295718 -2378 295954
rect -2934 295398 -2698 295634
rect -2614 295398 -2378 295634
rect -2934 259718 -2698 259954
rect -2614 259718 -2378 259954
rect -2934 259398 -2698 259634
rect -2614 259398 -2378 259634
rect -2934 223718 -2698 223954
rect -2614 223718 -2378 223954
rect -2934 223398 -2698 223634
rect -2614 223398 -2378 223634
rect -2934 187718 -2698 187954
rect -2614 187718 -2378 187954
rect -2934 187398 -2698 187634
rect -2614 187398 -2378 187634
rect -2934 151718 -2698 151954
rect -2614 151718 -2378 151954
rect -2934 151398 -2698 151634
rect -2614 151398 -2378 151634
rect -2934 115718 -2698 115954
rect -2614 115718 -2378 115954
rect -2934 115398 -2698 115634
rect -2614 115398 -2378 115634
rect -2934 79718 -2698 79954
rect -2614 79718 -2378 79954
rect -2934 79398 -2698 79634
rect -2614 79398 -2378 79634
rect -2934 43718 -2698 43954
rect -2614 43718 -2378 43954
rect -2934 43398 -2698 43634
rect -2614 43398 -2378 43634
rect -2934 7718 -2698 7954
rect -2614 7718 -2378 7954
rect -2934 7398 -2698 7634
rect -2614 7398 -2378 7634
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 6326 705562 6562 705798
rect 6646 705562 6882 705798
rect 6326 705242 6562 705478
rect 6646 705242 6882 705478
rect 6326 691718 6562 691954
rect 6646 691718 6882 691954
rect 6326 691398 6562 691634
rect 6646 691398 6882 691634
rect 6326 655718 6562 655954
rect 6646 655718 6882 655954
rect 6326 655398 6562 655634
rect 6646 655398 6882 655634
rect 6326 619718 6562 619954
rect 6646 619718 6882 619954
rect 6326 619398 6562 619634
rect 6646 619398 6882 619634
rect 6326 583718 6562 583954
rect 6646 583718 6882 583954
rect 6326 583398 6562 583634
rect 6646 583398 6882 583634
rect 6326 547718 6562 547954
rect 6646 547718 6882 547954
rect 6326 547398 6562 547634
rect 6646 547398 6882 547634
rect 6326 511718 6562 511954
rect 6646 511718 6882 511954
rect 6326 511398 6562 511634
rect 6646 511398 6882 511634
rect 6326 475718 6562 475954
rect 6646 475718 6882 475954
rect 6326 475398 6562 475634
rect 6646 475398 6882 475634
rect 6326 439718 6562 439954
rect 6646 439718 6882 439954
rect 6326 439398 6562 439634
rect 6646 439398 6882 439634
rect 6326 403718 6562 403954
rect 6646 403718 6882 403954
rect 6326 403398 6562 403634
rect 6646 403398 6882 403634
rect 6326 367718 6562 367954
rect 6646 367718 6882 367954
rect 6326 367398 6562 367634
rect 6646 367398 6882 367634
rect 6326 331718 6562 331954
rect 6646 331718 6882 331954
rect 6326 331398 6562 331634
rect 6646 331398 6882 331634
rect 6326 295718 6562 295954
rect 6646 295718 6882 295954
rect 6326 295398 6562 295634
rect 6646 295398 6882 295634
rect 6326 259718 6562 259954
rect 6646 259718 6882 259954
rect 6326 259398 6562 259634
rect 6646 259398 6882 259634
rect 6326 223718 6562 223954
rect 6646 223718 6882 223954
rect 6326 223398 6562 223634
rect 6646 223398 6882 223634
rect 6326 187718 6562 187954
rect 6646 187718 6882 187954
rect 6326 187398 6562 187634
rect 6646 187398 6882 187634
rect 6326 151718 6562 151954
rect 6646 151718 6882 151954
rect 6326 151398 6562 151634
rect 6646 151398 6882 151634
rect 6326 115718 6562 115954
rect 6646 115718 6882 115954
rect 6326 115398 6562 115634
rect 6646 115398 6882 115634
rect 6326 79718 6562 79954
rect 6646 79718 6882 79954
rect 6326 79398 6562 79634
rect 6646 79398 6882 79634
rect 6326 43718 6562 43954
rect 6646 43718 6882 43954
rect 6326 43398 6562 43634
rect 6646 43398 6882 43634
rect 6326 7718 6562 7954
rect 6646 7718 6882 7954
rect 6326 7398 6562 7634
rect 6646 7398 6882 7634
rect 6326 -1542 6562 -1306
rect 6646 -1542 6882 -1306
rect 6326 -1862 6562 -1626
rect 6646 -1862 6882 -1626
rect 10826 706522 11062 706758
rect 11146 706522 11382 706758
rect 10826 706202 11062 706438
rect 11146 706202 11382 706438
rect 10826 696218 11062 696454
rect 11146 696218 11382 696454
rect 10826 695898 11062 696134
rect 11146 695898 11382 696134
rect 10826 660218 11062 660454
rect 11146 660218 11382 660454
rect 10826 659898 11062 660134
rect 11146 659898 11382 660134
rect 10826 624218 11062 624454
rect 11146 624218 11382 624454
rect 10826 623898 11062 624134
rect 11146 623898 11382 624134
rect 10826 588218 11062 588454
rect 11146 588218 11382 588454
rect 10826 587898 11062 588134
rect 11146 587898 11382 588134
rect 10826 552218 11062 552454
rect 11146 552218 11382 552454
rect 10826 551898 11062 552134
rect 11146 551898 11382 552134
rect 10826 516218 11062 516454
rect 11146 516218 11382 516454
rect 10826 515898 11062 516134
rect 11146 515898 11382 516134
rect 10826 480218 11062 480454
rect 11146 480218 11382 480454
rect 10826 479898 11062 480134
rect 11146 479898 11382 480134
rect 10826 444218 11062 444454
rect 11146 444218 11382 444454
rect 10826 443898 11062 444134
rect 11146 443898 11382 444134
rect 10826 408218 11062 408454
rect 11146 408218 11382 408454
rect 10826 407898 11062 408134
rect 11146 407898 11382 408134
rect 10826 372218 11062 372454
rect 11146 372218 11382 372454
rect 10826 371898 11062 372134
rect 11146 371898 11382 372134
rect 10826 336218 11062 336454
rect 11146 336218 11382 336454
rect 10826 335898 11062 336134
rect 11146 335898 11382 336134
rect 10826 300218 11062 300454
rect 11146 300218 11382 300454
rect 10826 299898 11062 300134
rect 11146 299898 11382 300134
rect 10826 264218 11062 264454
rect 11146 264218 11382 264454
rect 10826 263898 11062 264134
rect 11146 263898 11382 264134
rect 10826 228218 11062 228454
rect 11146 228218 11382 228454
rect 10826 227898 11062 228134
rect 11146 227898 11382 228134
rect 10826 192218 11062 192454
rect 11146 192218 11382 192454
rect 10826 191898 11062 192134
rect 11146 191898 11382 192134
rect 10826 156218 11062 156454
rect 11146 156218 11382 156454
rect 10826 155898 11062 156134
rect 11146 155898 11382 156134
rect 10826 120218 11062 120454
rect 11146 120218 11382 120454
rect 10826 119898 11062 120134
rect 11146 119898 11382 120134
rect 10826 84218 11062 84454
rect 11146 84218 11382 84454
rect 10826 83898 11062 84134
rect 11146 83898 11382 84134
rect 10826 48218 11062 48454
rect 11146 48218 11382 48454
rect 10826 47898 11062 48134
rect 11146 47898 11382 48134
rect 10826 12218 11062 12454
rect 11146 12218 11382 12454
rect 10826 11898 11062 12134
rect 11146 11898 11382 12134
rect 10826 -2502 11062 -2266
rect 11146 -2502 11382 -2266
rect 10826 -2822 11062 -2586
rect 11146 -2822 11382 -2586
rect 15326 707482 15562 707718
rect 15646 707482 15882 707718
rect 15326 707162 15562 707398
rect 15646 707162 15882 707398
rect 15326 700718 15562 700954
rect 15646 700718 15882 700954
rect 15326 700398 15562 700634
rect 15646 700398 15882 700634
rect 15326 664718 15562 664954
rect 15646 664718 15882 664954
rect 15326 664398 15562 664634
rect 15646 664398 15882 664634
rect 15326 628718 15562 628954
rect 15646 628718 15882 628954
rect 15326 628398 15562 628634
rect 15646 628398 15882 628634
rect 15326 592718 15562 592954
rect 15646 592718 15882 592954
rect 15326 592398 15562 592634
rect 15646 592398 15882 592634
rect 15326 556718 15562 556954
rect 15646 556718 15882 556954
rect 15326 556398 15562 556634
rect 15646 556398 15882 556634
rect 15326 520718 15562 520954
rect 15646 520718 15882 520954
rect 15326 520398 15562 520634
rect 15646 520398 15882 520634
rect 15326 484718 15562 484954
rect 15646 484718 15882 484954
rect 15326 484398 15562 484634
rect 15646 484398 15882 484634
rect 15326 448718 15562 448954
rect 15646 448718 15882 448954
rect 15326 448398 15562 448634
rect 15646 448398 15882 448634
rect 15326 412718 15562 412954
rect 15646 412718 15882 412954
rect 15326 412398 15562 412634
rect 15646 412398 15882 412634
rect 15326 376718 15562 376954
rect 15646 376718 15882 376954
rect 15326 376398 15562 376634
rect 15646 376398 15882 376634
rect 15326 340718 15562 340954
rect 15646 340718 15882 340954
rect 15326 340398 15562 340634
rect 15646 340398 15882 340634
rect 15326 304718 15562 304954
rect 15646 304718 15882 304954
rect 15326 304398 15562 304634
rect 15646 304398 15882 304634
rect 15326 268718 15562 268954
rect 15646 268718 15882 268954
rect 15326 268398 15562 268634
rect 15646 268398 15882 268634
rect 15326 232718 15562 232954
rect 15646 232718 15882 232954
rect 15326 232398 15562 232634
rect 15646 232398 15882 232634
rect 15326 196718 15562 196954
rect 15646 196718 15882 196954
rect 15326 196398 15562 196634
rect 15646 196398 15882 196634
rect 15326 160718 15562 160954
rect 15646 160718 15882 160954
rect 15326 160398 15562 160634
rect 15646 160398 15882 160634
rect 15326 124718 15562 124954
rect 15646 124718 15882 124954
rect 15326 124398 15562 124634
rect 15646 124398 15882 124634
rect 15326 88718 15562 88954
rect 15646 88718 15882 88954
rect 15326 88398 15562 88634
rect 15646 88398 15882 88634
rect 15326 52718 15562 52954
rect 15646 52718 15882 52954
rect 15326 52398 15562 52634
rect 15646 52398 15882 52634
rect 15326 16718 15562 16954
rect 15646 16718 15882 16954
rect 15326 16398 15562 16634
rect 15646 16398 15882 16634
rect 15326 -3462 15562 -3226
rect 15646 -3462 15882 -3226
rect 15326 -3782 15562 -3546
rect 15646 -3782 15882 -3546
rect 19826 708442 20062 708678
rect 20146 708442 20382 708678
rect 19826 708122 20062 708358
rect 20146 708122 20382 708358
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -4422 20062 -4186
rect 20146 -4422 20382 -4186
rect 19826 -4742 20062 -4506
rect 20146 -4742 20382 -4506
rect 24326 709402 24562 709638
rect 24646 709402 24882 709638
rect 24326 709082 24562 709318
rect 24646 709082 24882 709318
rect 24326 673718 24562 673954
rect 24646 673718 24882 673954
rect 24326 673398 24562 673634
rect 24646 673398 24882 673634
rect 24326 637718 24562 637954
rect 24646 637718 24882 637954
rect 24326 637398 24562 637634
rect 24646 637398 24882 637634
rect 24326 601718 24562 601954
rect 24646 601718 24882 601954
rect 24326 601398 24562 601634
rect 24646 601398 24882 601634
rect 24326 565718 24562 565954
rect 24646 565718 24882 565954
rect 24326 565398 24562 565634
rect 24646 565398 24882 565634
rect 24326 529718 24562 529954
rect 24646 529718 24882 529954
rect 24326 529398 24562 529634
rect 24646 529398 24882 529634
rect 24326 493718 24562 493954
rect 24646 493718 24882 493954
rect 24326 493398 24562 493634
rect 24646 493398 24882 493634
rect 24326 457718 24562 457954
rect 24646 457718 24882 457954
rect 24326 457398 24562 457634
rect 24646 457398 24882 457634
rect 24326 421718 24562 421954
rect 24646 421718 24882 421954
rect 24326 421398 24562 421634
rect 24646 421398 24882 421634
rect 24326 385718 24562 385954
rect 24646 385718 24882 385954
rect 24326 385398 24562 385634
rect 24646 385398 24882 385634
rect 24326 349718 24562 349954
rect 24646 349718 24882 349954
rect 24326 349398 24562 349634
rect 24646 349398 24882 349634
rect 24326 313718 24562 313954
rect 24646 313718 24882 313954
rect 24326 313398 24562 313634
rect 24646 313398 24882 313634
rect 24326 277718 24562 277954
rect 24646 277718 24882 277954
rect 24326 277398 24562 277634
rect 24646 277398 24882 277634
rect 24326 241718 24562 241954
rect 24646 241718 24882 241954
rect 24326 241398 24562 241634
rect 24646 241398 24882 241634
rect 24326 205718 24562 205954
rect 24646 205718 24882 205954
rect 24326 205398 24562 205634
rect 24646 205398 24882 205634
rect 24326 169718 24562 169954
rect 24646 169718 24882 169954
rect 24326 169398 24562 169634
rect 24646 169398 24882 169634
rect 24326 133718 24562 133954
rect 24646 133718 24882 133954
rect 24326 133398 24562 133634
rect 24646 133398 24882 133634
rect 24326 97718 24562 97954
rect 24646 97718 24882 97954
rect 24326 97398 24562 97634
rect 24646 97398 24882 97634
rect 24326 61718 24562 61954
rect 24646 61718 24882 61954
rect 24326 61398 24562 61634
rect 24646 61398 24882 61634
rect 24326 25718 24562 25954
rect 24646 25718 24882 25954
rect 24326 25398 24562 25634
rect 24646 25398 24882 25634
rect 24326 -5382 24562 -5146
rect 24646 -5382 24882 -5146
rect 24326 -5702 24562 -5466
rect 24646 -5702 24882 -5466
rect 28826 710362 29062 710598
rect 29146 710362 29382 710598
rect 28826 710042 29062 710278
rect 29146 710042 29382 710278
rect 28826 678218 29062 678454
rect 29146 678218 29382 678454
rect 28826 677898 29062 678134
rect 29146 677898 29382 678134
rect 28826 642218 29062 642454
rect 29146 642218 29382 642454
rect 28826 641898 29062 642134
rect 29146 641898 29382 642134
rect 28826 606218 29062 606454
rect 29146 606218 29382 606454
rect 28826 605898 29062 606134
rect 29146 605898 29382 606134
rect 28826 570218 29062 570454
rect 29146 570218 29382 570454
rect 28826 569898 29062 570134
rect 29146 569898 29382 570134
rect 28826 534218 29062 534454
rect 29146 534218 29382 534454
rect 28826 533898 29062 534134
rect 29146 533898 29382 534134
rect 28826 498218 29062 498454
rect 29146 498218 29382 498454
rect 28826 497898 29062 498134
rect 29146 497898 29382 498134
rect 28826 462218 29062 462454
rect 29146 462218 29382 462454
rect 28826 461898 29062 462134
rect 29146 461898 29382 462134
rect 28826 426218 29062 426454
rect 29146 426218 29382 426454
rect 28826 425898 29062 426134
rect 29146 425898 29382 426134
rect 28826 390218 29062 390454
rect 29146 390218 29382 390454
rect 28826 389898 29062 390134
rect 29146 389898 29382 390134
rect 28826 354218 29062 354454
rect 29146 354218 29382 354454
rect 28826 353898 29062 354134
rect 29146 353898 29382 354134
rect 28826 318218 29062 318454
rect 29146 318218 29382 318454
rect 28826 317898 29062 318134
rect 29146 317898 29382 318134
rect 28826 282218 29062 282454
rect 29146 282218 29382 282454
rect 28826 281898 29062 282134
rect 29146 281898 29382 282134
rect 28826 246218 29062 246454
rect 29146 246218 29382 246454
rect 28826 245898 29062 246134
rect 29146 245898 29382 246134
rect 28826 210218 29062 210454
rect 29146 210218 29382 210454
rect 28826 209898 29062 210134
rect 29146 209898 29382 210134
rect 28826 174218 29062 174454
rect 29146 174218 29382 174454
rect 28826 173898 29062 174134
rect 29146 173898 29382 174134
rect 28826 138218 29062 138454
rect 29146 138218 29382 138454
rect 28826 137898 29062 138134
rect 29146 137898 29382 138134
rect 28826 102218 29062 102454
rect 29146 102218 29382 102454
rect 28826 101898 29062 102134
rect 29146 101898 29382 102134
rect 28826 66218 29062 66454
rect 29146 66218 29382 66454
rect 28826 65898 29062 66134
rect 29146 65898 29382 66134
rect 28826 30218 29062 30454
rect 29146 30218 29382 30454
rect 28826 29898 29062 30134
rect 29146 29898 29382 30134
rect 28826 -6342 29062 -6106
rect 29146 -6342 29382 -6106
rect 28826 -6662 29062 -6426
rect 29146 -6662 29382 -6426
rect 33326 711322 33562 711558
rect 33646 711322 33882 711558
rect 33326 711002 33562 711238
rect 33646 711002 33882 711238
rect 33326 682718 33562 682954
rect 33646 682718 33882 682954
rect 33326 682398 33562 682634
rect 33646 682398 33882 682634
rect 33326 646718 33562 646954
rect 33646 646718 33882 646954
rect 33326 646398 33562 646634
rect 33646 646398 33882 646634
rect 33326 610718 33562 610954
rect 33646 610718 33882 610954
rect 33326 610398 33562 610634
rect 33646 610398 33882 610634
rect 33326 574718 33562 574954
rect 33646 574718 33882 574954
rect 33326 574398 33562 574634
rect 33646 574398 33882 574634
rect 33326 538718 33562 538954
rect 33646 538718 33882 538954
rect 33326 538398 33562 538634
rect 33646 538398 33882 538634
rect 33326 502718 33562 502954
rect 33646 502718 33882 502954
rect 33326 502398 33562 502634
rect 33646 502398 33882 502634
rect 33326 466718 33562 466954
rect 33646 466718 33882 466954
rect 33326 466398 33562 466634
rect 33646 466398 33882 466634
rect 33326 430718 33562 430954
rect 33646 430718 33882 430954
rect 33326 430398 33562 430634
rect 33646 430398 33882 430634
rect 33326 394718 33562 394954
rect 33646 394718 33882 394954
rect 33326 394398 33562 394634
rect 33646 394398 33882 394634
rect 33326 358718 33562 358954
rect 33646 358718 33882 358954
rect 33326 358398 33562 358634
rect 33646 358398 33882 358634
rect 33326 322718 33562 322954
rect 33646 322718 33882 322954
rect 33326 322398 33562 322634
rect 33646 322398 33882 322634
rect 33326 286718 33562 286954
rect 33646 286718 33882 286954
rect 33326 286398 33562 286634
rect 33646 286398 33882 286634
rect 33326 250718 33562 250954
rect 33646 250718 33882 250954
rect 33326 250398 33562 250634
rect 33646 250398 33882 250634
rect 33326 214718 33562 214954
rect 33646 214718 33882 214954
rect 33326 214398 33562 214634
rect 33646 214398 33882 214634
rect 33326 178718 33562 178954
rect 33646 178718 33882 178954
rect 33326 178398 33562 178634
rect 33646 178398 33882 178634
rect 33326 142718 33562 142954
rect 33646 142718 33882 142954
rect 33326 142398 33562 142634
rect 33646 142398 33882 142634
rect 33326 106718 33562 106954
rect 33646 106718 33882 106954
rect 33326 106398 33562 106634
rect 33646 106398 33882 106634
rect 33326 70718 33562 70954
rect 33646 70718 33882 70954
rect 33326 70398 33562 70634
rect 33646 70398 33882 70634
rect 33326 34718 33562 34954
rect 33646 34718 33882 34954
rect 33326 34398 33562 34634
rect 33646 34398 33882 34634
rect 33326 -7302 33562 -7066
rect 33646 -7302 33882 -7066
rect 33326 -7622 33562 -7386
rect 33646 -7622 33882 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 42326 705562 42562 705798
rect 42646 705562 42882 705798
rect 42326 705242 42562 705478
rect 42646 705242 42882 705478
rect 42326 691718 42562 691954
rect 42646 691718 42882 691954
rect 42326 691398 42562 691634
rect 42646 691398 42882 691634
rect 42326 655718 42562 655954
rect 42646 655718 42882 655954
rect 42326 655398 42562 655634
rect 42646 655398 42882 655634
rect 42326 619718 42562 619954
rect 42646 619718 42882 619954
rect 42326 619398 42562 619634
rect 42646 619398 42882 619634
rect 42326 583718 42562 583954
rect 42646 583718 42882 583954
rect 42326 583398 42562 583634
rect 42646 583398 42882 583634
rect 42326 547718 42562 547954
rect 42646 547718 42882 547954
rect 42326 547398 42562 547634
rect 42646 547398 42882 547634
rect 42326 511718 42562 511954
rect 42646 511718 42882 511954
rect 42326 511398 42562 511634
rect 42646 511398 42882 511634
rect 42326 475718 42562 475954
rect 42646 475718 42882 475954
rect 42326 475398 42562 475634
rect 42646 475398 42882 475634
rect 42326 439718 42562 439954
rect 42646 439718 42882 439954
rect 42326 439398 42562 439634
rect 42646 439398 42882 439634
rect 42326 403718 42562 403954
rect 42646 403718 42882 403954
rect 42326 403398 42562 403634
rect 42646 403398 42882 403634
rect 42326 367718 42562 367954
rect 42646 367718 42882 367954
rect 42326 367398 42562 367634
rect 42646 367398 42882 367634
rect 42326 331718 42562 331954
rect 42646 331718 42882 331954
rect 42326 331398 42562 331634
rect 42646 331398 42882 331634
rect 42326 295718 42562 295954
rect 42646 295718 42882 295954
rect 42326 295398 42562 295634
rect 42646 295398 42882 295634
rect 42326 259718 42562 259954
rect 42646 259718 42882 259954
rect 42326 259398 42562 259634
rect 42646 259398 42882 259634
rect 42326 223718 42562 223954
rect 42646 223718 42882 223954
rect 42326 223398 42562 223634
rect 42646 223398 42882 223634
rect 42326 187718 42562 187954
rect 42646 187718 42882 187954
rect 42326 187398 42562 187634
rect 42646 187398 42882 187634
rect 42326 151718 42562 151954
rect 42646 151718 42882 151954
rect 42326 151398 42562 151634
rect 42646 151398 42882 151634
rect 42326 115718 42562 115954
rect 42646 115718 42882 115954
rect 42326 115398 42562 115634
rect 42646 115398 42882 115634
rect 42326 79718 42562 79954
rect 42646 79718 42882 79954
rect 42326 79398 42562 79634
rect 42646 79398 42882 79634
rect 42326 43718 42562 43954
rect 42646 43718 42882 43954
rect 42326 43398 42562 43634
rect 42646 43398 42882 43634
rect 42326 7718 42562 7954
rect 42646 7718 42882 7954
rect 42326 7398 42562 7634
rect 42646 7398 42882 7634
rect 42326 -1542 42562 -1306
rect 42646 -1542 42882 -1306
rect 42326 -1862 42562 -1626
rect 42646 -1862 42882 -1626
rect 46826 706522 47062 706758
rect 47146 706522 47382 706758
rect 46826 706202 47062 706438
rect 47146 706202 47382 706438
rect 46826 696218 47062 696454
rect 47146 696218 47382 696454
rect 46826 695898 47062 696134
rect 47146 695898 47382 696134
rect 46826 660218 47062 660454
rect 47146 660218 47382 660454
rect 46826 659898 47062 660134
rect 47146 659898 47382 660134
rect 46826 624218 47062 624454
rect 47146 624218 47382 624454
rect 46826 623898 47062 624134
rect 47146 623898 47382 624134
rect 46826 588218 47062 588454
rect 47146 588218 47382 588454
rect 46826 587898 47062 588134
rect 47146 587898 47382 588134
rect 46826 552218 47062 552454
rect 47146 552218 47382 552454
rect 46826 551898 47062 552134
rect 47146 551898 47382 552134
rect 46826 516218 47062 516454
rect 47146 516218 47382 516454
rect 46826 515898 47062 516134
rect 47146 515898 47382 516134
rect 46826 480218 47062 480454
rect 47146 480218 47382 480454
rect 46826 479898 47062 480134
rect 47146 479898 47382 480134
rect 46826 444218 47062 444454
rect 47146 444218 47382 444454
rect 46826 443898 47062 444134
rect 47146 443898 47382 444134
rect 46826 408218 47062 408454
rect 47146 408218 47382 408454
rect 46826 407898 47062 408134
rect 47146 407898 47382 408134
rect 46826 372218 47062 372454
rect 47146 372218 47382 372454
rect 46826 371898 47062 372134
rect 47146 371898 47382 372134
rect 46826 336218 47062 336454
rect 47146 336218 47382 336454
rect 46826 335898 47062 336134
rect 47146 335898 47382 336134
rect 46826 300218 47062 300454
rect 47146 300218 47382 300454
rect 46826 299898 47062 300134
rect 47146 299898 47382 300134
rect 46826 264218 47062 264454
rect 47146 264218 47382 264454
rect 46826 263898 47062 264134
rect 47146 263898 47382 264134
rect 46826 228218 47062 228454
rect 47146 228218 47382 228454
rect 46826 227898 47062 228134
rect 47146 227898 47382 228134
rect 46826 192218 47062 192454
rect 47146 192218 47382 192454
rect 46826 191898 47062 192134
rect 47146 191898 47382 192134
rect 46826 156218 47062 156454
rect 47146 156218 47382 156454
rect 46826 155898 47062 156134
rect 47146 155898 47382 156134
rect 46826 120218 47062 120454
rect 47146 120218 47382 120454
rect 46826 119898 47062 120134
rect 47146 119898 47382 120134
rect 46826 84218 47062 84454
rect 47146 84218 47382 84454
rect 46826 83898 47062 84134
rect 47146 83898 47382 84134
rect 46826 48218 47062 48454
rect 47146 48218 47382 48454
rect 46826 47898 47062 48134
rect 47146 47898 47382 48134
rect 46826 12218 47062 12454
rect 47146 12218 47382 12454
rect 46826 11898 47062 12134
rect 47146 11898 47382 12134
rect 46826 -2502 47062 -2266
rect 47146 -2502 47382 -2266
rect 46826 -2822 47062 -2586
rect 47146 -2822 47382 -2586
rect 51326 707482 51562 707718
rect 51646 707482 51882 707718
rect 51326 707162 51562 707398
rect 51646 707162 51882 707398
rect 51326 700718 51562 700954
rect 51646 700718 51882 700954
rect 51326 700398 51562 700634
rect 51646 700398 51882 700634
rect 51326 664718 51562 664954
rect 51646 664718 51882 664954
rect 51326 664398 51562 664634
rect 51646 664398 51882 664634
rect 51326 628718 51562 628954
rect 51646 628718 51882 628954
rect 51326 628398 51562 628634
rect 51646 628398 51882 628634
rect 51326 592718 51562 592954
rect 51646 592718 51882 592954
rect 51326 592398 51562 592634
rect 51646 592398 51882 592634
rect 51326 556718 51562 556954
rect 51646 556718 51882 556954
rect 51326 556398 51562 556634
rect 51646 556398 51882 556634
rect 51326 520718 51562 520954
rect 51646 520718 51882 520954
rect 51326 520398 51562 520634
rect 51646 520398 51882 520634
rect 51326 484718 51562 484954
rect 51646 484718 51882 484954
rect 51326 484398 51562 484634
rect 51646 484398 51882 484634
rect 51326 448718 51562 448954
rect 51646 448718 51882 448954
rect 51326 448398 51562 448634
rect 51646 448398 51882 448634
rect 51326 412718 51562 412954
rect 51646 412718 51882 412954
rect 51326 412398 51562 412634
rect 51646 412398 51882 412634
rect 51326 376718 51562 376954
rect 51646 376718 51882 376954
rect 51326 376398 51562 376634
rect 51646 376398 51882 376634
rect 51326 340718 51562 340954
rect 51646 340718 51882 340954
rect 51326 340398 51562 340634
rect 51646 340398 51882 340634
rect 51326 304718 51562 304954
rect 51646 304718 51882 304954
rect 51326 304398 51562 304634
rect 51646 304398 51882 304634
rect 51326 268718 51562 268954
rect 51646 268718 51882 268954
rect 51326 268398 51562 268634
rect 51646 268398 51882 268634
rect 51326 232718 51562 232954
rect 51646 232718 51882 232954
rect 51326 232398 51562 232634
rect 51646 232398 51882 232634
rect 51326 196718 51562 196954
rect 51646 196718 51882 196954
rect 51326 196398 51562 196634
rect 51646 196398 51882 196634
rect 51326 160718 51562 160954
rect 51646 160718 51882 160954
rect 51326 160398 51562 160634
rect 51646 160398 51882 160634
rect 51326 124718 51562 124954
rect 51646 124718 51882 124954
rect 51326 124398 51562 124634
rect 51646 124398 51882 124634
rect 51326 88718 51562 88954
rect 51646 88718 51882 88954
rect 51326 88398 51562 88634
rect 51646 88398 51882 88634
rect 51326 52718 51562 52954
rect 51646 52718 51882 52954
rect 51326 52398 51562 52634
rect 51646 52398 51882 52634
rect 51326 16718 51562 16954
rect 51646 16718 51882 16954
rect 51326 16398 51562 16634
rect 51646 16398 51882 16634
rect 51326 -3462 51562 -3226
rect 51646 -3462 51882 -3226
rect 51326 -3782 51562 -3546
rect 51646 -3782 51882 -3546
rect 55826 708442 56062 708678
rect 56146 708442 56382 708678
rect 55826 708122 56062 708358
rect 56146 708122 56382 708358
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -4422 56062 -4186
rect 56146 -4422 56382 -4186
rect 55826 -4742 56062 -4506
rect 56146 -4742 56382 -4506
rect 60326 709402 60562 709638
rect 60646 709402 60882 709638
rect 60326 709082 60562 709318
rect 60646 709082 60882 709318
rect 60326 673718 60562 673954
rect 60646 673718 60882 673954
rect 60326 673398 60562 673634
rect 60646 673398 60882 673634
rect 60326 637718 60562 637954
rect 60646 637718 60882 637954
rect 60326 637398 60562 637634
rect 60646 637398 60882 637634
rect 60326 601718 60562 601954
rect 60646 601718 60882 601954
rect 60326 601398 60562 601634
rect 60646 601398 60882 601634
rect 60326 565718 60562 565954
rect 60646 565718 60882 565954
rect 60326 565398 60562 565634
rect 60646 565398 60882 565634
rect 60326 529718 60562 529954
rect 60646 529718 60882 529954
rect 60326 529398 60562 529634
rect 60646 529398 60882 529634
rect 60326 493718 60562 493954
rect 60646 493718 60882 493954
rect 60326 493398 60562 493634
rect 60646 493398 60882 493634
rect 60326 457718 60562 457954
rect 60646 457718 60882 457954
rect 60326 457398 60562 457634
rect 60646 457398 60882 457634
rect 60326 421718 60562 421954
rect 60646 421718 60882 421954
rect 60326 421398 60562 421634
rect 60646 421398 60882 421634
rect 60326 385718 60562 385954
rect 60646 385718 60882 385954
rect 60326 385398 60562 385634
rect 60646 385398 60882 385634
rect 60326 349718 60562 349954
rect 60646 349718 60882 349954
rect 60326 349398 60562 349634
rect 60646 349398 60882 349634
rect 60326 313718 60562 313954
rect 60646 313718 60882 313954
rect 60326 313398 60562 313634
rect 60646 313398 60882 313634
rect 60326 277718 60562 277954
rect 60646 277718 60882 277954
rect 60326 277398 60562 277634
rect 60646 277398 60882 277634
rect 60326 241718 60562 241954
rect 60646 241718 60882 241954
rect 60326 241398 60562 241634
rect 60646 241398 60882 241634
rect 60326 205718 60562 205954
rect 60646 205718 60882 205954
rect 60326 205398 60562 205634
rect 60646 205398 60882 205634
rect 60326 169718 60562 169954
rect 60646 169718 60882 169954
rect 60326 169398 60562 169634
rect 60646 169398 60882 169634
rect 60326 133718 60562 133954
rect 60646 133718 60882 133954
rect 60326 133398 60562 133634
rect 60646 133398 60882 133634
rect 60326 97718 60562 97954
rect 60646 97718 60882 97954
rect 60326 97398 60562 97634
rect 60646 97398 60882 97634
rect 60326 61718 60562 61954
rect 60646 61718 60882 61954
rect 60326 61398 60562 61634
rect 60646 61398 60882 61634
rect 60326 25718 60562 25954
rect 60646 25718 60882 25954
rect 60326 25398 60562 25634
rect 60646 25398 60882 25634
rect 60326 -5382 60562 -5146
rect 60646 -5382 60882 -5146
rect 60326 -5702 60562 -5466
rect 60646 -5702 60882 -5466
rect 64826 710362 65062 710598
rect 65146 710362 65382 710598
rect 64826 710042 65062 710278
rect 65146 710042 65382 710278
rect 64826 678218 65062 678454
rect 65146 678218 65382 678454
rect 64826 677898 65062 678134
rect 65146 677898 65382 678134
rect 64826 642218 65062 642454
rect 65146 642218 65382 642454
rect 64826 641898 65062 642134
rect 65146 641898 65382 642134
rect 64826 606218 65062 606454
rect 65146 606218 65382 606454
rect 64826 605898 65062 606134
rect 65146 605898 65382 606134
rect 64826 570218 65062 570454
rect 65146 570218 65382 570454
rect 64826 569898 65062 570134
rect 65146 569898 65382 570134
rect 64826 534218 65062 534454
rect 65146 534218 65382 534454
rect 64826 533898 65062 534134
rect 65146 533898 65382 534134
rect 64826 498218 65062 498454
rect 65146 498218 65382 498454
rect 64826 497898 65062 498134
rect 65146 497898 65382 498134
rect 64826 462218 65062 462454
rect 65146 462218 65382 462454
rect 64826 461898 65062 462134
rect 65146 461898 65382 462134
rect 64826 426218 65062 426454
rect 65146 426218 65382 426454
rect 64826 425898 65062 426134
rect 65146 425898 65382 426134
rect 64826 390218 65062 390454
rect 65146 390218 65382 390454
rect 64826 389898 65062 390134
rect 65146 389898 65382 390134
rect 64826 354218 65062 354454
rect 65146 354218 65382 354454
rect 64826 353898 65062 354134
rect 65146 353898 65382 354134
rect 64826 318218 65062 318454
rect 65146 318218 65382 318454
rect 64826 317898 65062 318134
rect 65146 317898 65382 318134
rect 64826 282218 65062 282454
rect 65146 282218 65382 282454
rect 64826 281898 65062 282134
rect 65146 281898 65382 282134
rect 64826 246218 65062 246454
rect 65146 246218 65382 246454
rect 64826 245898 65062 246134
rect 65146 245898 65382 246134
rect 64826 210218 65062 210454
rect 65146 210218 65382 210454
rect 64826 209898 65062 210134
rect 65146 209898 65382 210134
rect 64826 174218 65062 174454
rect 65146 174218 65382 174454
rect 64826 173898 65062 174134
rect 65146 173898 65382 174134
rect 64826 138218 65062 138454
rect 65146 138218 65382 138454
rect 64826 137898 65062 138134
rect 65146 137898 65382 138134
rect 64826 102218 65062 102454
rect 65146 102218 65382 102454
rect 64826 101898 65062 102134
rect 65146 101898 65382 102134
rect 64826 66218 65062 66454
rect 65146 66218 65382 66454
rect 64826 65898 65062 66134
rect 65146 65898 65382 66134
rect 64826 30218 65062 30454
rect 65146 30218 65382 30454
rect 64826 29898 65062 30134
rect 65146 29898 65382 30134
rect 64826 -6342 65062 -6106
rect 65146 -6342 65382 -6106
rect 64826 -6662 65062 -6426
rect 65146 -6662 65382 -6426
rect 69326 711322 69562 711558
rect 69646 711322 69882 711558
rect 69326 711002 69562 711238
rect 69646 711002 69882 711238
rect 69326 682718 69562 682954
rect 69646 682718 69882 682954
rect 69326 682398 69562 682634
rect 69646 682398 69882 682634
rect 69326 646718 69562 646954
rect 69646 646718 69882 646954
rect 69326 646398 69562 646634
rect 69646 646398 69882 646634
rect 69326 610718 69562 610954
rect 69646 610718 69882 610954
rect 69326 610398 69562 610634
rect 69646 610398 69882 610634
rect 69326 574718 69562 574954
rect 69646 574718 69882 574954
rect 69326 574398 69562 574634
rect 69646 574398 69882 574634
rect 69326 538718 69562 538954
rect 69646 538718 69882 538954
rect 69326 538398 69562 538634
rect 69646 538398 69882 538634
rect 69326 502718 69562 502954
rect 69646 502718 69882 502954
rect 69326 502398 69562 502634
rect 69646 502398 69882 502634
rect 69326 466718 69562 466954
rect 69646 466718 69882 466954
rect 69326 466398 69562 466634
rect 69646 466398 69882 466634
rect 69326 430718 69562 430954
rect 69646 430718 69882 430954
rect 69326 430398 69562 430634
rect 69646 430398 69882 430634
rect 69326 394718 69562 394954
rect 69646 394718 69882 394954
rect 69326 394398 69562 394634
rect 69646 394398 69882 394634
rect 69326 358718 69562 358954
rect 69646 358718 69882 358954
rect 69326 358398 69562 358634
rect 69646 358398 69882 358634
rect 69326 322718 69562 322954
rect 69646 322718 69882 322954
rect 69326 322398 69562 322634
rect 69646 322398 69882 322634
rect 69326 286718 69562 286954
rect 69646 286718 69882 286954
rect 69326 286398 69562 286634
rect 69646 286398 69882 286634
rect 69326 250718 69562 250954
rect 69646 250718 69882 250954
rect 69326 250398 69562 250634
rect 69646 250398 69882 250634
rect 69326 214718 69562 214954
rect 69646 214718 69882 214954
rect 69326 214398 69562 214634
rect 69646 214398 69882 214634
rect 69326 178718 69562 178954
rect 69646 178718 69882 178954
rect 69326 178398 69562 178634
rect 69646 178398 69882 178634
rect 69326 142718 69562 142954
rect 69646 142718 69882 142954
rect 69326 142398 69562 142634
rect 69646 142398 69882 142634
rect 69326 106718 69562 106954
rect 69646 106718 69882 106954
rect 69326 106398 69562 106634
rect 69646 106398 69882 106634
rect 69326 70718 69562 70954
rect 69646 70718 69882 70954
rect 69326 70398 69562 70634
rect 69646 70398 69882 70634
rect 69326 34718 69562 34954
rect 69646 34718 69882 34954
rect 69326 34398 69562 34634
rect 69646 34398 69882 34634
rect 69326 -7302 69562 -7066
rect 69646 -7302 69882 -7066
rect 69326 -7622 69562 -7386
rect 69646 -7622 69882 -7386
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 73826 435218 74062 435454
rect 74146 435218 74382 435454
rect 73826 434898 74062 435134
rect 74146 434898 74382 435134
rect 73826 399218 74062 399454
rect 74146 399218 74382 399454
rect 73826 398898 74062 399134
rect 74146 398898 74382 399134
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 73826 291218 74062 291454
rect 74146 291218 74382 291454
rect 73826 290898 74062 291134
rect 74146 290898 74382 291134
rect 73826 255218 74062 255454
rect 74146 255218 74382 255454
rect 73826 254898 74062 255134
rect 74146 254898 74382 255134
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 73826 147218 74062 147454
rect 74146 147218 74382 147454
rect 73826 146898 74062 147134
rect 74146 146898 74382 147134
rect 73826 111218 74062 111454
rect 74146 111218 74382 111454
rect 73826 110898 74062 111134
rect 74146 110898 74382 111134
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 78326 705562 78562 705798
rect 78646 705562 78882 705798
rect 78326 705242 78562 705478
rect 78646 705242 78882 705478
rect 78326 691718 78562 691954
rect 78646 691718 78882 691954
rect 78326 691398 78562 691634
rect 78646 691398 78882 691634
rect 78326 655718 78562 655954
rect 78646 655718 78882 655954
rect 78326 655398 78562 655634
rect 78646 655398 78882 655634
rect 78326 619718 78562 619954
rect 78646 619718 78882 619954
rect 78326 619398 78562 619634
rect 78646 619398 78882 619634
rect 78326 583718 78562 583954
rect 78646 583718 78882 583954
rect 78326 583398 78562 583634
rect 78646 583398 78882 583634
rect 78326 547718 78562 547954
rect 78646 547718 78882 547954
rect 78326 547398 78562 547634
rect 78646 547398 78882 547634
rect 78326 511718 78562 511954
rect 78646 511718 78882 511954
rect 78326 511398 78562 511634
rect 78646 511398 78882 511634
rect 78326 475718 78562 475954
rect 78646 475718 78882 475954
rect 78326 475398 78562 475634
rect 78646 475398 78882 475634
rect 78326 439718 78562 439954
rect 78646 439718 78882 439954
rect 78326 439398 78562 439634
rect 78646 439398 78882 439634
rect 78326 403718 78562 403954
rect 78646 403718 78882 403954
rect 78326 403398 78562 403634
rect 78646 403398 78882 403634
rect 78326 367718 78562 367954
rect 78646 367718 78882 367954
rect 78326 367398 78562 367634
rect 78646 367398 78882 367634
rect 78326 331718 78562 331954
rect 78646 331718 78882 331954
rect 78326 331398 78562 331634
rect 78646 331398 78882 331634
rect 78326 295718 78562 295954
rect 78646 295718 78882 295954
rect 78326 295398 78562 295634
rect 78646 295398 78882 295634
rect 78326 259718 78562 259954
rect 78646 259718 78882 259954
rect 78326 259398 78562 259634
rect 78646 259398 78882 259634
rect 78326 223718 78562 223954
rect 78646 223718 78882 223954
rect 78326 223398 78562 223634
rect 78646 223398 78882 223634
rect 78326 187718 78562 187954
rect 78646 187718 78882 187954
rect 78326 187398 78562 187634
rect 78646 187398 78882 187634
rect 78326 151718 78562 151954
rect 78646 151718 78882 151954
rect 78326 151398 78562 151634
rect 78646 151398 78882 151634
rect 78326 115718 78562 115954
rect 78646 115718 78882 115954
rect 78326 115398 78562 115634
rect 78646 115398 78882 115634
rect 78326 79718 78562 79954
rect 78646 79718 78882 79954
rect 78326 79398 78562 79634
rect 78646 79398 78882 79634
rect 78326 43718 78562 43954
rect 78646 43718 78882 43954
rect 78326 43398 78562 43634
rect 78646 43398 78882 43634
rect 78326 7718 78562 7954
rect 78646 7718 78882 7954
rect 78326 7398 78562 7634
rect 78646 7398 78882 7634
rect 78326 -1542 78562 -1306
rect 78646 -1542 78882 -1306
rect 78326 -1862 78562 -1626
rect 78646 -1862 78882 -1626
rect 82826 706522 83062 706758
rect 83146 706522 83382 706758
rect 82826 706202 83062 706438
rect 83146 706202 83382 706438
rect 82826 696218 83062 696454
rect 83146 696218 83382 696454
rect 82826 695898 83062 696134
rect 83146 695898 83382 696134
rect 82826 660218 83062 660454
rect 83146 660218 83382 660454
rect 82826 659898 83062 660134
rect 83146 659898 83382 660134
rect 82826 624218 83062 624454
rect 83146 624218 83382 624454
rect 82826 623898 83062 624134
rect 83146 623898 83382 624134
rect 82826 588218 83062 588454
rect 83146 588218 83382 588454
rect 82826 587898 83062 588134
rect 83146 587898 83382 588134
rect 82826 552218 83062 552454
rect 83146 552218 83382 552454
rect 82826 551898 83062 552134
rect 83146 551898 83382 552134
rect 82826 516218 83062 516454
rect 83146 516218 83382 516454
rect 82826 515898 83062 516134
rect 83146 515898 83382 516134
rect 82826 480218 83062 480454
rect 83146 480218 83382 480454
rect 82826 479898 83062 480134
rect 83146 479898 83382 480134
rect 82826 444218 83062 444454
rect 83146 444218 83382 444454
rect 82826 443898 83062 444134
rect 83146 443898 83382 444134
rect 82826 408218 83062 408454
rect 83146 408218 83382 408454
rect 82826 407898 83062 408134
rect 83146 407898 83382 408134
rect 82826 372218 83062 372454
rect 83146 372218 83382 372454
rect 82826 371898 83062 372134
rect 83146 371898 83382 372134
rect 82826 336218 83062 336454
rect 83146 336218 83382 336454
rect 82826 335898 83062 336134
rect 83146 335898 83382 336134
rect 82826 300218 83062 300454
rect 83146 300218 83382 300454
rect 82826 299898 83062 300134
rect 83146 299898 83382 300134
rect 82826 264218 83062 264454
rect 83146 264218 83382 264454
rect 82826 263898 83062 264134
rect 83146 263898 83382 264134
rect 82826 228218 83062 228454
rect 83146 228218 83382 228454
rect 82826 227898 83062 228134
rect 83146 227898 83382 228134
rect 82826 192218 83062 192454
rect 83146 192218 83382 192454
rect 82826 191898 83062 192134
rect 83146 191898 83382 192134
rect 82826 156218 83062 156454
rect 83146 156218 83382 156454
rect 82826 155898 83062 156134
rect 83146 155898 83382 156134
rect 82826 120218 83062 120454
rect 83146 120218 83382 120454
rect 82826 119898 83062 120134
rect 83146 119898 83382 120134
rect 82826 84218 83062 84454
rect 83146 84218 83382 84454
rect 82826 83898 83062 84134
rect 83146 83898 83382 84134
rect 82826 48218 83062 48454
rect 83146 48218 83382 48454
rect 82826 47898 83062 48134
rect 83146 47898 83382 48134
rect 82826 12218 83062 12454
rect 83146 12218 83382 12454
rect 82826 11898 83062 12134
rect 83146 11898 83382 12134
rect 82826 -2502 83062 -2266
rect 83146 -2502 83382 -2266
rect 82826 -2822 83062 -2586
rect 83146 -2822 83382 -2586
rect 87326 707482 87562 707718
rect 87646 707482 87882 707718
rect 87326 707162 87562 707398
rect 87646 707162 87882 707398
rect 87326 700718 87562 700954
rect 87646 700718 87882 700954
rect 87326 700398 87562 700634
rect 87646 700398 87882 700634
rect 87326 664718 87562 664954
rect 87646 664718 87882 664954
rect 87326 664398 87562 664634
rect 87646 664398 87882 664634
rect 87326 628718 87562 628954
rect 87646 628718 87882 628954
rect 87326 628398 87562 628634
rect 87646 628398 87882 628634
rect 87326 592718 87562 592954
rect 87646 592718 87882 592954
rect 87326 592398 87562 592634
rect 87646 592398 87882 592634
rect 87326 556718 87562 556954
rect 87646 556718 87882 556954
rect 87326 556398 87562 556634
rect 87646 556398 87882 556634
rect 87326 520718 87562 520954
rect 87646 520718 87882 520954
rect 87326 520398 87562 520634
rect 87646 520398 87882 520634
rect 87326 484718 87562 484954
rect 87646 484718 87882 484954
rect 87326 484398 87562 484634
rect 87646 484398 87882 484634
rect 87326 448718 87562 448954
rect 87646 448718 87882 448954
rect 87326 448398 87562 448634
rect 87646 448398 87882 448634
rect 87326 412718 87562 412954
rect 87646 412718 87882 412954
rect 87326 412398 87562 412634
rect 87646 412398 87882 412634
rect 87326 376718 87562 376954
rect 87646 376718 87882 376954
rect 87326 376398 87562 376634
rect 87646 376398 87882 376634
rect 87326 340718 87562 340954
rect 87646 340718 87882 340954
rect 87326 340398 87562 340634
rect 87646 340398 87882 340634
rect 87326 304718 87562 304954
rect 87646 304718 87882 304954
rect 87326 304398 87562 304634
rect 87646 304398 87882 304634
rect 87326 268718 87562 268954
rect 87646 268718 87882 268954
rect 87326 268398 87562 268634
rect 87646 268398 87882 268634
rect 87326 232718 87562 232954
rect 87646 232718 87882 232954
rect 87326 232398 87562 232634
rect 87646 232398 87882 232634
rect 87326 196718 87562 196954
rect 87646 196718 87882 196954
rect 87326 196398 87562 196634
rect 87646 196398 87882 196634
rect 87326 160718 87562 160954
rect 87646 160718 87882 160954
rect 87326 160398 87562 160634
rect 87646 160398 87882 160634
rect 87326 124718 87562 124954
rect 87646 124718 87882 124954
rect 87326 124398 87562 124634
rect 87646 124398 87882 124634
rect 87326 88718 87562 88954
rect 87646 88718 87882 88954
rect 87326 88398 87562 88634
rect 87646 88398 87882 88634
rect 87326 52718 87562 52954
rect 87646 52718 87882 52954
rect 87326 52398 87562 52634
rect 87646 52398 87882 52634
rect 87326 16718 87562 16954
rect 87646 16718 87882 16954
rect 87326 16398 87562 16634
rect 87646 16398 87882 16634
rect 87326 -3462 87562 -3226
rect 87646 -3462 87882 -3226
rect 87326 -3782 87562 -3546
rect 87646 -3782 87882 -3546
rect 91826 708442 92062 708678
rect 92146 708442 92382 708678
rect 91826 708122 92062 708358
rect 92146 708122 92382 708358
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 91826 561218 92062 561454
rect 92146 561218 92382 561454
rect 91826 560898 92062 561134
rect 92146 560898 92382 561134
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 91826 453218 92062 453454
rect 92146 453218 92382 453454
rect 91826 452898 92062 453134
rect 92146 452898 92382 453134
rect 91826 417218 92062 417454
rect 92146 417218 92382 417454
rect 91826 416898 92062 417134
rect 92146 416898 92382 417134
rect 91826 381218 92062 381454
rect 92146 381218 92382 381454
rect 91826 380898 92062 381134
rect 92146 380898 92382 381134
rect 91826 345218 92062 345454
rect 92146 345218 92382 345454
rect 91826 344898 92062 345134
rect 92146 344898 92382 345134
rect 91826 309218 92062 309454
rect 92146 309218 92382 309454
rect 91826 308898 92062 309134
rect 92146 308898 92382 309134
rect 91826 273218 92062 273454
rect 92146 273218 92382 273454
rect 91826 272898 92062 273134
rect 92146 272898 92382 273134
rect 91826 237218 92062 237454
rect 92146 237218 92382 237454
rect 91826 236898 92062 237134
rect 92146 236898 92382 237134
rect 91826 201218 92062 201454
rect 92146 201218 92382 201454
rect 91826 200898 92062 201134
rect 92146 200898 92382 201134
rect 91826 165218 92062 165454
rect 92146 165218 92382 165454
rect 91826 164898 92062 165134
rect 92146 164898 92382 165134
rect 91826 129218 92062 129454
rect 92146 129218 92382 129454
rect 91826 128898 92062 129134
rect 92146 128898 92382 129134
rect 91826 93218 92062 93454
rect 92146 93218 92382 93454
rect 91826 92898 92062 93134
rect 92146 92898 92382 93134
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -4422 92062 -4186
rect 92146 -4422 92382 -4186
rect 91826 -4742 92062 -4506
rect 92146 -4742 92382 -4506
rect 96326 709402 96562 709638
rect 96646 709402 96882 709638
rect 96326 709082 96562 709318
rect 96646 709082 96882 709318
rect 96326 673718 96562 673954
rect 96646 673718 96882 673954
rect 96326 673398 96562 673634
rect 96646 673398 96882 673634
rect 96326 637718 96562 637954
rect 96646 637718 96882 637954
rect 96326 637398 96562 637634
rect 96646 637398 96882 637634
rect 96326 601718 96562 601954
rect 96646 601718 96882 601954
rect 96326 601398 96562 601634
rect 96646 601398 96882 601634
rect 96326 565718 96562 565954
rect 96646 565718 96882 565954
rect 96326 565398 96562 565634
rect 96646 565398 96882 565634
rect 96326 529718 96562 529954
rect 96646 529718 96882 529954
rect 96326 529398 96562 529634
rect 96646 529398 96882 529634
rect 96326 493718 96562 493954
rect 96646 493718 96882 493954
rect 96326 493398 96562 493634
rect 96646 493398 96882 493634
rect 96326 457718 96562 457954
rect 96646 457718 96882 457954
rect 96326 457398 96562 457634
rect 96646 457398 96882 457634
rect 96326 421718 96562 421954
rect 96646 421718 96882 421954
rect 96326 421398 96562 421634
rect 96646 421398 96882 421634
rect 96326 385718 96562 385954
rect 96646 385718 96882 385954
rect 96326 385398 96562 385634
rect 96646 385398 96882 385634
rect 96326 349718 96562 349954
rect 96646 349718 96882 349954
rect 96326 349398 96562 349634
rect 96646 349398 96882 349634
rect 96326 313718 96562 313954
rect 96646 313718 96882 313954
rect 96326 313398 96562 313634
rect 96646 313398 96882 313634
rect 96326 277718 96562 277954
rect 96646 277718 96882 277954
rect 96326 277398 96562 277634
rect 96646 277398 96882 277634
rect 96326 241718 96562 241954
rect 96646 241718 96882 241954
rect 96326 241398 96562 241634
rect 96646 241398 96882 241634
rect 96326 205718 96562 205954
rect 96646 205718 96882 205954
rect 96326 205398 96562 205634
rect 96646 205398 96882 205634
rect 96326 169718 96562 169954
rect 96646 169718 96882 169954
rect 96326 169398 96562 169634
rect 96646 169398 96882 169634
rect 96326 133718 96562 133954
rect 96646 133718 96882 133954
rect 96326 133398 96562 133634
rect 96646 133398 96882 133634
rect 96326 97718 96562 97954
rect 96646 97718 96882 97954
rect 96326 97398 96562 97634
rect 96646 97398 96882 97634
rect 96326 61718 96562 61954
rect 96646 61718 96882 61954
rect 96326 61398 96562 61634
rect 96646 61398 96882 61634
rect 96326 25718 96562 25954
rect 96646 25718 96882 25954
rect 96326 25398 96562 25634
rect 96646 25398 96882 25634
rect 96326 -5382 96562 -5146
rect 96646 -5382 96882 -5146
rect 96326 -5702 96562 -5466
rect 96646 -5702 96882 -5466
rect 100826 710362 101062 710598
rect 101146 710362 101382 710598
rect 100826 710042 101062 710278
rect 101146 710042 101382 710278
rect 100826 678218 101062 678454
rect 101146 678218 101382 678454
rect 100826 677898 101062 678134
rect 101146 677898 101382 678134
rect 100826 642218 101062 642454
rect 101146 642218 101382 642454
rect 100826 641898 101062 642134
rect 101146 641898 101382 642134
rect 100826 606218 101062 606454
rect 101146 606218 101382 606454
rect 100826 605898 101062 606134
rect 101146 605898 101382 606134
rect 100826 570218 101062 570454
rect 101146 570218 101382 570454
rect 100826 569898 101062 570134
rect 101146 569898 101382 570134
rect 100826 534218 101062 534454
rect 101146 534218 101382 534454
rect 100826 533898 101062 534134
rect 101146 533898 101382 534134
rect 100826 498218 101062 498454
rect 101146 498218 101382 498454
rect 100826 497898 101062 498134
rect 101146 497898 101382 498134
rect 100826 462218 101062 462454
rect 101146 462218 101382 462454
rect 100826 461898 101062 462134
rect 101146 461898 101382 462134
rect 100826 426218 101062 426454
rect 101146 426218 101382 426454
rect 100826 425898 101062 426134
rect 101146 425898 101382 426134
rect 100826 390218 101062 390454
rect 101146 390218 101382 390454
rect 100826 389898 101062 390134
rect 101146 389898 101382 390134
rect 100826 354218 101062 354454
rect 101146 354218 101382 354454
rect 100826 353898 101062 354134
rect 101146 353898 101382 354134
rect 100826 318218 101062 318454
rect 101146 318218 101382 318454
rect 100826 317898 101062 318134
rect 101146 317898 101382 318134
rect 100826 282218 101062 282454
rect 101146 282218 101382 282454
rect 100826 281898 101062 282134
rect 101146 281898 101382 282134
rect 100826 246218 101062 246454
rect 101146 246218 101382 246454
rect 100826 245898 101062 246134
rect 101146 245898 101382 246134
rect 100826 210218 101062 210454
rect 101146 210218 101382 210454
rect 100826 209898 101062 210134
rect 101146 209898 101382 210134
rect 100826 174218 101062 174454
rect 101146 174218 101382 174454
rect 100826 173898 101062 174134
rect 101146 173898 101382 174134
rect 100826 138218 101062 138454
rect 101146 138218 101382 138454
rect 100826 137898 101062 138134
rect 101146 137898 101382 138134
rect 100826 102218 101062 102454
rect 101146 102218 101382 102454
rect 100826 101898 101062 102134
rect 101146 101898 101382 102134
rect 100826 66218 101062 66454
rect 101146 66218 101382 66454
rect 100826 65898 101062 66134
rect 101146 65898 101382 66134
rect 100826 30218 101062 30454
rect 101146 30218 101382 30454
rect 100826 29898 101062 30134
rect 101146 29898 101382 30134
rect 100826 -6342 101062 -6106
rect 101146 -6342 101382 -6106
rect 100826 -6662 101062 -6426
rect 101146 -6662 101382 -6426
rect 105326 711322 105562 711558
rect 105646 711322 105882 711558
rect 105326 711002 105562 711238
rect 105646 711002 105882 711238
rect 105326 682718 105562 682954
rect 105646 682718 105882 682954
rect 105326 682398 105562 682634
rect 105646 682398 105882 682634
rect 105326 646718 105562 646954
rect 105646 646718 105882 646954
rect 105326 646398 105562 646634
rect 105646 646398 105882 646634
rect 105326 610718 105562 610954
rect 105646 610718 105882 610954
rect 105326 610398 105562 610634
rect 105646 610398 105882 610634
rect 105326 574718 105562 574954
rect 105646 574718 105882 574954
rect 105326 574398 105562 574634
rect 105646 574398 105882 574634
rect 105326 538718 105562 538954
rect 105646 538718 105882 538954
rect 105326 538398 105562 538634
rect 105646 538398 105882 538634
rect 105326 502718 105562 502954
rect 105646 502718 105882 502954
rect 105326 502398 105562 502634
rect 105646 502398 105882 502634
rect 105326 466718 105562 466954
rect 105646 466718 105882 466954
rect 105326 466398 105562 466634
rect 105646 466398 105882 466634
rect 105326 430718 105562 430954
rect 105646 430718 105882 430954
rect 105326 430398 105562 430634
rect 105646 430398 105882 430634
rect 105326 394718 105562 394954
rect 105646 394718 105882 394954
rect 105326 394398 105562 394634
rect 105646 394398 105882 394634
rect 105326 358718 105562 358954
rect 105646 358718 105882 358954
rect 105326 358398 105562 358634
rect 105646 358398 105882 358634
rect 105326 322718 105562 322954
rect 105646 322718 105882 322954
rect 105326 322398 105562 322634
rect 105646 322398 105882 322634
rect 105326 286718 105562 286954
rect 105646 286718 105882 286954
rect 105326 286398 105562 286634
rect 105646 286398 105882 286634
rect 105326 250718 105562 250954
rect 105646 250718 105882 250954
rect 105326 250398 105562 250634
rect 105646 250398 105882 250634
rect 105326 214718 105562 214954
rect 105646 214718 105882 214954
rect 105326 214398 105562 214634
rect 105646 214398 105882 214634
rect 105326 178718 105562 178954
rect 105646 178718 105882 178954
rect 105326 178398 105562 178634
rect 105646 178398 105882 178634
rect 105326 142718 105562 142954
rect 105646 142718 105882 142954
rect 105326 142398 105562 142634
rect 105646 142398 105882 142634
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 109826 435218 110062 435454
rect 110146 435218 110382 435454
rect 109826 434898 110062 435134
rect 110146 434898 110382 435134
rect 109826 399218 110062 399454
rect 110146 399218 110382 399454
rect 109826 398898 110062 399134
rect 110146 398898 110382 399134
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 109826 327218 110062 327454
rect 110146 327218 110382 327454
rect 109826 326898 110062 327134
rect 110146 326898 110382 327134
rect 109826 291218 110062 291454
rect 110146 291218 110382 291454
rect 109826 290898 110062 291134
rect 110146 290898 110382 291134
rect 114326 705562 114562 705798
rect 114646 705562 114882 705798
rect 114326 705242 114562 705478
rect 114646 705242 114882 705478
rect 114326 691718 114562 691954
rect 114646 691718 114882 691954
rect 114326 691398 114562 691634
rect 114646 691398 114882 691634
rect 114326 655718 114562 655954
rect 114646 655718 114882 655954
rect 114326 655398 114562 655634
rect 114646 655398 114882 655634
rect 114326 619718 114562 619954
rect 114646 619718 114882 619954
rect 114326 619398 114562 619634
rect 114646 619398 114882 619634
rect 114326 583718 114562 583954
rect 114646 583718 114882 583954
rect 114326 583398 114562 583634
rect 114646 583398 114882 583634
rect 114326 547718 114562 547954
rect 114646 547718 114882 547954
rect 114326 547398 114562 547634
rect 114646 547398 114882 547634
rect 114326 511718 114562 511954
rect 114646 511718 114882 511954
rect 114326 511398 114562 511634
rect 114646 511398 114882 511634
rect 114326 475718 114562 475954
rect 114646 475718 114882 475954
rect 114326 475398 114562 475634
rect 114646 475398 114882 475634
rect 114326 439718 114562 439954
rect 114646 439718 114882 439954
rect 114326 439398 114562 439634
rect 114646 439398 114882 439634
rect 114326 403718 114562 403954
rect 114646 403718 114882 403954
rect 114326 403398 114562 403634
rect 114646 403398 114882 403634
rect 114326 367718 114562 367954
rect 114646 367718 114882 367954
rect 114326 367398 114562 367634
rect 114646 367398 114882 367634
rect 114326 331718 114562 331954
rect 114646 331718 114882 331954
rect 114326 331398 114562 331634
rect 114646 331398 114882 331634
rect 114326 295718 114562 295954
rect 114646 295718 114882 295954
rect 114326 295398 114562 295634
rect 114646 295398 114882 295634
rect 109826 255218 110062 255454
rect 110146 255218 110382 255454
rect 109826 254898 110062 255134
rect 110146 254898 110382 255134
rect 109826 219218 110062 219454
rect 110146 219218 110382 219454
rect 109826 218898 110062 219134
rect 110146 218898 110382 219134
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 109826 147218 110062 147454
rect 110146 147218 110382 147454
rect 109826 146898 110062 147134
rect 110146 146898 110382 147134
rect 105326 106718 105562 106954
rect 105646 106718 105882 106954
rect 105326 106398 105562 106634
rect 105646 106398 105882 106634
rect 105326 70718 105562 70954
rect 105646 70718 105882 70954
rect 105326 70398 105562 70634
rect 105646 70398 105882 70634
rect 105326 34718 105562 34954
rect 105646 34718 105882 34954
rect 105326 34398 105562 34634
rect 105646 34398 105882 34634
rect 109826 111218 110062 111454
rect 110146 111218 110382 111454
rect 109826 110898 110062 111134
rect 110146 110898 110382 111134
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 118826 706522 119062 706758
rect 119146 706522 119382 706758
rect 118826 706202 119062 706438
rect 119146 706202 119382 706438
rect 118826 696218 119062 696454
rect 119146 696218 119382 696454
rect 118826 695898 119062 696134
rect 119146 695898 119382 696134
rect 118826 660218 119062 660454
rect 119146 660218 119382 660454
rect 118826 659898 119062 660134
rect 119146 659898 119382 660134
rect 118826 624218 119062 624454
rect 119146 624218 119382 624454
rect 118826 623898 119062 624134
rect 119146 623898 119382 624134
rect 118826 588218 119062 588454
rect 119146 588218 119382 588454
rect 118826 587898 119062 588134
rect 119146 587898 119382 588134
rect 118826 552218 119062 552454
rect 119146 552218 119382 552454
rect 118826 551898 119062 552134
rect 119146 551898 119382 552134
rect 118826 516218 119062 516454
rect 119146 516218 119382 516454
rect 118826 515898 119062 516134
rect 119146 515898 119382 516134
rect 118826 480218 119062 480454
rect 119146 480218 119382 480454
rect 118826 479898 119062 480134
rect 119146 479898 119382 480134
rect 118826 444218 119062 444454
rect 119146 444218 119382 444454
rect 118826 443898 119062 444134
rect 119146 443898 119382 444134
rect 118826 408218 119062 408454
rect 119146 408218 119382 408454
rect 118826 407898 119062 408134
rect 119146 407898 119382 408134
rect 118826 372218 119062 372454
rect 119146 372218 119382 372454
rect 118826 371898 119062 372134
rect 119146 371898 119382 372134
rect 118826 336218 119062 336454
rect 119146 336218 119382 336454
rect 118826 335898 119062 336134
rect 119146 335898 119382 336134
rect 118826 300218 119062 300454
rect 119146 300218 119382 300454
rect 118826 299898 119062 300134
rect 119146 299898 119382 300134
rect 118826 264218 119062 264454
rect 119146 264218 119382 264454
rect 118826 263898 119062 264134
rect 119146 263898 119382 264134
rect 114326 259718 114562 259954
rect 114646 259718 114882 259954
rect 114326 259398 114562 259634
rect 114646 259398 114882 259634
rect 114326 223718 114562 223954
rect 114646 223718 114882 223954
rect 114326 223398 114562 223634
rect 114646 223398 114882 223634
rect 114326 187718 114562 187954
rect 114646 187718 114882 187954
rect 114326 187398 114562 187634
rect 114646 187398 114882 187634
rect 114326 151718 114562 151954
rect 114646 151718 114882 151954
rect 114326 151398 114562 151634
rect 114646 151398 114882 151634
rect 114326 115718 114562 115954
rect 114646 115718 114882 115954
rect 114326 115398 114562 115634
rect 114646 115398 114882 115634
rect 114326 79718 114562 79954
rect 114646 79718 114882 79954
rect 114326 79398 114562 79634
rect 114646 79398 114882 79634
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 105326 -7302 105562 -7066
rect 105646 -7302 105882 -7066
rect 105326 -7622 105562 -7386
rect 105646 -7622 105882 -7386
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 123326 707482 123562 707718
rect 123646 707482 123882 707718
rect 123326 707162 123562 707398
rect 123646 707162 123882 707398
rect 123326 700718 123562 700954
rect 123646 700718 123882 700954
rect 123326 700398 123562 700634
rect 123646 700398 123882 700634
rect 123326 664718 123562 664954
rect 123646 664718 123882 664954
rect 123326 664398 123562 664634
rect 123646 664398 123882 664634
rect 123326 628718 123562 628954
rect 123646 628718 123882 628954
rect 123326 628398 123562 628634
rect 123646 628398 123882 628634
rect 123326 592718 123562 592954
rect 123646 592718 123882 592954
rect 123326 592398 123562 592634
rect 123646 592398 123882 592634
rect 123326 556718 123562 556954
rect 123646 556718 123882 556954
rect 123326 556398 123562 556634
rect 123646 556398 123882 556634
rect 123326 520718 123562 520954
rect 123646 520718 123882 520954
rect 123326 520398 123562 520634
rect 123646 520398 123882 520634
rect 123326 484718 123562 484954
rect 123646 484718 123882 484954
rect 123326 484398 123562 484634
rect 123646 484398 123882 484634
rect 123326 448718 123562 448954
rect 123646 448718 123882 448954
rect 123326 448398 123562 448634
rect 123646 448398 123882 448634
rect 123326 412718 123562 412954
rect 123646 412718 123882 412954
rect 123326 412398 123562 412634
rect 123646 412398 123882 412634
rect 123326 376718 123562 376954
rect 123646 376718 123882 376954
rect 123326 376398 123562 376634
rect 123646 376398 123882 376634
rect 123326 340718 123562 340954
rect 123646 340718 123882 340954
rect 123326 340398 123562 340634
rect 123646 340398 123882 340634
rect 123326 304718 123562 304954
rect 123646 304718 123882 304954
rect 123326 304398 123562 304634
rect 123646 304398 123882 304634
rect 123326 268718 123562 268954
rect 123646 268718 123882 268954
rect 123326 268398 123562 268634
rect 123646 268398 123882 268634
rect 118826 192218 119062 192454
rect 119146 192218 119382 192454
rect 118826 191898 119062 192134
rect 119146 191898 119382 192134
rect 118826 156218 119062 156454
rect 119146 156218 119382 156454
rect 118826 155898 119062 156134
rect 119146 155898 119382 156134
rect 114326 43718 114562 43954
rect 114646 43718 114882 43954
rect 114326 43398 114562 43634
rect 114646 43398 114882 43634
rect 127826 708442 128062 708678
rect 128146 708442 128382 708678
rect 127826 708122 128062 708358
rect 128146 708122 128382 708358
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 127826 453218 128062 453454
rect 128146 453218 128382 453454
rect 127826 452898 128062 453134
rect 128146 452898 128382 453134
rect 127826 417218 128062 417454
rect 128146 417218 128382 417454
rect 127826 416898 128062 417134
rect 128146 416898 128382 417134
rect 127826 381218 128062 381454
rect 128146 381218 128382 381454
rect 127826 380898 128062 381134
rect 128146 380898 128382 381134
rect 127826 345218 128062 345454
rect 128146 345218 128382 345454
rect 127826 344898 128062 345134
rect 128146 344898 128382 345134
rect 127826 309218 128062 309454
rect 128146 309218 128382 309454
rect 127826 308898 128062 309134
rect 128146 308898 128382 309134
rect 127826 273218 128062 273454
rect 128146 273218 128382 273454
rect 127826 272898 128062 273134
rect 128146 272898 128382 273134
rect 132326 709402 132562 709638
rect 132646 709402 132882 709638
rect 132326 709082 132562 709318
rect 132646 709082 132882 709318
rect 132326 673718 132562 673954
rect 132646 673718 132882 673954
rect 132326 673398 132562 673634
rect 132646 673398 132882 673634
rect 132326 637718 132562 637954
rect 132646 637718 132882 637954
rect 132326 637398 132562 637634
rect 132646 637398 132882 637634
rect 132326 601718 132562 601954
rect 132646 601718 132882 601954
rect 132326 601398 132562 601634
rect 132646 601398 132882 601634
rect 132326 565718 132562 565954
rect 132646 565718 132882 565954
rect 132326 565398 132562 565634
rect 132646 565398 132882 565634
rect 132326 529718 132562 529954
rect 132646 529718 132882 529954
rect 132326 529398 132562 529634
rect 132646 529398 132882 529634
rect 132326 493718 132562 493954
rect 132646 493718 132882 493954
rect 132326 493398 132562 493634
rect 132646 493398 132882 493634
rect 132326 457718 132562 457954
rect 132646 457718 132882 457954
rect 132326 457398 132562 457634
rect 132646 457398 132882 457634
rect 132326 421718 132562 421954
rect 132646 421718 132882 421954
rect 132326 421398 132562 421634
rect 132646 421398 132882 421634
rect 132326 385718 132562 385954
rect 132646 385718 132882 385954
rect 132326 385398 132562 385634
rect 132646 385398 132882 385634
rect 132326 349718 132562 349954
rect 132646 349718 132882 349954
rect 132326 349398 132562 349634
rect 132646 349398 132882 349634
rect 132326 313718 132562 313954
rect 132646 313718 132882 313954
rect 132326 313398 132562 313634
rect 132646 313398 132882 313634
rect 132326 277718 132562 277954
rect 132646 277718 132882 277954
rect 132326 277398 132562 277634
rect 132646 277398 132882 277634
rect 136826 710362 137062 710598
rect 137146 710362 137382 710598
rect 136826 710042 137062 710278
rect 137146 710042 137382 710278
rect 136826 678218 137062 678454
rect 137146 678218 137382 678454
rect 136826 677898 137062 678134
rect 137146 677898 137382 678134
rect 136826 642218 137062 642454
rect 137146 642218 137382 642454
rect 136826 641898 137062 642134
rect 137146 641898 137382 642134
rect 136826 606218 137062 606454
rect 137146 606218 137382 606454
rect 136826 605898 137062 606134
rect 137146 605898 137382 606134
rect 136826 570218 137062 570454
rect 137146 570218 137382 570454
rect 136826 569898 137062 570134
rect 137146 569898 137382 570134
rect 136826 534218 137062 534454
rect 137146 534218 137382 534454
rect 136826 533898 137062 534134
rect 137146 533898 137382 534134
rect 136826 498218 137062 498454
rect 137146 498218 137382 498454
rect 136826 497898 137062 498134
rect 137146 497898 137382 498134
rect 136826 462218 137062 462454
rect 137146 462218 137382 462454
rect 136826 461898 137062 462134
rect 137146 461898 137382 462134
rect 136826 426218 137062 426454
rect 137146 426218 137382 426454
rect 136826 425898 137062 426134
rect 137146 425898 137382 426134
rect 136826 390218 137062 390454
rect 137146 390218 137382 390454
rect 136826 389898 137062 390134
rect 137146 389898 137382 390134
rect 136826 354218 137062 354454
rect 137146 354218 137382 354454
rect 136826 353898 137062 354134
rect 137146 353898 137382 354134
rect 136826 318218 137062 318454
rect 137146 318218 137382 318454
rect 136826 317898 137062 318134
rect 137146 317898 137382 318134
rect 136826 282218 137062 282454
rect 137146 282218 137382 282454
rect 136826 281898 137062 282134
rect 137146 281898 137382 282134
rect 141326 711322 141562 711558
rect 141646 711322 141882 711558
rect 141326 711002 141562 711238
rect 141646 711002 141882 711238
rect 141326 682718 141562 682954
rect 141646 682718 141882 682954
rect 141326 682398 141562 682634
rect 141646 682398 141882 682634
rect 141326 646718 141562 646954
rect 141646 646718 141882 646954
rect 141326 646398 141562 646634
rect 141646 646398 141882 646634
rect 141326 610718 141562 610954
rect 141646 610718 141882 610954
rect 141326 610398 141562 610634
rect 141646 610398 141882 610634
rect 141326 574718 141562 574954
rect 141646 574718 141882 574954
rect 141326 574398 141562 574634
rect 141646 574398 141882 574634
rect 141326 538718 141562 538954
rect 141646 538718 141882 538954
rect 141326 538398 141562 538634
rect 141646 538398 141882 538634
rect 141326 502718 141562 502954
rect 141646 502718 141882 502954
rect 141326 502398 141562 502634
rect 141646 502398 141882 502634
rect 141326 466718 141562 466954
rect 141646 466718 141882 466954
rect 141326 466398 141562 466634
rect 141646 466398 141882 466634
rect 141326 430718 141562 430954
rect 141646 430718 141882 430954
rect 141326 430398 141562 430634
rect 141646 430398 141882 430634
rect 141326 394718 141562 394954
rect 141646 394718 141882 394954
rect 141326 394398 141562 394634
rect 141646 394398 141882 394634
rect 141326 358718 141562 358954
rect 141646 358718 141882 358954
rect 141326 358398 141562 358634
rect 141646 358398 141882 358634
rect 141326 322718 141562 322954
rect 141646 322718 141882 322954
rect 141326 322398 141562 322634
rect 141646 322398 141882 322634
rect 141326 286718 141562 286954
rect 141646 286718 141882 286954
rect 141326 286398 141562 286634
rect 141646 286398 141882 286634
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 150326 705562 150562 705798
rect 150646 705562 150882 705798
rect 150326 705242 150562 705478
rect 150646 705242 150882 705478
rect 150326 691718 150562 691954
rect 150646 691718 150882 691954
rect 150326 691398 150562 691634
rect 150646 691398 150882 691634
rect 150326 655718 150562 655954
rect 150646 655718 150882 655954
rect 150326 655398 150562 655634
rect 150646 655398 150882 655634
rect 150326 619718 150562 619954
rect 150646 619718 150882 619954
rect 150326 619398 150562 619634
rect 150646 619398 150882 619634
rect 150326 583718 150562 583954
rect 150646 583718 150882 583954
rect 150326 583398 150562 583634
rect 150646 583398 150882 583634
rect 150326 547718 150562 547954
rect 150646 547718 150882 547954
rect 150326 547398 150562 547634
rect 150646 547398 150882 547634
rect 150326 511718 150562 511954
rect 150646 511718 150882 511954
rect 150326 511398 150562 511634
rect 150646 511398 150882 511634
rect 150326 475718 150562 475954
rect 150646 475718 150882 475954
rect 150326 475398 150562 475634
rect 150646 475398 150882 475634
rect 150326 439718 150562 439954
rect 150646 439718 150882 439954
rect 150326 439398 150562 439634
rect 150646 439398 150882 439634
rect 150326 403718 150562 403954
rect 150646 403718 150882 403954
rect 150326 403398 150562 403634
rect 150646 403398 150882 403634
rect 150326 367718 150562 367954
rect 150646 367718 150882 367954
rect 150326 367398 150562 367634
rect 150646 367398 150882 367634
rect 150326 331718 150562 331954
rect 150646 331718 150882 331954
rect 150326 331398 150562 331634
rect 150646 331398 150882 331634
rect 150326 295718 150562 295954
rect 150646 295718 150882 295954
rect 150326 295398 150562 295634
rect 150646 295398 150882 295634
rect 154826 706522 155062 706758
rect 155146 706522 155382 706758
rect 154826 706202 155062 706438
rect 155146 706202 155382 706438
rect 154826 696218 155062 696454
rect 155146 696218 155382 696454
rect 154826 695898 155062 696134
rect 155146 695898 155382 696134
rect 154826 660218 155062 660454
rect 155146 660218 155382 660454
rect 154826 659898 155062 660134
rect 155146 659898 155382 660134
rect 154826 624218 155062 624454
rect 155146 624218 155382 624454
rect 154826 623898 155062 624134
rect 155146 623898 155382 624134
rect 154826 588218 155062 588454
rect 155146 588218 155382 588454
rect 154826 587898 155062 588134
rect 155146 587898 155382 588134
rect 154826 552218 155062 552454
rect 155146 552218 155382 552454
rect 154826 551898 155062 552134
rect 155146 551898 155382 552134
rect 154826 516218 155062 516454
rect 155146 516218 155382 516454
rect 154826 515898 155062 516134
rect 155146 515898 155382 516134
rect 154826 480218 155062 480454
rect 155146 480218 155382 480454
rect 154826 479898 155062 480134
rect 155146 479898 155382 480134
rect 154826 444218 155062 444454
rect 155146 444218 155382 444454
rect 154826 443898 155062 444134
rect 155146 443898 155382 444134
rect 154826 408218 155062 408454
rect 155146 408218 155382 408454
rect 154826 407898 155062 408134
rect 155146 407898 155382 408134
rect 154826 372218 155062 372454
rect 155146 372218 155382 372454
rect 154826 371898 155062 372134
rect 155146 371898 155382 372134
rect 154826 336218 155062 336454
rect 155146 336218 155382 336454
rect 154826 335898 155062 336134
rect 155146 335898 155382 336134
rect 154826 300218 155062 300454
rect 155146 300218 155382 300454
rect 154826 299898 155062 300134
rect 155146 299898 155382 300134
rect 154826 264218 155062 264454
rect 155146 264218 155382 264454
rect 154826 263898 155062 264134
rect 155146 263898 155382 264134
rect 159326 707482 159562 707718
rect 159646 707482 159882 707718
rect 159326 707162 159562 707398
rect 159646 707162 159882 707398
rect 159326 700718 159562 700954
rect 159646 700718 159882 700954
rect 159326 700398 159562 700634
rect 159646 700398 159882 700634
rect 159326 664718 159562 664954
rect 159646 664718 159882 664954
rect 159326 664398 159562 664634
rect 159646 664398 159882 664634
rect 159326 628718 159562 628954
rect 159646 628718 159882 628954
rect 159326 628398 159562 628634
rect 159646 628398 159882 628634
rect 159326 592718 159562 592954
rect 159646 592718 159882 592954
rect 159326 592398 159562 592634
rect 159646 592398 159882 592634
rect 159326 556718 159562 556954
rect 159646 556718 159882 556954
rect 159326 556398 159562 556634
rect 159646 556398 159882 556634
rect 159326 520718 159562 520954
rect 159646 520718 159882 520954
rect 159326 520398 159562 520634
rect 159646 520398 159882 520634
rect 159326 484718 159562 484954
rect 159646 484718 159882 484954
rect 159326 484398 159562 484634
rect 159646 484398 159882 484634
rect 159326 448718 159562 448954
rect 159646 448718 159882 448954
rect 159326 448398 159562 448634
rect 159646 448398 159882 448634
rect 159326 412718 159562 412954
rect 159646 412718 159882 412954
rect 159326 412398 159562 412634
rect 159646 412398 159882 412634
rect 159326 376718 159562 376954
rect 159646 376718 159882 376954
rect 159326 376398 159562 376634
rect 159646 376398 159882 376634
rect 159326 340718 159562 340954
rect 159646 340718 159882 340954
rect 159326 340398 159562 340634
rect 159646 340398 159882 340634
rect 159326 304718 159562 304954
rect 159646 304718 159882 304954
rect 159326 304398 159562 304634
rect 159646 304398 159882 304634
rect 159326 268718 159562 268954
rect 159646 268718 159882 268954
rect 159326 268398 159562 268634
rect 159646 268398 159882 268634
rect 163826 708442 164062 708678
rect 164146 708442 164382 708678
rect 163826 708122 164062 708358
rect 164146 708122 164382 708358
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 163826 453218 164062 453454
rect 164146 453218 164382 453454
rect 163826 452898 164062 453134
rect 164146 452898 164382 453134
rect 163826 417218 164062 417454
rect 164146 417218 164382 417454
rect 163826 416898 164062 417134
rect 164146 416898 164382 417134
rect 163826 381218 164062 381454
rect 164146 381218 164382 381454
rect 163826 380898 164062 381134
rect 164146 380898 164382 381134
rect 163826 345218 164062 345454
rect 164146 345218 164382 345454
rect 163826 344898 164062 345134
rect 164146 344898 164382 345134
rect 163826 309218 164062 309454
rect 164146 309218 164382 309454
rect 163826 308898 164062 309134
rect 164146 308898 164382 309134
rect 163826 273218 164062 273454
rect 164146 273218 164382 273454
rect 163826 272898 164062 273134
rect 164146 272898 164382 273134
rect 168326 709402 168562 709638
rect 168646 709402 168882 709638
rect 168326 709082 168562 709318
rect 168646 709082 168882 709318
rect 168326 673718 168562 673954
rect 168646 673718 168882 673954
rect 168326 673398 168562 673634
rect 168646 673398 168882 673634
rect 168326 637718 168562 637954
rect 168646 637718 168882 637954
rect 168326 637398 168562 637634
rect 168646 637398 168882 637634
rect 168326 601718 168562 601954
rect 168646 601718 168882 601954
rect 168326 601398 168562 601634
rect 168646 601398 168882 601634
rect 168326 565718 168562 565954
rect 168646 565718 168882 565954
rect 168326 565398 168562 565634
rect 168646 565398 168882 565634
rect 168326 529718 168562 529954
rect 168646 529718 168882 529954
rect 168326 529398 168562 529634
rect 168646 529398 168882 529634
rect 168326 493718 168562 493954
rect 168646 493718 168882 493954
rect 168326 493398 168562 493634
rect 168646 493398 168882 493634
rect 168326 457718 168562 457954
rect 168646 457718 168882 457954
rect 168326 457398 168562 457634
rect 168646 457398 168882 457634
rect 168326 421718 168562 421954
rect 168646 421718 168882 421954
rect 168326 421398 168562 421634
rect 168646 421398 168882 421634
rect 168326 385718 168562 385954
rect 168646 385718 168882 385954
rect 168326 385398 168562 385634
rect 168646 385398 168882 385634
rect 168326 349718 168562 349954
rect 168646 349718 168882 349954
rect 168326 349398 168562 349634
rect 168646 349398 168882 349634
rect 168326 313718 168562 313954
rect 168646 313718 168882 313954
rect 168326 313398 168562 313634
rect 168646 313398 168882 313634
rect 168326 277718 168562 277954
rect 168646 277718 168882 277954
rect 168326 277398 168562 277634
rect 168646 277398 168882 277634
rect 172826 710362 173062 710598
rect 173146 710362 173382 710598
rect 172826 710042 173062 710278
rect 173146 710042 173382 710278
rect 172826 678218 173062 678454
rect 173146 678218 173382 678454
rect 172826 677898 173062 678134
rect 173146 677898 173382 678134
rect 172826 642218 173062 642454
rect 173146 642218 173382 642454
rect 172826 641898 173062 642134
rect 173146 641898 173382 642134
rect 172826 606218 173062 606454
rect 173146 606218 173382 606454
rect 172826 605898 173062 606134
rect 173146 605898 173382 606134
rect 172826 570218 173062 570454
rect 173146 570218 173382 570454
rect 172826 569898 173062 570134
rect 173146 569898 173382 570134
rect 172826 534218 173062 534454
rect 173146 534218 173382 534454
rect 172826 533898 173062 534134
rect 173146 533898 173382 534134
rect 172826 498218 173062 498454
rect 173146 498218 173382 498454
rect 172826 497898 173062 498134
rect 173146 497898 173382 498134
rect 172826 462218 173062 462454
rect 173146 462218 173382 462454
rect 172826 461898 173062 462134
rect 173146 461898 173382 462134
rect 172826 426218 173062 426454
rect 173146 426218 173382 426454
rect 172826 425898 173062 426134
rect 173146 425898 173382 426134
rect 172826 390218 173062 390454
rect 173146 390218 173382 390454
rect 172826 389898 173062 390134
rect 173146 389898 173382 390134
rect 172826 354218 173062 354454
rect 173146 354218 173382 354454
rect 172826 353898 173062 354134
rect 173146 353898 173382 354134
rect 172826 318218 173062 318454
rect 173146 318218 173382 318454
rect 172826 317898 173062 318134
rect 173146 317898 173382 318134
rect 172826 282218 173062 282454
rect 173146 282218 173382 282454
rect 172826 281898 173062 282134
rect 173146 281898 173382 282134
rect 177326 711322 177562 711558
rect 177646 711322 177882 711558
rect 177326 711002 177562 711238
rect 177646 711002 177882 711238
rect 177326 682718 177562 682954
rect 177646 682718 177882 682954
rect 177326 682398 177562 682634
rect 177646 682398 177882 682634
rect 177326 646718 177562 646954
rect 177646 646718 177882 646954
rect 177326 646398 177562 646634
rect 177646 646398 177882 646634
rect 177326 610718 177562 610954
rect 177646 610718 177882 610954
rect 177326 610398 177562 610634
rect 177646 610398 177882 610634
rect 177326 574718 177562 574954
rect 177646 574718 177882 574954
rect 177326 574398 177562 574634
rect 177646 574398 177882 574634
rect 177326 538718 177562 538954
rect 177646 538718 177882 538954
rect 177326 538398 177562 538634
rect 177646 538398 177882 538634
rect 177326 502718 177562 502954
rect 177646 502718 177882 502954
rect 177326 502398 177562 502634
rect 177646 502398 177882 502634
rect 177326 466718 177562 466954
rect 177646 466718 177882 466954
rect 177326 466398 177562 466634
rect 177646 466398 177882 466634
rect 177326 430718 177562 430954
rect 177646 430718 177882 430954
rect 177326 430398 177562 430634
rect 177646 430398 177882 430634
rect 177326 394718 177562 394954
rect 177646 394718 177882 394954
rect 177326 394398 177562 394634
rect 177646 394398 177882 394634
rect 177326 358718 177562 358954
rect 177646 358718 177882 358954
rect 177326 358398 177562 358634
rect 177646 358398 177882 358634
rect 177326 322718 177562 322954
rect 177646 322718 177882 322954
rect 177326 322398 177562 322634
rect 177646 322398 177882 322634
rect 177326 286718 177562 286954
rect 177646 286718 177882 286954
rect 177326 286398 177562 286634
rect 177646 286398 177882 286634
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 186326 705562 186562 705798
rect 186646 705562 186882 705798
rect 186326 705242 186562 705478
rect 186646 705242 186882 705478
rect 186326 691718 186562 691954
rect 186646 691718 186882 691954
rect 186326 691398 186562 691634
rect 186646 691398 186882 691634
rect 186326 655718 186562 655954
rect 186646 655718 186882 655954
rect 186326 655398 186562 655634
rect 186646 655398 186882 655634
rect 186326 619718 186562 619954
rect 186646 619718 186882 619954
rect 186326 619398 186562 619634
rect 186646 619398 186882 619634
rect 186326 583718 186562 583954
rect 186646 583718 186882 583954
rect 186326 583398 186562 583634
rect 186646 583398 186882 583634
rect 186326 547718 186562 547954
rect 186646 547718 186882 547954
rect 186326 547398 186562 547634
rect 186646 547398 186882 547634
rect 186326 511718 186562 511954
rect 186646 511718 186882 511954
rect 186326 511398 186562 511634
rect 186646 511398 186882 511634
rect 186326 475718 186562 475954
rect 186646 475718 186882 475954
rect 186326 475398 186562 475634
rect 186646 475398 186882 475634
rect 186326 439718 186562 439954
rect 186646 439718 186882 439954
rect 186326 439398 186562 439634
rect 186646 439398 186882 439634
rect 186326 403718 186562 403954
rect 186646 403718 186882 403954
rect 186326 403398 186562 403634
rect 186646 403398 186882 403634
rect 186326 367718 186562 367954
rect 186646 367718 186882 367954
rect 186326 367398 186562 367634
rect 186646 367398 186882 367634
rect 186326 331718 186562 331954
rect 186646 331718 186882 331954
rect 186326 331398 186562 331634
rect 186646 331398 186882 331634
rect 186326 295718 186562 295954
rect 186646 295718 186882 295954
rect 186326 295398 186562 295634
rect 186646 295398 186882 295634
rect 190826 706522 191062 706758
rect 191146 706522 191382 706758
rect 190826 706202 191062 706438
rect 191146 706202 191382 706438
rect 190826 696218 191062 696454
rect 191146 696218 191382 696454
rect 190826 695898 191062 696134
rect 191146 695898 191382 696134
rect 190826 660218 191062 660454
rect 191146 660218 191382 660454
rect 190826 659898 191062 660134
rect 191146 659898 191382 660134
rect 190826 624218 191062 624454
rect 191146 624218 191382 624454
rect 190826 623898 191062 624134
rect 191146 623898 191382 624134
rect 190826 588218 191062 588454
rect 191146 588218 191382 588454
rect 190826 587898 191062 588134
rect 191146 587898 191382 588134
rect 190826 552218 191062 552454
rect 191146 552218 191382 552454
rect 190826 551898 191062 552134
rect 191146 551898 191382 552134
rect 190826 516218 191062 516454
rect 191146 516218 191382 516454
rect 190826 515898 191062 516134
rect 191146 515898 191382 516134
rect 190826 480218 191062 480454
rect 191146 480218 191382 480454
rect 190826 479898 191062 480134
rect 191146 479898 191382 480134
rect 190826 444218 191062 444454
rect 191146 444218 191382 444454
rect 190826 443898 191062 444134
rect 191146 443898 191382 444134
rect 190826 408218 191062 408454
rect 191146 408218 191382 408454
rect 190826 407898 191062 408134
rect 191146 407898 191382 408134
rect 190826 372218 191062 372454
rect 191146 372218 191382 372454
rect 190826 371898 191062 372134
rect 191146 371898 191382 372134
rect 190826 336218 191062 336454
rect 191146 336218 191382 336454
rect 190826 335898 191062 336134
rect 191146 335898 191382 336134
rect 190826 300218 191062 300454
rect 191146 300218 191382 300454
rect 190826 299898 191062 300134
rect 191146 299898 191382 300134
rect 124250 255218 124486 255454
rect 124250 254898 124486 255134
rect 154970 255218 155206 255454
rect 154970 254898 155206 255134
rect 139610 223718 139846 223954
rect 139610 223398 139846 223634
rect 170330 223718 170566 223954
rect 170330 223398 170566 223634
rect 124250 219218 124486 219454
rect 124250 218898 124486 219134
rect 154970 219218 155206 219454
rect 154970 218898 155206 219134
rect 185690 255218 185926 255454
rect 185690 254898 185926 255134
rect 185690 219218 185926 219454
rect 185690 218898 185926 219134
rect 123326 196718 123562 196954
rect 123646 196718 123882 196954
rect 123326 196398 123562 196634
rect 123646 196398 123882 196634
rect 123326 160718 123562 160954
rect 123646 160718 123882 160954
rect 123326 160398 123562 160634
rect 123646 160398 123882 160634
rect 124250 111218 124486 111454
rect 124250 110898 124486 111134
rect 118826 48218 119062 48454
rect 119146 48218 119382 48454
rect 118826 47898 119062 48134
rect 119146 47898 119382 48134
rect 114326 7718 114562 7954
rect 114646 7718 114882 7954
rect 114326 7398 114562 7634
rect 114646 7398 114882 7634
rect 114326 -1542 114562 -1306
rect 114646 -1542 114882 -1306
rect 114326 -1862 114562 -1626
rect 114646 -1862 114882 -1626
rect 118826 12218 119062 12454
rect 119146 12218 119382 12454
rect 118826 11898 119062 12134
rect 119146 11898 119382 12134
rect 118826 -2502 119062 -2266
rect 119146 -2502 119382 -2266
rect 118826 -2822 119062 -2586
rect 119146 -2822 119382 -2586
rect 123326 52718 123562 52954
rect 123646 52718 123882 52954
rect 123326 52398 123562 52634
rect 123646 52398 123882 52634
rect 123326 16718 123562 16954
rect 123646 16718 123882 16954
rect 123326 16398 123562 16634
rect 123646 16398 123882 16634
rect 123326 -3462 123562 -3226
rect 123646 -3462 123882 -3226
rect 123326 -3782 123562 -3546
rect 123646 -3782 123882 -3546
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -4422 128062 -4186
rect 128146 -4422 128382 -4186
rect 127826 -4742 128062 -4506
rect 128146 -4742 128382 -4506
rect 132326 61718 132562 61954
rect 132646 61718 132882 61954
rect 132326 61398 132562 61634
rect 132646 61398 132882 61634
rect 136826 66218 137062 66454
rect 137146 66218 137382 66454
rect 136826 65898 137062 66134
rect 137146 65898 137382 66134
rect 132326 25718 132562 25954
rect 132646 25718 132882 25954
rect 132326 25398 132562 25634
rect 132646 25398 132882 25634
rect 132326 -5382 132562 -5146
rect 132646 -5382 132882 -5146
rect 132326 -5702 132562 -5466
rect 132646 -5702 132882 -5466
rect 139610 115718 139846 115954
rect 139610 115398 139846 115634
rect 141326 178718 141562 178954
rect 141646 178718 141882 178954
rect 141326 178398 141562 178634
rect 141646 178398 141882 178634
rect 141326 142718 141562 142954
rect 141646 142718 141882 142954
rect 141326 142398 141562 142634
rect 141646 142398 141882 142634
rect 145826 183218 146062 183454
rect 146146 183218 146382 183454
rect 145826 182898 146062 183134
rect 146146 182898 146382 183134
rect 141326 70718 141562 70954
rect 141646 70718 141882 70954
rect 141326 70398 141562 70634
rect 141646 70398 141882 70634
rect 136826 30218 137062 30454
rect 137146 30218 137382 30454
rect 136826 29898 137062 30134
rect 137146 29898 137382 30134
rect 136826 -6342 137062 -6106
rect 137146 -6342 137382 -6106
rect 136826 -6662 137062 -6426
rect 137146 -6662 137382 -6426
rect 141326 34718 141562 34954
rect 141646 34718 141882 34954
rect 141326 34398 141562 34634
rect 141646 34398 141882 34634
rect 145826 147218 146062 147454
rect 146146 147218 146382 147454
rect 145826 146898 146062 147134
rect 146146 146898 146382 147134
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 150326 187718 150562 187954
rect 150646 187718 150882 187954
rect 150326 187398 150562 187634
rect 150646 187398 150882 187634
rect 150326 151718 150562 151954
rect 150646 151718 150882 151954
rect 150326 151398 150562 151634
rect 150646 151398 150882 151634
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 141326 -7302 141562 -7066
rect 141646 -7302 141882 -7066
rect 141326 -7622 141562 -7386
rect 141646 -7622 141882 -7386
rect 154826 192218 155062 192454
rect 155146 192218 155382 192454
rect 154826 191898 155062 192134
rect 155146 191898 155382 192134
rect 154826 156218 155062 156454
rect 155146 156218 155382 156454
rect 154826 155898 155062 156134
rect 155146 155898 155382 156134
rect 154970 111218 155206 111454
rect 154970 110898 155206 111134
rect 150326 43718 150562 43954
rect 150646 43718 150882 43954
rect 150326 43398 150562 43634
rect 150646 43398 150882 43634
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 159326 196718 159562 196954
rect 159646 196718 159882 196954
rect 159326 196398 159562 196634
rect 159646 196398 159882 196634
rect 159326 160718 159562 160954
rect 159646 160718 159882 160954
rect 159326 160398 159562 160634
rect 159646 160398 159882 160634
rect 159326 52718 159562 52954
rect 159646 52718 159882 52954
rect 159326 52398 159562 52634
rect 159646 52398 159882 52634
rect 154826 48218 155062 48454
rect 155146 48218 155382 48454
rect 154826 47898 155062 48134
rect 155146 47898 155382 48134
rect 150326 7718 150562 7954
rect 150646 7718 150882 7954
rect 150326 7398 150562 7634
rect 150646 7398 150882 7634
rect 150326 -1542 150562 -1306
rect 150646 -1542 150882 -1306
rect 150326 -1862 150562 -1626
rect 150646 -1862 150882 -1626
rect 154826 12218 155062 12454
rect 155146 12218 155382 12454
rect 154826 11898 155062 12134
rect 155146 11898 155382 12134
rect 154826 -2502 155062 -2266
rect 155146 -2502 155382 -2266
rect 154826 -2822 155062 -2586
rect 155146 -2822 155382 -2586
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 159326 16718 159562 16954
rect 159646 16718 159882 16954
rect 159326 16398 159562 16634
rect 159646 16398 159882 16634
rect 159326 -3462 159562 -3226
rect 159646 -3462 159882 -3226
rect 159326 -3782 159562 -3546
rect 159646 -3782 159882 -3546
rect 168326 61718 168562 61954
rect 168646 61718 168882 61954
rect 168326 61398 168562 61634
rect 168646 61398 168882 61634
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -4422 164062 -4186
rect 164146 -4422 164382 -4186
rect 163826 -4742 164062 -4506
rect 164146 -4742 164382 -4506
rect 170330 115718 170566 115954
rect 170330 115398 170566 115634
rect 172826 66218 173062 66454
rect 173146 66218 173382 66454
rect 172826 65898 173062 66134
rect 173146 65898 173382 66134
rect 168326 25718 168562 25954
rect 168646 25718 168882 25954
rect 168326 25398 168562 25634
rect 168646 25398 168882 25634
rect 168326 -5382 168562 -5146
rect 168646 -5382 168882 -5146
rect 168326 -5702 168562 -5466
rect 168646 -5702 168882 -5466
rect 177326 178718 177562 178954
rect 177646 178718 177882 178954
rect 177326 178398 177562 178634
rect 177646 178398 177882 178634
rect 177326 142718 177562 142954
rect 177646 142718 177882 142954
rect 177326 142398 177562 142634
rect 177646 142398 177882 142634
rect 177326 70718 177562 70954
rect 177646 70718 177882 70954
rect 177326 70398 177562 70634
rect 177646 70398 177882 70634
rect 172826 30218 173062 30454
rect 173146 30218 173382 30454
rect 172826 29898 173062 30134
rect 173146 29898 173382 30134
rect 172826 -6342 173062 -6106
rect 173146 -6342 173382 -6106
rect 172826 -6662 173062 -6426
rect 173146 -6662 173382 -6426
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 177326 34718 177562 34954
rect 177646 34718 177882 34954
rect 177326 34398 177562 34634
rect 177646 34398 177882 34634
rect 177326 -7302 177562 -7066
rect 177646 -7302 177882 -7066
rect 177326 -7622 177562 -7386
rect 177646 -7622 177882 -7386
rect 186326 187718 186562 187954
rect 186646 187718 186882 187954
rect 186326 187398 186562 187634
rect 186646 187398 186882 187634
rect 186326 151718 186562 151954
rect 186646 151718 186882 151954
rect 186326 151398 186562 151634
rect 186646 151398 186882 151634
rect 185690 111218 185926 111454
rect 185690 110898 185926 111134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 195326 707482 195562 707718
rect 195646 707482 195882 707718
rect 195326 707162 195562 707398
rect 195646 707162 195882 707398
rect 195326 700718 195562 700954
rect 195646 700718 195882 700954
rect 195326 700398 195562 700634
rect 195646 700398 195882 700634
rect 195326 664718 195562 664954
rect 195646 664718 195882 664954
rect 195326 664398 195562 664634
rect 195646 664398 195882 664634
rect 195326 628718 195562 628954
rect 195646 628718 195882 628954
rect 195326 628398 195562 628634
rect 195646 628398 195882 628634
rect 195326 592718 195562 592954
rect 195646 592718 195882 592954
rect 195326 592398 195562 592634
rect 195646 592398 195882 592634
rect 195326 556718 195562 556954
rect 195646 556718 195882 556954
rect 195326 556398 195562 556634
rect 195646 556398 195882 556634
rect 195326 520718 195562 520954
rect 195646 520718 195882 520954
rect 195326 520398 195562 520634
rect 195646 520398 195882 520634
rect 195326 484718 195562 484954
rect 195646 484718 195882 484954
rect 195326 484398 195562 484634
rect 195646 484398 195882 484634
rect 195326 448718 195562 448954
rect 195646 448718 195882 448954
rect 195326 448398 195562 448634
rect 195646 448398 195882 448634
rect 195326 412718 195562 412954
rect 195646 412718 195882 412954
rect 195326 412398 195562 412634
rect 195646 412398 195882 412634
rect 195326 376718 195562 376954
rect 195646 376718 195882 376954
rect 195326 376398 195562 376634
rect 195646 376398 195882 376634
rect 195326 340718 195562 340954
rect 195646 340718 195882 340954
rect 195326 340398 195562 340634
rect 195646 340398 195882 340634
rect 195326 304718 195562 304954
rect 195646 304718 195882 304954
rect 195326 304398 195562 304634
rect 195646 304398 195882 304634
rect 195326 268718 195562 268954
rect 195646 268718 195882 268954
rect 195326 268398 195562 268634
rect 195646 268398 195882 268634
rect 190826 264218 191062 264454
rect 191146 264218 191382 264454
rect 190826 263898 191062 264134
rect 191146 263898 191382 264134
rect 190826 192218 191062 192454
rect 191146 192218 191382 192454
rect 190826 191898 191062 192134
rect 191146 191898 191382 192134
rect 190826 156218 191062 156454
rect 191146 156218 191382 156454
rect 190826 155898 191062 156134
rect 191146 155898 191382 156134
rect 186326 43718 186562 43954
rect 186646 43718 186882 43954
rect 186326 43398 186562 43634
rect 186646 43398 186882 43634
rect 190826 48218 191062 48454
rect 191146 48218 191382 48454
rect 190826 47898 191062 48134
rect 191146 47898 191382 48134
rect 186326 7718 186562 7954
rect 186646 7718 186882 7954
rect 186326 7398 186562 7634
rect 186646 7398 186882 7634
rect 186326 -1542 186562 -1306
rect 186646 -1542 186882 -1306
rect 186326 -1862 186562 -1626
rect 186646 -1862 186882 -1626
rect 195326 232718 195562 232954
rect 195646 232718 195882 232954
rect 195326 232398 195562 232634
rect 195646 232398 195882 232634
rect 199826 708442 200062 708678
rect 200146 708442 200382 708678
rect 199826 708122 200062 708358
rect 200146 708122 200382 708358
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 199826 525218 200062 525454
rect 200146 525218 200382 525454
rect 199826 524898 200062 525134
rect 200146 524898 200382 525134
rect 199826 489218 200062 489454
rect 200146 489218 200382 489454
rect 199826 488898 200062 489134
rect 200146 488898 200382 489134
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 199826 417218 200062 417454
rect 200146 417218 200382 417454
rect 199826 416898 200062 417134
rect 200146 416898 200382 417134
rect 199826 381218 200062 381454
rect 200146 381218 200382 381454
rect 199826 380898 200062 381134
rect 200146 380898 200382 381134
rect 199826 345218 200062 345454
rect 200146 345218 200382 345454
rect 199826 344898 200062 345134
rect 200146 344898 200382 345134
rect 199826 309218 200062 309454
rect 200146 309218 200382 309454
rect 199826 308898 200062 309134
rect 200146 308898 200382 309134
rect 199826 273218 200062 273454
rect 200146 273218 200382 273454
rect 199826 272898 200062 273134
rect 200146 272898 200382 273134
rect 199826 237218 200062 237454
rect 200146 237218 200382 237454
rect 199826 236898 200062 237134
rect 200146 236898 200382 237134
rect 199826 201218 200062 201454
rect 200146 201218 200382 201454
rect 199826 200898 200062 201134
rect 200146 200898 200382 201134
rect 195326 196718 195562 196954
rect 195646 196718 195882 196954
rect 195326 196398 195562 196634
rect 195646 196398 195882 196634
rect 195326 160718 195562 160954
rect 195646 160718 195882 160954
rect 195326 160398 195562 160634
rect 195646 160398 195882 160634
rect 195326 124718 195562 124954
rect 195646 124718 195882 124954
rect 195326 124398 195562 124634
rect 195646 124398 195882 124634
rect 195326 88718 195562 88954
rect 195646 88718 195882 88954
rect 195326 88398 195562 88634
rect 195646 88398 195882 88634
rect 195326 52718 195562 52954
rect 195646 52718 195882 52954
rect 195326 52398 195562 52634
rect 195646 52398 195882 52634
rect 190826 12218 191062 12454
rect 191146 12218 191382 12454
rect 190826 11898 191062 12134
rect 191146 11898 191382 12134
rect 190826 -2502 191062 -2266
rect 191146 -2502 191382 -2266
rect 190826 -2822 191062 -2586
rect 191146 -2822 191382 -2586
rect 204326 709402 204562 709638
rect 204646 709402 204882 709638
rect 204326 709082 204562 709318
rect 204646 709082 204882 709318
rect 204326 673718 204562 673954
rect 204646 673718 204882 673954
rect 204326 673398 204562 673634
rect 204646 673398 204882 673634
rect 204326 637718 204562 637954
rect 204646 637718 204882 637954
rect 204326 637398 204562 637634
rect 204646 637398 204882 637634
rect 204326 601718 204562 601954
rect 204646 601718 204882 601954
rect 204326 601398 204562 601634
rect 204646 601398 204882 601634
rect 204326 565718 204562 565954
rect 204646 565718 204882 565954
rect 204326 565398 204562 565634
rect 204646 565398 204882 565634
rect 204326 529718 204562 529954
rect 204646 529718 204882 529954
rect 204326 529398 204562 529634
rect 204646 529398 204882 529634
rect 204326 493718 204562 493954
rect 204646 493718 204882 493954
rect 204326 493398 204562 493634
rect 204646 493398 204882 493634
rect 204326 457718 204562 457954
rect 204646 457718 204882 457954
rect 204326 457398 204562 457634
rect 204646 457398 204882 457634
rect 204326 421718 204562 421954
rect 204646 421718 204882 421954
rect 204326 421398 204562 421634
rect 204646 421398 204882 421634
rect 204326 385718 204562 385954
rect 204646 385718 204882 385954
rect 204326 385398 204562 385634
rect 204646 385398 204882 385634
rect 204326 349718 204562 349954
rect 204646 349718 204882 349954
rect 204326 349398 204562 349634
rect 204646 349398 204882 349634
rect 204326 313718 204562 313954
rect 204646 313718 204882 313954
rect 204326 313398 204562 313634
rect 204646 313398 204882 313634
rect 204326 277718 204562 277954
rect 204646 277718 204882 277954
rect 204326 277398 204562 277634
rect 204646 277398 204882 277634
rect 204326 241718 204562 241954
rect 204646 241718 204882 241954
rect 204326 241398 204562 241634
rect 204646 241398 204882 241634
rect 204326 205718 204562 205954
rect 204646 205718 204882 205954
rect 204326 205398 204562 205634
rect 204646 205398 204882 205634
rect 199826 165218 200062 165454
rect 200146 165218 200382 165454
rect 199826 164898 200062 165134
rect 200146 164898 200382 165134
rect 199826 129218 200062 129454
rect 200146 129218 200382 129454
rect 199826 128898 200062 129134
rect 200146 128898 200382 129134
rect 199826 93218 200062 93454
rect 200146 93218 200382 93454
rect 199826 92898 200062 93134
rect 200146 92898 200382 93134
rect 204326 169718 204562 169954
rect 204646 169718 204882 169954
rect 204326 169398 204562 169634
rect 204646 169398 204882 169634
rect 204326 133718 204562 133954
rect 204646 133718 204882 133954
rect 204326 133398 204562 133634
rect 204646 133398 204882 133634
rect 204326 97718 204562 97954
rect 204646 97718 204882 97954
rect 204326 97398 204562 97634
rect 204646 97398 204882 97634
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 195326 16718 195562 16954
rect 195646 16718 195882 16954
rect 195326 16398 195562 16634
rect 195646 16398 195882 16634
rect 195326 -3462 195562 -3226
rect 195646 -3462 195882 -3226
rect 195326 -3782 195562 -3546
rect 195646 -3782 195882 -3546
rect 204326 61718 204562 61954
rect 204646 61718 204882 61954
rect 204326 61398 204562 61634
rect 204646 61398 204882 61634
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -4422 200062 -4186
rect 200146 -4422 200382 -4186
rect 199826 -4742 200062 -4506
rect 200146 -4742 200382 -4506
rect 204326 25718 204562 25954
rect 204646 25718 204882 25954
rect 204326 25398 204562 25634
rect 204646 25398 204882 25634
rect 204326 -5382 204562 -5146
rect 204646 -5382 204882 -5146
rect 204326 -5702 204562 -5466
rect 204646 -5702 204882 -5466
rect 208826 710362 209062 710598
rect 209146 710362 209382 710598
rect 208826 710042 209062 710278
rect 209146 710042 209382 710278
rect 208826 678218 209062 678454
rect 209146 678218 209382 678454
rect 208826 677898 209062 678134
rect 209146 677898 209382 678134
rect 208826 642218 209062 642454
rect 209146 642218 209382 642454
rect 208826 641898 209062 642134
rect 209146 641898 209382 642134
rect 208826 606218 209062 606454
rect 209146 606218 209382 606454
rect 208826 605898 209062 606134
rect 209146 605898 209382 606134
rect 208826 570218 209062 570454
rect 209146 570218 209382 570454
rect 208826 569898 209062 570134
rect 209146 569898 209382 570134
rect 208826 534218 209062 534454
rect 209146 534218 209382 534454
rect 208826 533898 209062 534134
rect 209146 533898 209382 534134
rect 208826 498218 209062 498454
rect 209146 498218 209382 498454
rect 208826 497898 209062 498134
rect 209146 497898 209382 498134
rect 208826 462218 209062 462454
rect 209146 462218 209382 462454
rect 208826 461898 209062 462134
rect 209146 461898 209382 462134
rect 208826 426218 209062 426454
rect 209146 426218 209382 426454
rect 208826 425898 209062 426134
rect 209146 425898 209382 426134
rect 208826 390218 209062 390454
rect 209146 390218 209382 390454
rect 208826 389898 209062 390134
rect 209146 389898 209382 390134
rect 208826 354218 209062 354454
rect 209146 354218 209382 354454
rect 208826 353898 209062 354134
rect 209146 353898 209382 354134
rect 208826 318218 209062 318454
rect 209146 318218 209382 318454
rect 208826 317898 209062 318134
rect 209146 317898 209382 318134
rect 208826 282218 209062 282454
rect 209146 282218 209382 282454
rect 208826 281898 209062 282134
rect 209146 281898 209382 282134
rect 208826 246218 209062 246454
rect 209146 246218 209382 246454
rect 208826 245898 209062 246134
rect 209146 245898 209382 246134
rect 208826 210218 209062 210454
rect 209146 210218 209382 210454
rect 208826 209898 209062 210134
rect 209146 209898 209382 210134
rect 208826 174218 209062 174454
rect 209146 174218 209382 174454
rect 208826 173898 209062 174134
rect 209146 173898 209382 174134
rect 208826 138218 209062 138454
rect 209146 138218 209382 138454
rect 208826 137898 209062 138134
rect 209146 137898 209382 138134
rect 208826 102218 209062 102454
rect 209146 102218 209382 102454
rect 208826 101898 209062 102134
rect 209146 101898 209382 102134
rect 208826 66218 209062 66454
rect 209146 66218 209382 66454
rect 208826 65898 209062 66134
rect 209146 65898 209382 66134
rect 208826 30218 209062 30454
rect 209146 30218 209382 30454
rect 208826 29898 209062 30134
rect 209146 29898 209382 30134
rect 208826 -6342 209062 -6106
rect 209146 -6342 209382 -6106
rect 208826 -6662 209062 -6426
rect 209146 -6662 209382 -6426
rect 213326 711322 213562 711558
rect 213646 711322 213882 711558
rect 213326 711002 213562 711238
rect 213646 711002 213882 711238
rect 213326 682718 213562 682954
rect 213646 682718 213882 682954
rect 213326 682398 213562 682634
rect 213646 682398 213882 682634
rect 213326 646718 213562 646954
rect 213646 646718 213882 646954
rect 213326 646398 213562 646634
rect 213646 646398 213882 646634
rect 213326 610718 213562 610954
rect 213646 610718 213882 610954
rect 213326 610398 213562 610634
rect 213646 610398 213882 610634
rect 213326 574718 213562 574954
rect 213646 574718 213882 574954
rect 213326 574398 213562 574634
rect 213646 574398 213882 574634
rect 213326 538718 213562 538954
rect 213646 538718 213882 538954
rect 213326 538398 213562 538634
rect 213646 538398 213882 538634
rect 213326 502718 213562 502954
rect 213646 502718 213882 502954
rect 213326 502398 213562 502634
rect 213646 502398 213882 502634
rect 213326 466718 213562 466954
rect 213646 466718 213882 466954
rect 213326 466398 213562 466634
rect 213646 466398 213882 466634
rect 213326 430718 213562 430954
rect 213646 430718 213882 430954
rect 213326 430398 213562 430634
rect 213646 430398 213882 430634
rect 213326 394718 213562 394954
rect 213646 394718 213882 394954
rect 213326 394398 213562 394634
rect 213646 394398 213882 394634
rect 213326 358718 213562 358954
rect 213646 358718 213882 358954
rect 213326 358398 213562 358634
rect 213646 358398 213882 358634
rect 213326 322718 213562 322954
rect 213646 322718 213882 322954
rect 213326 322398 213562 322634
rect 213646 322398 213882 322634
rect 213326 286718 213562 286954
rect 213646 286718 213882 286954
rect 213326 286398 213562 286634
rect 213646 286398 213882 286634
rect 213326 250718 213562 250954
rect 213646 250718 213882 250954
rect 213326 250398 213562 250634
rect 213646 250398 213882 250634
rect 213326 214718 213562 214954
rect 213646 214718 213882 214954
rect 213326 214398 213562 214634
rect 213646 214398 213882 214634
rect 213326 178718 213562 178954
rect 213646 178718 213882 178954
rect 213326 178398 213562 178634
rect 213646 178398 213882 178634
rect 213326 142718 213562 142954
rect 213646 142718 213882 142954
rect 213326 142398 213562 142634
rect 213646 142398 213882 142634
rect 213326 106718 213562 106954
rect 213646 106718 213882 106954
rect 213326 106398 213562 106634
rect 213646 106398 213882 106634
rect 213326 70718 213562 70954
rect 213646 70718 213882 70954
rect 213326 70398 213562 70634
rect 213646 70398 213882 70634
rect 213326 34718 213562 34954
rect 213646 34718 213882 34954
rect 213326 34398 213562 34634
rect 213646 34398 213882 34634
rect 213326 -7302 213562 -7066
rect 213646 -7302 213882 -7066
rect 213326 -7622 213562 -7386
rect 213646 -7622 213882 -7386
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 217826 507218 218062 507454
rect 218146 507218 218382 507454
rect 217826 506898 218062 507134
rect 218146 506898 218382 507134
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 217826 435218 218062 435454
rect 218146 435218 218382 435454
rect 217826 434898 218062 435134
rect 218146 434898 218382 435134
rect 217826 399218 218062 399454
rect 218146 399218 218382 399454
rect 217826 398898 218062 399134
rect 218146 398898 218382 399134
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 217826 327218 218062 327454
rect 218146 327218 218382 327454
rect 217826 326898 218062 327134
rect 218146 326898 218382 327134
rect 217826 291218 218062 291454
rect 218146 291218 218382 291454
rect 217826 290898 218062 291134
rect 218146 290898 218382 291134
rect 217826 255218 218062 255454
rect 218146 255218 218382 255454
rect 217826 254898 218062 255134
rect 218146 254898 218382 255134
rect 217826 219218 218062 219454
rect 218146 219218 218382 219454
rect 217826 218898 218062 219134
rect 218146 218898 218382 219134
rect 217826 183218 218062 183454
rect 218146 183218 218382 183454
rect 217826 182898 218062 183134
rect 218146 182898 218382 183134
rect 217826 147218 218062 147454
rect 218146 147218 218382 147454
rect 217826 146898 218062 147134
rect 218146 146898 218382 147134
rect 217826 111218 218062 111454
rect 218146 111218 218382 111454
rect 217826 110898 218062 111134
rect 218146 110898 218382 111134
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 222326 705562 222562 705798
rect 222646 705562 222882 705798
rect 222326 705242 222562 705478
rect 222646 705242 222882 705478
rect 222326 691718 222562 691954
rect 222646 691718 222882 691954
rect 222326 691398 222562 691634
rect 222646 691398 222882 691634
rect 222326 655718 222562 655954
rect 222646 655718 222882 655954
rect 222326 655398 222562 655634
rect 222646 655398 222882 655634
rect 222326 619718 222562 619954
rect 222646 619718 222882 619954
rect 222326 619398 222562 619634
rect 222646 619398 222882 619634
rect 222326 583718 222562 583954
rect 222646 583718 222882 583954
rect 222326 583398 222562 583634
rect 222646 583398 222882 583634
rect 222326 547718 222562 547954
rect 222646 547718 222882 547954
rect 222326 547398 222562 547634
rect 222646 547398 222882 547634
rect 222326 511718 222562 511954
rect 222646 511718 222882 511954
rect 222326 511398 222562 511634
rect 222646 511398 222882 511634
rect 222326 475718 222562 475954
rect 222646 475718 222882 475954
rect 222326 475398 222562 475634
rect 222646 475398 222882 475634
rect 222326 439718 222562 439954
rect 222646 439718 222882 439954
rect 222326 439398 222562 439634
rect 222646 439398 222882 439634
rect 222326 403718 222562 403954
rect 222646 403718 222882 403954
rect 222326 403398 222562 403634
rect 222646 403398 222882 403634
rect 222326 367718 222562 367954
rect 222646 367718 222882 367954
rect 222326 367398 222562 367634
rect 222646 367398 222882 367634
rect 222326 331718 222562 331954
rect 222646 331718 222882 331954
rect 222326 331398 222562 331634
rect 222646 331398 222882 331634
rect 222326 295718 222562 295954
rect 222646 295718 222882 295954
rect 222326 295398 222562 295634
rect 222646 295398 222882 295634
rect 222326 259718 222562 259954
rect 222646 259718 222882 259954
rect 222326 259398 222562 259634
rect 222646 259398 222882 259634
rect 222326 223718 222562 223954
rect 222646 223718 222882 223954
rect 222326 223398 222562 223634
rect 222646 223398 222882 223634
rect 222326 187718 222562 187954
rect 222646 187718 222882 187954
rect 222326 187398 222562 187634
rect 222646 187398 222882 187634
rect 222326 151718 222562 151954
rect 222646 151718 222882 151954
rect 222326 151398 222562 151634
rect 222646 151398 222882 151634
rect 222326 115718 222562 115954
rect 222646 115718 222882 115954
rect 222326 115398 222562 115634
rect 222646 115398 222882 115634
rect 222326 79718 222562 79954
rect 222646 79718 222882 79954
rect 222326 79398 222562 79634
rect 222646 79398 222882 79634
rect 222326 43718 222562 43954
rect 222646 43718 222882 43954
rect 222326 43398 222562 43634
rect 222646 43398 222882 43634
rect 222326 7718 222562 7954
rect 222646 7718 222882 7954
rect 222326 7398 222562 7634
rect 222646 7398 222882 7634
rect 222326 -1542 222562 -1306
rect 222646 -1542 222882 -1306
rect 222326 -1862 222562 -1626
rect 222646 -1862 222882 -1626
rect 226826 706522 227062 706758
rect 227146 706522 227382 706758
rect 226826 706202 227062 706438
rect 227146 706202 227382 706438
rect 226826 696218 227062 696454
rect 227146 696218 227382 696454
rect 226826 695898 227062 696134
rect 227146 695898 227382 696134
rect 226826 660218 227062 660454
rect 227146 660218 227382 660454
rect 226826 659898 227062 660134
rect 227146 659898 227382 660134
rect 226826 624218 227062 624454
rect 227146 624218 227382 624454
rect 226826 623898 227062 624134
rect 227146 623898 227382 624134
rect 226826 588218 227062 588454
rect 227146 588218 227382 588454
rect 226826 587898 227062 588134
rect 227146 587898 227382 588134
rect 226826 552218 227062 552454
rect 227146 552218 227382 552454
rect 226826 551898 227062 552134
rect 227146 551898 227382 552134
rect 226826 516218 227062 516454
rect 227146 516218 227382 516454
rect 226826 515898 227062 516134
rect 227146 515898 227382 516134
rect 226826 480218 227062 480454
rect 227146 480218 227382 480454
rect 226826 479898 227062 480134
rect 227146 479898 227382 480134
rect 226826 444218 227062 444454
rect 227146 444218 227382 444454
rect 226826 443898 227062 444134
rect 227146 443898 227382 444134
rect 226826 408218 227062 408454
rect 227146 408218 227382 408454
rect 226826 407898 227062 408134
rect 227146 407898 227382 408134
rect 226826 372218 227062 372454
rect 227146 372218 227382 372454
rect 226826 371898 227062 372134
rect 227146 371898 227382 372134
rect 226826 336218 227062 336454
rect 227146 336218 227382 336454
rect 226826 335898 227062 336134
rect 227146 335898 227382 336134
rect 226826 300218 227062 300454
rect 227146 300218 227382 300454
rect 226826 299898 227062 300134
rect 227146 299898 227382 300134
rect 226826 264218 227062 264454
rect 227146 264218 227382 264454
rect 226826 263898 227062 264134
rect 227146 263898 227382 264134
rect 226826 228218 227062 228454
rect 227146 228218 227382 228454
rect 226826 227898 227062 228134
rect 227146 227898 227382 228134
rect 226826 192218 227062 192454
rect 227146 192218 227382 192454
rect 226826 191898 227062 192134
rect 227146 191898 227382 192134
rect 226826 156218 227062 156454
rect 227146 156218 227382 156454
rect 226826 155898 227062 156134
rect 227146 155898 227382 156134
rect 226826 120218 227062 120454
rect 227146 120218 227382 120454
rect 226826 119898 227062 120134
rect 227146 119898 227382 120134
rect 226826 84218 227062 84454
rect 227146 84218 227382 84454
rect 226826 83898 227062 84134
rect 227146 83898 227382 84134
rect 226826 48218 227062 48454
rect 227146 48218 227382 48454
rect 226826 47898 227062 48134
rect 227146 47898 227382 48134
rect 226826 12218 227062 12454
rect 227146 12218 227382 12454
rect 226826 11898 227062 12134
rect 227146 11898 227382 12134
rect 226826 -2502 227062 -2266
rect 227146 -2502 227382 -2266
rect 226826 -2822 227062 -2586
rect 227146 -2822 227382 -2586
rect 231326 707482 231562 707718
rect 231646 707482 231882 707718
rect 231326 707162 231562 707398
rect 231646 707162 231882 707398
rect 231326 700718 231562 700954
rect 231646 700718 231882 700954
rect 231326 700398 231562 700634
rect 231646 700398 231882 700634
rect 231326 664718 231562 664954
rect 231646 664718 231882 664954
rect 231326 664398 231562 664634
rect 231646 664398 231882 664634
rect 231326 628718 231562 628954
rect 231646 628718 231882 628954
rect 231326 628398 231562 628634
rect 231646 628398 231882 628634
rect 231326 592718 231562 592954
rect 231646 592718 231882 592954
rect 231326 592398 231562 592634
rect 231646 592398 231882 592634
rect 231326 556718 231562 556954
rect 231646 556718 231882 556954
rect 231326 556398 231562 556634
rect 231646 556398 231882 556634
rect 231326 520718 231562 520954
rect 231646 520718 231882 520954
rect 231326 520398 231562 520634
rect 231646 520398 231882 520634
rect 231326 484718 231562 484954
rect 231646 484718 231882 484954
rect 231326 484398 231562 484634
rect 231646 484398 231882 484634
rect 231326 448718 231562 448954
rect 231646 448718 231882 448954
rect 231326 448398 231562 448634
rect 231646 448398 231882 448634
rect 231326 412718 231562 412954
rect 231646 412718 231882 412954
rect 231326 412398 231562 412634
rect 231646 412398 231882 412634
rect 231326 376718 231562 376954
rect 231646 376718 231882 376954
rect 231326 376398 231562 376634
rect 231646 376398 231882 376634
rect 231326 340718 231562 340954
rect 231646 340718 231882 340954
rect 231326 340398 231562 340634
rect 231646 340398 231882 340634
rect 231326 304718 231562 304954
rect 231646 304718 231882 304954
rect 231326 304398 231562 304634
rect 231646 304398 231882 304634
rect 231326 268718 231562 268954
rect 231646 268718 231882 268954
rect 231326 268398 231562 268634
rect 231646 268398 231882 268634
rect 231326 232718 231562 232954
rect 231646 232718 231882 232954
rect 231326 232398 231562 232634
rect 231646 232398 231882 232634
rect 231326 196718 231562 196954
rect 231646 196718 231882 196954
rect 231326 196398 231562 196634
rect 231646 196398 231882 196634
rect 231326 160718 231562 160954
rect 231646 160718 231882 160954
rect 231326 160398 231562 160634
rect 231646 160398 231882 160634
rect 231326 124718 231562 124954
rect 231646 124718 231882 124954
rect 231326 124398 231562 124634
rect 231646 124398 231882 124634
rect 231326 88718 231562 88954
rect 231646 88718 231882 88954
rect 231326 88398 231562 88634
rect 231646 88398 231882 88634
rect 231326 52718 231562 52954
rect 231646 52718 231882 52954
rect 231326 52398 231562 52634
rect 231646 52398 231882 52634
rect 231326 16718 231562 16954
rect 231646 16718 231882 16954
rect 231326 16398 231562 16634
rect 231646 16398 231882 16634
rect 231326 -3462 231562 -3226
rect 231646 -3462 231882 -3226
rect 231326 -3782 231562 -3546
rect 231646 -3782 231882 -3546
rect 235826 708442 236062 708678
rect 236146 708442 236382 708678
rect 235826 708122 236062 708358
rect 236146 708122 236382 708358
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 235826 561218 236062 561454
rect 236146 561218 236382 561454
rect 235826 560898 236062 561134
rect 236146 560898 236382 561134
rect 235826 525218 236062 525454
rect 236146 525218 236382 525454
rect 235826 524898 236062 525134
rect 236146 524898 236382 525134
rect 235826 489218 236062 489454
rect 236146 489218 236382 489454
rect 235826 488898 236062 489134
rect 236146 488898 236382 489134
rect 235826 453218 236062 453454
rect 236146 453218 236382 453454
rect 235826 452898 236062 453134
rect 236146 452898 236382 453134
rect 235826 417218 236062 417454
rect 236146 417218 236382 417454
rect 235826 416898 236062 417134
rect 236146 416898 236382 417134
rect 235826 381218 236062 381454
rect 236146 381218 236382 381454
rect 235826 380898 236062 381134
rect 236146 380898 236382 381134
rect 235826 345218 236062 345454
rect 236146 345218 236382 345454
rect 235826 344898 236062 345134
rect 236146 344898 236382 345134
rect 235826 309218 236062 309454
rect 236146 309218 236382 309454
rect 235826 308898 236062 309134
rect 236146 308898 236382 309134
rect 235826 273218 236062 273454
rect 236146 273218 236382 273454
rect 235826 272898 236062 273134
rect 236146 272898 236382 273134
rect 235826 237218 236062 237454
rect 236146 237218 236382 237454
rect 235826 236898 236062 237134
rect 236146 236898 236382 237134
rect 235826 201218 236062 201454
rect 236146 201218 236382 201454
rect 235826 200898 236062 201134
rect 236146 200898 236382 201134
rect 235826 165218 236062 165454
rect 236146 165218 236382 165454
rect 235826 164898 236062 165134
rect 236146 164898 236382 165134
rect 235826 129218 236062 129454
rect 236146 129218 236382 129454
rect 235826 128898 236062 129134
rect 236146 128898 236382 129134
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -4422 236062 -4186
rect 236146 -4422 236382 -4186
rect 235826 -4742 236062 -4506
rect 236146 -4742 236382 -4506
rect 240326 709402 240562 709638
rect 240646 709402 240882 709638
rect 240326 709082 240562 709318
rect 240646 709082 240882 709318
rect 240326 673718 240562 673954
rect 240646 673718 240882 673954
rect 240326 673398 240562 673634
rect 240646 673398 240882 673634
rect 240326 637718 240562 637954
rect 240646 637718 240882 637954
rect 240326 637398 240562 637634
rect 240646 637398 240882 637634
rect 240326 601718 240562 601954
rect 240646 601718 240882 601954
rect 240326 601398 240562 601634
rect 240646 601398 240882 601634
rect 240326 565718 240562 565954
rect 240646 565718 240882 565954
rect 240326 565398 240562 565634
rect 240646 565398 240882 565634
rect 240326 529718 240562 529954
rect 240646 529718 240882 529954
rect 240326 529398 240562 529634
rect 240646 529398 240882 529634
rect 240326 493718 240562 493954
rect 240646 493718 240882 493954
rect 240326 493398 240562 493634
rect 240646 493398 240882 493634
rect 240326 457718 240562 457954
rect 240646 457718 240882 457954
rect 240326 457398 240562 457634
rect 240646 457398 240882 457634
rect 240326 421718 240562 421954
rect 240646 421718 240882 421954
rect 240326 421398 240562 421634
rect 240646 421398 240882 421634
rect 240326 385718 240562 385954
rect 240646 385718 240882 385954
rect 240326 385398 240562 385634
rect 240646 385398 240882 385634
rect 240326 349718 240562 349954
rect 240646 349718 240882 349954
rect 240326 349398 240562 349634
rect 240646 349398 240882 349634
rect 240326 313718 240562 313954
rect 240646 313718 240882 313954
rect 240326 313398 240562 313634
rect 240646 313398 240882 313634
rect 240326 277718 240562 277954
rect 240646 277718 240882 277954
rect 240326 277398 240562 277634
rect 240646 277398 240882 277634
rect 240326 241718 240562 241954
rect 240646 241718 240882 241954
rect 240326 241398 240562 241634
rect 240646 241398 240882 241634
rect 240326 205718 240562 205954
rect 240646 205718 240882 205954
rect 240326 205398 240562 205634
rect 240646 205398 240882 205634
rect 240326 169718 240562 169954
rect 240646 169718 240882 169954
rect 240326 169398 240562 169634
rect 240646 169398 240882 169634
rect 240326 133718 240562 133954
rect 240646 133718 240882 133954
rect 240326 133398 240562 133634
rect 240646 133398 240882 133634
rect 240326 97718 240562 97954
rect 240646 97718 240882 97954
rect 240326 97398 240562 97634
rect 240646 97398 240882 97634
rect 240326 61718 240562 61954
rect 240646 61718 240882 61954
rect 240326 61398 240562 61634
rect 240646 61398 240882 61634
rect 240326 25718 240562 25954
rect 240646 25718 240882 25954
rect 240326 25398 240562 25634
rect 240646 25398 240882 25634
rect 240326 -5382 240562 -5146
rect 240646 -5382 240882 -5146
rect 240326 -5702 240562 -5466
rect 240646 -5702 240882 -5466
rect 244826 710362 245062 710598
rect 245146 710362 245382 710598
rect 244826 710042 245062 710278
rect 245146 710042 245382 710278
rect 244826 678218 245062 678454
rect 245146 678218 245382 678454
rect 244826 677898 245062 678134
rect 245146 677898 245382 678134
rect 244826 642218 245062 642454
rect 245146 642218 245382 642454
rect 244826 641898 245062 642134
rect 245146 641898 245382 642134
rect 244826 606218 245062 606454
rect 245146 606218 245382 606454
rect 244826 605898 245062 606134
rect 245146 605898 245382 606134
rect 244826 570218 245062 570454
rect 245146 570218 245382 570454
rect 244826 569898 245062 570134
rect 245146 569898 245382 570134
rect 244826 534218 245062 534454
rect 245146 534218 245382 534454
rect 244826 533898 245062 534134
rect 245146 533898 245382 534134
rect 244826 498218 245062 498454
rect 245146 498218 245382 498454
rect 244826 497898 245062 498134
rect 245146 497898 245382 498134
rect 244826 462218 245062 462454
rect 245146 462218 245382 462454
rect 244826 461898 245062 462134
rect 245146 461898 245382 462134
rect 244826 426218 245062 426454
rect 245146 426218 245382 426454
rect 244826 425898 245062 426134
rect 245146 425898 245382 426134
rect 244826 390218 245062 390454
rect 245146 390218 245382 390454
rect 244826 389898 245062 390134
rect 245146 389898 245382 390134
rect 244826 354218 245062 354454
rect 245146 354218 245382 354454
rect 244826 353898 245062 354134
rect 245146 353898 245382 354134
rect 244826 318218 245062 318454
rect 245146 318218 245382 318454
rect 244826 317898 245062 318134
rect 245146 317898 245382 318134
rect 244826 282218 245062 282454
rect 245146 282218 245382 282454
rect 244826 281898 245062 282134
rect 245146 281898 245382 282134
rect 244826 246218 245062 246454
rect 245146 246218 245382 246454
rect 244826 245898 245062 246134
rect 245146 245898 245382 246134
rect 244826 210218 245062 210454
rect 245146 210218 245382 210454
rect 244826 209898 245062 210134
rect 245146 209898 245382 210134
rect 244826 174218 245062 174454
rect 245146 174218 245382 174454
rect 244826 173898 245062 174134
rect 245146 173898 245382 174134
rect 244826 138218 245062 138454
rect 245146 138218 245382 138454
rect 244826 137898 245062 138134
rect 245146 137898 245382 138134
rect 244826 102218 245062 102454
rect 245146 102218 245382 102454
rect 244826 101898 245062 102134
rect 245146 101898 245382 102134
rect 244826 66218 245062 66454
rect 245146 66218 245382 66454
rect 244826 65898 245062 66134
rect 245146 65898 245382 66134
rect 244826 30218 245062 30454
rect 245146 30218 245382 30454
rect 244826 29898 245062 30134
rect 245146 29898 245382 30134
rect 244826 -6342 245062 -6106
rect 245146 -6342 245382 -6106
rect 244826 -6662 245062 -6426
rect 245146 -6662 245382 -6426
rect 249326 711322 249562 711558
rect 249646 711322 249882 711558
rect 249326 711002 249562 711238
rect 249646 711002 249882 711238
rect 249326 682718 249562 682954
rect 249646 682718 249882 682954
rect 249326 682398 249562 682634
rect 249646 682398 249882 682634
rect 249326 646718 249562 646954
rect 249646 646718 249882 646954
rect 249326 646398 249562 646634
rect 249646 646398 249882 646634
rect 249326 610718 249562 610954
rect 249646 610718 249882 610954
rect 249326 610398 249562 610634
rect 249646 610398 249882 610634
rect 249326 574718 249562 574954
rect 249646 574718 249882 574954
rect 249326 574398 249562 574634
rect 249646 574398 249882 574634
rect 249326 538718 249562 538954
rect 249646 538718 249882 538954
rect 249326 538398 249562 538634
rect 249646 538398 249882 538634
rect 249326 502718 249562 502954
rect 249646 502718 249882 502954
rect 249326 502398 249562 502634
rect 249646 502398 249882 502634
rect 249326 466718 249562 466954
rect 249646 466718 249882 466954
rect 249326 466398 249562 466634
rect 249646 466398 249882 466634
rect 249326 430718 249562 430954
rect 249646 430718 249882 430954
rect 249326 430398 249562 430634
rect 249646 430398 249882 430634
rect 249326 394718 249562 394954
rect 249646 394718 249882 394954
rect 249326 394398 249562 394634
rect 249646 394398 249882 394634
rect 249326 358718 249562 358954
rect 249646 358718 249882 358954
rect 249326 358398 249562 358634
rect 249646 358398 249882 358634
rect 249326 322718 249562 322954
rect 249646 322718 249882 322954
rect 249326 322398 249562 322634
rect 249646 322398 249882 322634
rect 249326 286718 249562 286954
rect 249646 286718 249882 286954
rect 249326 286398 249562 286634
rect 249646 286398 249882 286634
rect 249326 250718 249562 250954
rect 249646 250718 249882 250954
rect 249326 250398 249562 250634
rect 249646 250398 249882 250634
rect 249326 214718 249562 214954
rect 249646 214718 249882 214954
rect 249326 214398 249562 214634
rect 249646 214398 249882 214634
rect 249326 178718 249562 178954
rect 249646 178718 249882 178954
rect 249326 178398 249562 178634
rect 249646 178398 249882 178634
rect 249326 142718 249562 142954
rect 249646 142718 249882 142954
rect 249326 142398 249562 142634
rect 249646 142398 249882 142634
rect 249326 106718 249562 106954
rect 249646 106718 249882 106954
rect 249326 106398 249562 106634
rect 249646 106398 249882 106634
rect 249326 70718 249562 70954
rect 249646 70718 249882 70954
rect 249326 70398 249562 70634
rect 249646 70398 249882 70634
rect 249326 34718 249562 34954
rect 249646 34718 249882 34954
rect 249326 34398 249562 34634
rect 249646 34398 249882 34634
rect 249326 -7302 249562 -7066
rect 249646 -7302 249882 -7066
rect 249326 -7622 249562 -7386
rect 249646 -7622 249882 -7386
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 253826 507218 254062 507454
rect 254146 507218 254382 507454
rect 253826 506898 254062 507134
rect 254146 506898 254382 507134
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 253826 435218 254062 435454
rect 254146 435218 254382 435454
rect 253826 434898 254062 435134
rect 254146 434898 254382 435134
rect 253826 399218 254062 399454
rect 254146 399218 254382 399454
rect 253826 398898 254062 399134
rect 254146 398898 254382 399134
rect 253826 363218 254062 363454
rect 254146 363218 254382 363454
rect 253826 362898 254062 363134
rect 254146 362898 254382 363134
rect 253826 327218 254062 327454
rect 254146 327218 254382 327454
rect 253826 326898 254062 327134
rect 254146 326898 254382 327134
rect 253826 291218 254062 291454
rect 254146 291218 254382 291454
rect 253826 290898 254062 291134
rect 254146 290898 254382 291134
rect 253826 255218 254062 255454
rect 254146 255218 254382 255454
rect 253826 254898 254062 255134
rect 254146 254898 254382 255134
rect 253826 219218 254062 219454
rect 254146 219218 254382 219454
rect 253826 218898 254062 219134
rect 254146 218898 254382 219134
rect 253826 183218 254062 183454
rect 254146 183218 254382 183454
rect 253826 182898 254062 183134
rect 254146 182898 254382 183134
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 258326 705562 258562 705798
rect 258646 705562 258882 705798
rect 258326 705242 258562 705478
rect 258646 705242 258882 705478
rect 258326 691718 258562 691954
rect 258646 691718 258882 691954
rect 258326 691398 258562 691634
rect 258646 691398 258882 691634
rect 258326 655718 258562 655954
rect 258646 655718 258882 655954
rect 258326 655398 258562 655634
rect 258646 655398 258882 655634
rect 258326 619718 258562 619954
rect 258646 619718 258882 619954
rect 258326 619398 258562 619634
rect 258646 619398 258882 619634
rect 258326 583718 258562 583954
rect 258646 583718 258882 583954
rect 258326 583398 258562 583634
rect 258646 583398 258882 583634
rect 258326 547718 258562 547954
rect 258646 547718 258882 547954
rect 258326 547398 258562 547634
rect 258646 547398 258882 547634
rect 258326 511718 258562 511954
rect 258646 511718 258882 511954
rect 258326 511398 258562 511634
rect 258646 511398 258882 511634
rect 258326 475718 258562 475954
rect 258646 475718 258882 475954
rect 258326 475398 258562 475634
rect 258646 475398 258882 475634
rect 258326 439718 258562 439954
rect 258646 439718 258882 439954
rect 258326 439398 258562 439634
rect 258646 439398 258882 439634
rect 258326 403718 258562 403954
rect 258646 403718 258882 403954
rect 258326 403398 258562 403634
rect 258646 403398 258882 403634
rect 258326 367718 258562 367954
rect 258646 367718 258882 367954
rect 258326 367398 258562 367634
rect 258646 367398 258882 367634
rect 258326 331718 258562 331954
rect 258646 331718 258882 331954
rect 258326 331398 258562 331634
rect 258646 331398 258882 331634
rect 258326 295718 258562 295954
rect 258646 295718 258882 295954
rect 258326 295398 258562 295634
rect 258646 295398 258882 295634
rect 258326 259718 258562 259954
rect 258646 259718 258882 259954
rect 258326 259398 258562 259634
rect 258646 259398 258882 259634
rect 258326 223718 258562 223954
rect 258646 223718 258882 223954
rect 258326 223398 258562 223634
rect 258646 223398 258882 223634
rect 258326 187718 258562 187954
rect 258646 187718 258882 187954
rect 258326 187398 258562 187634
rect 258646 187398 258882 187634
rect 258326 151718 258562 151954
rect 258646 151718 258882 151954
rect 258326 151398 258562 151634
rect 258646 151398 258882 151634
rect 258326 115718 258562 115954
rect 258646 115718 258882 115954
rect 258326 115398 258562 115634
rect 258646 115398 258882 115634
rect 258326 79718 258562 79954
rect 258646 79718 258882 79954
rect 258326 79398 258562 79634
rect 258646 79398 258882 79634
rect 258326 43718 258562 43954
rect 258646 43718 258882 43954
rect 258326 43398 258562 43634
rect 258646 43398 258882 43634
rect 258326 7718 258562 7954
rect 258646 7718 258882 7954
rect 258326 7398 258562 7634
rect 258646 7398 258882 7634
rect 258326 -1542 258562 -1306
rect 258646 -1542 258882 -1306
rect 258326 -1862 258562 -1626
rect 258646 -1862 258882 -1626
rect 262826 706522 263062 706758
rect 263146 706522 263382 706758
rect 262826 706202 263062 706438
rect 263146 706202 263382 706438
rect 262826 696218 263062 696454
rect 263146 696218 263382 696454
rect 262826 695898 263062 696134
rect 263146 695898 263382 696134
rect 262826 660218 263062 660454
rect 263146 660218 263382 660454
rect 262826 659898 263062 660134
rect 263146 659898 263382 660134
rect 262826 624218 263062 624454
rect 263146 624218 263382 624454
rect 262826 623898 263062 624134
rect 263146 623898 263382 624134
rect 262826 588218 263062 588454
rect 263146 588218 263382 588454
rect 262826 587898 263062 588134
rect 263146 587898 263382 588134
rect 262826 552218 263062 552454
rect 263146 552218 263382 552454
rect 262826 551898 263062 552134
rect 263146 551898 263382 552134
rect 262826 516218 263062 516454
rect 263146 516218 263382 516454
rect 262826 515898 263062 516134
rect 263146 515898 263382 516134
rect 262826 480218 263062 480454
rect 263146 480218 263382 480454
rect 262826 479898 263062 480134
rect 263146 479898 263382 480134
rect 262826 444218 263062 444454
rect 263146 444218 263382 444454
rect 262826 443898 263062 444134
rect 263146 443898 263382 444134
rect 262826 408218 263062 408454
rect 263146 408218 263382 408454
rect 262826 407898 263062 408134
rect 263146 407898 263382 408134
rect 262826 372218 263062 372454
rect 263146 372218 263382 372454
rect 262826 371898 263062 372134
rect 263146 371898 263382 372134
rect 262826 336218 263062 336454
rect 263146 336218 263382 336454
rect 262826 335898 263062 336134
rect 263146 335898 263382 336134
rect 262826 300218 263062 300454
rect 263146 300218 263382 300454
rect 262826 299898 263062 300134
rect 263146 299898 263382 300134
rect 262826 264218 263062 264454
rect 263146 264218 263382 264454
rect 262826 263898 263062 264134
rect 263146 263898 263382 264134
rect 262826 228218 263062 228454
rect 263146 228218 263382 228454
rect 262826 227898 263062 228134
rect 263146 227898 263382 228134
rect 262826 192218 263062 192454
rect 263146 192218 263382 192454
rect 262826 191898 263062 192134
rect 263146 191898 263382 192134
rect 262826 156218 263062 156454
rect 263146 156218 263382 156454
rect 262826 155898 263062 156134
rect 263146 155898 263382 156134
rect 262826 120218 263062 120454
rect 263146 120218 263382 120454
rect 262826 119898 263062 120134
rect 263146 119898 263382 120134
rect 262826 84218 263062 84454
rect 263146 84218 263382 84454
rect 262826 83898 263062 84134
rect 263146 83898 263382 84134
rect 262826 48218 263062 48454
rect 263146 48218 263382 48454
rect 262826 47898 263062 48134
rect 263146 47898 263382 48134
rect 262826 12218 263062 12454
rect 263146 12218 263382 12454
rect 262826 11898 263062 12134
rect 263146 11898 263382 12134
rect 262826 -2502 263062 -2266
rect 263146 -2502 263382 -2266
rect 262826 -2822 263062 -2586
rect 263146 -2822 263382 -2586
rect 267326 707482 267562 707718
rect 267646 707482 267882 707718
rect 267326 707162 267562 707398
rect 267646 707162 267882 707398
rect 267326 700718 267562 700954
rect 267646 700718 267882 700954
rect 267326 700398 267562 700634
rect 267646 700398 267882 700634
rect 267326 664718 267562 664954
rect 267646 664718 267882 664954
rect 267326 664398 267562 664634
rect 267646 664398 267882 664634
rect 267326 628718 267562 628954
rect 267646 628718 267882 628954
rect 267326 628398 267562 628634
rect 267646 628398 267882 628634
rect 267326 592718 267562 592954
rect 267646 592718 267882 592954
rect 267326 592398 267562 592634
rect 267646 592398 267882 592634
rect 267326 556718 267562 556954
rect 267646 556718 267882 556954
rect 267326 556398 267562 556634
rect 267646 556398 267882 556634
rect 267326 520718 267562 520954
rect 267646 520718 267882 520954
rect 267326 520398 267562 520634
rect 267646 520398 267882 520634
rect 267326 484718 267562 484954
rect 267646 484718 267882 484954
rect 267326 484398 267562 484634
rect 267646 484398 267882 484634
rect 267326 448718 267562 448954
rect 267646 448718 267882 448954
rect 267326 448398 267562 448634
rect 267646 448398 267882 448634
rect 267326 412718 267562 412954
rect 267646 412718 267882 412954
rect 267326 412398 267562 412634
rect 267646 412398 267882 412634
rect 267326 376718 267562 376954
rect 267646 376718 267882 376954
rect 267326 376398 267562 376634
rect 267646 376398 267882 376634
rect 267326 340718 267562 340954
rect 267646 340718 267882 340954
rect 267326 340398 267562 340634
rect 267646 340398 267882 340634
rect 267326 304718 267562 304954
rect 267646 304718 267882 304954
rect 267326 304398 267562 304634
rect 267646 304398 267882 304634
rect 267326 268718 267562 268954
rect 267646 268718 267882 268954
rect 267326 268398 267562 268634
rect 267646 268398 267882 268634
rect 267326 232718 267562 232954
rect 267646 232718 267882 232954
rect 267326 232398 267562 232634
rect 267646 232398 267882 232634
rect 267326 196718 267562 196954
rect 267646 196718 267882 196954
rect 267326 196398 267562 196634
rect 267646 196398 267882 196634
rect 267326 160718 267562 160954
rect 267646 160718 267882 160954
rect 267326 160398 267562 160634
rect 267646 160398 267882 160634
rect 267326 124718 267562 124954
rect 267646 124718 267882 124954
rect 267326 124398 267562 124634
rect 267646 124398 267882 124634
rect 267326 88718 267562 88954
rect 267646 88718 267882 88954
rect 267326 88398 267562 88634
rect 267646 88398 267882 88634
rect 267326 52718 267562 52954
rect 267646 52718 267882 52954
rect 267326 52398 267562 52634
rect 267646 52398 267882 52634
rect 267326 16718 267562 16954
rect 267646 16718 267882 16954
rect 267326 16398 267562 16634
rect 267646 16398 267882 16634
rect 267326 -3462 267562 -3226
rect 267646 -3462 267882 -3226
rect 267326 -3782 267562 -3546
rect 267646 -3782 267882 -3546
rect 271826 708442 272062 708678
rect 272146 708442 272382 708678
rect 271826 708122 272062 708358
rect 272146 708122 272382 708358
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 271826 525218 272062 525454
rect 272146 525218 272382 525454
rect 271826 524898 272062 525134
rect 272146 524898 272382 525134
rect 271826 489218 272062 489454
rect 272146 489218 272382 489454
rect 271826 488898 272062 489134
rect 272146 488898 272382 489134
rect 271826 453218 272062 453454
rect 272146 453218 272382 453454
rect 271826 452898 272062 453134
rect 272146 452898 272382 453134
rect 271826 417218 272062 417454
rect 272146 417218 272382 417454
rect 271826 416898 272062 417134
rect 272146 416898 272382 417134
rect 271826 381218 272062 381454
rect 272146 381218 272382 381454
rect 271826 380898 272062 381134
rect 272146 380898 272382 381134
rect 271826 345218 272062 345454
rect 272146 345218 272382 345454
rect 271826 344898 272062 345134
rect 272146 344898 272382 345134
rect 271826 309218 272062 309454
rect 272146 309218 272382 309454
rect 271826 308898 272062 309134
rect 272146 308898 272382 309134
rect 271826 273218 272062 273454
rect 272146 273218 272382 273454
rect 271826 272898 272062 273134
rect 272146 272898 272382 273134
rect 271826 237218 272062 237454
rect 272146 237218 272382 237454
rect 271826 236898 272062 237134
rect 272146 236898 272382 237134
rect 271826 201218 272062 201454
rect 272146 201218 272382 201454
rect 271826 200898 272062 201134
rect 272146 200898 272382 201134
rect 271826 165218 272062 165454
rect 272146 165218 272382 165454
rect 271826 164898 272062 165134
rect 272146 164898 272382 165134
rect 271826 129218 272062 129454
rect 272146 129218 272382 129454
rect 271826 128898 272062 129134
rect 272146 128898 272382 129134
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -4422 272062 -4186
rect 272146 -4422 272382 -4186
rect 271826 -4742 272062 -4506
rect 272146 -4742 272382 -4506
rect 276326 709402 276562 709638
rect 276646 709402 276882 709638
rect 276326 709082 276562 709318
rect 276646 709082 276882 709318
rect 276326 673718 276562 673954
rect 276646 673718 276882 673954
rect 276326 673398 276562 673634
rect 276646 673398 276882 673634
rect 276326 637718 276562 637954
rect 276646 637718 276882 637954
rect 276326 637398 276562 637634
rect 276646 637398 276882 637634
rect 276326 601718 276562 601954
rect 276646 601718 276882 601954
rect 276326 601398 276562 601634
rect 276646 601398 276882 601634
rect 276326 565718 276562 565954
rect 276646 565718 276882 565954
rect 276326 565398 276562 565634
rect 276646 565398 276882 565634
rect 276326 529718 276562 529954
rect 276646 529718 276882 529954
rect 276326 529398 276562 529634
rect 276646 529398 276882 529634
rect 276326 493718 276562 493954
rect 276646 493718 276882 493954
rect 276326 493398 276562 493634
rect 276646 493398 276882 493634
rect 276326 457718 276562 457954
rect 276646 457718 276882 457954
rect 276326 457398 276562 457634
rect 276646 457398 276882 457634
rect 276326 421718 276562 421954
rect 276646 421718 276882 421954
rect 276326 421398 276562 421634
rect 276646 421398 276882 421634
rect 276326 385718 276562 385954
rect 276646 385718 276882 385954
rect 276326 385398 276562 385634
rect 276646 385398 276882 385634
rect 276326 349718 276562 349954
rect 276646 349718 276882 349954
rect 276326 349398 276562 349634
rect 276646 349398 276882 349634
rect 276326 313718 276562 313954
rect 276646 313718 276882 313954
rect 276326 313398 276562 313634
rect 276646 313398 276882 313634
rect 276326 277718 276562 277954
rect 276646 277718 276882 277954
rect 276326 277398 276562 277634
rect 276646 277398 276882 277634
rect 276326 241718 276562 241954
rect 276646 241718 276882 241954
rect 276326 241398 276562 241634
rect 276646 241398 276882 241634
rect 276326 205718 276562 205954
rect 276646 205718 276882 205954
rect 276326 205398 276562 205634
rect 276646 205398 276882 205634
rect 276326 169718 276562 169954
rect 276646 169718 276882 169954
rect 276326 169398 276562 169634
rect 276646 169398 276882 169634
rect 276326 133718 276562 133954
rect 276646 133718 276882 133954
rect 276326 133398 276562 133634
rect 276646 133398 276882 133634
rect 276326 97718 276562 97954
rect 276646 97718 276882 97954
rect 276326 97398 276562 97634
rect 276646 97398 276882 97634
rect 276326 61718 276562 61954
rect 276646 61718 276882 61954
rect 276326 61398 276562 61634
rect 276646 61398 276882 61634
rect 276326 25718 276562 25954
rect 276646 25718 276882 25954
rect 276326 25398 276562 25634
rect 276646 25398 276882 25634
rect 276326 -5382 276562 -5146
rect 276646 -5382 276882 -5146
rect 276326 -5702 276562 -5466
rect 276646 -5702 276882 -5466
rect 280826 710362 281062 710598
rect 281146 710362 281382 710598
rect 280826 710042 281062 710278
rect 281146 710042 281382 710278
rect 280826 678218 281062 678454
rect 281146 678218 281382 678454
rect 280826 677898 281062 678134
rect 281146 677898 281382 678134
rect 280826 642218 281062 642454
rect 281146 642218 281382 642454
rect 280826 641898 281062 642134
rect 281146 641898 281382 642134
rect 280826 606218 281062 606454
rect 281146 606218 281382 606454
rect 280826 605898 281062 606134
rect 281146 605898 281382 606134
rect 280826 570218 281062 570454
rect 281146 570218 281382 570454
rect 280826 569898 281062 570134
rect 281146 569898 281382 570134
rect 280826 534218 281062 534454
rect 281146 534218 281382 534454
rect 280826 533898 281062 534134
rect 281146 533898 281382 534134
rect 280826 498218 281062 498454
rect 281146 498218 281382 498454
rect 280826 497898 281062 498134
rect 281146 497898 281382 498134
rect 280826 462218 281062 462454
rect 281146 462218 281382 462454
rect 280826 461898 281062 462134
rect 281146 461898 281382 462134
rect 280826 426218 281062 426454
rect 281146 426218 281382 426454
rect 280826 425898 281062 426134
rect 281146 425898 281382 426134
rect 280826 390218 281062 390454
rect 281146 390218 281382 390454
rect 280826 389898 281062 390134
rect 281146 389898 281382 390134
rect 280826 354218 281062 354454
rect 281146 354218 281382 354454
rect 280826 353898 281062 354134
rect 281146 353898 281382 354134
rect 280826 318218 281062 318454
rect 281146 318218 281382 318454
rect 280826 317898 281062 318134
rect 281146 317898 281382 318134
rect 280826 282218 281062 282454
rect 281146 282218 281382 282454
rect 280826 281898 281062 282134
rect 281146 281898 281382 282134
rect 280826 246218 281062 246454
rect 281146 246218 281382 246454
rect 280826 245898 281062 246134
rect 281146 245898 281382 246134
rect 280826 210218 281062 210454
rect 281146 210218 281382 210454
rect 280826 209898 281062 210134
rect 281146 209898 281382 210134
rect 280826 174218 281062 174454
rect 281146 174218 281382 174454
rect 280826 173898 281062 174134
rect 281146 173898 281382 174134
rect 280826 138218 281062 138454
rect 281146 138218 281382 138454
rect 280826 137898 281062 138134
rect 281146 137898 281382 138134
rect 280826 102218 281062 102454
rect 281146 102218 281382 102454
rect 280826 101898 281062 102134
rect 281146 101898 281382 102134
rect 280826 66218 281062 66454
rect 281146 66218 281382 66454
rect 280826 65898 281062 66134
rect 281146 65898 281382 66134
rect 280826 30218 281062 30454
rect 281146 30218 281382 30454
rect 280826 29898 281062 30134
rect 281146 29898 281382 30134
rect 280826 -6342 281062 -6106
rect 281146 -6342 281382 -6106
rect 280826 -6662 281062 -6426
rect 281146 -6662 281382 -6426
rect 285326 711322 285562 711558
rect 285646 711322 285882 711558
rect 285326 711002 285562 711238
rect 285646 711002 285882 711238
rect 285326 682718 285562 682954
rect 285646 682718 285882 682954
rect 285326 682398 285562 682634
rect 285646 682398 285882 682634
rect 285326 646718 285562 646954
rect 285646 646718 285882 646954
rect 285326 646398 285562 646634
rect 285646 646398 285882 646634
rect 285326 610718 285562 610954
rect 285646 610718 285882 610954
rect 285326 610398 285562 610634
rect 285646 610398 285882 610634
rect 285326 574718 285562 574954
rect 285646 574718 285882 574954
rect 285326 574398 285562 574634
rect 285646 574398 285882 574634
rect 285326 538718 285562 538954
rect 285646 538718 285882 538954
rect 285326 538398 285562 538634
rect 285646 538398 285882 538634
rect 285326 502718 285562 502954
rect 285646 502718 285882 502954
rect 285326 502398 285562 502634
rect 285646 502398 285882 502634
rect 285326 466718 285562 466954
rect 285646 466718 285882 466954
rect 285326 466398 285562 466634
rect 285646 466398 285882 466634
rect 285326 430718 285562 430954
rect 285646 430718 285882 430954
rect 285326 430398 285562 430634
rect 285646 430398 285882 430634
rect 285326 394718 285562 394954
rect 285646 394718 285882 394954
rect 285326 394398 285562 394634
rect 285646 394398 285882 394634
rect 285326 358718 285562 358954
rect 285646 358718 285882 358954
rect 285326 358398 285562 358634
rect 285646 358398 285882 358634
rect 285326 322718 285562 322954
rect 285646 322718 285882 322954
rect 285326 322398 285562 322634
rect 285646 322398 285882 322634
rect 285326 286718 285562 286954
rect 285646 286718 285882 286954
rect 285326 286398 285562 286634
rect 285646 286398 285882 286634
rect 285326 250718 285562 250954
rect 285646 250718 285882 250954
rect 285326 250398 285562 250634
rect 285646 250398 285882 250634
rect 285326 214718 285562 214954
rect 285646 214718 285882 214954
rect 285326 214398 285562 214634
rect 285646 214398 285882 214634
rect 285326 178718 285562 178954
rect 285646 178718 285882 178954
rect 285326 178398 285562 178634
rect 285646 178398 285882 178634
rect 285326 142718 285562 142954
rect 285646 142718 285882 142954
rect 285326 142398 285562 142634
rect 285646 142398 285882 142634
rect 285326 106718 285562 106954
rect 285646 106718 285882 106954
rect 285326 106398 285562 106634
rect 285646 106398 285882 106634
rect 285326 70718 285562 70954
rect 285646 70718 285882 70954
rect 285326 70398 285562 70634
rect 285646 70398 285882 70634
rect 285326 34718 285562 34954
rect 285646 34718 285882 34954
rect 285326 34398 285562 34634
rect 285646 34398 285882 34634
rect 285326 -7302 285562 -7066
rect 285646 -7302 285882 -7066
rect 285326 -7622 285562 -7386
rect 285646 -7622 285882 -7386
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 289826 435218 290062 435454
rect 290146 435218 290382 435454
rect 289826 434898 290062 435134
rect 290146 434898 290382 435134
rect 289826 399218 290062 399454
rect 290146 399218 290382 399454
rect 289826 398898 290062 399134
rect 290146 398898 290382 399134
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 289826 327218 290062 327454
rect 290146 327218 290382 327454
rect 289826 326898 290062 327134
rect 290146 326898 290382 327134
rect 289826 291218 290062 291454
rect 290146 291218 290382 291454
rect 289826 290898 290062 291134
rect 290146 290898 290382 291134
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 289826 219218 290062 219454
rect 290146 219218 290382 219454
rect 289826 218898 290062 219134
rect 290146 218898 290382 219134
rect 289826 183218 290062 183454
rect 290146 183218 290382 183454
rect 289826 182898 290062 183134
rect 290146 182898 290382 183134
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 294326 705562 294562 705798
rect 294646 705562 294882 705798
rect 294326 705242 294562 705478
rect 294646 705242 294882 705478
rect 294326 691718 294562 691954
rect 294646 691718 294882 691954
rect 294326 691398 294562 691634
rect 294646 691398 294882 691634
rect 294326 655718 294562 655954
rect 294646 655718 294882 655954
rect 294326 655398 294562 655634
rect 294646 655398 294882 655634
rect 294326 619718 294562 619954
rect 294646 619718 294882 619954
rect 294326 619398 294562 619634
rect 294646 619398 294882 619634
rect 294326 583718 294562 583954
rect 294646 583718 294882 583954
rect 294326 583398 294562 583634
rect 294646 583398 294882 583634
rect 294326 547718 294562 547954
rect 294646 547718 294882 547954
rect 294326 547398 294562 547634
rect 294646 547398 294882 547634
rect 294326 511718 294562 511954
rect 294646 511718 294882 511954
rect 294326 511398 294562 511634
rect 294646 511398 294882 511634
rect 294326 475718 294562 475954
rect 294646 475718 294882 475954
rect 294326 475398 294562 475634
rect 294646 475398 294882 475634
rect 294326 439718 294562 439954
rect 294646 439718 294882 439954
rect 294326 439398 294562 439634
rect 294646 439398 294882 439634
rect 294326 403718 294562 403954
rect 294646 403718 294882 403954
rect 294326 403398 294562 403634
rect 294646 403398 294882 403634
rect 294326 367718 294562 367954
rect 294646 367718 294882 367954
rect 294326 367398 294562 367634
rect 294646 367398 294882 367634
rect 294326 331718 294562 331954
rect 294646 331718 294882 331954
rect 294326 331398 294562 331634
rect 294646 331398 294882 331634
rect 294326 295718 294562 295954
rect 294646 295718 294882 295954
rect 294326 295398 294562 295634
rect 294646 295398 294882 295634
rect 294326 259718 294562 259954
rect 294646 259718 294882 259954
rect 294326 259398 294562 259634
rect 294646 259398 294882 259634
rect 294326 223718 294562 223954
rect 294646 223718 294882 223954
rect 294326 223398 294562 223634
rect 294646 223398 294882 223634
rect 294326 187718 294562 187954
rect 294646 187718 294882 187954
rect 294326 187398 294562 187634
rect 294646 187398 294882 187634
rect 294326 151718 294562 151954
rect 294646 151718 294882 151954
rect 294326 151398 294562 151634
rect 294646 151398 294882 151634
rect 294326 115718 294562 115954
rect 294646 115718 294882 115954
rect 294326 115398 294562 115634
rect 294646 115398 294882 115634
rect 294326 79718 294562 79954
rect 294646 79718 294882 79954
rect 294326 79398 294562 79634
rect 294646 79398 294882 79634
rect 294326 43718 294562 43954
rect 294646 43718 294882 43954
rect 294326 43398 294562 43634
rect 294646 43398 294882 43634
rect 294326 7718 294562 7954
rect 294646 7718 294882 7954
rect 294326 7398 294562 7634
rect 294646 7398 294882 7634
rect 294326 -1542 294562 -1306
rect 294646 -1542 294882 -1306
rect 294326 -1862 294562 -1626
rect 294646 -1862 294882 -1626
rect 298826 706522 299062 706758
rect 299146 706522 299382 706758
rect 298826 706202 299062 706438
rect 299146 706202 299382 706438
rect 298826 696218 299062 696454
rect 299146 696218 299382 696454
rect 298826 695898 299062 696134
rect 299146 695898 299382 696134
rect 298826 660218 299062 660454
rect 299146 660218 299382 660454
rect 298826 659898 299062 660134
rect 299146 659898 299382 660134
rect 298826 624218 299062 624454
rect 299146 624218 299382 624454
rect 298826 623898 299062 624134
rect 299146 623898 299382 624134
rect 298826 588218 299062 588454
rect 299146 588218 299382 588454
rect 298826 587898 299062 588134
rect 299146 587898 299382 588134
rect 298826 552218 299062 552454
rect 299146 552218 299382 552454
rect 298826 551898 299062 552134
rect 299146 551898 299382 552134
rect 298826 516218 299062 516454
rect 299146 516218 299382 516454
rect 298826 515898 299062 516134
rect 299146 515898 299382 516134
rect 298826 480218 299062 480454
rect 299146 480218 299382 480454
rect 298826 479898 299062 480134
rect 299146 479898 299382 480134
rect 298826 444218 299062 444454
rect 299146 444218 299382 444454
rect 298826 443898 299062 444134
rect 299146 443898 299382 444134
rect 298826 408218 299062 408454
rect 299146 408218 299382 408454
rect 298826 407898 299062 408134
rect 299146 407898 299382 408134
rect 298826 372218 299062 372454
rect 299146 372218 299382 372454
rect 298826 371898 299062 372134
rect 299146 371898 299382 372134
rect 298826 336218 299062 336454
rect 299146 336218 299382 336454
rect 298826 335898 299062 336134
rect 299146 335898 299382 336134
rect 298826 300218 299062 300454
rect 299146 300218 299382 300454
rect 298826 299898 299062 300134
rect 299146 299898 299382 300134
rect 298826 264218 299062 264454
rect 299146 264218 299382 264454
rect 298826 263898 299062 264134
rect 299146 263898 299382 264134
rect 298826 228218 299062 228454
rect 299146 228218 299382 228454
rect 298826 227898 299062 228134
rect 299146 227898 299382 228134
rect 298826 192218 299062 192454
rect 299146 192218 299382 192454
rect 298826 191898 299062 192134
rect 299146 191898 299382 192134
rect 298826 156218 299062 156454
rect 299146 156218 299382 156454
rect 298826 155898 299062 156134
rect 299146 155898 299382 156134
rect 298826 120218 299062 120454
rect 299146 120218 299382 120454
rect 298826 119898 299062 120134
rect 299146 119898 299382 120134
rect 298826 84218 299062 84454
rect 299146 84218 299382 84454
rect 298826 83898 299062 84134
rect 299146 83898 299382 84134
rect 298826 48218 299062 48454
rect 299146 48218 299382 48454
rect 298826 47898 299062 48134
rect 299146 47898 299382 48134
rect 298826 12218 299062 12454
rect 299146 12218 299382 12454
rect 298826 11898 299062 12134
rect 299146 11898 299382 12134
rect 298826 -2502 299062 -2266
rect 299146 -2502 299382 -2266
rect 298826 -2822 299062 -2586
rect 299146 -2822 299382 -2586
rect 303326 707482 303562 707718
rect 303646 707482 303882 707718
rect 303326 707162 303562 707398
rect 303646 707162 303882 707398
rect 303326 700718 303562 700954
rect 303646 700718 303882 700954
rect 303326 700398 303562 700634
rect 303646 700398 303882 700634
rect 303326 664718 303562 664954
rect 303646 664718 303882 664954
rect 303326 664398 303562 664634
rect 303646 664398 303882 664634
rect 303326 628718 303562 628954
rect 303646 628718 303882 628954
rect 303326 628398 303562 628634
rect 303646 628398 303882 628634
rect 303326 592718 303562 592954
rect 303646 592718 303882 592954
rect 303326 592398 303562 592634
rect 303646 592398 303882 592634
rect 303326 556718 303562 556954
rect 303646 556718 303882 556954
rect 303326 556398 303562 556634
rect 303646 556398 303882 556634
rect 303326 520718 303562 520954
rect 303646 520718 303882 520954
rect 303326 520398 303562 520634
rect 303646 520398 303882 520634
rect 303326 484718 303562 484954
rect 303646 484718 303882 484954
rect 303326 484398 303562 484634
rect 303646 484398 303882 484634
rect 303326 448718 303562 448954
rect 303646 448718 303882 448954
rect 303326 448398 303562 448634
rect 303646 448398 303882 448634
rect 303326 412718 303562 412954
rect 303646 412718 303882 412954
rect 303326 412398 303562 412634
rect 303646 412398 303882 412634
rect 303326 376718 303562 376954
rect 303646 376718 303882 376954
rect 303326 376398 303562 376634
rect 303646 376398 303882 376634
rect 303326 340718 303562 340954
rect 303646 340718 303882 340954
rect 303326 340398 303562 340634
rect 303646 340398 303882 340634
rect 303326 304718 303562 304954
rect 303646 304718 303882 304954
rect 303326 304398 303562 304634
rect 303646 304398 303882 304634
rect 303326 268718 303562 268954
rect 303646 268718 303882 268954
rect 303326 268398 303562 268634
rect 303646 268398 303882 268634
rect 303326 232718 303562 232954
rect 303646 232718 303882 232954
rect 303326 232398 303562 232634
rect 303646 232398 303882 232634
rect 303326 196718 303562 196954
rect 303646 196718 303882 196954
rect 303326 196398 303562 196634
rect 303646 196398 303882 196634
rect 303326 160718 303562 160954
rect 303646 160718 303882 160954
rect 303326 160398 303562 160634
rect 303646 160398 303882 160634
rect 303326 124718 303562 124954
rect 303646 124718 303882 124954
rect 303326 124398 303562 124634
rect 303646 124398 303882 124634
rect 303326 88718 303562 88954
rect 303646 88718 303882 88954
rect 303326 88398 303562 88634
rect 303646 88398 303882 88634
rect 303326 52718 303562 52954
rect 303646 52718 303882 52954
rect 303326 52398 303562 52634
rect 303646 52398 303882 52634
rect 303326 16718 303562 16954
rect 303646 16718 303882 16954
rect 303326 16398 303562 16634
rect 303646 16398 303882 16634
rect 303326 -3462 303562 -3226
rect 303646 -3462 303882 -3226
rect 303326 -3782 303562 -3546
rect 303646 -3782 303882 -3546
rect 307826 708442 308062 708678
rect 308146 708442 308382 708678
rect 307826 708122 308062 708358
rect 308146 708122 308382 708358
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 307826 525218 308062 525454
rect 308146 525218 308382 525454
rect 307826 524898 308062 525134
rect 308146 524898 308382 525134
rect 307826 489218 308062 489454
rect 308146 489218 308382 489454
rect 307826 488898 308062 489134
rect 308146 488898 308382 489134
rect 307826 453218 308062 453454
rect 308146 453218 308382 453454
rect 307826 452898 308062 453134
rect 308146 452898 308382 453134
rect 307826 417218 308062 417454
rect 308146 417218 308382 417454
rect 307826 416898 308062 417134
rect 308146 416898 308382 417134
rect 307826 381218 308062 381454
rect 308146 381218 308382 381454
rect 307826 380898 308062 381134
rect 308146 380898 308382 381134
rect 307826 345218 308062 345454
rect 308146 345218 308382 345454
rect 307826 344898 308062 345134
rect 308146 344898 308382 345134
rect 307826 309218 308062 309454
rect 308146 309218 308382 309454
rect 307826 308898 308062 309134
rect 308146 308898 308382 309134
rect 307826 273218 308062 273454
rect 308146 273218 308382 273454
rect 307826 272898 308062 273134
rect 308146 272898 308382 273134
rect 307826 237218 308062 237454
rect 308146 237218 308382 237454
rect 307826 236898 308062 237134
rect 308146 236898 308382 237134
rect 307826 201218 308062 201454
rect 308146 201218 308382 201454
rect 307826 200898 308062 201134
rect 308146 200898 308382 201134
rect 307826 165218 308062 165454
rect 308146 165218 308382 165454
rect 307826 164898 308062 165134
rect 308146 164898 308382 165134
rect 307826 129218 308062 129454
rect 308146 129218 308382 129454
rect 307826 128898 308062 129134
rect 308146 128898 308382 129134
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -4422 308062 -4186
rect 308146 -4422 308382 -4186
rect 307826 -4742 308062 -4506
rect 308146 -4742 308382 -4506
rect 312326 709402 312562 709638
rect 312646 709402 312882 709638
rect 312326 709082 312562 709318
rect 312646 709082 312882 709318
rect 312326 673718 312562 673954
rect 312646 673718 312882 673954
rect 312326 673398 312562 673634
rect 312646 673398 312882 673634
rect 312326 637718 312562 637954
rect 312646 637718 312882 637954
rect 312326 637398 312562 637634
rect 312646 637398 312882 637634
rect 312326 601718 312562 601954
rect 312646 601718 312882 601954
rect 312326 601398 312562 601634
rect 312646 601398 312882 601634
rect 312326 565718 312562 565954
rect 312646 565718 312882 565954
rect 312326 565398 312562 565634
rect 312646 565398 312882 565634
rect 312326 529718 312562 529954
rect 312646 529718 312882 529954
rect 312326 529398 312562 529634
rect 312646 529398 312882 529634
rect 312326 493718 312562 493954
rect 312646 493718 312882 493954
rect 312326 493398 312562 493634
rect 312646 493398 312882 493634
rect 312326 457718 312562 457954
rect 312646 457718 312882 457954
rect 312326 457398 312562 457634
rect 312646 457398 312882 457634
rect 312326 421718 312562 421954
rect 312646 421718 312882 421954
rect 312326 421398 312562 421634
rect 312646 421398 312882 421634
rect 312326 385718 312562 385954
rect 312646 385718 312882 385954
rect 312326 385398 312562 385634
rect 312646 385398 312882 385634
rect 312326 349718 312562 349954
rect 312646 349718 312882 349954
rect 312326 349398 312562 349634
rect 312646 349398 312882 349634
rect 312326 313718 312562 313954
rect 312646 313718 312882 313954
rect 312326 313398 312562 313634
rect 312646 313398 312882 313634
rect 312326 277718 312562 277954
rect 312646 277718 312882 277954
rect 312326 277398 312562 277634
rect 312646 277398 312882 277634
rect 312326 241718 312562 241954
rect 312646 241718 312882 241954
rect 312326 241398 312562 241634
rect 312646 241398 312882 241634
rect 312326 205718 312562 205954
rect 312646 205718 312882 205954
rect 312326 205398 312562 205634
rect 312646 205398 312882 205634
rect 312326 169718 312562 169954
rect 312646 169718 312882 169954
rect 312326 169398 312562 169634
rect 312646 169398 312882 169634
rect 312326 133718 312562 133954
rect 312646 133718 312882 133954
rect 312326 133398 312562 133634
rect 312646 133398 312882 133634
rect 312326 97718 312562 97954
rect 312646 97718 312882 97954
rect 312326 97398 312562 97634
rect 312646 97398 312882 97634
rect 312326 61718 312562 61954
rect 312646 61718 312882 61954
rect 312326 61398 312562 61634
rect 312646 61398 312882 61634
rect 312326 25718 312562 25954
rect 312646 25718 312882 25954
rect 312326 25398 312562 25634
rect 312646 25398 312882 25634
rect 312326 -5382 312562 -5146
rect 312646 -5382 312882 -5146
rect 312326 -5702 312562 -5466
rect 312646 -5702 312882 -5466
rect 316826 710362 317062 710598
rect 317146 710362 317382 710598
rect 316826 710042 317062 710278
rect 317146 710042 317382 710278
rect 316826 678218 317062 678454
rect 317146 678218 317382 678454
rect 316826 677898 317062 678134
rect 317146 677898 317382 678134
rect 316826 642218 317062 642454
rect 317146 642218 317382 642454
rect 316826 641898 317062 642134
rect 317146 641898 317382 642134
rect 316826 606218 317062 606454
rect 317146 606218 317382 606454
rect 316826 605898 317062 606134
rect 317146 605898 317382 606134
rect 316826 570218 317062 570454
rect 317146 570218 317382 570454
rect 316826 569898 317062 570134
rect 317146 569898 317382 570134
rect 316826 534218 317062 534454
rect 317146 534218 317382 534454
rect 316826 533898 317062 534134
rect 317146 533898 317382 534134
rect 316826 498218 317062 498454
rect 317146 498218 317382 498454
rect 316826 497898 317062 498134
rect 317146 497898 317382 498134
rect 316826 462218 317062 462454
rect 317146 462218 317382 462454
rect 316826 461898 317062 462134
rect 317146 461898 317382 462134
rect 316826 426218 317062 426454
rect 317146 426218 317382 426454
rect 316826 425898 317062 426134
rect 317146 425898 317382 426134
rect 316826 390218 317062 390454
rect 317146 390218 317382 390454
rect 316826 389898 317062 390134
rect 317146 389898 317382 390134
rect 316826 354218 317062 354454
rect 317146 354218 317382 354454
rect 316826 353898 317062 354134
rect 317146 353898 317382 354134
rect 316826 318218 317062 318454
rect 317146 318218 317382 318454
rect 316826 317898 317062 318134
rect 317146 317898 317382 318134
rect 316826 282218 317062 282454
rect 317146 282218 317382 282454
rect 316826 281898 317062 282134
rect 317146 281898 317382 282134
rect 316826 246218 317062 246454
rect 317146 246218 317382 246454
rect 316826 245898 317062 246134
rect 317146 245898 317382 246134
rect 316826 210218 317062 210454
rect 317146 210218 317382 210454
rect 316826 209898 317062 210134
rect 317146 209898 317382 210134
rect 316826 174218 317062 174454
rect 317146 174218 317382 174454
rect 316826 173898 317062 174134
rect 317146 173898 317382 174134
rect 316826 138218 317062 138454
rect 317146 138218 317382 138454
rect 316826 137898 317062 138134
rect 317146 137898 317382 138134
rect 316826 102218 317062 102454
rect 317146 102218 317382 102454
rect 316826 101898 317062 102134
rect 317146 101898 317382 102134
rect 316826 66218 317062 66454
rect 317146 66218 317382 66454
rect 316826 65898 317062 66134
rect 317146 65898 317382 66134
rect 316826 30218 317062 30454
rect 317146 30218 317382 30454
rect 316826 29898 317062 30134
rect 317146 29898 317382 30134
rect 316826 -6342 317062 -6106
rect 317146 -6342 317382 -6106
rect 316826 -6662 317062 -6426
rect 317146 -6662 317382 -6426
rect 321326 711322 321562 711558
rect 321646 711322 321882 711558
rect 321326 711002 321562 711238
rect 321646 711002 321882 711238
rect 321326 682718 321562 682954
rect 321646 682718 321882 682954
rect 321326 682398 321562 682634
rect 321646 682398 321882 682634
rect 321326 646718 321562 646954
rect 321646 646718 321882 646954
rect 321326 646398 321562 646634
rect 321646 646398 321882 646634
rect 321326 610718 321562 610954
rect 321646 610718 321882 610954
rect 321326 610398 321562 610634
rect 321646 610398 321882 610634
rect 321326 574718 321562 574954
rect 321646 574718 321882 574954
rect 321326 574398 321562 574634
rect 321646 574398 321882 574634
rect 321326 538718 321562 538954
rect 321646 538718 321882 538954
rect 321326 538398 321562 538634
rect 321646 538398 321882 538634
rect 321326 502718 321562 502954
rect 321646 502718 321882 502954
rect 321326 502398 321562 502634
rect 321646 502398 321882 502634
rect 321326 466718 321562 466954
rect 321646 466718 321882 466954
rect 321326 466398 321562 466634
rect 321646 466398 321882 466634
rect 321326 430718 321562 430954
rect 321646 430718 321882 430954
rect 321326 430398 321562 430634
rect 321646 430398 321882 430634
rect 321326 394718 321562 394954
rect 321646 394718 321882 394954
rect 321326 394398 321562 394634
rect 321646 394398 321882 394634
rect 321326 358718 321562 358954
rect 321646 358718 321882 358954
rect 321326 358398 321562 358634
rect 321646 358398 321882 358634
rect 321326 322718 321562 322954
rect 321646 322718 321882 322954
rect 321326 322398 321562 322634
rect 321646 322398 321882 322634
rect 321326 286718 321562 286954
rect 321646 286718 321882 286954
rect 321326 286398 321562 286634
rect 321646 286398 321882 286634
rect 321326 250718 321562 250954
rect 321646 250718 321882 250954
rect 321326 250398 321562 250634
rect 321646 250398 321882 250634
rect 321326 214718 321562 214954
rect 321646 214718 321882 214954
rect 321326 214398 321562 214634
rect 321646 214398 321882 214634
rect 321326 178718 321562 178954
rect 321646 178718 321882 178954
rect 321326 178398 321562 178634
rect 321646 178398 321882 178634
rect 321326 142718 321562 142954
rect 321646 142718 321882 142954
rect 321326 142398 321562 142634
rect 321646 142398 321882 142634
rect 321326 106718 321562 106954
rect 321646 106718 321882 106954
rect 321326 106398 321562 106634
rect 321646 106398 321882 106634
rect 321326 70718 321562 70954
rect 321646 70718 321882 70954
rect 321326 70398 321562 70634
rect 321646 70398 321882 70634
rect 321326 34718 321562 34954
rect 321646 34718 321882 34954
rect 321326 34398 321562 34634
rect 321646 34398 321882 34634
rect 321326 -7302 321562 -7066
rect 321646 -7302 321882 -7066
rect 321326 -7622 321562 -7386
rect 321646 -7622 321882 -7386
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 325826 435218 326062 435454
rect 326146 435218 326382 435454
rect 325826 434898 326062 435134
rect 326146 434898 326382 435134
rect 325826 399218 326062 399454
rect 326146 399218 326382 399454
rect 325826 398898 326062 399134
rect 326146 398898 326382 399134
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 325826 327218 326062 327454
rect 326146 327218 326382 327454
rect 325826 326898 326062 327134
rect 326146 326898 326382 327134
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 325826 219218 326062 219454
rect 326146 219218 326382 219454
rect 325826 218898 326062 219134
rect 326146 218898 326382 219134
rect 325826 183218 326062 183454
rect 326146 183218 326382 183454
rect 325826 182898 326062 183134
rect 326146 182898 326382 183134
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 330326 705562 330562 705798
rect 330646 705562 330882 705798
rect 330326 705242 330562 705478
rect 330646 705242 330882 705478
rect 330326 691718 330562 691954
rect 330646 691718 330882 691954
rect 330326 691398 330562 691634
rect 330646 691398 330882 691634
rect 330326 655718 330562 655954
rect 330646 655718 330882 655954
rect 330326 655398 330562 655634
rect 330646 655398 330882 655634
rect 330326 619718 330562 619954
rect 330646 619718 330882 619954
rect 330326 619398 330562 619634
rect 330646 619398 330882 619634
rect 330326 583718 330562 583954
rect 330646 583718 330882 583954
rect 330326 583398 330562 583634
rect 330646 583398 330882 583634
rect 330326 547718 330562 547954
rect 330646 547718 330882 547954
rect 330326 547398 330562 547634
rect 330646 547398 330882 547634
rect 330326 511718 330562 511954
rect 330646 511718 330882 511954
rect 330326 511398 330562 511634
rect 330646 511398 330882 511634
rect 330326 475718 330562 475954
rect 330646 475718 330882 475954
rect 330326 475398 330562 475634
rect 330646 475398 330882 475634
rect 330326 439718 330562 439954
rect 330646 439718 330882 439954
rect 330326 439398 330562 439634
rect 330646 439398 330882 439634
rect 330326 403718 330562 403954
rect 330646 403718 330882 403954
rect 330326 403398 330562 403634
rect 330646 403398 330882 403634
rect 330326 367718 330562 367954
rect 330646 367718 330882 367954
rect 330326 367398 330562 367634
rect 330646 367398 330882 367634
rect 330326 331718 330562 331954
rect 330646 331718 330882 331954
rect 330326 331398 330562 331634
rect 330646 331398 330882 331634
rect 330326 295718 330562 295954
rect 330646 295718 330882 295954
rect 330326 295398 330562 295634
rect 330646 295398 330882 295634
rect 330326 259718 330562 259954
rect 330646 259718 330882 259954
rect 330326 259398 330562 259634
rect 330646 259398 330882 259634
rect 330326 223718 330562 223954
rect 330646 223718 330882 223954
rect 330326 223398 330562 223634
rect 330646 223398 330882 223634
rect 330326 187718 330562 187954
rect 330646 187718 330882 187954
rect 330326 187398 330562 187634
rect 330646 187398 330882 187634
rect 330326 151718 330562 151954
rect 330646 151718 330882 151954
rect 330326 151398 330562 151634
rect 330646 151398 330882 151634
rect 330326 115718 330562 115954
rect 330646 115718 330882 115954
rect 330326 115398 330562 115634
rect 330646 115398 330882 115634
rect 330326 79718 330562 79954
rect 330646 79718 330882 79954
rect 330326 79398 330562 79634
rect 330646 79398 330882 79634
rect 330326 43718 330562 43954
rect 330646 43718 330882 43954
rect 330326 43398 330562 43634
rect 330646 43398 330882 43634
rect 330326 7718 330562 7954
rect 330646 7718 330882 7954
rect 330326 7398 330562 7634
rect 330646 7398 330882 7634
rect 330326 -1542 330562 -1306
rect 330646 -1542 330882 -1306
rect 330326 -1862 330562 -1626
rect 330646 -1862 330882 -1626
rect 334826 706522 335062 706758
rect 335146 706522 335382 706758
rect 334826 706202 335062 706438
rect 335146 706202 335382 706438
rect 334826 696218 335062 696454
rect 335146 696218 335382 696454
rect 334826 695898 335062 696134
rect 335146 695898 335382 696134
rect 334826 660218 335062 660454
rect 335146 660218 335382 660454
rect 334826 659898 335062 660134
rect 335146 659898 335382 660134
rect 334826 624218 335062 624454
rect 335146 624218 335382 624454
rect 334826 623898 335062 624134
rect 335146 623898 335382 624134
rect 334826 588218 335062 588454
rect 335146 588218 335382 588454
rect 334826 587898 335062 588134
rect 335146 587898 335382 588134
rect 334826 552218 335062 552454
rect 335146 552218 335382 552454
rect 334826 551898 335062 552134
rect 335146 551898 335382 552134
rect 334826 516218 335062 516454
rect 335146 516218 335382 516454
rect 334826 515898 335062 516134
rect 335146 515898 335382 516134
rect 334826 480218 335062 480454
rect 335146 480218 335382 480454
rect 334826 479898 335062 480134
rect 335146 479898 335382 480134
rect 334826 444218 335062 444454
rect 335146 444218 335382 444454
rect 334826 443898 335062 444134
rect 335146 443898 335382 444134
rect 334826 408218 335062 408454
rect 335146 408218 335382 408454
rect 334826 407898 335062 408134
rect 335146 407898 335382 408134
rect 334826 372218 335062 372454
rect 335146 372218 335382 372454
rect 334826 371898 335062 372134
rect 335146 371898 335382 372134
rect 334826 336218 335062 336454
rect 335146 336218 335382 336454
rect 334826 335898 335062 336134
rect 335146 335898 335382 336134
rect 334826 300218 335062 300454
rect 335146 300218 335382 300454
rect 334826 299898 335062 300134
rect 335146 299898 335382 300134
rect 334826 264218 335062 264454
rect 335146 264218 335382 264454
rect 334826 263898 335062 264134
rect 335146 263898 335382 264134
rect 334826 228218 335062 228454
rect 335146 228218 335382 228454
rect 334826 227898 335062 228134
rect 335146 227898 335382 228134
rect 334826 192218 335062 192454
rect 335146 192218 335382 192454
rect 334826 191898 335062 192134
rect 335146 191898 335382 192134
rect 334826 156218 335062 156454
rect 335146 156218 335382 156454
rect 334826 155898 335062 156134
rect 335146 155898 335382 156134
rect 334826 120218 335062 120454
rect 335146 120218 335382 120454
rect 334826 119898 335062 120134
rect 335146 119898 335382 120134
rect 334826 84218 335062 84454
rect 335146 84218 335382 84454
rect 334826 83898 335062 84134
rect 335146 83898 335382 84134
rect 334826 48218 335062 48454
rect 335146 48218 335382 48454
rect 334826 47898 335062 48134
rect 335146 47898 335382 48134
rect 334826 12218 335062 12454
rect 335146 12218 335382 12454
rect 334826 11898 335062 12134
rect 335146 11898 335382 12134
rect 334826 -2502 335062 -2266
rect 335146 -2502 335382 -2266
rect 334826 -2822 335062 -2586
rect 335146 -2822 335382 -2586
rect 339326 707482 339562 707718
rect 339646 707482 339882 707718
rect 339326 707162 339562 707398
rect 339646 707162 339882 707398
rect 339326 700718 339562 700954
rect 339646 700718 339882 700954
rect 339326 700398 339562 700634
rect 339646 700398 339882 700634
rect 339326 664718 339562 664954
rect 339646 664718 339882 664954
rect 339326 664398 339562 664634
rect 339646 664398 339882 664634
rect 339326 628718 339562 628954
rect 339646 628718 339882 628954
rect 339326 628398 339562 628634
rect 339646 628398 339882 628634
rect 339326 592718 339562 592954
rect 339646 592718 339882 592954
rect 339326 592398 339562 592634
rect 339646 592398 339882 592634
rect 339326 556718 339562 556954
rect 339646 556718 339882 556954
rect 339326 556398 339562 556634
rect 339646 556398 339882 556634
rect 339326 520718 339562 520954
rect 339646 520718 339882 520954
rect 339326 520398 339562 520634
rect 339646 520398 339882 520634
rect 339326 484718 339562 484954
rect 339646 484718 339882 484954
rect 339326 484398 339562 484634
rect 339646 484398 339882 484634
rect 339326 448718 339562 448954
rect 339646 448718 339882 448954
rect 339326 448398 339562 448634
rect 339646 448398 339882 448634
rect 339326 412718 339562 412954
rect 339646 412718 339882 412954
rect 339326 412398 339562 412634
rect 339646 412398 339882 412634
rect 339326 376718 339562 376954
rect 339646 376718 339882 376954
rect 339326 376398 339562 376634
rect 339646 376398 339882 376634
rect 339326 340718 339562 340954
rect 339646 340718 339882 340954
rect 339326 340398 339562 340634
rect 339646 340398 339882 340634
rect 339326 304718 339562 304954
rect 339646 304718 339882 304954
rect 339326 304398 339562 304634
rect 339646 304398 339882 304634
rect 339326 268718 339562 268954
rect 339646 268718 339882 268954
rect 339326 268398 339562 268634
rect 339646 268398 339882 268634
rect 339326 232718 339562 232954
rect 339646 232718 339882 232954
rect 339326 232398 339562 232634
rect 339646 232398 339882 232634
rect 339326 196718 339562 196954
rect 339646 196718 339882 196954
rect 339326 196398 339562 196634
rect 339646 196398 339882 196634
rect 339326 160718 339562 160954
rect 339646 160718 339882 160954
rect 339326 160398 339562 160634
rect 339646 160398 339882 160634
rect 339326 124718 339562 124954
rect 339646 124718 339882 124954
rect 339326 124398 339562 124634
rect 339646 124398 339882 124634
rect 339326 88718 339562 88954
rect 339646 88718 339882 88954
rect 339326 88398 339562 88634
rect 339646 88398 339882 88634
rect 339326 52718 339562 52954
rect 339646 52718 339882 52954
rect 339326 52398 339562 52634
rect 339646 52398 339882 52634
rect 339326 16718 339562 16954
rect 339646 16718 339882 16954
rect 339326 16398 339562 16634
rect 339646 16398 339882 16634
rect 339326 -3462 339562 -3226
rect 339646 -3462 339882 -3226
rect 339326 -3782 339562 -3546
rect 339646 -3782 339882 -3546
rect 343826 708442 344062 708678
rect 344146 708442 344382 708678
rect 343826 708122 344062 708358
rect 344146 708122 344382 708358
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 343826 561218 344062 561454
rect 344146 561218 344382 561454
rect 343826 560898 344062 561134
rect 344146 560898 344382 561134
rect 343826 525218 344062 525454
rect 344146 525218 344382 525454
rect 343826 524898 344062 525134
rect 344146 524898 344382 525134
rect 343826 489218 344062 489454
rect 344146 489218 344382 489454
rect 343826 488898 344062 489134
rect 344146 488898 344382 489134
rect 343826 453218 344062 453454
rect 344146 453218 344382 453454
rect 343826 452898 344062 453134
rect 344146 452898 344382 453134
rect 343826 417218 344062 417454
rect 344146 417218 344382 417454
rect 343826 416898 344062 417134
rect 344146 416898 344382 417134
rect 343826 381218 344062 381454
rect 344146 381218 344382 381454
rect 343826 380898 344062 381134
rect 344146 380898 344382 381134
rect 343826 345218 344062 345454
rect 344146 345218 344382 345454
rect 343826 344898 344062 345134
rect 344146 344898 344382 345134
rect 343826 309218 344062 309454
rect 344146 309218 344382 309454
rect 343826 308898 344062 309134
rect 344146 308898 344382 309134
rect 343826 273218 344062 273454
rect 344146 273218 344382 273454
rect 343826 272898 344062 273134
rect 344146 272898 344382 273134
rect 343826 237218 344062 237454
rect 344146 237218 344382 237454
rect 343826 236898 344062 237134
rect 344146 236898 344382 237134
rect 343826 201218 344062 201454
rect 344146 201218 344382 201454
rect 343826 200898 344062 201134
rect 344146 200898 344382 201134
rect 343826 165218 344062 165454
rect 344146 165218 344382 165454
rect 343826 164898 344062 165134
rect 344146 164898 344382 165134
rect 343826 129218 344062 129454
rect 344146 129218 344382 129454
rect 343826 128898 344062 129134
rect 344146 128898 344382 129134
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -4422 344062 -4186
rect 344146 -4422 344382 -4186
rect 343826 -4742 344062 -4506
rect 344146 -4742 344382 -4506
rect 348326 709402 348562 709638
rect 348646 709402 348882 709638
rect 348326 709082 348562 709318
rect 348646 709082 348882 709318
rect 348326 673718 348562 673954
rect 348646 673718 348882 673954
rect 348326 673398 348562 673634
rect 348646 673398 348882 673634
rect 348326 637718 348562 637954
rect 348646 637718 348882 637954
rect 348326 637398 348562 637634
rect 348646 637398 348882 637634
rect 348326 601718 348562 601954
rect 348646 601718 348882 601954
rect 348326 601398 348562 601634
rect 348646 601398 348882 601634
rect 348326 565718 348562 565954
rect 348646 565718 348882 565954
rect 348326 565398 348562 565634
rect 348646 565398 348882 565634
rect 348326 529718 348562 529954
rect 348646 529718 348882 529954
rect 348326 529398 348562 529634
rect 348646 529398 348882 529634
rect 348326 493718 348562 493954
rect 348646 493718 348882 493954
rect 348326 493398 348562 493634
rect 348646 493398 348882 493634
rect 348326 457718 348562 457954
rect 348646 457718 348882 457954
rect 348326 457398 348562 457634
rect 348646 457398 348882 457634
rect 348326 421718 348562 421954
rect 348646 421718 348882 421954
rect 348326 421398 348562 421634
rect 348646 421398 348882 421634
rect 348326 385718 348562 385954
rect 348646 385718 348882 385954
rect 348326 385398 348562 385634
rect 348646 385398 348882 385634
rect 348326 349718 348562 349954
rect 348646 349718 348882 349954
rect 348326 349398 348562 349634
rect 348646 349398 348882 349634
rect 348326 313718 348562 313954
rect 348646 313718 348882 313954
rect 348326 313398 348562 313634
rect 348646 313398 348882 313634
rect 348326 277718 348562 277954
rect 348646 277718 348882 277954
rect 348326 277398 348562 277634
rect 348646 277398 348882 277634
rect 348326 241718 348562 241954
rect 348646 241718 348882 241954
rect 348326 241398 348562 241634
rect 348646 241398 348882 241634
rect 348326 205718 348562 205954
rect 348646 205718 348882 205954
rect 348326 205398 348562 205634
rect 348646 205398 348882 205634
rect 348326 169718 348562 169954
rect 348646 169718 348882 169954
rect 348326 169398 348562 169634
rect 348646 169398 348882 169634
rect 348326 133718 348562 133954
rect 348646 133718 348882 133954
rect 348326 133398 348562 133634
rect 348646 133398 348882 133634
rect 348326 97718 348562 97954
rect 348646 97718 348882 97954
rect 348326 97398 348562 97634
rect 348646 97398 348882 97634
rect 348326 61718 348562 61954
rect 348646 61718 348882 61954
rect 348326 61398 348562 61634
rect 348646 61398 348882 61634
rect 348326 25718 348562 25954
rect 348646 25718 348882 25954
rect 348326 25398 348562 25634
rect 348646 25398 348882 25634
rect 348326 -5382 348562 -5146
rect 348646 -5382 348882 -5146
rect 348326 -5702 348562 -5466
rect 348646 -5702 348882 -5466
rect 352826 710362 353062 710598
rect 353146 710362 353382 710598
rect 352826 710042 353062 710278
rect 353146 710042 353382 710278
rect 352826 678218 353062 678454
rect 353146 678218 353382 678454
rect 352826 677898 353062 678134
rect 353146 677898 353382 678134
rect 352826 642218 353062 642454
rect 353146 642218 353382 642454
rect 352826 641898 353062 642134
rect 353146 641898 353382 642134
rect 352826 606218 353062 606454
rect 353146 606218 353382 606454
rect 352826 605898 353062 606134
rect 353146 605898 353382 606134
rect 352826 570218 353062 570454
rect 353146 570218 353382 570454
rect 352826 569898 353062 570134
rect 353146 569898 353382 570134
rect 352826 534218 353062 534454
rect 353146 534218 353382 534454
rect 352826 533898 353062 534134
rect 353146 533898 353382 534134
rect 352826 498218 353062 498454
rect 353146 498218 353382 498454
rect 352826 497898 353062 498134
rect 353146 497898 353382 498134
rect 352826 462218 353062 462454
rect 353146 462218 353382 462454
rect 352826 461898 353062 462134
rect 353146 461898 353382 462134
rect 352826 426218 353062 426454
rect 353146 426218 353382 426454
rect 352826 425898 353062 426134
rect 353146 425898 353382 426134
rect 352826 390218 353062 390454
rect 353146 390218 353382 390454
rect 352826 389898 353062 390134
rect 353146 389898 353382 390134
rect 352826 354218 353062 354454
rect 353146 354218 353382 354454
rect 352826 353898 353062 354134
rect 353146 353898 353382 354134
rect 352826 318218 353062 318454
rect 353146 318218 353382 318454
rect 352826 317898 353062 318134
rect 353146 317898 353382 318134
rect 352826 282218 353062 282454
rect 353146 282218 353382 282454
rect 352826 281898 353062 282134
rect 353146 281898 353382 282134
rect 352826 246218 353062 246454
rect 353146 246218 353382 246454
rect 352826 245898 353062 246134
rect 353146 245898 353382 246134
rect 352826 210218 353062 210454
rect 353146 210218 353382 210454
rect 352826 209898 353062 210134
rect 353146 209898 353382 210134
rect 352826 174218 353062 174454
rect 353146 174218 353382 174454
rect 352826 173898 353062 174134
rect 353146 173898 353382 174134
rect 352826 138218 353062 138454
rect 353146 138218 353382 138454
rect 352826 137898 353062 138134
rect 353146 137898 353382 138134
rect 352826 102218 353062 102454
rect 353146 102218 353382 102454
rect 352826 101898 353062 102134
rect 353146 101898 353382 102134
rect 352826 66218 353062 66454
rect 353146 66218 353382 66454
rect 352826 65898 353062 66134
rect 353146 65898 353382 66134
rect 352826 30218 353062 30454
rect 353146 30218 353382 30454
rect 352826 29898 353062 30134
rect 353146 29898 353382 30134
rect 352826 -6342 353062 -6106
rect 353146 -6342 353382 -6106
rect 352826 -6662 353062 -6426
rect 353146 -6662 353382 -6426
rect 357326 711322 357562 711558
rect 357646 711322 357882 711558
rect 357326 711002 357562 711238
rect 357646 711002 357882 711238
rect 357326 682718 357562 682954
rect 357646 682718 357882 682954
rect 357326 682398 357562 682634
rect 357646 682398 357882 682634
rect 357326 646718 357562 646954
rect 357646 646718 357882 646954
rect 357326 646398 357562 646634
rect 357646 646398 357882 646634
rect 357326 610718 357562 610954
rect 357646 610718 357882 610954
rect 357326 610398 357562 610634
rect 357646 610398 357882 610634
rect 357326 574718 357562 574954
rect 357646 574718 357882 574954
rect 357326 574398 357562 574634
rect 357646 574398 357882 574634
rect 357326 538718 357562 538954
rect 357646 538718 357882 538954
rect 357326 538398 357562 538634
rect 357646 538398 357882 538634
rect 357326 502718 357562 502954
rect 357646 502718 357882 502954
rect 357326 502398 357562 502634
rect 357646 502398 357882 502634
rect 357326 466718 357562 466954
rect 357646 466718 357882 466954
rect 357326 466398 357562 466634
rect 357646 466398 357882 466634
rect 357326 430718 357562 430954
rect 357646 430718 357882 430954
rect 357326 430398 357562 430634
rect 357646 430398 357882 430634
rect 357326 394718 357562 394954
rect 357646 394718 357882 394954
rect 357326 394398 357562 394634
rect 357646 394398 357882 394634
rect 357326 358718 357562 358954
rect 357646 358718 357882 358954
rect 357326 358398 357562 358634
rect 357646 358398 357882 358634
rect 357326 322718 357562 322954
rect 357646 322718 357882 322954
rect 357326 322398 357562 322634
rect 357646 322398 357882 322634
rect 357326 286718 357562 286954
rect 357646 286718 357882 286954
rect 357326 286398 357562 286634
rect 357646 286398 357882 286634
rect 357326 250718 357562 250954
rect 357646 250718 357882 250954
rect 357326 250398 357562 250634
rect 357646 250398 357882 250634
rect 357326 214718 357562 214954
rect 357646 214718 357882 214954
rect 357326 214398 357562 214634
rect 357646 214398 357882 214634
rect 357326 178718 357562 178954
rect 357646 178718 357882 178954
rect 357326 178398 357562 178634
rect 357646 178398 357882 178634
rect 357326 142718 357562 142954
rect 357646 142718 357882 142954
rect 357326 142398 357562 142634
rect 357646 142398 357882 142634
rect 357326 106718 357562 106954
rect 357646 106718 357882 106954
rect 357326 106398 357562 106634
rect 357646 106398 357882 106634
rect 357326 70718 357562 70954
rect 357646 70718 357882 70954
rect 357326 70398 357562 70634
rect 357646 70398 357882 70634
rect 357326 34718 357562 34954
rect 357646 34718 357882 34954
rect 357326 34398 357562 34634
rect 357646 34398 357882 34634
rect 357326 -7302 357562 -7066
rect 357646 -7302 357882 -7066
rect 357326 -7622 357562 -7386
rect 357646 -7622 357882 -7386
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 366326 705562 366562 705798
rect 366646 705562 366882 705798
rect 366326 705242 366562 705478
rect 366646 705242 366882 705478
rect 366326 691718 366562 691954
rect 366646 691718 366882 691954
rect 366326 691398 366562 691634
rect 366646 691398 366882 691634
rect 366326 655718 366562 655954
rect 366646 655718 366882 655954
rect 366326 655398 366562 655634
rect 366646 655398 366882 655634
rect 366326 619718 366562 619954
rect 366646 619718 366882 619954
rect 366326 619398 366562 619634
rect 366646 619398 366882 619634
rect 366326 583718 366562 583954
rect 366646 583718 366882 583954
rect 366326 583398 366562 583634
rect 366646 583398 366882 583634
rect 366326 547718 366562 547954
rect 366646 547718 366882 547954
rect 366326 547398 366562 547634
rect 366646 547398 366882 547634
rect 366326 511718 366562 511954
rect 366646 511718 366882 511954
rect 366326 511398 366562 511634
rect 366646 511398 366882 511634
rect 366326 475718 366562 475954
rect 366646 475718 366882 475954
rect 366326 475398 366562 475634
rect 366646 475398 366882 475634
rect 366326 439718 366562 439954
rect 366646 439718 366882 439954
rect 366326 439398 366562 439634
rect 366646 439398 366882 439634
rect 366326 403718 366562 403954
rect 366646 403718 366882 403954
rect 366326 403398 366562 403634
rect 366646 403398 366882 403634
rect 366326 367718 366562 367954
rect 366646 367718 366882 367954
rect 366326 367398 366562 367634
rect 366646 367398 366882 367634
rect 366326 331718 366562 331954
rect 366646 331718 366882 331954
rect 366326 331398 366562 331634
rect 366646 331398 366882 331634
rect 366326 295718 366562 295954
rect 366646 295718 366882 295954
rect 366326 295398 366562 295634
rect 366646 295398 366882 295634
rect 366326 259718 366562 259954
rect 366646 259718 366882 259954
rect 366326 259398 366562 259634
rect 366646 259398 366882 259634
rect 366326 223718 366562 223954
rect 366646 223718 366882 223954
rect 366326 223398 366562 223634
rect 366646 223398 366882 223634
rect 366326 187718 366562 187954
rect 366646 187718 366882 187954
rect 366326 187398 366562 187634
rect 366646 187398 366882 187634
rect 366326 151718 366562 151954
rect 366646 151718 366882 151954
rect 366326 151398 366562 151634
rect 366646 151398 366882 151634
rect 366326 115718 366562 115954
rect 366646 115718 366882 115954
rect 366326 115398 366562 115634
rect 366646 115398 366882 115634
rect 366326 79718 366562 79954
rect 366646 79718 366882 79954
rect 366326 79398 366562 79634
rect 366646 79398 366882 79634
rect 366326 43718 366562 43954
rect 366646 43718 366882 43954
rect 366326 43398 366562 43634
rect 366646 43398 366882 43634
rect 366326 7718 366562 7954
rect 366646 7718 366882 7954
rect 366326 7398 366562 7634
rect 366646 7398 366882 7634
rect 366326 -1542 366562 -1306
rect 366646 -1542 366882 -1306
rect 366326 -1862 366562 -1626
rect 366646 -1862 366882 -1626
rect 370826 706522 371062 706758
rect 371146 706522 371382 706758
rect 370826 706202 371062 706438
rect 371146 706202 371382 706438
rect 370826 696218 371062 696454
rect 371146 696218 371382 696454
rect 370826 695898 371062 696134
rect 371146 695898 371382 696134
rect 370826 660218 371062 660454
rect 371146 660218 371382 660454
rect 370826 659898 371062 660134
rect 371146 659898 371382 660134
rect 370826 624218 371062 624454
rect 371146 624218 371382 624454
rect 370826 623898 371062 624134
rect 371146 623898 371382 624134
rect 370826 588218 371062 588454
rect 371146 588218 371382 588454
rect 370826 587898 371062 588134
rect 371146 587898 371382 588134
rect 370826 552218 371062 552454
rect 371146 552218 371382 552454
rect 370826 551898 371062 552134
rect 371146 551898 371382 552134
rect 370826 516218 371062 516454
rect 371146 516218 371382 516454
rect 370826 515898 371062 516134
rect 371146 515898 371382 516134
rect 370826 480218 371062 480454
rect 371146 480218 371382 480454
rect 370826 479898 371062 480134
rect 371146 479898 371382 480134
rect 370826 444218 371062 444454
rect 371146 444218 371382 444454
rect 370826 443898 371062 444134
rect 371146 443898 371382 444134
rect 370826 408218 371062 408454
rect 371146 408218 371382 408454
rect 370826 407898 371062 408134
rect 371146 407898 371382 408134
rect 370826 372218 371062 372454
rect 371146 372218 371382 372454
rect 370826 371898 371062 372134
rect 371146 371898 371382 372134
rect 370826 336218 371062 336454
rect 371146 336218 371382 336454
rect 370826 335898 371062 336134
rect 371146 335898 371382 336134
rect 370826 300218 371062 300454
rect 371146 300218 371382 300454
rect 370826 299898 371062 300134
rect 371146 299898 371382 300134
rect 370826 264218 371062 264454
rect 371146 264218 371382 264454
rect 370826 263898 371062 264134
rect 371146 263898 371382 264134
rect 370826 228218 371062 228454
rect 371146 228218 371382 228454
rect 370826 227898 371062 228134
rect 371146 227898 371382 228134
rect 370826 192218 371062 192454
rect 371146 192218 371382 192454
rect 370826 191898 371062 192134
rect 371146 191898 371382 192134
rect 370826 156218 371062 156454
rect 371146 156218 371382 156454
rect 370826 155898 371062 156134
rect 371146 155898 371382 156134
rect 370826 120218 371062 120454
rect 371146 120218 371382 120454
rect 370826 119898 371062 120134
rect 371146 119898 371382 120134
rect 370826 84218 371062 84454
rect 371146 84218 371382 84454
rect 370826 83898 371062 84134
rect 371146 83898 371382 84134
rect 370826 48218 371062 48454
rect 371146 48218 371382 48454
rect 370826 47898 371062 48134
rect 371146 47898 371382 48134
rect 370826 12218 371062 12454
rect 371146 12218 371382 12454
rect 370826 11898 371062 12134
rect 371146 11898 371382 12134
rect 370826 -2502 371062 -2266
rect 371146 -2502 371382 -2266
rect 370826 -2822 371062 -2586
rect 371146 -2822 371382 -2586
rect 375326 707482 375562 707718
rect 375646 707482 375882 707718
rect 375326 707162 375562 707398
rect 375646 707162 375882 707398
rect 375326 700718 375562 700954
rect 375646 700718 375882 700954
rect 375326 700398 375562 700634
rect 375646 700398 375882 700634
rect 375326 664718 375562 664954
rect 375646 664718 375882 664954
rect 375326 664398 375562 664634
rect 375646 664398 375882 664634
rect 375326 628718 375562 628954
rect 375646 628718 375882 628954
rect 375326 628398 375562 628634
rect 375646 628398 375882 628634
rect 375326 592718 375562 592954
rect 375646 592718 375882 592954
rect 375326 592398 375562 592634
rect 375646 592398 375882 592634
rect 375326 556718 375562 556954
rect 375646 556718 375882 556954
rect 375326 556398 375562 556634
rect 375646 556398 375882 556634
rect 375326 520718 375562 520954
rect 375646 520718 375882 520954
rect 375326 520398 375562 520634
rect 375646 520398 375882 520634
rect 375326 484718 375562 484954
rect 375646 484718 375882 484954
rect 375326 484398 375562 484634
rect 375646 484398 375882 484634
rect 375326 448718 375562 448954
rect 375646 448718 375882 448954
rect 375326 448398 375562 448634
rect 375646 448398 375882 448634
rect 375326 412718 375562 412954
rect 375646 412718 375882 412954
rect 375326 412398 375562 412634
rect 375646 412398 375882 412634
rect 375326 376718 375562 376954
rect 375646 376718 375882 376954
rect 375326 376398 375562 376634
rect 375646 376398 375882 376634
rect 375326 340718 375562 340954
rect 375646 340718 375882 340954
rect 375326 340398 375562 340634
rect 375646 340398 375882 340634
rect 375326 304718 375562 304954
rect 375646 304718 375882 304954
rect 375326 304398 375562 304634
rect 375646 304398 375882 304634
rect 375326 268718 375562 268954
rect 375646 268718 375882 268954
rect 375326 268398 375562 268634
rect 375646 268398 375882 268634
rect 375326 232718 375562 232954
rect 375646 232718 375882 232954
rect 375326 232398 375562 232634
rect 375646 232398 375882 232634
rect 375326 196718 375562 196954
rect 375646 196718 375882 196954
rect 375326 196398 375562 196634
rect 375646 196398 375882 196634
rect 375326 160718 375562 160954
rect 375646 160718 375882 160954
rect 375326 160398 375562 160634
rect 375646 160398 375882 160634
rect 375326 124718 375562 124954
rect 375646 124718 375882 124954
rect 375326 124398 375562 124634
rect 375646 124398 375882 124634
rect 375326 88718 375562 88954
rect 375646 88718 375882 88954
rect 375326 88398 375562 88634
rect 375646 88398 375882 88634
rect 375326 52718 375562 52954
rect 375646 52718 375882 52954
rect 375326 52398 375562 52634
rect 375646 52398 375882 52634
rect 375326 16718 375562 16954
rect 375646 16718 375882 16954
rect 375326 16398 375562 16634
rect 375646 16398 375882 16634
rect 375326 -3462 375562 -3226
rect 375646 -3462 375882 -3226
rect 375326 -3782 375562 -3546
rect 375646 -3782 375882 -3546
rect 379826 708442 380062 708678
rect 380146 708442 380382 708678
rect 379826 708122 380062 708358
rect 380146 708122 380382 708358
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 379826 417218 380062 417454
rect 380146 417218 380382 417454
rect 379826 416898 380062 417134
rect 380146 416898 380382 417134
rect 379826 381218 380062 381454
rect 380146 381218 380382 381454
rect 379826 380898 380062 381134
rect 380146 380898 380382 381134
rect 379826 345218 380062 345454
rect 380146 345218 380382 345454
rect 379826 344898 380062 345134
rect 380146 344898 380382 345134
rect 379826 309218 380062 309454
rect 380146 309218 380382 309454
rect 379826 308898 380062 309134
rect 380146 308898 380382 309134
rect 379826 273218 380062 273454
rect 380146 273218 380382 273454
rect 379826 272898 380062 273134
rect 380146 272898 380382 273134
rect 379826 237218 380062 237454
rect 380146 237218 380382 237454
rect 379826 236898 380062 237134
rect 380146 236898 380382 237134
rect 379826 201218 380062 201454
rect 380146 201218 380382 201454
rect 379826 200898 380062 201134
rect 380146 200898 380382 201134
rect 379826 165218 380062 165454
rect 380146 165218 380382 165454
rect 379826 164898 380062 165134
rect 380146 164898 380382 165134
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -4422 380062 -4186
rect 380146 -4422 380382 -4186
rect 379826 -4742 380062 -4506
rect 380146 -4742 380382 -4506
rect 384326 709402 384562 709638
rect 384646 709402 384882 709638
rect 384326 709082 384562 709318
rect 384646 709082 384882 709318
rect 384326 673718 384562 673954
rect 384646 673718 384882 673954
rect 384326 673398 384562 673634
rect 384646 673398 384882 673634
rect 384326 637718 384562 637954
rect 384646 637718 384882 637954
rect 384326 637398 384562 637634
rect 384646 637398 384882 637634
rect 384326 601718 384562 601954
rect 384646 601718 384882 601954
rect 384326 601398 384562 601634
rect 384646 601398 384882 601634
rect 384326 565718 384562 565954
rect 384646 565718 384882 565954
rect 384326 565398 384562 565634
rect 384646 565398 384882 565634
rect 384326 529718 384562 529954
rect 384646 529718 384882 529954
rect 384326 529398 384562 529634
rect 384646 529398 384882 529634
rect 384326 493718 384562 493954
rect 384646 493718 384882 493954
rect 384326 493398 384562 493634
rect 384646 493398 384882 493634
rect 384326 457718 384562 457954
rect 384646 457718 384882 457954
rect 384326 457398 384562 457634
rect 384646 457398 384882 457634
rect 384326 421718 384562 421954
rect 384646 421718 384882 421954
rect 384326 421398 384562 421634
rect 384646 421398 384882 421634
rect 384326 385718 384562 385954
rect 384646 385718 384882 385954
rect 384326 385398 384562 385634
rect 384646 385398 384882 385634
rect 384326 349718 384562 349954
rect 384646 349718 384882 349954
rect 384326 349398 384562 349634
rect 384646 349398 384882 349634
rect 384326 313718 384562 313954
rect 384646 313718 384882 313954
rect 384326 313398 384562 313634
rect 384646 313398 384882 313634
rect 384326 277718 384562 277954
rect 384646 277718 384882 277954
rect 384326 277398 384562 277634
rect 384646 277398 384882 277634
rect 384326 241718 384562 241954
rect 384646 241718 384882 241954
rect 384326 241398 384562 241634
rect 384646 241398 384882 241634
rect 384326 205718 384562 205954
rect 384646 205718 384882 205954
rect 384326 205398 384562 205634
rect 384646 205398 384882 205634
rect 384326 169718 384562 169954
rect 384646 169718 384882 169954
rect 384326 169398 384562 169634
rect 384646 169398 384882 169634
rect 384326 133718 384562 133954
rect 384646 133718 384882 133954
rect 384326 133398 384562 133634
rect 384646 133398 384882 133634
rect 384326 97718 384562 97954
rect 384646 97718 384882 97954
rect 384326 97398 384562 97634
rect 384646 97398 384882 97634
rect 384326 61718 384562 61954
rect 384646 61718 384882 61954
rect 384326 61398 384562 61634
rect 384646 61398 384882 61634
rect 384326 25718 384562 25954
rect 384646 25718 384882 25954
rect 384326 25398 384562 25634
rect 384646 25398 384882 25634
rect 384326 -5382 384562 -5146
rect 384646 -5382 384882 -5146
rect 384326 -5702 384562 -5466
rect 384646 -5702 384882 -5466
rect 388826 710362 389062 710598
rect 389146 710362 389382 710598
rect 388826 710042 389062 710278
rect 389146 710042 389382 710278
rect 388826 678218 389062 678454
rect 389146 678218 389382 678454
rect 388826 677898 389062 678134
rect 389146 677898 389382 678134
rect 388826 642218 389062 642454
rect 389146 642218 389382 642454
rect 388826 641898 389062 642134
rect 389146 641898 389382 642134
rect 388826 606218 389062 606454
rect 389146 606218 389382 606454
rect 388826 605898 389062 606134
rect 389146 605898 389382 606134
rect 388826 570218 389062 570454
rect 389146 570218 389382 570454
rect 388826 569898 389062 570134
rect 389146 569898 389382 570134
rect 388826 534218 389062 534454
rect 389146 534218 389382 534454
rect 388826 533898 389062 534134
rect 389146 533898 389382 534134
rect 388826 498218 389062 498454
rect 389146 498218 389382 498454
rect 388826 497898 389062 498134
rect 389146 497898 389382 498134
rect 388826 462218 389062 462454
rect 389146 462218 389382 462454
rect 388826 461898 389062 462134
rect 389146 461898 389382 462134
rect 388826 426218 389062 426454
rect 389146 426218 389382 426454
rect 388826 425898 389062 426134
rect 389146 425898 389382 426134
rect 388826 390218 389062 390454
rect 389146 390218 389382 390454
rect 388826 389898 389062 390134
rect 389146 389898 389382 390134
rect 388826 354218 389062 354454
rect 389146 354218 389382 354454
rect 388826 353898 389062 354134
rect 389146 353898 389382 354134
rect 388826 318218 389062 318454
rect 389146 318218 389382 318454
rect 388826 317898 389062 318134
rect 389146 317898 389382 318134
rect 388826 282218 389062 282454
rect 389146 282218 389382 282454
rect 388826 281898 389062 282134
rect 389146 281898 389382 282134
rect 388826 246218 389062 246454
rect 389146 246218 389382 246454
rect 388826 245898 389062 246134
rect 389146 245898 389382 246134
rect 388826 210218 389062 210454
rect 389146 210218 389382 210454
rect 388826 209898 389062 210134
rect 389146 209898 389382 210134
rect 388826 174218 389062 174454
rect 389146 174218 389382 174454
rect 388826 173898 389062 174134
rect 389146 173898 389382 174134
rect 388826 138218 389062 138454
rect 389146 138218 389382 138454
rect 388826 137898 389062 138134
rect 389146 137898 389382 138134
rect 388826 102218 389062 102454
rect 389146 102218 389382 102454
rect 388826 101898 389062 102134
rect 389146 101898 389382 102134
rect 388826 66218 389062 66454
rect 389146 66218 389382 66454
rect 388826 65898 389062 66134
rect 389146 65898 389382 66134
rect 388826 30218 389062 30454
rect 389146 30218 389382 30454
rect 388826 29898 389062 30134
rect 389146 29898 389382 30134
rect 388826 -6342 389062 -6106
rect 389146 -6342 389382 -6106
rect 388826 -6662 389062 -6426
rect 389146 -6662 389382 -6426
rect 393326 711322 393562 711558
rect 393646 711322 393882 711558
rect 393326 711002 393562 711238
rect 393646 711002 393882 711238
rect 393326 682718 393562 682954
rect 393646 682718 393882 682954
rect 393326 682398 393562 682634
rect 393646 682398 393882 682634
rect 393326 646718 393562 646954
rect 393646 646718 393882 646954
rect 393326 646398 393562 646634
rect 393646 646398 393882 646634
rect 393326 610718 393562 610954
rect 393646 610718 393882 610954
rect 393326 610398 393562 610634
rect 393646 610398 393882 610634
rect 393326 574718 393562 574954
rect 393646 574718 393882 574954
rect 393326 574398 393562 574634
rect 393646 574398 393882 574634
rect 393326 538718 393562 538954
rect 393646 538718 393882 538954
rect 393326 538398 393562 538634
rect 393646 538398 393882 538634
rect 393326 502718 393562 502954
rect 393646 502718 393882 502954
rect 393326 502398 393562 502634
rect 393646 502398 393882 502634
rect 393326 466718 393562 466954
rect 393646 466718 393882 466954
rect 393326 466398 393562 466634
rect 393646 466398 393882 466634
rect 393326 430718 393562 430954
rect 393646 430718 393882 430954
rect 393326 430398 393562 430634
rect 393646 430398 393882 430634
rect 393326 394718 393562 394954
rect 393646 394718 393882 394954
rect 393326 394398 393562 394634
rect 393646 394398 393882 394634
rect 393326 358718 393562 358954
rect 393646 358718 393882 358954
rect 393326 358398 393562 358634
rect 393646 358398 393882 358634
rect 393326 322718 393562 322954
rect 393646 322718 393882 322954
rect 393326 322398 393562 322634
rect 393646 322398 393882 322634
rect 393326 286718 393562 286954
rect 393646 286718 393882 286954
rect 393326 286398 393562 286634
rect 393646 286398 393882 286634
rect 393326 250718 393562 250954
rect 393646 250718 393882 250954
rect 393326 250398 393562 250634
rect 393646 250398 393882 250634
rect 393326 214718 393562 214954
rect 393646 214718 393882 214954
rect 393326 214398 393562 214634
rect 393646 214398 393882 214634
rect 393326 178718 393562 178954
rect 393646 178718 393882 178954
rect 393326 178398 393562 178634
rect 393646 178398 393882 178634
rect 393326 142718 393562 142954
rect 393646 142718 393882 142954
rect 393326 142398 393562 142634
rect 393646 142398 393882 142634
rect 393326 106718 393562 106954
rect 393646 106718 393882 106954
rect 393326 106398 393562 106634
rect 393646 106398 393882 106634
rect 393326 70718 393562 70954
rect 393646 70718 393882 70954
rect 393326 70398 393562 70634
rect 393646 70398 393882 70634
rect 393326 34718 393562 34954
rect 393646 34718 393882 34954
rect 393326 34398 393562 34634
rect 393646 34398 393882 34634
rect 393326 -7302 393562 -7066
rect 393646 -7302 393882 -7066
rect 393326 -7622 393562 -7386
rect 393646 -7622 393882 -7386
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 402326 705562 402562 705798
rect 402646 705562 402882 705798
rect 402326 705242 402562 705478
rect 402646 705242 402882 705478
rect 402326 691718 402562 691954
rect 402646 691718 402882 691954
rect 402326 691398 402562 691634
rect 402646 691398 402882 691634
rect 402326 655718 402562 655954
rect 402646 655718 402882 655954
rect 402326 655398 402562 655634
rect 402646 655398 402882 655634
rect 402326 619718 402562 619954
rect 402646 619718 402882 619954
rect 402326 619398 402562 619634
rect 402646 619398 402882 619634
rect 402326 583718 402562 583954
rect 402646 583718 402882 583954
rect 402326 583398 402562 583634
rect 402646 583398 402882 583634
rect 402326 547718 402562 547954
rect 402646 547718 402882 547954
rect 402326 547398 402562 547634
rect 402646 547398 402882 547634
rect 402326 511718 402562 511954
rect 402646 511718 402882 511954
rect 402326 511398 402562 511634
rect 402646 511398 402882 511634
rect 402326 475718 402562 475954
rect 402646 475718 402882 475954
rect 402326 475398 402562 475634
rect 402646 475398 402882 475634
rect 402326 439718 402562 439954
rect 402646 439718 402882 439954
rect 402326 439398 402562 439634
rect 402646 439398 402882 439634
rect 402326 403718 402562 403954
rect 402646 403718 402882 403954
rect 402326 403398 402562 403634
rect 402646 403398 402882 403634
rect 402326 367718 402562 367954
rect 402646 367718 402882 367954
rect 402326 367398 402562 367634
rect 402646 367398 402882 367634
rect 402326 331718 402562 331954
rect 402646 331718 402882 331954
rect 402326 331398 402562 331634
rect 402646 331398 402882 331634
rect 402326 295718 402562 295954
rect 402646 295718 402882 295954
rect 402326 295398 402562 295634
rect 402646 295398 402882 295634
rect 402326 259718 402562 259954
rect 402646 259718 402882 259954
rect 402326 259398 402562 259634
rect 402646 259398 402882 259634
rect 402326 223718 402562 223954
rect 402646 223718 402882 223954
rect 402326 223398 402562 223634
rect 402646 223398 402882 223634
rect 402326 187718 402562 187954
rect 402646 187718 402882 187954
rect 402326 187398 402562 187634
rect 402646 187398 402882 187634
rect 402326 151718 402562 151954
rect 402646 151718 402882 151954
rect 402326 151398 402562 151634
rect 402646 151398 402882 151634
rect 402326 115718 402562 115954
rect 402646 115718 402882 115954
rect 402326 115398 402562 115634
rect 402646 115398 402882 115634
rect 402326 79718 402562 79954
rect 402646 79718 402882 79954
rect 402326 79398 402562 79634
rect 402646 79398 402882 79634
rect 402326 43718 402562 43954
rect 402646 43718 402882 43954
rect 402326 43398 402562 43634
rect 402646 43398 402882 43634
rect 402326 7718 402562 7954
rect 402646 7718 402882 7954
rect 402326 7398 402562 7634
rect 402646 7398 402882 7634
rect 402326 -1542 402562 -1306
rect 402646 -1542 402882 -1306
rect 402326 -1862 402562 -1626
rect 402646 -1862 402882 -1626
rect 406826 706522 407062 706758
rect 407146 706522 407382 706758
rect 406826 706202 407062 706438
rect 407146 706202 407382 706438
rect 406826 696218 407062 696454
rect 407146 696218 407382 696454
rect 406826 695898 407062 696134
rect 407146 695898 407382 696134
rect 406826 660218 407062 660454
rect 407146 660218 407382 660454
rect 406826 659898 407062 660134
rect 407146 659898 407382 660134
rect 406826 624218 407062 624454
rect 407146 624218 407382 624454
rect 406826 623898 407062 624134
rect 407146 623898 407382 624134
rect 406826 588218 407062 588454
rect 407146 588218 407382 588454
rect 406826 587898 407062 588134
rect 407146 587898 407382 588134
rect 406826 552218 407062 552454
rect 407146 552218 407382 552454
rect 406826 551898 407062 552134
rect 407146 551898 407382 552134
rect 406826 516218 407062 516454
rect 407146 516218 407382 516454
rect 406826 515898 407062 516134
rect 407146 515898 407382 516134
rect 406826 480218 407062 480454
rect 407146 480218 407382 480454
rect 406826 479898 407062 480134
rect 407146 479898 407382 480134
rect 406826 444218 407062 444454
rect 407146 444218 407382 444454
rect 406826 443898 407062 444134
rect 407146 443898 407382 444134
rect 406826 408218 407062 408454
rect 407146 408218 407382 408454
rect 406826 407898 407062 408134
rect 407146 407898 407382 408134
rect 406826 372218 407062 372454
rect 407146 372218 407382 372454
rect 406826 371898 407062 372134
rect 407146 371898 407382 372134
rect 406826 336218 407062 336454
rect 407146 336218 407382 336454
rect 406826 335898 407062 336134
rect 407146 335898 407382 336134
rect 406826 300218 407062 300454
rect 407146 300218 407382 300454
rect 406826 299898 407062 300134
rect 407146 299898 407382 300134
rect 406826 264218 407062 264454
rect 407146 264218 407382 264454
rect 406826 263898 407062 264134
rect 407146 263898 407382 264134
rect 406826 228218 407062 228454
rect 407146 228218 407382 228454
rect 406826 227898 407062 228134
rect 407146 227898 407382 228134
rect 406826 192218 407062 192454
rect 407146 192218 407382 192454
rect 406826 191898 407062 192134
rect 407146 191898 407382 192134
rect 406826 156218 407062 156454
rect 407146 156218 407382 156454
rect 406826 155898 407062 156134
rect 407146 155898 407382 156134
rect 406826 120218 407062 120454
rect 407146 120218 407382 120454
rect 406826 119898 407062 120134
rect 407146 119898 407382 120134
rect 406826 84218 407062 84454
rect 407146 84218 407382 84454
rect 406826 83898 407062 84134
rect 407146 83898 407382 84134
rect 406826 48218 407062 48454
rect 407146 48218 407382 48454
rect 406826 47898 407062 48134
rect 407146 47898 407382 48134
rect 406826 12218 407062 12454
rect 407146 12218 407382 12454
rect 406826 11898 407062 12134
rect 407146 11898 407382 12134
rect 406826 -2502 407062 -2266
rect 407146 -2502 407382 -2266
rect 406826 -2822 407062 -2586
rect 407146 -2822 407382 -2586
rect 411326 707482 411562 707718
rect 411646 707482 411882 707718
rect 411326 707162 411562 707398
rect 411646 707162 411882 707398
rect 411326 700718 411562 700954
rect 411646 700718 411882 700954
rect 411326 700398 411562 700634
rect 411646 700398 411882 700634
rect 411326 664718 411562 664954
rect 411646 664718 411882 664954
rect 411326 664398 411562 664634
rect 411646 664398 411882 664634
rect 411326 628718 411562 628954
rect 411646 628718 411882 628954
rect 411326 628398 411562 628634
rect 411646 628398 411882 628634
rect 411326 592718 411562 592954
rect 411646 592718 411882 592954
rect 411326 592398 411562 592634
rect 411646 592398 411882 592634
rect 411326 556718 411562 556954
rect 411646 556718 411882 556954
rect 411326 556398 411562 556634
rect 411646 556398 411882 556634
rect 411326 520718 411562 520954
rect 411646 520718 411882 520954
rect 411326 520398 411562 520634
rect 411646 520398 411882 520634
rect 411326 484718 411562 484954
rect 411646 484718 411882 484954
rect 411326 484398 411562 484634
rect 411646 484398 411882 484634
rect 411326 448718 411562 448954
rect 411646 448718 411882 448954
rect 411326 448398 411562 448634
rect 411646 448398 411882 448634
rect 411326 412718 411562 412954
rect 411646 412718 411882 412954
rect 411326 412398 411562 412634
rect 411646 412398 411882 412634
rect 411326 376718 411562 376954
rect 411646 376718 411882 376954
rect 411326 376398 411562 376634
rect 411646 376398 411882 376634
rect 411326 340718 411562 340954
rect 411646 340718 411882 340954
rect 411326 340398 411562 340634
rect 411646 340398 411882 340634
rect 411326 304718 411562 304954
rect 411646 304718 411882 304954
rect 411326 304398 411562 304634
rect 411646 304398 411882 304634
rect 411326 268718 411562 268954
rect 411646 268718 411882 268954
rect 411326 268398 411562 268634
rect 411646 268398 411882 268634
rect 411326 232718 411562 232954
rect 411646 232718 411882 232954
rect 411326 232398 411562 232634
rect 411646 232398 411882 232634
rect 411326 196718 411562 196954
rect 411646 196718 411882 196954
rect 411326 196398 411562 196634
rect 411646 196398 411882 196634
rect 411326 160718 411562 160954
rect 411646 160718 411882 160954
rect 411326 160398 411562 160634
rect 411646 160398 411882 160634
rect 411326 124718 411562 124954
rect 411646 124718 411882 124954
rect 411326 124398 411562 124634
rect 411646 124398 411882 124634
rect 411326 88718 411562 88954
rect 411646 88718 411882 88954
rect 411326 88398 411562 88634
rect 411646 88398 411882 88634
rect 411326 52718 411562 52954
rect 411646 52718 411882 52954
rect 411326 52398 411562 52634
rect 411646 52398 411882 52634
rect 411326 16718 411562 16954
rect 411646 16718 411882 16954
rect 411326 16398 411562 16634
rect 411646 16398 411882 16634
rect 411326 -3462 411562 -3226
rect 411646 -3462 411882 -3226
rect 411326 -3782 411562 -3546
rect 411646 -3782 411882 -3546
rect 415826 708442 416062 708678
rect 416146 708442 416382 708678
rect 415826 708122 416062 708358
rect 416146 708122 416382 708358
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 415826 381218 416062 381454
rect 416146 381218 416382 381454
rect 415826 380898 416062 381134
rect 416146 380898 416382 381134
rect 415826 345218 416062 345454
rect 416146 345218 416382 345454
rect 415826 344898 416062 345134
rect 416146 344898 416382 345134
rect 415826 309218 416062 309454
rect 416146 309218 416382 309454
rect 415826 308898 416062 309134
rect 416146 308898 416382 309134
rect 415826 273218 416062 273454
rect 416146 273218 416382 273454
rect 415826 272898 416062 273134
rect 416146 272898 416382 273134
rect 415826 237218 416062 237454
rect 416146 237218 416382 237454
rect 415826 236898 416062 237134
rect 416146 236898 416382 237134
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -4422 416062 -4186
rect 416146 -4422 416382 -4186
rect 415826 -4742 416062 -4506
rect 416146 -4742 416382 -4506
rect 420326 709402 420562 709638
rect 420646 709402 420882 709638
rect 420326 709082 420562 709318
rect 420646 709082 420882 709318
rect 420326 673718 420562 673954
rect 420646 673718 420882 673954
rect 420326 673398 420562 673634
rect 420646 673398 420882 673634
rect 420326 637718 420562 637954
rect 420646 637718 420882 637954
rect 420326 637398 420562 637634
rect 420646 637398 420882 637634
rect 420326 601718 420562 601954
rect 420646 601718 420882 601954
rect 420326 601398 420562 601634
rect 420646 601398 420882 601634
rect 420326 565718 420562 565954
rect 420646 565718 420882 565954
rect 420326 565398 420562 565634
rect 420646 565398 420882 565634
rect 420326 529718 420562 529954
rect 420646 529718 420882 529954
rect 420326 529398 420562 529634
rect 420646 529398 420882 529634
rect 420326 493718 420562 493954
rect 420646 493718 420882 493954
rect 420326 493398 420562 493634
rect 420646 493398 420882 493634
rect 420326 457718 420562 457954
rect 420646 457718 420882 457954
rect 420326 457398 420562 457634
rect 420646 457398 420882 457634
rect 420326 421718 420562 421954
rect 420646 421718 420882 421954
rect 420326 421398 420562 421634
rect 420646 421398 420882 421634
rect 420326 385718 420562 385954
rect 420646 385718 420882 385954
rect 420326 385398 420562 385634
rect 420646 385398 420882 385634
rect 420326 349718 420562 349954
rect 420646 349718 420882 349954
rect 420326 349398 420562 349634
rect 420646 349398 420882 349634
rect 420326 313718 420562 313954
rect 420646 313718 420882 313954
rect 420326 313398 420562 313634
rect 420646 313398 420882 313634
rect 420326 277718 420562 277954
rect 420646 277718 420882 277954
rect 420326 277398 420562 277634
rect 420646 277398 420882 277634
rect 420326 241718 420562 241954
rect 420646 241718 420882 241954
rect 420326 241398 420562 241634
rect 420646 241398 420882 241634
rect 420326 205718 420562 205954
rect 420646 205718 420882 205954
rect 420326 205398 420562 205634
rect 420646 205398 420882 205634
rect 420326 169718 420562 169954
rect 420646 169718 420882 169954
rect 420326 169398 420562 169634
rect 420646 169398 420882 169634
rect 420326 133718 420562 133954
rect 420646 133718 420882 133954
rect 420326 133398 420562 133634
rect 420646 133398 420882 133634
rect 420326 97718 420562 97954
rect 420646 97718 420882 97954
rect 420326 97398 420562 97634
rect 420646 97398 420882 97634
rect 420326 61718 420562 61954
rect 420646 61718 420882 61954
rect 420326 61398 420562 61634
rect 420646 61398 420882 61634
rect 420326 25718 420562 25954
rect 420646 25718 420882 25954
rect 420326 25398 420562 25634
rect 420646 25398 420882 25634
rect 420326 -5382 420562 -5146
rect 420646 -5382 420882 -5146
rect 420326 -5702 420562 -5466
rect 420646 -5702 420882 -5466
rect 424826 710362 425062 710598
rect 425146 710362 425382 710598
rect 424826 710042 425062 710278
rect 425146 710042 425382 710278
rect 424826 678218 425062 678454
rect 425146 678218 425382 678454
rect 424826 677898 425062 678134
rect 425146 677898 425382 678134
rect 424826 642218 425062 642454
rect 425146 642218 425382 642454
rect 424826 641898 425062 642134
rect 425146 641898 425382 642134
rect 424826 606218 425062 606454
rect 425146 606218 425382 606454
rect 424826 605898 425062 606134
rect 425146 605898 425382 606134
rect 424826 570218 425062 570454
rect 425146 570218 425382 570454
rect 424826 569898 425062 570134
rect 425146 569898 425382 570134
rect 424826 534218 425062 534454
rect 425146 534218 425382 534454
rect 424826 533898 425062 534134
rect 425146 533898 425382 534134
rect 424826 498218 425062 498454
rect 425146 498218 425382 498454
rect 424826 497898 425062 498134
rect 425146 497898 425382 498134
rect 424826 462218 425062 462454
rect 425146 462218 425382 462454
rect 424826 461898 425062 462134
rect 425146 461898 425382 462134
rect 424826 426218 425062 426454
rect 425146 426218 425382 426454
rect 424826 425898 425062 426134
rect 425146 425898 425382 426134
rect 424826 390218 425062 390454
rect 425146 390218 425382 390454
rect 424826 389898 425062 390134
rect 425146 389898 425382 390134
rect 424826 354218 425062 354454
rect 425146 354218 425382 354454
rect 424826 353898 425062 354134
rect 425146 353898 425382 354134
rect 424826 318218 425062 318454
rect 425146 318218 425382 318454
rect 424826 317898 425062 318134
rect 425146 317898 425382 318134
rect 424826 282218 425062 282454
rect 425146 282218 425382 282454
rect 424826 281898 425062 282134
rect 425146 281898 425382 282134
rect 424826 246218 425062 246454
rect 425146 246218 425382 246454
rect 424826 245898 425062 246134
rect 425146 245898 425382 246134
rect 424826 210218 425062 210454
rect 425146 210218 425382 210454
rect 424826 209898 425062 210134
rect 425146 209898 425382 210134
rect 424826 174218 425062 174454
rect 425146 174218 425382 174454
rect 424826 173898 425062 174134
rect 425146 173898 425382 174134
rect 424826 138218 425062 138454
rect 425146 138218 425382 138454
rect 424826 137898 425062 138134
rect 425146 137898 425382 138134
rect 424826 102218 425062 102454
rect 425146 102218 425382 102454
rect 424826 101898 425062 102134
rect 425146 101898 425382 102134
rect 424826 66218 425062 66454
rect 425146 66218 425382 66454
rect 424826 65898 425062 66134
rect 425146 65898 425382 66134
rect 424826 30218 425062 30454
rect 425146 30218 425382 30454
rect 424826 29898 425062 30134
rect 425146 29898 425382 30134
rect 424826 -6342 425062 -6106
rect 425146 -6342 425382 -6106
rect 424826 -6662 425062 -6426
rect 425146 -6662 425382 -6426
rect 429326 711322 429562 711558
rect 429646 711322 429882 711558
rect 429326 711002 429562 711238
rect 429646 711002 429882 711238
rect 429326 682718 429562 682954
rect 429646 682718 429882 682954
rect 429326 682398 429562 682634
rect 429646 682398 429882 682634
rect 429326 646718 429562 646954
rect 429646 646718 429882 646954
rect 429326 646398 429562 646634
rect 429646 646398 429882 646634
rect 429326 610718 429562 610954
rect 429646 610718 429882 610954
rect 429326 610398 429562 610634
rect 429646 610398 429882 610634
rect 429326 574718 429562 574954
rect 429646 574718 429882 574954
rect 429326 574398 429562 574634
rect 429646 574398 429882 574634
rect 429326 538718 429562 538954
rect 429646 538718 429882 538954
rect 429326 538398 429562 538634
rect 429646 538398 429882 538634
rect 429326 502718 429562 502954
rect 429646 502718 429882 502954
rect 429326 502398 429562 502634
rect 429646 502398 429882 502634
rect 429326 466718 429562 466954
rect 429646 466718 429882 466954
rect 429326 466398 429562 466634
rect 429646 466398 429882 466634
rect 429326 430718 429562 430954
rect 429646 430718 429882 430954
rect 429326 430398 429562 430634
rect 429646 430398 429882 430634
rect 429326 394718 429562 394954
rect 429646 394718 429882 394954
rect 429326 394398 429562 394634
rect 429646 394398 429882 394634
rect 429326 358718 429562 358954
rect 429646 358718 429882 358954
rect 429326 358398 429562 358634
rect 429646 358398 429882 358634
rect 429326 322718 429562 322954
rect 429646 322718 429882 322954
rect 429326 322398 429562 322634
rect 429646 322398 429882 322634
rect 429326 286718 429562 286954
rect 429646 286718 429882 286954
rect 429326 286398 429562 286634
rect 429646 286398 429882 286634
rect 429326 250718 429562 250954
rect 429646 250718 429882 250954
rect 429326 250398 429562 250634
rect 429646 250398 429882 250634
rect 429326 214718 429562 214954
rect 429646 214718 429882 214954
rect 429326 214398 429562 214634
rect 429646 214398 429882 214634
rect 429326 178718 429562 178954
rect 429646 178718 429882 178954
rect 429326 178398 429562 178634
rect 429646 178398 429882 178634
rect 429326 142718 429562 142954
rect 429646 142718 429882 142954
rect 429326 142398 429562 142634
rect 429646 142398 429882 142634
rect 429326 106718 429562 106954
rect 429646 106718 429882 106954
rect 429326 106398 429562 106634
rect 429646 106398 429882 106634
rect 429326 70718 429562 70954
rect 429646 70718 429882 70954
rect 429326 70398 429562 70634
rect 429646 70398 429882 70634
rect 429326 34718 429562 34954
rect 429646 34718 429882 34954
rect 429326 34398 429562 34634
rect 429646 34398 429882 34634
rect 429326 -7302 429562 -7066
rect 429646 -7302 429882 -7066
rect 429326 -7622 429562 -7386
rect 429646 -7622 429882 -7386
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 438326 705562 438562 705798
rect 438646 705562 438882 705798
rect 438326 705242 438562 705478
rect 438646 705242 438882 705478
rect 438326 691718 438562 691954
rect 438646 691718 438882 691954
rect 438326 691398 438562 691634
rect 438646 691398 438882 691634
rect 438326 655718 438562 655954
rect 438646 655718 438882 655954
rect 438326 655398 438562 655634
rect 438646 655398 438882 655634
rect 438326 619718 438562 619954
rect 438646 619718 438882 619954
rect 438326 619398 438562 619634
rect 438646 619398 438882 619634
rect 438326 583718 438562 583954
rect 438646 583718 438882 583954
rect 438326 583398 438562 583634
rect 438646 583398 438882 583634
rect 438326 547718 438562 547954
rect 438646 547718 438882 547954
rect 438326 547398 438562 547634
rect 438646 547398 438882 547634
rect 438326 511718 438562 511954
rect 438646 511718 438882 511954
rect 438326 511398 438562 511634
rect 438646 511398 438882 511634
rect 438326 475718 438562 475954
rect 438646 475718 438882 475954
rect 438326 475398 438562 475634
rect 438646 475398 438882 475634
rect 438326 439718 438562 439954
rect 438646 439718 438882 439954
rect 438326 439398 438562 439634
rect 438646 439398 438882 439634
rect 438326 403718 438562 403954
rect 438646 403718 438882 403954
rect 438326 403398 438562 403634
rect 438646 403398 438882 403634
rect 438326 367718 438562 367954
rect 438646 367718 438882 367954
rect 438326 367398 438562 367634
rect 438646 367398 438882 367634
rect 438326 331718 438562 331954
rect 438646 331718 438882 331954
rect 438326 331398 438562 331634
rect 438646 331398 438882 331634
rect 438326 295718 438562 295954
rect 438646 295718 438882 295954
rect 438326 295398 438562 295634
rect 438646 295398 438882 295634
rect 438326 259718 438562 259954
rect 438646 259718 438882 259954
rect 438326 259398 438562 259634
rect 438646 259398 438882 259634
rect 438326 223718 438562 223954
rect 438646 223718 438882 223954
rect 438326 223398 438562 223634
rect 438646 223398 438882 223634
rect 438326 187718 438562 187954
rect 438646 187718 438882 187954
rect 438326 187398 438562 187634
rect 438646 187398 438882 187634
rect 438326 151718 438562 151954
rect 438646 151718 438882 151954
rect 438326 151398 438562 151634
rect 438646 151398 438882 151634
rect 438326 115718 438562 115954
rect 438646 115718 438882 115954
rect 438326 115398 438562 115634
rect 438646 115398 438882 115634
rect 438326 79718 438562 79954
rect 438646 79718 438882 79954
rect 438326 79398 438562 79634
rect 438646 79398 438882 79634
rect 438326 43718 438562 43954
rect 438646 43718 438882 43954
rect 438326 43398 438562 43634
rect 438646 43398 438882 43634
rect 438326 7718 438562 7954
rect 438646 7718 438882 7954
rect 438326 7398 438562 7634
rect 438646 7398 438882 7634
rect 438326 -1542 438562 -1306
rect 438646 -1542 438882 -1306
rect 438326 -1862 438562 -1626
rect 438646 -1862 438882 -1626
rect 442826 706522 443062 706758
rect 443146 706522 443382 706758
rect 442826 706202 443062 706438
rect 443146 706202 443382 706438
rect 442826 696218 443062 696454
rect 443146 696218 443382 696454
rect 442826 695898 443062 696134
rect 443146 695898 443382 696134
rect 442826 660218 443062 660454
rect 443146 660218 443382 660454
rect 442826 659898 443062 660134
rect 443146 659898 443382 660134
rect 442826 624218 443062 624454
rect 443146 624218 443382 624454
rect 442826 623898 443062 624134
rect 443146 623898 443382 624134
rect 442826 588218 443062 588454
rect 443146 588218 443382 588454
rect 442826 587898 443062 588134
rect 443146 587898 443382 588134
rect 442826 552218 443062 552454
rect 443146 552218 443382 552454
rect 442826 551898 443062 552134
rect 443146 551898 443382 552134
rect 442826 516218 443062 516454
rect 443146 516218 443382 516454
rect 442826 515898 443062 516134
rect 443146 515898 443382 516134
rect 442826 480218 443062 480454
rect 443146 480218 443382 480454
rect 442826 479898 443062 480134
rect 443146 479898 443382 480134
rect 442826 444218 443062 444454
rect 443146 444218 443382 444454
rect 442826 443898 443062 444134
rect 443146 443898 443382 444134
rect 442826 408218 443062 408454
rect 443146 408218 443382 408454
rect 442826 407898 443062 408134
rect 443146 407898 443382 408134
rect 442826 372218 443062 372454
rect 443146 372218 443382 372454
rect 442826 371898 443062 372134
rect 443146 371898 443382 372134
rect 442826 336218 443062 336454
rect 443146 336218 443382 336454
rect 442826 335898 443062 336134
rect 443146 335898 443382 336134
rect 442826 300218 443062 300454
rect 443146 300218 443382 300454
rect 442826 299898 443062 300134
rect 443146 299898 443382 300134
rect 442826 264218 443062 264454
rect 443146 264218 443382 264454
rect 442826 263898 443062 264134
rect 443146 263898 443382 264134
rect 442826 228218 443062 228454
rect 443146 228218 443382 228454
rect 442826 227898 443062 228134
rect 443146 227898 443382 228134
rect 442826 192218 443062 192454
rect 443146 192218 443382 192454
rect 442826 191898 443062 192134
rect 443146 191898 443382 192134
rect 442826 156218 443062 156454
rect 443146 156218 443382 156454
rect 442826 155898 443062 156134
rect 443146 155898 443382 156134
rect 442826 120218 443062 120454
rect 443146 120218 443382 120454
rect 442826 119898 443062 120134
rect 443146 119898 443382 120134
rect 442826 84218 443062 84454
rect 443146 84218 443382 84454
rect 442826 83898 443062 84134
rect 443146 83898 443382 84134
rect 442826 48218 443062 48454
rect 443146 48218 443382 48454
rect 442826 47898 443062 48134
rect 443146 47898 443382 48134
rect 442826 12218 443062 12454
rect 443146 12218 443382 12454
rect 442826 11898 443062 12134
rect 443146 11898 443382 12134
rect 442826 -2502 443062 -2266
rect 443146 -2502 443382 -2266
rect 442826 -2822 443062 -2586
rect 443146 -2822 443382 -2586
rect 447326 707482 447562 707718
rect 447646 707482 447882 707718
rect 447326 707162 447562 707398
rect 447646 707162 447882 707398
rect 447326 700718 447562 700954
rect 447646 700718 447882 700954
rect 447326 700398 447562 700634
rect 447646 700398 447882 700634
rect 447326 664718 447562 664954
rect 447646 664718 447882 664954
rect 447326 664398 447562 664634
rect 447646 664398 447882 664634
rect 447326 628718 447562 628954
rect 447646 628718 447882 628954
rect 447326 628398 447562 628634
rect 447646 628398 447882 628634
rect 447326 592718 447562 592954
rect 447646 592718 447882 592954
rect 447326 592398 447562 592634
rect 447646 592398 447882 592634
rect 447326 556718 447562 556954
rect 447646 556718 447882 556954
rect 447326 556398 447562 556634
rect 447646 556398 447882 556634
rect 447326 520718 447562 520954
rect 447646 520718 447882 520954
rect 447326 520398 447562 520634
rect 447646 520398 447882 520634
rect 447326 484718 447562 484954
rect 447646 484718 447882 484954
rect 447326 484398 447562 484634
rect 447646 484398 447882 484634
rect 447326 448718 447562 448954
rect 447646 448718 447882 448954
rect 447326 448398 447562 448634
rect 447646 448398 447882 448634
rect 447326 412718 447562 412954
rect 447646 412718 447882 412954
rect 447326 412398 447562 412634
rect 447646 412398 447882 412634
rect 447326 376718 447562 376954
rect 447646 376718 447882 376954
rect 447326 376398 447562 376634
rect 447646 376398 447882 376634
rect 447326 340718 447562 340954
rect 447646 340718 447882 340954
rect 447326 340398 447562 340634
rect 447646 340398 447882 340634
rect 447326 304718 447562 304954
rect 447646 304718 447882 304954
rect 447326 304398 447562 304634
rect 447646 304398 447882 304634
rect 447326 268718 447562 268954
rect 447646 268718 447882 268954
rect 447326 268398 447562 268634
rect 447646 268398 447882 268634
rect 447326 232718 447562 232954
rect 447646 232718 447882 232954
rect 447326 232398 447562 232634
rect 447646 232398 447882 232634
rect 447326 196718 447562 196954
rect 447646 196718 447882 196954
rect 447326 196398 447562 196634
rect 447646 196398 447882 196634
rect 447326 160718 447562 160954
rect 447646 160718 447882 160954
rect 447326 160398 447562 160634
rect 447646 160398 447882 160634
rect 447326 124718 447562 124954
rect 447646 124718 447882 124954
rect 447326 124398 447562 124634
rect 447646 124398 447882 124634
rect 447326 88718 447562 88954
rect 447646 88718 447882 88954
rect 447326 88398 447562 88634
rect 447646 88398 447882 88634
rect 447326 52718 447562 52954
rect 447646 52718 447882 52954
rect 447326 52398 447562 52634
rect 447646 52398 447882 52634
rect 447326 16718 447562 16954
rect 447646 16718 447882 16954
rect 447326 16398 447562 16634
rect 447646 16398 447882 16634
rect 447326 -3462 447562 -3226
rect 447646 -3462 447882 -3226
rect 447326 -3782 447562 -3546
rect 447646 -3782 447882 -3546
rect 451826 708442 452062 708678
rect 452146 708442 452382 708678
rect 451826 708122 452062 708358
rect 452146 708122 452382 708358
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 451826 309218 452062 309454
rect 452146 309218 452382 309454
rect 451826 308898 452062 309134
rect 452146 308898 452382 309134
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -4422 452062 -4186
rect 452146 -4422 452382 -4186
rect 451826 -4742 452062 -4506
rect 452146 -4742 452382 -4506
rect 456326 709402 456562 709638
rect 456646 709402 456882 709638
rect 456326 709082 456562 709318
rect 456646 709082 456882 709318
rect 456326 673718 456562 673954
rect 456646 673718 456882 673954
rect 456326 673398 456562 673634
rect 456646 673398 456882 673634
rect 456326 637718 456562 637954
rect 456646 637718 456882 637954
rect 456326 637398 456562 637634
rect 456646 637398 456882 637634
rect 456326 601718 456562 601954
rect 456646 601718 456882 601954
rect 456326 601398 456562 601634
rect 456646 601398 456882 601634
rect 456326 565718 456562 565954
rect 456646 565718 456882 565954
rect 456326 565398 456562 565634
rect 456646 565398 456882 565634
rect 456326 529718 456562 529954
rect 456646 529718 456882 529954
rect 456326 529398 456562 529634
rect 456646 529398 456882 529634
rect 456326 493718 456562 493954
rect 456646 493718 456882 493954
rect 456326 493398 456562 493634
rect 456646 493398 456882 493634
rect 456326 457718 456562 457954
rect 456646 457718 456882 457954
rect 456326 457398 456562 457634
rect 456646 457398 456882 457634
rect 456326 421718 456562 421954
rect 456646 421718 456882 421954
rect 456326 421398 456562 421634
rect 456646 421398 456882 421634
rect 456326 385718 456562 385954
rect 456646 385718 456882 385954
rect 456326 385398 456562 385634
rect 456646 385398 456882 385634
rect 456326 349718 456562 349954
rect 456646 349718 456882 349954
rect 456326 349398 456562 349634
rect 456646 349398 456882 349634
rect 456326 313718 456562 313954
rect 456646 313718 456882 313954
rect 456326 313398 456562 313634
rect 456646 313398 456882 313634
rect 456326 277718 456562 277954
rect 456646 277718 456882 277954
rect 456326 277398 456562 277634
rect 456646 277398 456882 277634
rect 456326 241718 456562 241954
rect 456646 241718 456882 241954
rect 456326 241398 456562 241634
rect 456646 241398 456882 241634
rect 456326 205718 456562 205954
rect 456646 205718 456882 205954
rect 456326 205398 456562 205634
rect 456646 205398 456882 205634
rect 456326 169718 456562 169954
rect 456646 169718 456882 169954
rect 456326 169398 456562 169634
rect 456646 169398 456882 169634
rect 456326 133718 456562 133954
rect 456646 133718 456882 133954
rect 456326 133398 456562 133634
rect 456646 133398 456882 133634
rect 456326 97718 456562 97954
rect 456646 97718 456882 97954
rect 456326 97398 456562 97634
rect 456646 97398 456882 97634
rect 456326 61718 456562 61954
rect 456646 61718 456882 61954
rect 456326 61398 456562 61634
rect 456646 61398 456882 61634
rect 456326 25718 456562 25954
rect 456646 25718 456882 25954
rect 456326 25398 456562 25634
rect 456646 25398 456882 25634
rect 456326 -5382 456562 -5146
rect 456646 -5382 456882 -5146
rect 456326 -5702 456562 -5466
rect 456646 -5702 456882 -5466
rect 460826 710362 461062 710598
rect 461146 710362 461382 710598
rect 460826 710042 461062 710278
rect 461146 710042 461382 710278
rect 460826 678218 461062 678454
rect 461146 678218 461382 678454
rect 460826 677898 461062 678134
rect 461146 677898 461382 678134
rect 460826 642218 461062 642454
rect 461146 642218 461382 642454
rect 460826 641898 461062 642134
rect 461146 641898 461382 642134
rect 460826 606218 461062 606454
rect 461146 606218 461382 606454
rect 460826 605898 461062 606134
rect 461146 605898 461382 606134
rect 460826 570218 461062 570454
rect 461146 570218 461382 570454
rect 460826 569898 461062 570134
rect 461146 569898 461382 570134
rect 460826 534218 461062 534454
rect 461146 534218 461382 534454
rect 460826 533898 461062 534134
rect 461146 533898 461382 534134
rect 460826 498218 461062 498454
rect 461146 498218 461382 498454
rect 460826 497898 461062 498134
rect 461146 497898 461382 498134
rect 460826 462218 461062 462454
rect 461146 462218 461382 462454
rect 460826 461898 461062 462134
rect 461146 461898 461382 462134
rect 460826 426218 461062 426454
rect 461146 426218 461382 426454
rect 460826 425898 461062 426134
rect 461146 425898 461382 426134
rect 460826 390218 461062 390454
rect 461146 390218 461382 390454
rect 460826 389898 461062 390134
rect 461146 389898 461382 390134
rect 460826 354218 461062 354454
rect 461146 354218 461382 354454
rect 460826 353898 461062 354134
rect 461146 353898 461382 354134
rect 460826 318218 461062 318454
rect 461146 318218 461382 318454
rect 460826 317898 461062 318134
rect 461146 317898 461382 318134
rect 460826 282218 461062 282454
rect 461146 282218 461382 282454
rect 460826 281898 461062 282134
rect 461146 281898 461382 282134
rect 460826 246218 461062 246454
rect 461146 246218 461382 246454
rect 460826 245898 461062 246134
rect 461146 245898 461382 246134
rect 460826 210218 461062 210454
rect 461146 210218 461382 210454
rect 460826 209898 461062 210134
rect 461146 209898 461382 210134
rect 460826 174218 461062 174454
rect 461146 174218 461382 174454
rect 460826 173898 461062 174134
rect 461146 173898 461382 174134
rect 460826 138218 461062 138454
rect 461146 138218 461382 138454
rect 460826 137898 461062 138134
rect 461146 137898 461382 138134
rect 460826 102218 461062 102454
rect 461146 102218 461382 102454
rect 460826 101898 461062 102134
rect 461146 101898 461382 102134
rect 460826 66218 461062 66454
rect 461146 66218 461382 66454
rect 460826 65898 461062 66134
rect 461146 65898 461382 66134
rect 460826 30218 461062 30454
rect 461146 30218 461382 30454
rect 460826 29898 461062 30134
rect 461146 29898 461382 30134
rect 460826 -6342 461062 -6106
rect 461146 -6342 461382 -6106
rect 460826 -6662 461062 -6426
rect 461146 -6662 461382 -6426
rect 465326 711322 465562 711558
rect 465646 711322 465882 711558
rect 465326 711002 465562 711238
rect 465646 711002 465882 711238
rect 465326 682718 465562 682954
rect 465646 682718 465882 682954
rect 465326 682398 465562 682634
rect 465646 682398 465882 682634
rect 465326 646718 465562 646954
rect 465646 646718 465882 646954
rect 465326 646398 465562 646634
rect 465646 646398 465882 646634
rect 465326 610718 465562 610954
rect 465646 610718 465882 610954
rect 465326 610398 465562 610634
rect 465646 610398 465882 610634
rect 465326 574718 465562 574954
rect 465646 574718 465882 574954
rect 465326 574398 465562 574634
rect 465646 574398 465882 574634
rect 465326 538718 465562 538954
rect 465646 538718 465882 538954
rect 465326 538398 465562 538634
rect 465646 538398 465882 538634
rect 465326 502718 465562 502954
rect 465646 502718 465882 502954
rect 465326 502398 465562 502634
rect 465646 502398 465882 502634
rect 465326 466718 465562 466954
rect 465646 466718 465882 466954
rect 465326 466398 465562 466634
rect 465646 466398 465882 466634
rect 465326 430718 465562 430954
rect 465646 430718 465882 430954
rect 465326 430398 465562 430634
rect 465646 430398 465882 430634
rect 465326 394718 465562 394954
rect 465646 394718 465882 394954
rect 465326 394398 465562 394634
rect 465646 394398 465882 394634
rect 465326 358718 465562 358954
rect 465646 358718 465882 358954
rect 465326 358398 465562 358634
rect 465646 358398 465882 358634
rect 465326 322718 465562 322954
rect 465646 322718 465882 322954
rect 465326 322398 465562 322634
rect 465646 322398 465882 322634
rect 465326 286718 465562 286954
rect 465646 286718 465882 286954
rect 465326 286398 465562 286634
rect 465646 286398 465882 286634
rect 465326 250718 465562 250954
rect 465646 250718 465882 250954
rect 465326 250398 465562 250634
rect 465646 250398 465882 250634
rect 465326 214718 465562 214954
rect 465646 214718 465882 214954
rect 465326 214398 465562 214634
rect 465646 214398 465882 214634
rect 465326 178718 465562 178954
rect 465646 178718 465882 178954
rect 465326 178398 465562 178634
rect 465646 178398 465882 178634
rect 465326 142718 465562 142954
rect 465646 142718 465882 142954
rect 465326 142398 465562 142634
rect 465646 142398 465882 142634
rect 465326 106718 465562 106954
rect 465646 106718 465882 106954
rect 465326 106398 465562 106634
rect 465646 106398 465882 106634
rect 465326 70718 465562 70954
rect 465646 70718 465882 70954
rect 465326 70398 465562 70634
rect 465646 70398 465882 70634
rect 465326 34718 465562 34954
rect 465646 34718 465882 34954
rect 465326 34398 465562 34634
rect 465646 34398 465882 34634
rect 465326 -7302 465562 -7066
rect 465646 -7302 465882 -7066
rect 465326 -7622 465562 -7386
rect 465646 -7622 465882 -7386
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 474326 705562 474562 705798
rect 474646 705562 474882 705798
rect 474326 705242 474562 705478
rect 474646 705242 474882 705478
rect 474326 691718 474562 691954
rect 474646 691718 474882 691954
rect 474326 691398 474562 691634
rect 474646 691398 474882 691634
rect 474326 655718 474562 655954
rect 474646 655718 474882 655954
rect 474326 655398 474562 655634
rect 474646 655398 474882 655634
rect 474326 619718 474562 619954
rect 474646 619718 474882 619954
rect 474326 619398 474562 619634
rect 474646 619398 474882 619634
rect 474326 583718 474562 583954
rect 474646 583718 474882 583954
rect 474326 583398 474562 583634
rect 474646 583398 474882 583634
rect 474326 547718 474562 547954
rect 474646 547718 474882 547954
rect 474326 547398 474562 547634
rect 474646 547398 474882 547634
rect 474326 511718 474562 511954
rect 474646 511718 474882 511954
rect 474326 511398 474562 511634
rect 474646 511398 474882 511634
rect 474326 475718 474562 475954
rect 474646 475718 474882 475954
rect 474326 475398 474562 475634
rect 474646 475398 474882 475634
rect 474326 439718 474562 439954
rect 474646 439718 474882 439954
rect 474326 439398 474562 439634
rect 474646 439398 474882 439634
rect 474326 403718 474562 403954
rect 474646 403718 474882 403954
rect 474326 403398 474562 403634
rect 474646 403398 474882 403634
rect 474326 367718 474562 367954
rect 474646 367718 474882 367954
rect 474326 367398 474562 367634
rect 474646 367398 474882 367634
rect 474326 331718 474562 331954
rect 474646 331718 474882 331954
rect 474326 331398 474562 331634
rect 474646 331398 474882 331634
rect 474326 295718 474562 295954
rect 474646 295718 474882 295954
rect 474326 295398 474562 295634
rect 474646 295398 474882 295634
rect 474326 259718 474562 259954
rect 474646 259718 474882 259954
rect 474326 259398 474562 259634
rect 474646 259398 474882 259634
rect 474326 223718 474562 223954
rect 474646 223718 474882 223954
rect 474326 223398 474562 223634
rect 474646 223398 474882 223634
rect 474326 187718 474562 187954
rect 474646 187718 474882 187954
rect 474326 187398 474562 187634
rect 474646 187398 474882 187634
rect 474326 151718 474562 151954
rect 474646 151718 474882 151954
rect 474326 151398 474562 151634
rect 474646 151398 474882 151634
rect 474326 115718 474562 115954
rect 474646 115718 474882 115954
rect 474326 115398 474562 115634
rect 474646 115398 474882 115634
rect 474326 79718 474562 79954
rect 474646 79718 474882 79954
rect 474326 79398 474562 79634
rect 474646 79398 474882 79634
rect 474326 43718 474562 43954
rect 474646 43718 474882 43954
rect 474326 43398 474562 43634
rect 474646 43398 474882 43634
rect 474326 7718 474562 7954
rect 474646 7718 474882 7954
rect 474326 7398 474562 7634
rect 474646 7398 474882 7634
rect 474326 -1542 474562 -1306
rect 474646 -1542 474882 -1306
rect 474326 -1862 474562 -1626
rect 474646 -1862 474882 -1626
rect 478826 706522 479062 706758
rect 479146 706522 479382 706758
rect 478826 706202 479062 706438
rect 479146 706202 479382 706438
rect 478826 696218 479062 696454
rect 479146 696218 479382 696454
rect 478826 695898 479062 696134
rect 479146 695898 479382 696134
rect 478826 660218 479062 660454
rect 479146 660218 479382 660454
rect 478826 659898 479062 660134
rect 479146 659898 479382 660134
rect 478826 624218 479062 624454
rect 479146 624218 479382 624454
rect 478826 623898 479062 624134
rect 479146 623898 479382 624134
rect 478826 588218 479062 588454
rect 479146 588218 479382 588454
rect 478826 587898 479062 588134
rect 479146 587898 479382 588134
rect 478826 552218 479062 552454
rect 479146 552218 479382 552454
rect 478826 551898 479062 552134
rect 479146 551898 479382 552134
rect 478826 516218 479062 516454
rect 479146 516218 479382 516454
rect 478826 515898 479062 516134
rect 479146 515898 479382 516134
rect 478826 480218 479062 480454
rect 479146 480218 479382 480454
rect 478826 479898 479062 480134
rect 479146 479898 479382 480134
rect 478826 444218 479062 444454
rect 479146 444218 479382 444454
rect 478826 443898 479062 444134
rect 479146 443898 479382 444134
rect 478826 408218 479062 408454
rect 479146 408218 479382 408454
rect 478826 407898 479062 408134
rect 479146 407898 479382 408134
rect 478826 372218 479062 372454
rect 479146 372218 479382 372454
rect 478826 371898 479062 372134
rect 479146 371898 479382 372134
rect 478826 336218 479062 336454
rect 479146 336218 479382 336454
rect 478826 335898 479062 336134
rect 479146 335898 479382 336134
rect 478826 300218 479062 300454
rect 479146 300218 479382 300454
rect 478826 299898 479062 300134
rect 479146 299898 479382 300134
rect 478826 264218 479062 264454
rect 479146 264218 479382 264454
rect 478826 263898 479062 264134
rect 479146 263898 479382 264134
rect 478826 228218 479062 228454
rect 479146 228218 479382 228454
rect 478826 227898 479062 228134
rect 479146 227898 479382 228134
rect 478826 192218 479062 192454
rect 479146 192218 479382 192454
rect 478826 191898 479062 192134
rect 479146 191898 479382 192134
rect 478826 156218 479062 156454
rect 479146 156218 479382 156454
rect 478826 155898 479062 156134
rect 479146 155898 479382 156134
rect 478826 120218 479062 120454
rect 479146 120218 479382 120454
rect 478826 119898 479062 120134
rect 479146 119898 479382 120134
rect 478826 84218 479062 84454
rect 479146 84218 479382 84454
rect 478826 83898 479062 84134
rect 479146 83898 479382 84134
rect 478826 48218 479062 48454
rect 479146 48218 479382 48454
rect 478826 47898 479062 48134
rect 479146 47898 479382 48134
rect 478826 12218 479062 12454
rect 479146 12218 479382 12454
rect 478826 11898 479062 12134
rect 479146 11898 479382 12134
rect 478826 -2502 479062 -2266
rect 479146 -2502 479382 -2266
rect 478826 -2822 479062 -2586
rect 479146 -2822 479382 -2586
rect 483326 707482 483562 707718
rect 483646 707482 483882 707718
rect 483326 707162 483562 707398
rect 483646 707162 483882 707398
rect 483326 700718 483562 700954
rect 483646 700718 483882 700954
rect 483326 700398 483562 700634
rect 483646 700398 483882 700634
rect 483326 664718 483562 664954
rect 483646 664718 483882 664954
rect 483326 664398 483562 664634
rect 483646 664398 483882 664634
rect 483326 628718 483562 628954
rect 483646 628718 483882 628954
rect 483326 628398 483562 628634
rect 483646 628398 483882 628634
rect 483326 592718 483562 592954
rect 483646 592718 483882 592954
rect 483326 592398 483562 592634
rect 483646 592398 483882 592634
rect 483326 556718 483562 556954
rect 483646 556718 483882 556954
rect 483326 556398 483562 556634
rect 483646 556398 483882 556634
rect 483326 520718 483562 520954
rect 483646 520718 483882 520954
rect 483326 520398 483562 520634
rect 483646 520398 483882 520634
rect 483326 484718 483562 484954
rect 483646 484718 483882 484954
rect 483326 484398 483562 484634
rect 483646 484398 483882 484634
rect 483326 448718 483562 448954
rect 483646 448718 483882 448954
rect 483326 448398 483562 448634
rect 483646 448398 483882 448634
rect 483326 412718 483562 412954
rect 483646 412718 483882 412954
rect 483326 412398 483562 412634
rect 483646 412398 483882 412634
rect 483326 376718 483562 376954
rect 483646 376718 483882 376954
rect 483326 376398 483562 376634
rect 483646 376398 483882 376634
rect 483326 340718 483562 340954
rect 483646 340718 483882 340954
rect 483326 340398 483562 340634
rect 483646 340398 483882 340634
rect 483326 304718 483562 304954
rect 483646 304718 483882 304954
rect 483326 304398 483562 304634
rect 483646 304398 483882 304634
rect 483326 268718 483562 268954
rect 483646 268718 483882 268954
rect 483326 268398 483562 268634
rect 483646 268398 483882 268634
rect 483326 232718 483562 232954
rect 483646 232718 483882 232954
rect 483326 232398 483562 232634
rect 483646 232398 483882 232634
rect 483326 196718 483562 196954
rect 483646 196718 483882 196954
rect 483326 196398 483562 196634
rect 483646 196398 483882 196634
rect 483326 160718 483562 160954
rect 483646 160718 483882 160954
rect 483326 160398 483562 160634
rect 483646 160398 483882 160634
rect 483326 124718 483562 124954
rect 483646 124718 483882 124954
rect 483326 124398 483562 124634
rect 483646 124398 483882 124634
rect 483326 88718 483562 88954
rect 483646 88718 483882 88954
rect 483326 88398 483562 88634
rect 483646 88398 483882 88634
rect 483326 52718 483562 52954
rect 483646 52718 483882 52954
rect 483326 52398 483562 52634
rect 483646 52398 483882 52634
rect 483326 16718 483562 16954
rect 483646 16718 483882 16954
rect 483326 16398 483562 16634
rect 483646 16398 483882 16634
rect 483326 -3462 483562 -3226
rect 483646 -3462 483882 -3226
rect 483326 -3782 483562 -3546
rect 483646 -3782 483882 -3546
rect 487826 708442 488062 708678
rect 488146 708442 488382 708678
rect 487826 708122 488062 708358
rect 488146 708122 488382 708358
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -4422 488062 -4186
rect 488146 -4422 488382 -4186
rect 487826 -4742 488062 -4506
rect 488146 -4742 488382 -4506
rect 492326 709402 492562 709638
rect 492646 709402 492882 709638
rect 492326 709082 492562 709318
rect 492646 709082 492882 709318
rect 492326 673718 492562 673954
rect 492646 673718 492882 673954
rect 492326 673398 492562 673634
rect 492646 673398 492882 673634
rect 492326 637718 492562 637954
rect 492646 637718 492882 637954
rect 492326 637398 492562 637634
rect 492646 637398 492882 637634
rect 492326 601718 492562 601954
rect 492646 601718 492882 601954
rect 492326 601398 492562 601634
rect 492646 601398 492882 601634
rect 492326 565718 492562 565954
rect 492646 565718 492882 565954
rect 492326 565398 492562 565634
rect 492646 565398 492882 565634
rect 492326 529718 492562 529954
rect 492646 529718 492882 529954
rect 492326 529398 492562 529634
rect 492646 529398 492882 529634
rect 492326 493718 492562 493954
rect 492646 493718 492882 493954
rect 492326 493398 492562 493634
rect 492646 493398 492882 493634
rect 492326 457718 492562 457954
rect 492646 457718 492882 457954
rect 492326 457398 492562 457634
rect 492646 457398 492882 457634
rect 492326 421718 492562 421954
rect 492646 421718 492882 421954
rect 492326 421398 492562 421634
rect 492646 421398 492882 421634
rect 492326 385718 492562 385954
rect 492646 385718 492882 385954
rect 492326 385398 492562 385634
rect 492646 385398 492882 385634
rect 492326 349718 492562 349954
rect 492646 349718 492882 349954
rect 492326 349398 492562 349634
rect 492646 349398 492882 349634
rect 492326 313718 492562 313954
rect 492646 313718 492882 313954
rect 492326 313398 492562 313634
rect 492646 313398 492882 313634
rect 492326 277718 492562 277954
rect 492646 277718 492882 277954
rect 492326 277398 492562 277634
rect 492646 277398 492882 277634
rect 492326 241718 492562 241954
rect 492646 241718 492882 241954
rect 492326 241398 492562 241634
rect 492646 241398 492882 241634
rect 492326 205718 492562 205954
rect 492646 205718 492882 205954
rect 492326 205398 492562 205634
rect 492646 205398 492882 205634
rect 492326 169718 492562 169954
rect 492646 169718 492882 169954
rect 492326 169398 492562 169634
rect 492646 169398 492882 169634
rect 492326 133718 492562 133954
rect 492646 133718 492882 133954
rect 492326 133398 492562 133634
rect 492646 133398 492882 133634
rect 492326 97718 492562 97954
rect 492646 97718 492882 97954
rect 492326 97398 492562 97634
rect 492646 97398 492882 97634
rect 492326 61718 492562 61954
rect 492646 61718 492882 61954
rect 492326 61398 492562 61634
rect 492646 61398 492882 61634
rect 492326 25718 492562 25954
rect 492646 25718 492882 25954
rect 492326 25398 492562 25634
rect 492646 25398 492882 25634
rect 492326 -5382 492562 -5146
rect 492646 -5382 492882 -5146
rect 492326 -5702 492562 -5466
rect 492646 -5702 492882 -5466
rect 496826 710362 497062 710598
rect 497146 710362 497382 710598
rect 496826 710042 497062 710278
rect 497146 710042 497382 710278
rect 496826 678218 497062 678454
rect 497146 678218 497382 678454
rect 496826 677898 497062 678134
rect 497146 677898 497382 678134
rect 496826 642218 497062 642454
rect 497146 642218 497382 642454
rect 496826 641898 497062 642134
rect 497146 641898 497382 642134
rect 496826 606218 497062 606454
rect 497146 606218 497382 606454
rect 496826 605898 497062 606134
rect 497146 605898 497382 606134
rect 496826 570218 497062 570454
rect 497146 570218 497382 570454
rect 496826 569898 497062 570134
rect 497146 569898 497382 570134
rect 496826 534218 497062 534454
rect 497146 534218 497382 534454
rect 496826 533898 497062 534134
rect 497146 533898 497382 534134
rect 496826 498218 497062 498454
rect 497146 498218 497382 498454
rect 496826 497898 497062 498134
rect 497146 497898 497382 498134
rect 496826 462218 497062 462454
rect 497146 462218 497382 462454
rect 496826 461898 497062 462134
rect 497146 461898 497382 462134
rect 496826 426218 497062 426454
rect 497146 426218 497382 426454
rect 496826 425898 497062 426134
rect 497146 425898 497382 426134
rect 496826 390218 497062 390454
rect 497146 390218 497382 390454
rect 496826 389898 497062 390134
rect 497146 389898 497382 390134
rect 496826 354218 497062 354454
rect 497146 354218 497382 354454
rect 496826 353898 497062 354134
rect 497146 353898 497382 354134
rect 496826 318218 497062 318454
rect 497146 318218 497382 318454
rect 496826 317898 497062 318134
rect 497146 317898 497382 318134
rect 496826 282218 497062 282454
rect 497146 282218 497382 282454
rect 496826 281898 497062 282134
rect 497146 281898 497382 282134
rect 496826 246218 497062 246454
rect 497146 246218 497382 246454
rect 496826 245898 497062 246134
rect 497146 245898 497382 246134
rect 496826 210218 497062 210454
rect 497146 210218 497382 210454
rect 496826 209898 497062 210134
rect 497146 209898 497382 210134
rect 496826 174218 497062 174454
rect 497146 174218 497382 174454
rect 496826 173898 497062 174134
rect 497146 173898 497382 174134
rect 496826 138218 497062 138454
rect 497146 138218 497382 138454
rect 496826 137898 497062 138134
rect 497146 137898 497382 138134
rect 496826 102218 497062 102454
rect 497146 102218 497382 102454
rect 496826 101898 497062 102134
rect 497146 101898 497382 102134
rect 496826 66218 497062 66454
rect 497146 66218 497382 66454
rect 496826 65898 497062 66134
rect 497146 65898 497382 66134
rect 496826 30218 497062 30454
rect 497146 30218 497382 30454
rect 496826 29898 497062 30134
rect 497146 29898 497382 30134
rect 496826 -6342 497062 -6106
rect 497146 -6342 497382 -6106
rect 496826 -6662 497062 -6426
rect 497146 -6662 497382 -6426
rect 501326 711322 501562 711558
rect 501646 711322 501882 711558
rect 501326 711002 501562 711238
rect 501646 711002 501882 711238
rect 501326 682718 501562 682954
rect 501646 682718 501882 682954
rect 501326 682398 501562 682634
rect 501646 682398 501882 682634
rect 501326 646718 501562 646954
rect 501646 646718 501882 646954
rect 501326 646398 501562 646634
rect 501646 646398 501882 646634
rect 501326 610718 501562 610954
rect 501646 610718 501882 610954
rect 501326 610398 501562 610634
rect 501646 610398 501882 610634
rect 501326 574718 501562 574954
rect 501646 574718 501882 574954
rect 501326 574398 501562 574634
rect 501646 574398 501882 574634
rect 501326 538718 501562 538954
rect 501646 538718 501882 538954
rect 501326 538398 501562 538634
rect 501646 538398 501882 538634
rect 501326 502718 501562 502954
rect 501646 502718 501882 502954
rect 501326 502398 501562 502634
rect 501646 502398 501882 502634
rect 501326 466718 501562 466954
rect 501646 466718 501882 466954
rect 501326 466398 501562 466634
rect 501646 466398 501882 466634
rect 501326 430718 501562 430954
rect 501646 430718 501882 430954
rect 501326 430398 501562 430634
rect 501646 430398 501882 430634
rect 501326 394718 501562 394954
rect 501646 394718 501882 394954
rect 501326 394398 501562 394634
rect 501646 394398 501882 394634
rect 501326 358718 501562 358954
rect 501646 358718 501882 358954
rect 501326 358398 501562 358634
rect 501646 358398 501882 358634
rect 501326 322718 501562 322954
rect 501646 322718 501882 322954
rect 501326 322398 501562 322634
rect 501646 322398 501882 322634
rect 501326 286718 501562 286954
rect 501646 286718 501882 286954
rect 501326 286398 501562 286634
rect 501646 286398 501882 286634
rect 501326 250718 501562 250954
rect 501646 250718 501882 250954
rect 501326 250398 501562 250634
rect 501646 250398 501882 250634
rect 501326 214718 501562 214954
rect 501646 214718 501882 214954
rect 501326 214398 501562 214634
rect 501646 214398 501882 214634
rect 501326 178718 501562 178954
rect 501646 178718 501882 178954
rect 501326 178398 501562 178634
rect 501646 178398 501882 178634
rect 501326 142718 501562 142954
rect 501646 142718 501882 142954
rect 501326 142398 501562 142634
rect 501646 142398 501882 142634
rect 501326 106718 501562 106954
rect 501646 106718 501882 106954
rect 501326 106398 501562 106634
rect 501646 106398 501882 106634
rect 501326 70718 501562 70954
rect 501646 70718 501882 70954
rect 501326 70398 501562 70634
rect 501646 70398 501882 70634
rect 501326 34718 501562 34954
rect 501646 34718 501882 34954
rect 501326 34398 501562 34634
rect 501646 34398 501882 34634
rect 501326 -7302 501562 -7066
rect 501646 -7302 501882 -7066
rect 501326 -7622 501562 -7386
rect 501646 -7622 501882 -7386
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 510326 705562 510562 705798
rect 510646 705562 510882 705798
rect 510326 705242 510562 705478
rect 510646 705242 510882 705478
rect 510326 691718 510562 691954
rect 510646 691718 510882 691954
rect 510326 691398 510562 691634
rect 510646 691398 510882 691634
rect 510326 655718 510562 655954
rect 510646 655718 510882 655954
rect 510326 655398 510562 655634
rect 510646 655398 510882 655634
rect 510326 619718 510562 619954
rect 510646 619718 510882 619954
rect 510326 619398 510562 619634
rect 510646 619398 510882 619634
rect 510326 583718 510562 583954
rect 510646 583718 510882 583954
rect 510326 583398 510562 583634
rect 510646 583398 510882 583634
rect 510326 547718 510562 547954
rect 510646 547718 510882 547954
rect 510326 547398 510562 547634
rect 510646 547398 510882 547634
rect 510326 511718 510562 511954
rect 510646 511718 510882 511954
rect 510326 511398 510562 511634
rect 510646 511398 510882 511634
rect 510326 475718 510562 475954
rect 510646 475718 510882 475954
rect 510326 475398 510562 475634
rect 510646 475398 510882 475634
rect 510326 439718 510562 439954
rect 510646 439718 510882 439954
rect 510326 439398 510562 439634
rect 510646 439398 510882 439634
rect 510326 403718 510562 403954
rect 510646 403718 510882 403954
rect 510326 403398 510562 403634
rect 510646 403398 510882 403634
rect 510326 367718 510562 367954
rect 510646 367718 510882 367954
rect 510326 367398 510562 367634
rect 510646 367398 510882 367634
rect 510326 331718 510562 331954
rect 510646 331718 510882 331954
rect 510326 331398 510562 331634
rect 510646 331398 510882 331634
rect 510326 295718 510562 295954
rect 510646 295718 510882 295954
rect 510326 295398 510562 295634
rect 510646 295398 510882 295634
rect 510326 259718 510562 259954
rect 510646 259718 510882 259954
rect 510326 259398 510562 259634
rect 510646 259398 510882 259634
rect 510326 223718 510562 223954
rect 510646 223718 510882 223954
rect 510326 223398 510562 223634
rect 510646 223398 510882 223634
rect 510326 187718 510562 187954
rect 510646 187718 510882 187954
rect 510326 187398 510562 187634
rect 510646 187398 510882 187634
rect 510326 151718 510562 151954
rect 510646 151718 510882 151954
rect 510326 151398 510562 151634
rect 510646 151398 510882 151634
rect 510326 115718 510562 115954
rect 510646 115718 510882 115954
rect 510326 115398 510562 115634
rect 510646 115398 510882 115634
rect 510326 79718 510562 79954
rect 510646 79718 510882 79954
rect 510326 79398 510562 79634
rect 510646 79398 510882 79634
rect 510326 43718 510562 43954
rect 510646 43718 510882 43954
rect 510326 43398 510562 43634
rect 510646 43398 510882 43634
rect 510326 7718 510562 7954
rect 510646 7718 510882 7954
rect 510326 7398 510562 7634
rect 510646 7398 510882 7634
rect 510326 -1542 510562 -1306
rect 510646 -1542 510882 -1306
rect 510326 -1862 510562 -1626
rect 510646 -1862 510882 -1626
rect 514826 706522 515062 706758
rect 515146 706522 515382 706758
rect 514826 706202 515062 706438
rect 515146 706202 515382 706438
rect 514826 696218 515062 696454
rect 515146 696218 515382 696454
rect 514826 695898 515062 696134
rect 515146 695898 515382 696134
rect 514826 660218 515062 660454
rect 515146 660218 515382 660454
rect 514826 659898 515062 660134
rect 515146 659898 515382 660134
rect 514826 624218 515062 624454
rect 515146 624218 515382 624454
rect 514826 623898 515062 624134
rect 515146 623898 515382 624134
rect 514826 588218 515062 588454
rect 515146 588218 515382 588454
rect 514826 587898 515062 588134
rect 515146 587898 515382 588134
rect 514826 552218 515062 552454
rect 515146 552218 515382 552454
rect 514826 551898 515062 552134
rect 515146 551898 515382 552134
rect 514826 516218 515062 516454
rect 515146 516218 515382 516454
rect 514826 515898 515062 516134
rect 515146 515898 515382 516134
rect 514826 480218 515062 480454
rect 515146 480218 515382 480454
rect 514826 479898 515062 480134
rect 515146 479898 515382 480134
rect 514826 444218 515062 444454
rect 515146 444218 515382 444454
rect 514826 443898 515062 444134
rect 515146 443898 515382 444134
rect 514826 408218 515062 408454
rect 515146 408218 515382 408454
rect 514826 407898 515062 408134
rect 515146 407898 515382 408134
rect 514826 372218 515062 372454
rect 515146 372218 515382 372454
rect 514826 371898 515062 372134
rect 515146 371898 515382 372134
rect 514826 336218 515062 336454
rect 515146 336218 515382 336454
rect 514826 335898 515062 336134
rect 515146 335898 515382 336134
rect 514826 300218 515062 300454
rect 515146 300218 515382 300454
rect 514826 299898 515062 300134
rect 515146 299898 515382 300134
rect 514826 264218 515062 264454
rect 515146 264218 515382 264454
rect 514826 263898 515062 264134
rect 515146 263898 515382 264134
rect 514826 228218 515062 228454
rect 515146 228218 515382 228454
rect 514826 227898 515062 228134
rect 515146 227898 515382 228134
rect 514826 192218 515062 192454
rect 515146 192218 515382 192454
rect 514826 191898 515062 192134
rect 515146 191898 515382 192134
rect 514826 156218 515062 156454
rect 515146 156218 515382 156454
rect 514826 155898 515062 156134
rect 515146 155898 515382 156134
rect 514826 120218 515062 120454
rect 515146 120218 515382 120454
rect 514826 119898 515062 120134
rect 515146 119898 515382 120134
rect 514826 84218 515062 84454
rect 515146 84218 515382 84454
rect 514826 83898 515062 84134
rect 515146 83898 515382 84134
rect 514826 48218 515062 48454
rect 515146 48218 515382 48454
rect 514826 47898 515062 48134
rect 515146 47898 515382 48134
rect 514826 12218 515062 12454
rect 515146 12218 515382 12454
rect 514826 11898 515062 12134
rect 515146 11898 515382 12134
rect 514826 -2502 515062 -2266
rect 515146 -2502 515382 -2266
rect 514826 -2822 515062 -2586
rect 515146 -2822 515382 -2586
rect 519326 707482 519562 707718
rect 519646 707482 519882 707718
rect 519326 707162 519562 707398
rect 519646 707162 519882 707398
rect 519326 700718 519562 700954
rect 519646 700718 519882 700954
rect 519326 700398 519562 700634
rect 519646 700398 519882 700634
rect 519326 664718 519562 664954
rect 519646 664718 519882 664954
rect 519326 664398 519562 664634
rect 519646 664398 519882 664634
rect 519326 628718 519562 628954
rect 519646 628718 519882 628954
rect 519326 628398 519562 628634
rect 519646 628398 519882 628634
rect 519326 592718 519562 592954
rect 519646 592718 519882 592954
rect 519326 592398 519562 592634
rect 519646 592398 519882 592634
rect 519326 556718 519562 556954
rect 519646 556718 519882 556954
rect 519326 556398 519562 556634
rect 519646 556398 519882 556634
rect 519326 520718 519562 520954
rect 519646 520718 519882 520954
rect 519326 520398 519562 520634
rect 519646 520398 519882 520634
rect 519326 484718 519562 484954
rect 519646 484718 519882 484954
rect 519326 484398 519562 484634
rect 519646 484398 519882 484634
rect 519326 448718 519562 448954
rect 519646 448718 519882 448954
rect 519326 448398 519562 448634
rect 519646 448398 519882 448634
rect 519326 412718 519562 412954
rect 519646 412718 519882 412954
rect 519326 412398 519562 412634
rect 519646 412398 519882 412634
rect 519326 376718 519562 376954
rect 519646 376718 519882 376954
rect 519326 376398 519562 376634
rect 519646 376398 519882 376634
rect 519326 340718 519562 340954
rect 519646 340718 519882 340954
rect 519326 340398 519562 340634
rect 519646 340398 519882 340634
rect 519326 304718 519562 304954
rect 519646 304718 519882 304954
rect 519326 304398 519562 304634
rect 519646 304398 519882 304634
rect 519326 268718 519562 268954
rect 519646 268718 519882 268954
rect 519326 268398 519562 268634
rect 519646 268398 519882 268634
rect 519326 232718 519562 232954
rect 519646 232718 519882 232954
rect 519326 232398 519562 232634
rect 519646 232398 519882 232634
rect 519326 196718 519562 196954
rect 519646 196718 519882 196954
rect 519326 196398 519562 196634
rect 519646 196398 519882 196634
rect 519326 160718 519562 160954
rect 519646 160718 519882 160954
rect 519326 160398 519562 160634
rect 519646 160398 519882 160634
rect 519326 124718 519562 124954
rect 519646 124718 519882 124954
rect 519326 124398 519562 124634
rect 519646 124398 519882 124634
rect 519326 88718 519562 88954
rect 519646 88718 519882 88954
rect 519326 88398 519562 88634
rect 519646 88398 519882 88634
rect 519326 52718 519562 52954
rect 519646 52718 519882 52954
rect 519326 52398 519562 52634
rect 519646 52398 519882 52634
rect 519326 16718 519562 16954
rect 519646 16718 519882 16954
rect 519326 16398 519562 16634
rect 519646 16398 519882 16634
rect 519326 -3462 519562 -3226
rect 519646 -3462 519882 -3226
rect 519326 -3782 519562 -3546
rect 519646 -3782 519882 -3546
rect 523826 708442 524062 708678
rect 524146 708442 524382 708678
rect 523826 708122 524062 708358
rect 524146 708122 524382 708358
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -4422 524062 -4186
rect 524146 -4422 524382 -4186
rect 523826 -4742 524062 -4506
rect 524146 -4742 524382 -4506
rect 528326 709402 528562 709638
rect 528646 709402 528882 709638
rect 528326 709082 528562 709318
rect 528646 709082 528882 709318
rect 528326 673718 528562 673954
rect 528646 673718 528882 673954
rect 528326 673398 528562 673634
rect 528646 673398 528882 673634
rect 528326 637718 528562 637954
rect 528646 637718 528882 637954
rect 528326 637398 528562 637634
rect 528646 637398 528882 637634
rect 528326 601718 528562 601954
rect 528646 601718 528882 601954
rect 528326 601398 528562 601634
rect 528646 601398 528882 601634
rect 528326 565718 528562 565954
rect 528646 565718 528882 565954
rect 528326 565398 528562 565634
rect 528646 565398 528882 565634
rect 528326 529718 528562 529954
rect 528646 529718 528882 529954
rect 528326 529398 528562 529634
rect 528646 529398 528882 529634
rect 528326 493718 528562 493954
rect 528646 493718 528882 493954
rect 528326 493398 528562 493634
rect 528646 493398 528882 493634
rect 528326 457718 528562 457954
rect 528646 457718 528882 457954
rect 528326 457398 528562 457634
rect 528646 457398 528882 457634
rect 528326 421718 528562 421954
rect 528646 421718 528882 421954
rect 528326 421398 528562 421634
rect 528646 421398 528882 421634
rect 528326 385718 528562 385954
rect 528646 385718 528882 385954
rect 528326 385398 528562 385634
rect 528646 385398 528882 385634
rect 528326 349718 528562 349954
rect 528646 349718 528882 349954
rect 528326 349398 528562 349634
rect 528646 349398 528882 349634
rect 528326 313718 528562 313954
rect 528646 313718 528882 313954
rect 528326 313398 528562 313634
rect 528646 313398 528882 313634
rect 528326 277718 528562 277954
rect 528646 277718 528882 277954
rect 528326 277398 528562 277634
rect 528646 277398 528882 277634
rect 528326 241718 528562 241954
rect 528646 241718 528882 241954
rect 528326 241398 528562 241634
rect 528646 241398 528882 241634
rect 528326 205718 528562 205954
rect 528646 205718 528882 205954
rect 528326 205398 528562 205634
rect 528646 205398 528882 205634
rect 528326 169718 528562 169954
rect 528646 169718 528882 169954
rect 528326 169398 528562 169634
rect 528646 169398 528882 169634
rect 528326 133718 528562 133954
rect 528646 133718 528882 133954
rect 528326 133398 528562 133634
rect 528646 133398 528882 133634
rect 528326 97718 528562 97954
rect 528646 97718 528882 97954
rect 528326 97398 528562 97634
rect 528646 97398 528882 97634
rect 528326 61718 528562 61954
rect 528646 61718 528882 61954
rect 528326 61398 528562 61634
rect 528646 61398 528882 61634
rect 528326 25718 528562 25954
rect 528646 25718 528882 25954
rect 528326 25398 528562 25634
rect 528646 25398 528882 25634
rect 528326 -5382 528562 -5146
rect 528646 -5382 528882 -5146
rect 528326 -5702 528562 -5466
rect 528646 -5702 528882 -5466
rect 532826 710362 533062 710598
rect 533146 710362 533382 710598
rect 532826 710042 533062 710278
rect 533146 710042 533382 710278
rect 532826 678218 533062 678454
rect 533146 678218 533382 678454
rect 532826 677898 533062 678134
rect 533146 677898 533382 678134
rect 532826 642218 533062 642454
rect 533146 642218 533382 642454
rect 532826 641898 533062 642134
rect 533146 641898 533382 642134
rect 532826 606218 533062 606454
rect 533146 606218 533382 606454
rect 532826 605898 533062 606134
rect 533146 605898 533382 606134
rect 532826 570218 533062 570454
rect 533146 570218 533382 570454
rect 532826 569898 533062 570134
rect 533146 569898 533382 570134
rect 532826 534218 533062 534454
rect 533146 534218 533382 534454
rect 532826 533898 533062 534134
rect 533146 533898 533382 534134
rect 532826 498218 533062 498454
rect 533146 498218 533382 498454
rect 532826 497898 533062 498134
rect 533146 497898 533382 498134
rect 532826 462218 533062 462454
rect 533146 462218 533382 462454
rect 532826 461898 533062 462134
rect 533146 461898 533382 462134
rect 532826 426218 533062 426454
rect 533146 426218 533382 426454
rect 532826 425898 533062 426134
rect 533146 425898 533382 426134
rect 532826 390218 533062 390454
rect 533146 390218 533382 390454
rect 532826 389898 533062 390134
rect 533146 389898 533382 390134
rect 532826 354218 533062 354454
rect 533146 354218 533382 354454
rect 532826 353898 533062 354134
rect 533146 353898 533382 354134
rect 532826 318218 533062 318454
rect 533146 318218 533382 318454
rect 532826 317898 533062 318134
rect 533146 317898 533382 318134
rect 532826 282218 533062 282454
rect 533146 282218 533382 282454
rect 532826 281898 533062 282134
rect 533146 281898 533382 282134
rect 532826 246218 533062 246454
rect 533146 246218 533382 246454
rect 532826 245898 533062 246134
rect 533146 245898 533382 246134
rect 532826 210218 533062 210454
rect 533146 210218 533382 210454
rect 532826 209898 533062 210134
rect 533146 209898 533382 210134
rect 532826 174218 533062 174454
rect 533146 174218 533382 174454
rect 532826 173898 533062 174134
rect 533146 173898 533382 174134
rect 532826 138218 533062 138454
rect 533146 138218 533382 138454
rect 532826 137898 533062 138134
rect 533146 137898 533382 138134
rect 532826 102218 533062 102454
rect 533146 102218 533382 102454
rect 532826 101898 533062 102134
rect 533146 101898 533382 102134
rect 532826 66218 533062 66454
rect 533146 66218 533382 66454
rect 532826 65898 533062 66134
rect 533146 65898 533382 66134
rect 532826 30218 533062 30454
rect 533146 30218 533382 30454
rect 532826 29898 533062 30134
rect 533146 29898 533382 30134
rect 532826 -6342 533062 -6106
rect 533146 -6342 533382 -6106
rect 532826 -6662 533062 -6426
rect 533146 -6662 533382 -6426
rect 537326 711322 537562 711558
rect 537646 711322 537882 711558
rect 537326 711002 537562 711238
rect 537646 711002 537882 711238
rect 537326 682718 537562 682954
rect 537646 682718 537882 682954
rect 537326 682398 537562 682634
rect 537646 682398 537882 682634
rect 537326 646718 537562 646954
rect 537646 646718 537882 646954
rect 537326 646398 537562 646634
rect 537646 646398 537882 646634
rect 537326 610718 537562 610954
rect 537646 610718 537882 610954
rect 537326 610398 537562 610634
rect 537646 610398 537882 610634
rect 537326 574718 537562 574954
rect 537646 574718 537882 574954
rect 537326 574398 537562 574634
rect 537646 574398 537882 574634
rect 537326 538718 537562 538954
rect 537646 538718 537882 538954
rect 537326 538398 537562 538634
rect 537646 538398 537882 538634
rect 537326 502718 537562 502954
rect 537646 502718 537882 502954
rect 537326 502398 537562 502634
rect 537646 502398 537882 502634
rect 537326 466718 537562 466954
rect 537646 466718 537882 466954
rect 537326 466398 537562 466634
rect 537646 466398 537882 466634
rect 537326 430718 537562 430954
rect 537646 430718 537882 430954
rect 537326 430398 537562 430634
rect 537646 430398 537882 430634
rect 537326 394718 537562 394954
rect 537646 394718 537882 394954
rect 537326 394398 537562 394634
rect 537646 394398 537882 394634
rect 537326 358718 537562 358954
rect 537646 358718 537882 358954
rect 537326 358398 537562 358634
rect 537646 358398 537882 358634
rect 537326 322718 537562 322954
rect 537646 322718 537882 322954
rect 537326 322398 537562 322634
rect 537646 322398 537882 322634
rect 537326 286718 537562 286954
rect 537646 286718 537882 286954
rect 537326 286398 537562 286634
rect 537646 286398 537882 286634
rect 537326 250718 537562 250954
rect 537646 250718 537882 250954
rect 537326 250398 537562 250634
rect 537646 250398 537882 250634
rect 537326 214718 537562 214954
rect 537646 214718 537882 214954
rect 537326 214398 537562 214634
rect 537646 214398 537882 214634
rect 537326 178718 537562 178954
rect 537646 178718 537882 178954
rect 537326 178398 537562 178634
rect 537646 178398 537882 178634
rect 537326 142718 537562 142954
rect 537646 142718 537882 142954
rect 537326 142398 537562 142634
rect 537646 142398 537882 142634
rect 537326 106718 537562 106954
rect 537646 106718 537882 106954
rect 537326 106398 537562 106634
rect 537646 106398 537882 106634
rect 537326 70718 537562 70954
rect 537646 70718 537882 70954
rect 537326 70398 537562 70634
rect 537646 70398 537882 70634
rect 537326 34718 537562 34954
rect 537646 34718 537882 34954
rect 537326 34398 537562 34634
rect 537646 34398 537882 34634
rect 537326 -7302 537562 -7066
rect 537646 -7302 537882 -7066
rect 537326 -7622 537562 -7386
rect 537646 -7622 537882 -7386
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 546326 705562 546562 705798
rect 546646 705562 546882 705798
rect 546326 705242 546562 705478
rect 546646 705242 546882 705478
rect 546326 691718 546562 691954
rect 546646 691718 546882 691954
rect 546326 691398 546562 691634
rect 546646 691398 546882 691634
rect 546326 655718 546562 655954
rect 546646 655718 546882 655954
rect 546326 655398 546562 655634
rect 546646 655398 546882 655634
rect 546326 619718 546562 619954
rect 546646 619718 546882 619954
rect 546326 619398 546562 619634
rect 546646 619398 546882 619634
rect 546326 583718 546562 583954
rect 546646 583718 546882 583954
rect 546326 583398 546562 583634
rect 546646 583398 546882 583634
rect 546326 547718 546562 547954
rect 546646 547718 546882 547954
rect 546326 547398 546562 547634
rect 546646 547398 546882 547634
rect 546326 511718 546562 511954
rect 546646 511718 546882 511954
rect 546326 511398 546562 511634
rect 546646 511398 546882 511634
rect 546326 475718 546562 475954
rect 546646 475718 546882 475954
rect 546326 475398 546562 475634
rect 546646 475398 546882 475634
rect 546326 439718 546562 439954
rect 546646 439718 546882 439954
rect 546326 439398 546562 439634
rect 546646 439398 546882 439634
rect 546326 403718 546562 403954
rect 546646 403718 546882 403954
rect 546326 403398 546562 403634
rect 546646 403398 546882 403634
rect 546326 367718 546562 367954
rect 546646 367718 546882 367954
rect 546326 367398 546562 367634
rect 546646 367398 546882 367634
rect 546326 331718 546562 331954
rect 546646 331718 546882 331954
rect 546326 331398 546562 331634
rect 546646 331398 546882 331634
rect 546326 295718 546562 295954
rect 546646 295718 546882 295954
rect 546326 295398 546562 295634
rect 546646 295398 546882 295634
rect 546326 259718 546562 259954
rect 546646 259718 546882 259954
rect 546326 259398 546562 259634
rect 546646 259398 546882 259634
rect 546326 223718 546562 223954
rect 546646 223718 546882 223954
rect 546326 223398 546562 223634
rect 546646 223398 546882 223634
rect 546326 187718 546562 187954
rect 546646 187718 546882 187954
rect 546326 187398 546562 187634
rect 546646 187398 546882 187634
rect 546326 151718 546562 151954
rect 546646 151718 546882 151954
rect 546326 151398 546562 151634
rect 546646 151398 546882 151634
rect 546326 115718 546562 115954
rect 546646 115718 546882 115954
rect 546326 115398 546562 115634
rect 546646 115398 546882 115634
rect 546326 79718 546562 79954
rect 546646 79718 546882 79954
rect 546326 79398 546562 79634
rect 546646 79398 546882 79634
rect 546326 43718 546562 43954
rect 546646 43718 546882 43954
rect 546326 43398 546562 43634
rect 546646 43398 546882 43634
rect 546326 7718 546562 7954
rect 546646 7718 546882 7954
rect 546326 7398 546562 7634
rect 546646 7398 546882 7634
rect 546326 -1542 546562 -1306
rect 546646 -1542 546882 -1306
rect 546326 -1862 546562 -1626
rect 546646 -1862 546882 -1626
rect 550826 706522 551062 706758
rect 551146 706522 551382 706758
rect 550826 706202 551062 706438
rect 551146 706202 551382 706438
rect 550826 696218 551062 696454
rect 551146 696218 551382 696454
rect 550826 695898 551062 696134
rect 551146 695898 551382 696134
rect 550826 660218 551062 660454
rect 551146 660218 551382 660454
rect 550826 659898 551062 660134
rect 551146 659898 551382 660134
rect 550826 624218 551062 624454
rect 551146 624218 551382 624454
rect 550826 623898 551062 624134
rect 551146 623898 551382 624134
rect 550826 588218 551062 588454
rect 551146 588218 551382 588454
rect 550826 587898 551062 588134
rect 551146 587898 551382 588134
rect 550826 552218 551062 552454
rect 551146 552218 551382 552454
rect 550826 551898 551062 552134
rect 551146 551898 551382 552134
rect 550826 516218 551062 516454
rect 551146 516218 551382 516454
rect 550826 515898 551062 516134
rect 551146 515898 551382 516134
rect 550826 480218 551062 480454
rect 551146 480218 551382 480454
rect 550826 479898 551062 480134
rect 551146 479898 551382 480134
rect 550826 444218 551062 444454
rect 551146 444218 551382 444454
rect 550826 443898 551062 444134
rect 551146 443898 551382 444134
rect 550826 408218 551062 408454
rect 551146 408218 551382 408454
rect 550826 407898 551062 408134
rect 551146 407898 551382 408134
rect 550826 372218 551062 372454
rect 551146 372218 551382 372454
rect 550826 371898 551062 372134
rect 551146 371898 551382 372134
rect 550826 336218 551062 336454
rect 551146 336218 551382 336454
rect 550826 335898 551062 336134
rect 551146 335898 551382 336134
rect 550826 300218 551062 300454
rect 551146 300218 551382 300454
rect 550826 299898 551062 300134
rect 551146 299898 551382 300134
rect 550826 264218 551062 264454
rect 551146 264218 551382 264454
rect 550826 263898 551062 264134
rect 551146 263898 551382 264134
rect 550826 228218 551062 228454
rect 551146 228218 551382 228454
rect 550826 227898 551062 228134
rect 551146 227898 551382 228134
rect 550826 192218 551062 192454
rect 551146 192218 551382 192454
rect 550826 191898 551062 192134
rect 551146 191898 551382 192134
rect 550826 156218 551062 156454
rect 551146 156218 551382 156454
rect 550826 155898 551062 156134
rect 551146 155898 551382 156134
rect 550826 120218 551062 120454
rect 551146 120218 551382 120454
rect 550826 119898 551062 120134
rect 551146 119898 551382 120134
rect 550826 84218 551062 84454
rect 551146 84218 551382 84454
rect 550826 83898 551062 84134
rect 551146 83898 551382 84134
rect 550826 48218 551062 48454
rect 551146 48218 551382 48454
rect 550826 47898 551062 48134
rect 551146 47898 551382 48134
rect 550826 12218 551062 12454
rect 551146 12218 551382 12454
rect 550826 11898 551062 12134
rect 551146 11898 551382 12134
rect 550826 -2502 551062 -2266
rect 551146 -2502 551382 -2266
rect 550826 -2822 551062 -2586
rect 551146 -2822 551382 -2586
rect 555326 707482 555562 707718
rect 555646 707482 555882 707718
rect 555326 707162 555562 707398
rect 555646 707162 555882 707398
rect 555326 700718 555562 700954
rect 555646 700718 555882 700954
rect 555326 700398 555562 700634
rect 555646 700398 555882 700634
rect 555326 664718 555562 664954
rect 555646 664718 555882 664954
rect 555326 664398 555562 664634
rect 555646 664398 555882 664634
rect 555326 628718 555562 628954
rect 555646 628718 555882 628954
rect 555326 628398 555562 628634
rect 555646 628398 555882 628634
rect 555326 592718 555562 592954
rect 555646 592718 555882 592954
rect 555326 592398 555562 592634
rect 555646 592398 555882 592634
rect 555326 556718 555562 556954
rect 555646 556718 555882 556954
rect 555326 556398 555562 556634
rect 555646 556398 555882 556634
rect 555326 520718 555562 520954
rect 555646 520718 555882 520954
rect 555326 520398 555562 520634
rect 555646 520398 555882 520634
rect 555326 484718 555562 484954
rect 555646 484718 555882 484954
rect 555326 484398 555562 484634
rect 555646 484398 555882 484634
rect 555326 448718 555562 448954
rect 555646 448718 555882 448954
rect 555326 448398 555562 448634
rect 555646 448398 555882 448634
rect 555326 412718 555562 412954
rect 555646 412718 555882 412954
rect 555326 412398 555562 412634
rect 555646 412398 555882 412634
rect 555326 376718 555562 376954
rect 555646 376718 555882 376954
rect 555326 376398 555562 376634
rect 555646 376398 555882 376634
rect 555326 340718 555562 340954
rect 555646 340718 555882 340954
rect 555326 340398 555562 340634
rect 555646 340398 555882 340634
rect 555326 304718 555562 304954
rect 555646 304718 555882 304954
rect 555326 304398 555562 304634
rect 555646 304398 555882 304634
rect 555326 268718 555562 268954
rect 555646 268718 555882 268954
rect 555326 268398 555562 268634
rect 555646 268398 555882 268634
rect 555326 232718 555562 232954
rect 555646 232718 555882 232954
rect 555326 232398 555562 232634
rect 555646 232398 555882 232634
rect 555326 196718 555562 196954
rect 555646 196718 555882 196954
rect 555326 196398 555562 196634
rect 555646 196398 555882 196634
rect 555326 160718 555562 160954
rect 555646 160718 555882 160954
rect 555326 160398 555562 160634
rect 555646 160398 555882 160634
rect 555326 124718 555562 124954
rect 555646 124718 555882 124954
rect 555326 124398 555562 124634
rect 555646 124398 555882 124634
rect 555326 88718 555562 88954
rect 555646 88718 555882 88954
rect 555326 88398 555562 88634
rect 555646 88398 555882 88634
rect 555326 52718 555562 52954
rect 555646 52718 555882 52954
rect 555326 52398 555562 52634
rect 555646 52398 555882 52634
rect 555326 16718 555562 16954
rect 555646 16718 555882 16954
rect 555326 16398 555562 16634
rect 555646 16398 555882 16634
rect 555326 -3462 555562 -3226
rect 555646 -3462 555882 -3226
rect 555326 -3782 555562 -3546
rect 555646 -3782 555882 -3546
rect 559826 708442 560062 708678
rect 560146 708442 560382 708678
rect 559826 708122 560062 708358
rect 560146 708122 560382 708358
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -4422 560062 -4186
rect 560146 -4422 560382 -4186
rect 559826 -4742 560062 -4506
rect 560146 -4742 560382 -4506
rect 564326 709402 564562 709638
rect 564646 709402 564882 709638
rect 564326 709082 564562 709318
rect 564646 709082 564882 709318
rect 564326 673718 564562 673954
rect 564646 673718 564882 673954
rect 564326 673398 564562 673634
rect 564646 673398 564882 673634
rect 564326 637718 564562 637954
rect 564646 637718 564882 637954
rect 564326 637398 564562 637634
rect 564646 637398 564882 637634
rect 564326 601718 564562 601954
rect 564646 601718 564882 601954
rect 564326 601398 564562 601634
rect 564646 601398 564882 601634
rect 564326 565718 564562 565954
rect 564646 565718 564882 565954
rect 564326 565398 564562 565634
rect 564646 565398 564882 565634
rect 564326 529718 564562 529954
rect 564646 529718 564882 529954
rect 564326 529398 564562 529634
rect 564646 529398 564882 529634
rect 564326 493718 564562 493954
rect 564646 493718 564882 493954
rect 564326 493398 564562 493634
rect 564646 493398 564882 493634
rect 564326 457718 564562 457954
rect 564646 457718 564882 457954
rect 564326 457398 564562 457634
rect 564646 457398 564882 457634
rect 564326 421718 564562 421954
rect 564646 421718 564882 421954
rect 564326 421398 564562 421634
rect 564646 421398 564882 421634
rect 564326 385718 564562 385954
rect 564646 385718 564882 385954
rect 564326 385398 564562 385634
rect 564646 385398 564882 385634
rect 564326 349718 564562 349954
rect 564646 349718 564882 349954
rect 564326 349398 564562 349634
rect 564646 349398 564882 349634
rect 564326 313718 564562 313954
rect 564646 313718 564882 313954
rect 564326 313398 564562 313634
rect 564646 313398 564882 313634
rect 564326 277718 564562 277954
rect 564646 277718 564882 277954
rect 564326 277398 564562 277634
rect 564646 277398 564882 277634
rect 564326 241718 564562 241954
rect 564646 241718 564882 241954
rect 564326 241398 564562 241634
rect 564646 241398 564882 241634
rect 564326 205718 564562 205954
rect 564646 205718 564882 205954
rect 564326 205398 564562 205634
rect 564646 205398 564882 205634
rect 564326 169718 564562 169954
rect 564646 169718 564882 169954
rect 564326 169398 564562 169634
rect 564646 169398 564882 169634
rect 564326 133718 564562 133954
rect 564646 133718 564882 133954
rect 564326 133398 564562 133634
rect 564646 133398 564882 133634
rect 564326 97718 564562 97954
rect 564646 97718 564882 97954
rect 564326 97398 564562 97634
rect 564646 97398 564882 97634
rect 564326 61718 564562 61954
rect 564646 61718 564882 61954
rect 564326 61398 564562 61634
rect 564646 61398 564882 61634
rect 564326 25718 564562 25954
rect 564646 25718 564882 25954
rect 564326 25398 564562 25634
rect 564646 25398 564882 25634
rect 564326 -5382 564562 -5146
rect 564646 -5382 564882 -5146
rect 564326 -5702 564562 -5466
rect 564646 -5702 564882 -5466
rect 568826 710362 569062 710598
rect 569146 710362 569382 710598
rect 568826 710042 569062 710278
rect 569146 710042 569382 710278
rect 568826 678218 569062 678454
rect 569146 678218 569382 678454
rect 568826 677898 569062 678134
rect 569146 677898 569382 678134
rect 568826 642218 569062 642454
rect 569146 642218 569382 642454
rect 568826 641898 569062 642134
rect 569146 641898 569382 642134
rect 568826 606218 569062 606454
rect 569146 606218 569382 606454
rect 568826 605898 569062 606134
rect 569146 605898 569382 606134
rect 568826 570218 569062 570454
rect 569146 570218 569382 570454
rect 568826 569898 569062 570134
rect 569146 569898 569382 570134
rect 568826 534218 569062 534454
rect 569146 534218 569382 534454
rect 568826 533898 569062 534134
rect 569146 533898 569382 534134
rect 568826 498218 569062 498454
rect 569146 498218 569382 498454
rect 568826 497898 569062 498134
rect 569146 497898 569382 498134
rect 568826 462218 569062 462454
rect 569146 462218 569382 462454
rect 568826 461898 569062 462134
rect 569146 461898 569382 462134
rect 568826 426218 569062 426454
rect 569146 426218 569382 426454
rect 568826 425898 569062 426134
rect 569146 425898 569382 426134
rect 568826 390218 569062 390454
rect 569146 390218 569382 390454
rect 568826 389898 569062 390134
rect 569146 389898 569382 390134
rect 568826 354218 569062 354454
rect 569146 354218 569382 354454
rect 568826 353898 569062 354134
rect 569146 353898 569382 354134
rect 568826 318218 569062 318454
rect 569146 318218 569382 318454
rect 568826 317898 569062 318134
rect 569146 317898 569382 318134
rect 568826 282218 569062 282454
rect 569146 282218 569382 282454
rect 568826 281898 569062 282134
rect 569146 281898 569382 282134
rect 568826 246218 569062 246454
rect 569146 246218 569382 246454
rect 568826 245898 569062 246134
rect 569146 245898 569382 246134
rect 568826 210218 569062 210454
rect 569146 210218 569382 210454
rect 568826 209898 569062 210134
rect 569146 209898 569382 210134
rect 568826 174218 569062 174454
rect 569146 174218 569382 174454
rect 568826 173898 569062 174134
rect 569146 173898 569382 174134
rect 568826 138218 569062 138454
rect 569146 138218 569382 138454
rect 568826 137898 569062 138134
rect 569146 137898 569382 138134
rect 568826 102218 569062 102454
rect 569146 102218 569382 102454
rect 568826 101898 569062 102134
rect 569146 101898 569382 102134
rect 568826 66218 569062 66454
rect 569146 66218 569382 66454
rect 568826 65898 569062 66134
rect 569146 65898 569382 66134
rect 568826 30218 569062 30454
rect 569146 30218 569382 30454
rect 568826 29898 569062 30134
rect 569146 29898 569382 30134
rect 568826 -6342 569062 -6106
rect 569146 -6342 569382 -6106
rect 568826 -6662 569062 -6426
rect 569146 -6662 569382 -6426
rect 573326 711322 573562 711558
rect 573646 711322 573882 711558
rect 573326 711002 573562 711238
rect 573646 711002 573882 711238
rect 573326 682718 573562 682954
rect 573646 682718 573882 682954
rect 573326 682398 573562 682634
rect 573646 682398 573882 682634
rect 573326 646718 573562 646954
rect 573646 646718 573882 646954
rect 573326 646398 573562 646634
rect 573646 646398 573882 646634
rect 573326 610718 573562 610954
rect 573646 610718 573882 610954
rect 573326 610398 573562 610634
rect 573646 610398 573882 610634
rect 573326 574718 573562 574954
rect 573646 574718 573882 574954
rect 573326 574398 573562 574634
rect 573646 574398 573882 574634
rect 573326 538718 573562 538954
rect 573646 538718 573882 538954
rect 573326 538398 573562 538634
rect 573646 538398 573882 538634
rect 573326 502718 573562 502954
rect 573646 502718 573882 502954
rect 573326 502398 573562 502634
rect 573646 502398 573882 502634
rect 573326 466718 573562 466954
rect 573646 466718 573882 466954
rect 573326 466398 573562 466634
rect 573646 466398 573882 466634
rect 573326 430718 573562 430954
rect 573646 430718 573882 430954
rect 573326 430398 573562 430634
rect 573646 430398 573882 430634
rect 573326 394718 573562 394954
rect 573646 394718 573882 394954
rect 573326 394398 573562 394634
rect 573646 394398 573882 394634
rect 573326 358718 573562 358954
rect 573646 358718 573882 358954
rect 573326 358398 573562 358634
rect 573646 358398 573882 358634
rect 573326 322718 573562 322954
rect 573646 322718 573882 322954
rect 573326 322398 573562 322634
rect 573646 322398 573882 322634
rect 573326 286718 573562 286954
rect 573646 286718 573882 286954
rect 573326 286398 573562 286634
rect 573646 286398 573882 286634
rect 573326 250718 573562 250954
rect 573646 250718 573882 250954
rect 573326 250398 573562 250634
rect 573646 250398 573882 250634
rect 573326 214718 573562 214954
rect 573646 214718 573882 214954
rect 573326 214398 573562 214634
rect 573646 214398 573882 214634
rect 573326 178718 573562 178954
rect 573646 178718 573882 178954
rect 573326 178398 573562 178634
rect 573646 178398 573882 178634
rect 573326 142718 573562 142954
rect 573646 142718 573882 142954
rect 573326 142398 573562 142634
rect 573646 142398 573882 142634
rect 573326 106718 573562 106954
rect 573646 106718 573882 106954
rect 573326 106398 573562 106634
rect 573646 106398 573882 106634
rect 573326 70718 573562 70954
rect 573646 70718 573882 70954
rect 573326 70398 573562 70634
rect 573646 70398 573882 70634
rect 573326 34718 573562 34954
rect 573646 34718 573882 34954
rect 573326 34398 573562 34634
rect 573646 34398 573882 34634
rect 573326 -7302 573562 -7066
rect 573646 -7302 573882 -7066
rect 573326 -7622 573562 -7386
rect 573646 -7622 573882 -7386
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 582326 705562 582562 705798
rect 582646 705562 582882 705798
rect 582326 705242 582562 705478
rect 582646 705242 582882 705478
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 582326 691718 582562 691954
rect 582646 691718 582882 691954
rect 582326 691398 582562 691634
rect 582646 691398 582882 691634
rect 582326 655718 582562 655954
rect 582646 655718 582882 655954
rect 582326 655398 582562 655634
rect 582646 655398 582882 655634
rect 582326 619718 582562 619954
rect 582646 619718 582882 619954
rect 582326 619398 582562 619634
rect 582646 619398 582882 619634
rect 582326 583718 582562 583954
rect 582646 583718 582882 583954
rect 582326 583398 582562 583634
rect 582646 583398 582882 583634
rect 582326 547718 582562 547954
rect 582646 547718 582882 547954
rect 582326 547398 582562 547634
rect 582646 547398 582882 547634
rect 582326 511718 582562 511954
rect 582646 511718 582882 511954
rect 582326 511398 582562 511634
rect 582646 511398 582882 511634
rect 582326 475718 582562 475954
rect 582646 475718 582882 475954
rect 582326 475398 582562 475634
rect 582646 475398 582882 475634
rect 582326 439718 582562 439954
rect 582646 439718 582882 439954
rect 582326 439398 582562 439634
rect 582646 439398 582882 439634
rect 582326 403718 582562 403954
rect 582646 403718 582882 403954
rect 582326 403398 582562 403634
rect 582646 403398 582882 403634
rect 582326 367718 582562 367954
rect 582646 367718 582882 367954
rect 582326 367398 582562 367634
rect 582646 367398 582882 367634
rect 582326 331718 582562 331954
rect 582646 331718 582882 331954
rect 582326 331398 582562 331634
rect 582646 331398 582882 331634
rect 582326 295718 582562 295954
rect 582646 295718 582882 295954
rect 582326 295398 582562 295634
rect 582646 295398 582882 295634
rect 582326 259718 582562 259954
rect 582646 259718 582882 259954
rect 582326 259398 582562 259634
rect 582646 259398 582882 259634
rect 582326 223718 582562 223954
rect 582646 223718 582882 223954
rect 582326 223398 582562 223634
rect 582646 223398 582882 223634
rect 582326 187718 582562 187954
rect 582646 187718 582882 187954
rect 582326 187398 582562 187634
rect 582646 187398 582882 187634
rect 582326 151718 582562 151954
rect 582646 151718 582882 151954
rect 582326 151398 582562 151634
rect 582646 151398 582882 151634
rect 582326 115718 582562 115954
rect 582646 115718 582882 115954
rect 582326 115398 582562 115634
rect 582646 115398 582882 115634
rect 582326 79718 582562 79954
rect 582646 79718 582882 79954
rect 582326 79398 582562 79634
rect 582646 79398 582882 79634
rect 582326 43718 582562 43954
rect 582646 43718 582882 43954
rect 582326 43398 582562 43634
rect 582646 43398 582882 43634
rect 582326 7718 582562 7954
rect 582646 7718 582882 7954
rect 582326 7398 582562 7634
rect 582646 7398 582882 7634
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 691718 586538 691954
rect 586622 691718 586858 691954
rect 586302 691398 586538 691634
rect 586622 691398 586858 691634
rect 586302 655718 586538 655954
rect 586622 655718 586858 655954
rect 586302 655398 586538 655634
rect 586622 655398 586858 655634
rect 586302 619718 586538 619954
rect 586622 619718 586858 619954
rect 586302 619398 586538 619634
rect 586622 619398 586858 619634
rect 586302 583718 586538 583954
rect 586622 583718 586858 583954
rect 586302 583398 586538 583634
rect 586622 583398 586858 583634
rect 586302 547718 586538 547954
rect 586622 547718 586858 547954
rect 586302 547398 586538 547634
rect 586622 547398 586858 547634
rect 586302 511718 586538 511954
rect 586622 511718 586858 511954
rect 586302 511398 586538 511634
rect 586622 511398 586858 511634
rect 586302 475718 586538 475954
rect 586622 475718 586858 475954
rect 586302 475398 586538 475634
rect 586622 475398 586858 475634
rect 586302 439718 586538 439954
rect 586622 439718 586858 439954
rect 586302 439398 586538 439634
rect 586622 439398 586858 439634
rect 586302 403718 586538 403954
rect 586622 403718 586858 403954
rect 586302 403398 586538 403634
rect 586622 403398 586858 403634
rect 586302 367718 586538 367954
rect 586622 367718 586858 367954
rect 586302 367398 586538 367634
rect 586622 367398 586858 367634
rect 586302 331718 586538 331954
rect 586622 331718 586858 331954
rect 586302 331398 586538 331634
rect 586622 331398 586858 331634
rect 586302 295718 586538 295954
rect 586622 295718 586858 295954
rect 586302 295398 586538 295634
rect 586622 295398 586858 295634
rect 586302 259718 586538 259954
rect 586622 259718 586858 259954
rect 586302 259398 586538 259634
rect 586622 259398 586858 259634
rect 586302 223718 586538 223954
rect 586622 223718 586858 223954
rect 586302 223398 586538 223634
rect 586622 223398 586858 223634
rect 586302 187718 586538 187954
rect 586622 187718 586858 187954
rect 586302 187398 586538 187634
rect 586622 187398 586858 187634
rect 586302 151718 586538 151954
rect 586622 151718 586858 151954
rect 586302 151398 586538 151634
rect 586622 151398 586858 151634
rect 586302 115718 586538 115954
rect 586622 115718 586858 115954
rect 586302 115398 586538 115634
rect 586622 115398 586858 115634
rect 586302 79718 586538 79954
rect 586622 79718 586858 79954
rect 586302 79398 586538 79634
rect 586622 79398 586858 79634
rect 586302 43718 586538 43954
rect 586622 43718 586858 43954
rect 586302 43398 586538 43634
rect 586622 43398 586858 43634
rect 586302 7718 586538 7954
rect 586622 7718 586858 7954
rect 586302 7398 586538 7634
rect 586622 7398 586858 7634
rect 582326 -1542 582562 -1306
rect 582646 -1542 582882 -1306
rect 582326 -1862 582562 -1626
rect 582646 -1862 582882 -1626
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 696218 587498 696454
rect 587582 696218 587818 696454
rect 587262 695898 587498 696134
rect 587582 695898 587818 696134
rect 587262 660218 587498 660454
rect 587582 660218 587818 660454
rect 587262 659898 587498 660134
rect 587582 659898 587818 660134
rect 587262 624218 587498 624454
rect 587582 624218 587818 624454
rect 587262 623898 587498 624134
rect 587582 623898 587818 624134
rect 587262 588218 587498 588454
rect 587582 588218 587818 588454
rect 587262 587898 587498 588134
rect 587582 587898 587818 588134
rect 587262 552218 587498 552454
rect 587582 552218 587818 552454
rect 587262 551898 587498 552134
rect 587582 551898 587818 552134
rect 587262 516218 587498 516454
rect 587582 516218 587818 516454
rect 587262 515898 587498 516134
rect 587582 515898 587818 516134
rect 587262 480218 587498 480454
rect 587582 480218 587818 480454
rect 587262 479898 587498 480134
rect 587582 479898 587818 480134
rect 587262 444218 587498 444454
rect 587582 444218 587818 444454
rect 587262 443898 587498 444134
rect 587582 443898 587818 444134
rect 587262 408218 587498 408454
rect 587582 408218 587818 408454
rect 587262 407898 587498 408134
rect 587582 407898 587818 408134
rect 587262 372218 587498 372454
rect 587582 372218 587818 372454
rect 587262 371898 587498 372134
rect 587582 371898 587818 372134
rect 587262 336218 587498 336454
rect 587582 336218 587818 336454
rect 587262 335898 587498 336134
rect 587582 335898 587818 336134
rect 587262 300218 587498 300454
rect 587582 300218 587818 300454
rect 587262 299898 587498 300134
rect 587582 299898 587818 300134
rect 587262 264218 587498 264454
rect 587582 264218 587818 264454
rect 587262 263898 587498 264134
rect 587582 263898 587818 264134
rect 587262 228218 587498 228454
rect 587582 228218 587818 228454
rect 587262 227898 587498 228134
rect 587582 227898 587818 228134
rect 587262 192218 587498 192454
rect 587582 192218 587818 192454
rect 587262 191898 587498 192134
rect 587582 191898 587818 192134
rect 587262 156218 587498 156454
rect 587582 156218 587818 156454
rect 587262 155898 587498 156134
rect 587582 155898 587818 156134
rect 587262 120218 587498 120454
rect 587582 120218 587818 120454
rect 587262 119898 587498 120134
rect 587582 119898 587818 120134
rect 587262 84218 587498 84454
rect 587582 84218 587818 84454
rect 587262 83898 587498 84134
rect 587582 83898 587818 84134
rect 587262 48218 587498 48454
rect 587582 48218 587818 48454
rect 587262 47898 587498 48134
rect 587582 47898 587818 48134
rect 587262 12218 587498 12454
rect 587582 12218 587818 12454
rect 587262 11898 587498 12134
rect 587582 11898 587818 12134
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 700718 588458 700954
rect 588542 700718 588778 700954
rect 588222 700398 588458 700634
rect 588542 700398 588778 700634
rect 588222 664718 588458 664954
rect 588542 664718 588778 664954
rect 588222 664398 588458 664634
rect 588542 664398 588778 664634
rect 588222 628718 588458 628954
rect 588542 628718 588778 628954
rect 588222 628398 588458 628634
rect 588542 628398 588778 628634
rect 588222 592718 588458 592954
rect 588542 592718 588778 592954
rect 588222 592398 588458 592634
rect 588542 592398 588778 592634
rect 588222 556718 588458 556954
rect 588542 556718 588778 556954
rect 588222 556398 588458 556634
rect 588542 556398 588778 556634
rect 588222 520718 588458 520954
rect 588542 520718 588778 520954
rect 588222 520398 588458 520634
rect 588542 520398 588778 520634
rect 588222 484718 588458 484954
rect 588542 484718 588778 484954
rect 588222 484398 588458 484634
rect 588542 484398 588778 484634
rect 588222 448718 588458 448954
rect 588542 448718 588778 448954
rect 588222 448398 588458 448634
rect 588542 448398 588778 448634
rect 588222 412718 588458 412954
rect 588542 412718 588778 412954
rect 588222 412398 588458 412634
rect 588542 412398 588778 412634
rect 588222 376718 588458 376954
rect 588542 376718 588778 376954
rect 588222 376398 588458 376634
rect 588542 376398 588778 376634
rect 588222 340718 588458 340954
rect 588542 340718 588778 340954
rect 588222 340398 588458 340634
rect 588542 340398 588778 340634
rect 588222 304718 588458 304954
rect 588542 304718 588778 304954
rect 588222 304398 588458 304634
rect 588542 304398 588778 304634
rect 588222 268718 588458 268954
rect 588542 268718 588778 268954
rect 588222 268398 588458 268634
rect 588542 268398 588778 268634
rect 588222 232718 588458 232954
rect 588542 232718 588778 232954
rect 588222 232398 588458 232634
rect 588542 232398 588778 232634
rect 588222 196718 588458 196954
rect 588542 196718 588778 196954
rect 588222 196398 588458 196634
rect 588542 196398 588778 196634
rect 588222 160718 588458 160954
rect 588542 160718 588778 160954
rect 588222 160398 588458 160634
rect 588542 160398 588778 160634
rect 588222 124718 588458 124954
rect 588542 124718 588778 124954
rect 588222 124398 588458 124634
rect 588542 124398 588778 124634
rect 588222 88718 588458 88954
rect 588542 88718 588778 88954
rect 588222 88398 588458 88634
rect 588542 88398 588778 88634
rect 588222 52718 588458 52954
rect 588542 52718 588778 52954
rect 588222 52398 588458 52634
rect 588542 52398 588778 52634
rect 588222 16718 588458 16954
rect 588542 16718 588778 16954
rect 588222 16398 588458 16634
rect 588542 16398 588778 16634
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 669218 589418 669454
rect 589502 669218 589738 669454
rect 589182 668898 589418 669134
rect 589502 668898 589738 669134
rect 589182 633218 589418 633454
rect 589502 633218 589738 633454
rect 589182 632898 589418 633134
rect 589502 632898 589738 633134
rect 589182 597218 589418 597454
rect 589502 597218 589738 597454
rect 589182 596898 589418 597134
rect 589502 596898 589738 597134
rect 589182 561218 589418 561454
rect 589502 561218 589738 561454
rect 589182 560898 589418 561134
rect 589502 560898 589738 561134
rect 589182 525218 589418 525454
rect 589502 525218 589738 525454
rect 589182 524898 589418 525134
rect 589502 524898 589738 525134
rect 589182 489218 589418 489454
rect 589502 489218 589738 489454
rect 589182 488898 589418 489134
rect 589502 488898 589738 489134
rect 589182 453218 589418 453454
rect 589502 453218 589738 453454
rect 589182 452898 589418 453134
rect 589502 452898 589738 453134
rect 589182 417218 589418 417454
rect 589502 417218 589738 417454
rect 589182 416898 589418 417134
rect 589502 416898 589738 417134
rect 589182 381218 589418 381454
rect 589502 381218 589738 381454
rect 589182 380898 589418 381134
rect 589502 380898 589738 381134
rect 589182 345218 589418 345454
rect 589502 345218 589738 345454
rect 589182 344898 589418 345134
rect 589502 344898 589738 345134
rect 589182 309218 589418 309454
rect 589502 309218 589738 309454
rect 589182 308898 589418 309134
rect 589502 308898 589738 309134
rect 589182 273218 589418 273454
rect 589502 273218 589738 273454
rect 589182 272898 589418 273134
rect 589502 272898 589738 273134
rect 589182 237218 589418 237454
rect 589502 237218 589738 237454
rect 589182 236898 589418 237134
rect 589502 236898 589738 237134
rect 589182 201218 589418 201454
rect 589502 201218 589738 201454
rect 589182 200898 589418 201134
rect 589502 200898 589738 201134
rect 589182 165218 589418 165454
rect 589502 165218 589738 165454
rect 589182 164898 589418 165134
rect 589502 164898 589738 165134
rect 589182 129218 589418 129454
rect 589502 129218 589738 129454
rect 589182 128898 589418 129134
rect 589502 128898 589738 129134
rect 589182 93218 589418 93454
rect 589502 93218 589738 93454
rect 589182 92898 589418 93134
rect 589502 92898 589738 93134
rect 589182 57218 589418 57454
rect 589502 57218 589738 57454
rect 589182 56898 589418 57134
rect 589502 56898 589738 57134
rect 589182 21218 589418 21454
rect 589502 21218 589738 21454
rect 589182 20898 589418 21134
rect 589502 20898 589738 21134
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 673718 590378 673954
rect 590462 673718 590698 673954
rect 590142 673398 590378 673634
rect 590462 673398 590698 673634
rect 590142 637718 590378 637954
rect 590462 637718 590698 637954
rect 590142 637398 590378 637634
rect 590462 637398 590698 637634
rect 590142 601718 590378 601954
rect 590462 601718 590698 601954
rect 590142 601398 590378 601634
rect 590462 601398 590698 601634
rect 590142 565718 590378 565954
rect 590462 565718 590698 565954
rect 590142 565398 590378 565634
rect 590462 565398 590698 565634
rect 590142 529718 590378 529954
rect 590462 529718 590698 529954
rect 590142 529398 590378 529634
rect 590462 529398 590698 529634
rect 590142 493718 590378 493954
rect 590462 493718 590698 493954
rect 590142 493398 590378 493634
rect 590462 493398 590698 493634
rect 590142 457718 590378 457954
rect 590462 457718 590698 457954
rect 590142 457398 590378 457634
rect 590462 457398 590698 457634
rect 590142 421718 590378 421954
rect 590462 421718 590698 421954
rect 590142 421398 590378 421634
rect 590462 421398 590698 421634
rect 590142 385718 590378 385954
rect 590462 385718 590698 385954
rect 590142 385398 590378 385634
rect 590462 385398 590698 385634
rect 590142 349718 590378 349954
rect 590462 349718 590698 349954
rect 590142 349398 590378 349634
rect 590462 349398 590698 349634
rect 590142 313718 590378 313954
rect 590462 313718 590698 313954
rect 590142 313398 590378 313634
rect 590462 313398 590698 313634
rect 590142 277718 590378 277954
rect 590462 277718 590698 277954
rect 590142 277398 590378 277634
rect 590462 277398 590698 277634
rect 590142 241718 590378 241954
rect 590462 241718 590698 241954
rect 590142 241398 590378 241634
rect 590462 241398 590698 241634
rect 590142 205718 590378 205954
rect 590462 205718 590698 205954
rect 590142 205398 590378 205634
rect 590462 205398 590698 205634
rect 590142 169718 590378 169954
rect 590462 169718 590698 169954
rect 590142 169398 590378 169634
rect 590462 169398 590698 169634
rect 590142 133718 590378 133954
rect 590462 133718 590698 133954
rect 590142 133398 590378 133634
rect 590462 133398 590698 133634
rect 590142 97718 590378 97954
rect 590462 97718 590698 97954
rect 590142 97398 590378 97634
rect 590462 97398 590698 97634
rect 590142 61718 590378 61954
rect 590462 61718 590698 61954
rect 590142 61398 590378 61634
rect 590462 61398 590698 61634
rect 590142 25718 590378 25954
rect 590462 25718 590698 25954
rect 590142 25398 590378 25634
rect 590462 25398 590698 25634
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 678218 591338 678454
rect 591422 678218 591658 678454
rect 591102 677898 591338 678134
rect 591422 677898 591658 678134
rect 591102 642218 591338 642454
rect 591422 642218 591658 642454
rect 591102 641898 591338 642134
rect 591422 641898 591658 642134
rect 591102 606218 591338 606454
rect 591422 606218 591658 606454
rect 591102 605898 591338 606134
rect 591422 605898 591658 606134
rect 591102 570218 591338 570454
rect 591422 570218 591658 570454
rect 591102 569898 591338 570134
rect 591422 569898 591658 570134
rect 591102 534218 591338 534454
rect 591422 534218 591658 534454
rect 591102 533898 591338 534134
rect 591422 533898 591658 534134
rect 591102 498218 591338 498454
rect 591422 498218 591658 498454
rect 591102 497898 591338 498134
rect 591422 497898 591658 498134
rect 591102 462218 591338 462454
rect 591422 462218 591658 462454
rect 591102 461898 591338 462134
rect 591422 461898 591658 462134
rect 591102 426218 591338 426454
rect 591422 426218 591658 426454
rect 591102 425898 591338 426134
rect 591422 425898 591658 426134
rect 591102 390218 591338 390454
rect 591422 390218 591658 390454
rect 591102 389898 591338 390134
rect 591422 389898 591658 390134
rect 591102 354218 591338 354454
rect 591422 354218 591658 354454
rect 591102 353898 591338 354134
rect 591422 353898 591658 354134
rect 591102 318218 591338 318454
rect 591422 318218 591658 318454
rect 591102 317898 591338 318134
rect 591422 317898 591658 318134
rect 591102 282218 591338 282454
rect 591422 282218 591658 282454
rect 591102 281898 591338 282134
rect 591422 281898 591658 282134
rect 591102 246218 591338 246454
rect 591422 246218 591658 246454
rect 591102 245898 591338 246134
rect 591422 245898 591658 246134
rect 591102 210218 591338 210454
rect 591422 210218 591658 210454
rect 591102 209898 591338 210134
rect 591422 209898 591658 210134
rect 591102 174218 591338 174454
rect 591422 174218 591658 174454
rect 591102 173898 591338 174134
rect 591422 173898 591658 174134
rect 591102 138218 591338 138454
rect 591422 138218 591658 138454
rect 591102 137898 591338 138134
rect 591422 137898 591658 138134
rect 591102 102218 591338 102454
rect 591422 102218 591658 102454
rect 591102 101898 591338 102134
rect 591422 101898 591658 102134
rect 591102 66218 591338 66454
rect 591422 66218 591658 66454
rect 591102 65898 591338 66134
rect 591422 65898 591658 66134
rect 591102 30218 591338 30454
rect 591422 30218 591658 30454
rect 591102 29898 591338 30134
rect 591422 29898 591658 30134
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 682718 592298 682954
rect 592382 682718 592618 682954
rect 592062 682398 592298 682634
rect 592382 682398 592618 682634
rect 592062 646718 592298 646954
rect 592382 646718 592618 646954
rect 592062 646398 592298 646634
rect 592382 646398 592618 646634
rect 592062 610718 592298 610954
rect 592382 610718 592618 610954
rect 592062 610398 592298 610634
rect 592382 610398 592618 610634
rect 592062 574718 592298 574954
rect 592382 574718 592618 574954
rect 592062 574398 592298 574634
rect 592382 574398 592618 574634
rect 592062 538718 592298 538954
rect 592382 538718 592618 538954
rect 592062 538398 592298 538634
rect 592382 538398 592618 538634
rect 592062 502718 592298 502954
rect 592382 502718 592618 502954
rect 592062 502398 592298 502634
rect 592382 502398 592618 502634
rect 592062 466718 592298 466954
rect 592382 466718 592618 466954
rect 592062 466398 592298 466634
rect 592382 466398 592618 466634
rect 592062 430718 592298 430954
rect 592382 430718 592618 430954
rect 592062 430398 592298 430634
rect 592382 430398 592618 430634
rect 592062 394718 592298 394954
rect 592382 394718 592618 394954
rect 592062 394398 592298 394634
rect 592382 394398 592618 394634
rect 592062 358718 592298 358954
rect 592382 358718 592618 358954
rect 592062 358398 592298 358634
rect 592382 358398 592618 358634
rect 592062 322718 592298 322954
rect 592382 322718 592618 322954
rect 592062 322398 592298 322634
rect 592382 322398 592618 322634
rect 592062 286718 592298 286954
rect 592382 286718 592618 286954
rect 592062 286398 592298 286634
rect 592382 286398 592618 286634
rect 592062 250718 592298 250954
rect 592382 250718 592618 250954
rect 592062 250398 592298 250634
rect 592382 250398 592618 250634
rect 592062 214718 592298 214954
rect 592382 214718 592618 214954
rect 592062 214398 592298 214634
rect 592382 214398 592618 214634
rect 592062 178718 592298 178954
rect 592382 178718 592618 178954
rect 592062 178398 592298 178634
rect 592382 178398 592618 178634
rect 592062 142718 592298 142954
rect 592382 142718 592618 142954
rect 592062 142398 592298 142634
rect 592382 142398 592618 142634
rect 592062 106718 592298 106954
rect 592382 106718 592618 106954
rect 592062 106398 592298 106634
rect 592382 106398 592618 106634
rect 592062 70718 592298 70954
rect 592382 70718 592618 70954
rect 592062 70398 592298 70634
rect 592382 70398 592618 70634
rect 592062 34718 592298 34954
rect 592382 34718 592618 34954
rect 592062 34398 592298 34634
rect 592382 34398 592618 34634
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 33326 711558
rect 33562 711322 33646 711558
rect 33882 711322 69326 711558
rect 69562 711322 69646 711558
rect 69882 711322 105326 711558
rect 105562 711322 105646 711558
rect 105882 711322 141326 711558
rect 141562 711322 141646 711558
rect 141882 711322 177326 711558
rect 177562 711322 177646 711558
rect 177882 711322 213326 711558
rect 213562 711322 213646 711558
rect 213882 711322 249326 711558
rect 249562 711322 249646 711558
rect 249882 711322 285326 711558
rect 285562 711322 285646 711558
rect 285882 711322 321326 711558
rect 321562 711322 321646 711558
rect 321882 711322 357326 711558
rect 357562 711322 357646 711558
rect 357882 711322 393326 711558
rect 393562 711322 393646 711558
rect 393882 711322 429326 711558
rect 429562 711322 429646 711558
rect 429882 711322 465326 711558
rect 465562 711322 465646 711558
rect 465882 711322 501326 711558
rect 501562 711322 501646 711558
rect 501882 711322 537326 711558
rect 537562 711322 537646 711558
rect 537882 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 33326 711238
rect 33562 711002 33646 711238
rect 33882 711002 69326 711238
rect 69562 711002 69646 711238
rect 69882 711002 105326 711238
rect 105562 711002 105646 711238
rect 105882 711002 141326 711238
rect 141562 711002 141646 711238
rect 141882 711002 177326 711238
rect 177562 711002 177646 711238
rect 177882 711002 213326 711238
rect 213562 711002 213646 711238
rect 213882 711002 249326 711238
rect 249562 711002 249646 711238
rect 249882 711002 285326 711238
rect 285562 711002 285646 711238
rect 285882 711002 321326 711238
rect 321562 711002 321646 711238
rect 321882 711002 357326 711238
rect 357562 711002 357646 711238
rect 357882 711002 393326 711238
rect 393562 711002 393646 711238
rect 393882 711002 429326 711238
rect 429562 711002 429646 711238
rect 429882 711002 465326 711238
rect 465562 711002 465646 711238
rect 465882 711002 501326 711238
rect 501562 711002 501646 711238
rect 501882 711002 537326 711238
rect 537562 711002 537646 711238
rect 537882 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 28826 710598
rect 29062 710362 29146 710598
rect 29382 710362 64826 710598
rect 65062 710362 65146 710598
rect 65382 710362 100826 710598
rect 101062 710362 101146 710598
rect 101382 710362 136826 710598
rect 137062 710362 137146 710598
rect 137382 710362 172826 710598
rect 173062 710362 173146 710598
rect 173382 710362 208826 710598
rect 209062 710362 209146 710598
rect 209382 710362 244826 710598
rect 245062 710362 245146 710598
rect 245382 710362 280826 710598
rect 281062 710362 281146 710598
rect 281382 710362 316826 710598
rect 317062 710362 317146 710598
rect 317382 710362 352826 710598
rect 353062 710362 353146 710598
rect 353382 710362 388826 710598
rect 389062 710362 389146 710598
rect 389382 710362 424826 710598
rect 425062 710362 425146 710598
rect 425382 710362 460826 710598
rect 461062 710362 461146 710598
rect 461382 710362 496826 710598
rect 497062 710362 497146 710598
rect 497382 710362 532826 710598
rect 533062 710362 533146 710598
rect 533382 710362 568826 710598
rect 569062 710362 569146 710598
rect 569382 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 28826 710278
rect 29062 710042 29146 710278
rect 29382 710042 64826 710278
rect 65062 710042 65146 710278
rect 65382 710042 100826 710278
rect 101062 710042 101146 710278
rect 101382 710042 136826 710278
rect 137062 710042 137146 710278
rect 137382 710042 172826 710278
rect 173062 710042 173146 710278
rect 173382 710042 208826 710278
rect 209062 710042 209146 710278
rect 209382 710042 244826 710278
rect 245062 710042 245146 710278
rect 245382 710042 280826 710278
rect 281062 710042 281146 710278
rect 281382 710042 316826 710278
rect 317062 710042 317146 710278
rect 317382 710042 352826 710278
rect 353062 710042 353146 710278
rect 353382 710042 388826 710278
rect 389062 710042 389146 710278
rect 389382 710042 424826 710278
rect 425062 710042 425146 710278
rect 425382 710042 460826 710278
rect 461062 710042 461146 710278
rect 461382 710042 496826 710278
rect 497062 710042 497146 710278
rect 497382 710042 532826 710278
rect 533062 710042 533146 710278
rect 533382 710042 568826 710278
rect 569062 710042 569146 710278
rect 569382 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 24326 709638
rect 24562 709402 24646 709638
rect 24882 709402 60326 709638
rect 60562 709402 60646 709638
rect 60882 709402 96326 709638
rect 96562 709402 96646 709638
rect 96882 709402 132326 709638
rect 132562 709402 132646 709638
rect 132882 709402 168326 709638
rect 168562 709402 168646 709638
rect 168882 709402 204326 709638
rect 204562 709402 204646 709638
rect 204882 709402 240326 709638
rect 240562 709402 240646 709638
rect 240882 709402 276326 709638
rect 276562 709402 276646 709638
rect 276882 709402 312326 709638
rect 312562 709402 312646 709638
rect 312882 709402 348326 709638
rect 348562 709402 348646 709638
rect 348882 709402 384326 709638
rect 384562 709402 384646 709638
rect 384882 709402 420326 709638
rect 420562 709402 420646 709638
rect 420882 709402 456326 709638
rect 456562 709402 456646 709638
rect 456882 709402 492326 709638
rect 492562 709402 492646 709638
rect 492882 709402 528326 709638
rect 528562 709402 528646 709638
rect 528882 709402 564326 709638
rect 564562 709402 564646 709638
rect 564882 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 24326 709318
rect 24562 709082 24646 709318
rect 24882 709082 60326 709318
rect 60562 709082 60646 709318
rect 60882 709082 96326 709318
rect 96562 709082 96646 709318
rect 96882 709082 132326 709318
rect 132562 709082 132646 709318
rect 132882 709082 168326 709318
rect 168562 709082 168646 709318
rect 168882 709082 204326 709318
rect 204562 709082 204646 709318
rect 204882 709082 240326 709318
rect 240562 709082 240646 709318
rect 240882 709082 276326 709318
rect 276562 709082 276646 709318
rect 276882 709082 312326 709318
rect 312562 709082 312646 709318
rect 312882 709082 348326 709318
rect 348562 709082 348646 709318
rect 348882 709082 384326 709318
rect 384562 709082 384646 709318
rect 384882 709082 420326 709318
rect 420562 709082 420646 709318
rect 420882 709082 456326 709318
rect 456562 709082 456646 709318
rect 456882 709082 492326 709318
rect 492562 709082 492646 709318
rect 492882 709082 528326 709318
rect 528562 709082 528646 709318
rect 528882 709082 564326 709318
rect 564562 709082 564646 709318
rect 564882 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 19826 708678
rect 20062 708442 20146 708678
rect 20382 708442 55826 708678
rect 56062 708442 56146 708678
rect 56382 708442 91826 708678
rect 92062 708442 92146 708678
rect 92382 708442 127826 708678
rect 128062 708442 128146 708678
rect 128382 708442 163826 708678
rect 164062 708442 164146 708678
rect 164382 708442 199826 708678
rect 200062 708442 200146 708678
rect 200382 708442 235826 708678
rect 236062 708442 236146 708678
rect 236382 708442 271826 708678
rect 272062 708442 272146 708678
rect 272382 708442 307826 708678
rect 308062 708442 308146 708678
rect 308382 708442 343826 708678
rect 344062 708442 344146 708678
rect 344382 708442 379826 708678
rect 380062 708442 380146 708678
rect 380382 708442 415826 708678
rect 416062 708442 416146 708678
rect 416382 708442 451826 708678
rect 452062 708442 452146 708678
rect 452382 708442 487826 708678
rect 488062 708442 488146 708678
rect 488382 708442 523826 708678
rect 524062 708442 524146 708678
rect 524382 708442 559826 708678
rect 560062 708442 560146 708678
rect 560382 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 19826 708358
rect 20062 708122 20146 708358
rect 20382 708122 55826 708358
rect 56062 708122 56146 708358
rect 56382 708122 91826 708358
rect 92062 708122 92146 708358
rect 92382 708122 127826 708358
rect 128062 708122 128146 708358
rect 128382 708122 163826 708358
rect 164062 708122 164146 708358
rect 164382 708122 199826 708358
rect 200062 708122 200146 708358
rect 200382 708122 235826 708358
rect 236062 708122 236146 708358
rect 236382 708122 271826 708358
rect 272062 708122 272146 708358
rect 272382 708122 307826 708358
rect 308062 708122 308146 708358
rect 308382 708122 343826 708358
rect 344062 708122 344146 708358
rect 344382 708122 379826 708358
rect 380062 708122 380146 708358
rect 380382 708122 415826 708358
rect 416062 708122 416146 708358
rect 416382 708122 451826 708358
rect 452062 708122 452146 708358
rect 452382 708122 487826 708358
rect 488062 708122 488146 708358
rect 488382 708122 523826 708358
rect 524062 708122 524146 708358
rect 524382 708122 559826 708358
rect 560062 708122 560146 708358
rect 560382 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 46826 706758
rect 47062 706522 47146 706758
rect 47382 706522 82826 706758
rect 83062 706522 83146 706758
rect 83382 706522 118826 706758
rect 119062 706522 119146 706758
rect 119382 706522 154826 706758
rect 155062 706522 155146 706758
rect 155382 706522 190826 706758
rect 191062 706522 191146 706758
rect 191382 706522 226826 706758
rect 227062 706522 227146 706758
rect 227382 706522 262826 706758
rect 263062 706522 263146 706758
rect 263382 706522 298826 706758
rect 299062 706522 299146 706758
rect 299382 706522 334826 706758
rect 335062 706522 335146 706758
rect 335382 706522 370826 706758
rect 371062 706522 371146 706758
rect 371382 706522 406826 706758
rect 407062 706522 407146 706758
rect 407382 706522 442826 706758
rect 443062 706522 443146 706758
rect 443382 706522 478826 706758
rect 479062 706522 479146 706758
rect 479382 706522 514826 706758
rect 515062 706522 515146 706758
rect 515382 706522 550826 706758
rect 551062 706522 551146 706758
rect 551382 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 46826 706438
rect 47062 706202 47146 706438
rect 47382 706202 82826 706438
rect 83062 706202 83146 706438
rect 83382 706202 118826 706438
rect 119062 706202 119146 706438
rect 119382 706202 154826 706438
rect 155062 706202 155146 706438
rect 155382 706202 190826 706438
rect 191062 706202 191146 706438
rect 191382 706202 226826 706438
rect 227062 706202 227146 706438
rect 227382 706202 262826 706438
rect 263062 706202 263146 706438
rect 263382 706202 298826 706438
rect 299062 706202 299146 706438
rect 299382 706202 334826 706438
rect 335062 706202 335146 706438
rect 335382 706202 370826 706438
rect 371062 706202 371146 706438
rect 371382 706202 406826 706438
rect 407062 706202 407146 706438
rect 407382 706202 442826 706438
rect 443062 706202 443146 706438
rect 443382 706202 478826 706438
rect 479062 706202 479146 706438
rect 479382 706202 514826 706438
rect 515062 706202 515146 706438
rect 515382 706202 550826 706438
rect 551062 706202 551146 706438
rect 551382 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 42326 705798
rect 42562 705562 42646 705798
rect 42882 705562 78326 705798
rect 78562 705562 78646 705798
rect 78882 705562 114326 705798
rect 114562 705562 114646 705798
rect 114882 705562 150326 705798
rect 150562 705562 150646 705798
rect 150882 705562 186326 705798
rect 186562 705562 186646 705798
rect 186882 705562 222326 705798
rect 222562 705562 222646 705798
rect 222882 705562 258326 705798
rect 258562 705562 258646 705798
rect 258882 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 330326 705798
rect 330562 705562 330646 705798
rect 330882 705562 366326 705798
rect 366562 705562 366646 705798
rect 366882 705562 402326 705798
rect 402562 705562 402646 705798
rect 402882 705562 438326 705798
rect 438562 705562 438646 705798
rect 438882 705562 474326 705798
rect 474562 705562 474646 705798
rect 474882 705562 510326 705798
rect 510562 705562 510646 705798
rect 510882 705562 546326 705798
rect 546562 705562 546646 705798
rect 546882 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 42326 705478
rect 42562 705242 42646 705478
rect 42882 705242 78326 705478
rect 78562 705242 78646 705478
rect 78882 705242 114326 705478
rect 114562 705242 114646 705478
rect 114882 705242 150326 705478
rect 150562 705242 150646 705478
rect 150882 705242 186326 705478
rect 186562 705242 186646 705478
rect 186882 705242 222326 705478
rect 222562 705242 222646 705478
rect 222882 705242 258326 705478
rect 258562 705242 258646 705478
rect 258882 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 330326 705478
rect 330562 705242 330646 705478
rect 330882 705242 366326 705478
rect 366562 705242 366646 705478
rect 366882 705242 402326 705478
rect 402562 705242 402646 705478
rect 402882 705242 438326 705478
rect 438562 705242 438646 705478
rect 438882 705242 474326 705478
rect 474562 705242 474646 705478
rect 474882 705242 510326 705478
rect 510562 705242 510646 705478
rect 510882 705242 546326 705478
rect 546562 705242 546646 705478
rect 546882 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 700954 592650 700986
rect -8726 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 592650 700954
rect -8726 700634 592650 700718
rect -8726 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 592650 700634
rect -8726 700366 592650 700398
rect -8726 696454 592650 696486
rect -8726 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 592650 696454
rect -8726 696134 592650 696218
rect -8726 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 592650 696134
rect -8726 695866 592650 695898
rect -8726 691954 592650 691986
rect -8726 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 592650 691954
rect -8726 691634 592650 691718
rect -8726 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 592650 691634
rect -8726 691366 592650 691398
rect -8726 687454 592650 687486
rect -8726 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 592650 687454
rect -8726 687134 592650 687218
rect -8726 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 592650 687134
rect -8726 686866 592650 686898
rect -8726 682954 592650 682986
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect -8726 682634 592650 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect -8726 682366 592650 682398
rect -8726 678454 592650 678486
rect -8726 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 424826 678454
rect 425062 678218 425146 678454
rect 425382 678218 460826 678454
rect 461062 678218 461146 678454
rect 461382 678218 496826 678454
rect 497062 678218 497146 678454
rect 497382 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 592650 678454
rect -8726 678134 592650 678218
rect -8726 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 424826 678134
rect 425062 677898 425146 678134
rect 425382 677898 460826 678134
rect 461062 677898 461146 678134
rect 461382 677898 496826 678134
rect 497062 677898 497146 678134
rect 497382 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 592650 678134
rect -8726 677866 592650 677898
rect -8726 673954 592650 673986
rect -8726 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 96326 673954
rect 96562 673718 96646 673954
rect 96882 673718 132326 673954
rect 132562 673718 132646 673954
rect 132882 673718 168326 673954
rect 168562 673718 168646 673954
rect 168882 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 240326 673954
rect 240562 673718 240646 673954
rect 240882 673718 276326 673954
rect 276562 673718 276646 673954
rect 276882 673718 312326 673954
rect 312562 673718 312646 673954
rect 312882 673718 348326 673954
rect 348562 673718 348646 673954
rect 348882 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 420326 673954
rect 420562 673718 420646 673954
rect 420882 673718 456326 673954
rect 456562 673718 456646 673954
rect 456882 673718 492326 673954
rect 492562 673718 492646 673954
rect 492882 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 592650 673954
rect -8726 673634 592650 673718
rect -8726 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 96326 673634
rect 96562 673398 96646 673634
rect 96882 673398 132326 673634
rect 132562 673398 132646 673634
rect 132882 673398 168326 673634
rect 168562 673398 168646 673634
rect 168882 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 240326 673634
rect 240562 673398 240646 673634
rect 240882 673398 276326 673634
rect 276562 673398 276646 673634
rect 276882 673398 312326 673634
rect 312562 673398 312646 673634
rect 312882 673398 348326 673634
rect 348562 673398 348646 673634
rect 348882 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 420326 673634
rect 420562 673398 420646 673634
rect 420882 673398 456326 673634
rect 456562 673398 456646 673634
rect 456882 673398 492326 673634
rect 492562 673398 492646 673634
rect 492882 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 592650 673634
rect -8726 673366 592650 673398
rect -8726 669454 592650 669486
rect -8726 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 592650 669454
rect -8726 669134 592650 669218
rect -8726 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 592650 669134
rect -8726 668866 592650 668898
rect -8726 664954 592650 664986
rect -8726 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 87326 664954
rect 87562 664718 87646 664954
rect 87882 664718 123326 664954
rect 123562 664718 123646 664954
rect 123882 664718 159326 664954
rect 159562 664718 159646 664954
rect 159882 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 231326 664954
rect 231562 664718 231646 664954
rect 231882 664718 267326 664954
rect 267562 664718 267646 664954
rect 267882 664718 303326 664954
rect 303562 664718 303646 664954
rect 303882 664718 339326 664954
rect 339562 664718 339646 664954
rect 339882 664718 375326 664954
rect 375562 664718 375646 664954
rect 375882 664718 411326 664954
rect 411562 664718 411646 664954
rect 411882 664718 447326 664954
rect 447562 664718 447646 664954
rect 447882 664718 483326 664954
rect 483562 664718 483646 664954
rect 483882 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 592650 664954
rect -8726 664634 592650 664718
rect -8726 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 87326 664634
rect 87562 664398 87646 664634
rect 87882 664398 123326 664634
rect 123562 664398 123646 664634
rect 123882 664398 159326 664634
rect 159562 664398 159646 664634
rect 159882 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 231326 664634
rect 231562 664398 231646 664634
rect 231882 664398 267326 664634
rect 267562 664398 267646 664634
rect 267882 664398 303326 664634
rect 303562 664398 303646 664634
rect 303882 664398 339326 664634
rect 339562 664398 339646 664634
rect 339882 664398 375326 664634
rect 375562 664398 375646 664634
rect 375882 664398 411326 664634
rect 411562 664398 411646 664634
rect 411882 664398 447326 664634
rect 447562 664398 447646 664634
rect 447882 664398 483326 664634
rect 483562 664398 483646 664634
rect 483882 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 592650 664634
rect -8726 664366 592650 664398
rect -8726 660454 592650 660486
rect -8726 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 82826 660454
rect 83062 660218 83146 660454
rect 83382 660218 118826 660454
rect 119062 660218 119146 660454
rect 119382 660218 154826 660454
rect 155062 660218 155146 660454
rect 155382 660218 190826 660454
rect 191062 660218 191146 660454
rect 191382 660218 226826 660454
rect 227062 660218 227146 660454
rect 227382 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 298826 660454
rect 299062 660218 299146 660454
rect 299382 660218 334826 660454
rect 335062 660218 335146 660454
rect 335382 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 442826 660454
rect 443062 660218 443146 660454
rect 443382 660218 478826 660454
rect 479062 660218 479146 660454
rect 479382 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 592650 660454
rect -8726 660134 592650 660218
rect -8726 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 82826 660134
rect 83062 659898 83146 660134
rect 83382 659898 118826 660134
rect 119062 659898 119146 660134
rect 119382 659898 154826 660134
rect 155062 659898 155146 660134
rect 155382 659898 190826 660134
rect 191062 659898 191146 660134
rect 191382 659898 226826 660134
rect 227062 659898 227146 660134
rect 227382 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 298826 660134
rect 299062 659898 299146 660134
rect 299382 659898 334826 660134
rect 335062 659898 335146 660134
rect 335382 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 442826 660134
rect 443062 659898 443146 660134
rect 443382 659898 478826 660134
rect 479062 659898 479146 660134
rect 479382 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 592650 660134
rect -8726 659866 592650 659898
rect -8726 655954 592650 655986
rect -8726 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 78326 655954
rect 78562 655718 78646 655954
rect 78882 655718 114326 655954
rect 114562 655718 114646 655954
rect 114882 655718 150326 655954
rect 150562 655718 150646 655954
rect 150882 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 222326 655954
rect 222562 655718 222646 655954
rect 222882 655718 258326 655954
rect 258562 655718 258646 655954
rect 258882 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 330326 655954
rect 330562 655718 330646 655954
rect 330882 655718 366326 655954
rect 366562 655718 366646 655954
rect 366882 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 438326 655954
rect 438562 655718 438646 655954
rect 438882 655718 474326 655954
rect 474562 655718 474646 655954
rect 474882 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 592650 655954
rect -8726 655634 592650 655718
rect -8726 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 78326 655634
rect 78562 655398 78646 655634
rect 78882 655398 114326 655634
rect 114562 655398 114646 655634
rect 114882 655398 150326 655634
rect 150562 655398 150646 655634
rect 150882 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 222326 655634
rect 222562 655398 222646 655634
rect 222882 655398 258326 655634
rect 258562 655398 258646 655634
rect 258882 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 330326 655634
rect 330562 655398 330646 655634
rect 330882 655398 366326 655634
rect 366562 655398 366646 655634
rect 366882 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 438326 655634
rect 438562 655398 438646 655634
rect 438882 655398 474326 655634
rect 474562 655398 474646 655634
rect 474882 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 592650 655634
rect -8726 655366 592650 655398
rect -8726 651454 592650 651486
rect -8726 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 592650 651454
rect -8726 651134 592650 651218
rect -8726 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 592650 651134
rect -8726 650866 592650 650898
rect -8726 646954 592650 646986
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 69326 646954
rect 69562 646718 69646 646954
rect 69882 646718 105326 646954
rect 105562 646718 105646 646954
rect 105882 646718 141326 646954
rect 141562 646718 141646 646954
rect 141882 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 213326 646954
rect 213562 646718 213646 646954
rect 213882 646718 249326 646954
rect 249562 646718 249646 646954
rect 249882 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 321326 646954
rect 321562 646718 321646 646954
rect 321882 646718 357326 646954
rect 357562 646718 357646 646954
rect 357882 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 429326 646954
rect 429562 646718 429646 646954
rect 429882 646718 465326 646954
rect 465562 646718 465646 646954
rect 465882 646718 501326 646954
rect 501562 646718 501646 646954
rect 501882 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect -8726 646634 592650 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 69326 646634
rect 69562 646398 69646 646634
rect 69882 646398 105326 646634
rect 105562 646398 105646 646634
rect 105882 646398 141326 646634
rect 141562 646398 141646 646634
rect 141882 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 213326 646634
rect 213562 646398 213646 646634
rect 213882 646398 249326 646634
rect 249562 646398 249646 646634
rect 249882 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 321326 646634
rect 321562 646398 321646 646634
rect 321882 646398 357326 646634
rect 357562 646398 357646 646634
rect 357882 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 429326 646634
rect 429562 646398 429646 646634
rect 429882 646398 465326 646634
rect 465562 646398 465646 646634
rect 465882 646398 501326 646634
rect 501562 646398 501646 646634
rect 501882 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect -8726 646366 592650 646398
rect -8726 642454 592650 642486
rect -8726 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 64826 642454
rect 65062 642218 65146 642454
rect 65382 642218 100826 642454
rect 101062 642218 101146 642454
rect 101382 642218 136826 642454
rect 137062 642218 137146 642454
rect 137382 642218 172826 642454
rect 173062 642218 173146 642454
rect 173382 642218 208826 642454
rect 209062 642218 209146 642454
rect 209382 642218 244826 642454
rect 245062 642218 245146 642454
rect 245382 642218 280826 642454
rect 281062 642218 281146 642454
rect 281382 642218 316826 642454
rect 317062 642218 317146 642454
rect 317382 642218 352826 642454
rect 353062 642218 353146 642454
rect 353382 642218 388826 642454
rect 389062 642218 389146 642454
rect 389382 642218 424826 642454
rect 425062 642218 425146 642454
rect 425382 642218 460826 642454
rect 461062 642218 461146 642454
rect 461382 642218 496826 642454
rect 497062 642218 497146 642454
rect 497382 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 592650 642454
rect -8726 642134 592650 642218
rect -8726 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 64826 642134
rect 65062 641898 65146 642134
rect 65382 641898 100826 642134
rect 101062 641898 101146 642134
rect 101382 641898 136826 642134
rect 137062 641898 137146 642134
rect 137382 641898 172826 642134
rect 173062 641898 173146 642134
rect 173382 641898 208826 642134
rect 209062 641898 209146 642134
rect 209382 641898 244826 642134
rect 245062 641898 245146 642134
rect 245382 641898 280826 642134
rect 281062 641898 281146 642134
rect 281382 641898 316826 642134
rect 317062 641898 317146 642134
rect 317382 641898 352826 642134
rect 353062 641898 353146 642134
rect 353382 641898 388826 642134
rect 389062 641898 389146 642134
rect 389382 641898 424826 642134
rect 425062 641898 425146 642134
rect 425382 641898 460826 642134
rect 461062 641898 461146 642134
rect 461382 641898 496826 642134
rect 497062 641898 497146 642134
rect 497382 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 592650 642134
rect -8726 641866 592650 641898
rect -8726 637954 592650 637986
rect -8726 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 60326 637954
rect 60562 637718 60646 637954
rect 60882 637718 96326 637954
rect 96562 637718 96646 637954
rect 96882 637718 132326 637954
rect 132562 637718 132646 637954
rect 132882 637718 168326 637954
rect 168562 637718 168646 637954
rect 168882 637718 204326 637954
rect 204562 637718 204646 637954
rect 204882 637718 240326 637954
rect 240562 637718 240646 637954
rect 240882 637718 276326 637954
rect 276562 637718 276646 637954
rect 276882 637718 312326 637954
rect 312562 637718 312646 637954
rect 312882 637718 348326 637954
rect 348562 637718 348646 637954
rect 348882 637718 384326 637954
rect 384562 637718 384646 637954
rect 384882 637718 420326 637954
rect 420562 637718 420646 637954
rect 420882 637718 456326 637954
rect 456562 637718 456646 637954
rect 456882 637718 492326 637954
rect 492562 637718 492646 637954
rect 492882 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 592650 637954
rect -8726 637634 592650 637718
rect -8726 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 60326 637634
rect 60562 637398 60646 637634
rect 60882 637398 96326 637634
rect 96562 637398 96646 637634
rect 96882 637398 132326 637634
rect 132562 637398 132646 637634
rect 132882 637398 168326 637634
rect 168562 637398 168646 637634
rect 168882 637398 204326 637634
rect 204562 637398 204646 637634
rect 204882 637398 240326 637634
rect 240562 637398 240646 637634
rect 240882 637398 276326 637634
rect 276562 637398 276646 637634
rect 276882 637398 312326 637634
rect 312562 637398 312646 637634
rect 312882 637398 348326 637634
rect 348562 637398 348646 637634
rect 348882 637398 384326 637634
rect 384562 637398 384646 637634
rect 384882 637398 420326 637634
rect 420562 637398 420646 637634
rect 420882 637398 456326 637634
rect 456562 637398 456646 637634
rect 456882 637398 492326 637634
rect 492562 637398 492646 637634
rect 492882 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 592650 637634
rect -8726 637366 592650 637398
rect -8726 633454 592650 633486
rect -8726 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 592650 633454
rect -8726 633134 592650 633218
rect -8726 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 592650 633134
rect -8726 632866 592650 632898
rect -8726 628954 592650 628986
rect -8726 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 51326 628954
rect 51562 628718 51646 628954
rect 51882 628718 87326 628954
rect 87562 628718 87646 628954
rect 87882 628718 123326 628954
rect 123562 628718 123646 628954
rect 123882 628718 159326 628954
rect 159562 628718 159646 628954
rect 159882 628718 195326 628954
rect 195562 628718 195646 628954
rect 195882 628718 231326 628954
rect 231562 628718 231646 628954
rect 231882 628718 267326 628954
rect 267562 628718 267646 628954
rect 267882 628718 303326 628954
rect 303562 628718 303646 628954
rect 303882 628718 339326 628954
rect 339562 628718 339646 628954
rect 339882 628718 375326 628954
rect 375562 628718 375646 628954
rect 375882 628718 411326 628954
rect 411562 628718 411646 628954
rect 411882 628718 447326 628954
rect 447562 628718 447646 628954
rect 447882 628718 483326 628954
rect 483562 628718 483646 628954
rect 483882 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 592650 628954
rect -8726 628634 592650 628718
rect -8726 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 51326 628634
rect 51562 628398 51646 628634
rect 51882 628398 87326 628634
rect 87562 628398 87646 628634
rect 87882 628398 123326 628634
rect 123562 628398 123646 628634
rect 123882 628398 159326 628634
rect 159562 628398 159646 628634
rect 159882 628398 195326 628634
rect 195562 628398 195646 628634
rect 195882 628398 231326 628634
rect 231562 628398 231646 628634
rect 231882 628398 267326 628634
rect 267562 628398 267646 628634
rect 267882 628398 303326 628634
rect 303562 628398 303646 628634
rect 303882 628398 339326 628634
rect 339562 628398 339646 628634
rect 339882 628398 375326 628634
rect 375562 628398 375646 628634
rect 375882 628398 411326 628634
rect 411562 628398 411646 628634
rect 411882 628398 447326 628634
rect 447562 628398 447646 628634
rect 447882 628398 483326 628634
rect 483562 628398 483646 628634
rect 483882 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 592650 628634
rect -8726 628366 592650 628398
rect -8726 624454 592650 624486
rect -8726 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 82826 624454
rect 83062 624218 83146 624454
rect 83382 624218 118826 624454
rect 119062 624218 119146 624454
rect 119382 624218 154826 624454
rect 155062 624218 155146 624454
rect 155382 624218 190826 624454
rect 191062 624218 191146 624454
rect 191382 624218 226826 624454
rect 227062 624218 227146 624454
rect 227382 624218 262826 624454
rect 263062 624218 263146 624454
rect 263382 624218 298826 624454
rect 299062 624218 299146 624454
rect 299382 624218 334826 624454
rect 335062 624218 335146 624454
rect 335382 624218 370826 624454
rect 371062 624218 371146 624454
rect 371382 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 442826 624454
rect 443062 624218 443146 624454
rect 443382 624218 478826 624454
rect 479062 624218 479146 624454
rect 479382 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 592650 624454
rect -8726 624134 592650 624218
rect -8726 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 82826 624134
rect 83062 623898 83146 624134
rect 83382 623898 118826 624134
rect 119062 623898 119146 624134
rect 119382 623898 154826 624134
rect 155062 623898 155146 624134
rect 155382 623898 190826 624134
rect 191062 623898 191146 624134
rect 191382 623898 226826 624134
rect 227062 623898 227146 624134
rect 227382 623898 262826 624134
rect 263062 623898 263146 624134
rect 263382 623898 298826 624134
rect 299062 623898 299146 624134
rect 299382 623898 334826 624134
rect 335062 623898 335146 624134
rect 335382 623898 370826 624134
rect 371062 623898 371146 624134
rect 371382 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 442826 624134
rect 443062 623898 443146 624134
rect 443382 623898 478826 624134
rect 479062 623898 479146 624134
rect 479382 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 592650 624134
rect -8726 623866 592650 623898
rect -8726 619954 592650 619986
rect -8726 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 78326 619954
rect 78562 619718 78646 619954
rect 78882 619718 114326 619954
rect 114562 619718 114646 619954
rect 114882 619718 150326 619954
rect 150562 619718 150646 619954
rect 150882 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 222326 619954
rect 222562 619718 222646 619954
rect 222882 619718 258326 619954
rect 258562 619718 258646 619954
rect 258882 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 330326 619954
rect 330562 619718 330646 619954
rect 330882 619718 366326 619954
rect 366562 619718 366646 619954
rect 366882 619718 402326 619954
rect 402562 619718 402646 619954
rect 402882 619718 438326 619954
rect 438562 619718 438646 619954
rect 438882 619718 474326 619954
rect 474562 619718 474646 619954
rect 474882 619718 510326 619954
rect 510562 619718 510646 619954
rect 510882 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 592650 619954
rect -8726 619634 592650 619718
rect -8726 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 78326 619634
rect 78562 619398 78646 619634
rect 78882 619398 114326 619634
rect 114562 619398 114646 619634
rect 114882 619398 150326 619634
rect 150562 619398 150646 619634
rect 150882 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 222326 619634
rect 222562 619398 222646 619634
rect 222882 619398 258326 619634
rect 258562 619398 258646 619634
rect 258882 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 330326 619634
rect 330562 619398 330646 619634
rect 330882 619398 366326 619634
rect 366562 619398 366646 619634
rect 366882 619398 402326 619634
rect 402562 619398 402646 619634
rect 402882 619398 438326 619634
rect 438562 619398 438646 619634
rect 438882 619398 474326 619634
rect 474562 619398 474646 619634
rect 474882 619398 510326 619634
rect 510562 619398 510646 619634
rect 510882 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 592650 619634
rect -8726 619366 592650 619398
rect -8726 615454 592650 615486
rect -8726 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 592650 615454
rect -8726 615134 592650 615218
rect -8726 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 592650 615134
rect -8726 614866 592650 614898
rect -8726 610954 592650 610986
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 69326 610954
rect 69562 610718 69646 610954
rect 69882 610718 105326 610954
rect 105562 610718 105646 610954
rect 105882 610718 141326 610954
rect 141562 610718 141646 610954
rect 141882 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 213326 610954
rect 213562 610718 213646 610954
rect 213882 610718 249326 610954
rect 249562 610718 249646 610954
rect 249882 610718 285326 610954
rect 285562 610718 285646 610954
rect 285882 610718 321326 610954
rect 321562 610718 321646 610954
rect 321882 610718 357326 610954
rect 357562 610718 357646 610954
rect 357882 610718 393326 610954
rect 393562 610718 393646 610954
rect 393882 610718 429326 610954
rect 429562 610718 429646 610954
rect 429882 610718 465326 610954
rect 465562 610718 465646 610954
rect 465882 610718 501326 610954
rect 501562 610718 501646 610954
rect 501882 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect -8726 610634 592650 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 69326 610634
rect 69562 610398 69646 610634
rect 69882 610398 105326 610634
rect 105562 610398 105646 610634
rect 105882 610398 141326 610634
rect 141562 610398 141646 610634
rect 141882 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 213326 610634
rect 213562 610398 213646 610634
rect 213882 610398 249326 610634
rect 249562 610398 249646 610634
rect 249882 610398 285326 610634
rect 285562 610398 285646 610634
rect 285882 610398 321326 610634
rect 321562 610398 321646 610634
rect 321882 610398 357326 610634
rect 357562 610398 357646 610634
rect 357882 610398 393326 610634
rect 393562 610398 393646 610634
rect 393882 610398 429326 610634
rect 429562 610398 429646 610634
rect 429882 610398 465326 610634
rect 465562 610398 465646 610634
rect 465882 610398 501326 610634
rect 501562 610398 501646 610634
rect 501882 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect -8726 610366 592650 610398
rect -8726 606454 592650 606486
rect -8726 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 64826 606454
rect 65062 606218 65146 606454
rect 65382 606218 100826 606454
rect 101062 606218 101146 606454
rect 101382 606218 136826 606454
rect 137062 606218 137146 606454
rect 137382 606218 172826 606454
rect 173062 606218 173146 606454
rect 173382 606218 208826 606454
rect 209062 606218 209146 606454
rect 209382 606218 244826 606454
rect 245062 606218 245146 606454
rect 245382 606218 280826 606454
rect 281062 606218 281146 606454
rect 281382 606218 316826 606454
rect 317062 606218 317146 606454
rect 317382 606218 352826 606454
rect 353062 606218 353146 606454
rect 353382 606218 388826 606454
rect 389062 606218 389146 606454
rect 389382 606218 424826 606454
rect 425062 606218 425146 606454
rect 425382 606218 460826 606454
rect 461062 606218 461146 606454
rect 461382 606218 496826 606454
rect 497062 606218 497146 606454
rect 497382 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 592650 606454
rect -8726 606134 592650 606218
rect -8726 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 64826 606134
rect 65062 605898 65146 606134
rect 65382 605898 100826 606134
rect 101062 605898 101146 606134
rect 101382 605898 136826 606134
rect 137062 605898 137146 606134
rect 137382 605898 172826 606134
rect 173062 605898 173146 606134
rect 173382 605898 208826 606134
rect 209062 605898 209146 606134
rect 209382 605898 244826 606134
rect 245062 605898 245146 606134
rect 245382 605898 280826 606134
rect 281062 605898 281146 606134
rect 281382 605898 316826 606134
rect 317062 605898 317146 606134
rect 317382 605898 352826 606134
rect 353062 605898 353146 606134
rect 353382 605898 388826 606134
rect 389062 605898 389146 606134
rect 389382 605898 424826 606134
rect 425062 605898 425146 606134
rect 425382 605898 460826 606134
rect 461062 605898 461146 606134
rect 461382 605898 496826 606134
rect 497062 605898 497146 606134
rect 497382 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 592650 606134
rect -8726 605866 592650 605898
rect -8726 601954 592650 601986
rect -8726 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 60326 601954
rect 60562 601718 60646 601954
rect 60882 601718 96326 601954
rect 96562 601718 96646 601954
rect 96882 601718 132326 601954
rect 132562 601718 132646 601954
rect 132882 601718 168326 601954
rect 168562 601718 168646 601954
rect 168882 601718 204326 601954
rect 204562 601718 204646 601954
rect 204882 601718 240326 601954
rect 240562 601718 240646 601954
rect 240882 601718 276326 601954
rect 276562 601718 276646 601954
rect 276882 601718 312326 601954
rect 312562 601718 312646 601954
rect 312882 601718 348326 601954
rect 348562 601718 348646 601954
rect 348882 601718 384326 601954
rect 384562 601718 384646 601954
rect 384882 601718 420326 601954
rect 420562 601718 420646 601954
rect 420882 601718 456326 601954
rect 456562 601718 456646 601954
rect 456882 601718 492326 601954
rect 492562 601718 492646 601954
rect 492882 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 592650 601954
rect -8726 601634 592650 601718
rect -8726 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 60326 601634
rect 60562 601398 60646 601634
rect 60882 601398 96326 601634
rect 96562 601398 96646 601634
rect 96882 601398 132326 601634
rect 132562 601398 132646 601634
rect 132882 601398 168326 601634
rect 168562 601398 168646 601634
rect 168882 601398 204326 601634
rect 204562 601398 204646 601634
rect 204882 601398 240326 601634
rect 240562 601398 240646 601634
rect 240882 601398 276326 601634
rect 276562 601398 276646 601634
rect 276882 601398 312326 601634
rect 312562 601398 312646 601634
rect 312882 601398 348326 601634
rect 348562 601398 348646 601634
rect 348882 601398 384326 601634
rect 384562 601398 384646 601634
rect 384882 601398 420326 601634
rect 420562 601398 420646 601634
rect 420882 601398 456326 601634
rect 456562 601398 456646 601634
rect 456882 601398 492326 601634
rect 492562 601398 492646 601634
rect 492882 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 592650 601634
rect -8726 601366 592650 601398
rect -8726 597454 592650 597486
rect -8726 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 592650 597454
rect -8726 597134 592650 597218
rect -8726 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 592650 597134
rect -8726 596866 592650 596898
rect -8726 592954 592650 592986
rect -8726 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 51326 592954
rect 51562 592718 51646 592954
rect 51882 592718 87326 592954
rect 87562 592718 87646 592954
rect 87882 592718 123326 592954
rect 123562 592718 123646 592954
rect 123882 592718 159326 592954
rect 159562 592718 159646 592954
rect 159882 592718 195326 592954
rect 195562 592718 195646 592954
rect 195882 592718 231326 592954
rect 231562 592718 231646 592954
rect 231882 592718 267326 592954
rect 267562 592718 267646 592954
rect 267882 592718 303326 592954
rect 303562 592718 303646 592954
rect 303882 592718 339326 592954
rect 339562 592718 339646 592954
rect 339882 592718 375326 592954
rect 375562 592718 375646 592954
rect 375882 592718 411326 592954
rect 411562 592718 411646 592954
rect 411882 592718 447326 592954
rect 447562 592718 447646 592954
rect 447882 592718 483326 592954
rect 483562 592718 483646 592954
rect 483882 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 592650 592954
rect -8726 592634 592650 592718
rect -8726 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 51326 592634
rect 51562 592398 51646 592634
rect 51882 592398 87326 592634
rect 87562 592398 87646 592634
rect 87882 592398 123326 592634
rect 123562 592398 123646 592634
rect 123882 592398 159326 592634
rect 159562 592398 159646 592634
rect 159882 592398 195326 592634
rect 195562 592398 195646 592634
rect 195882 592398 231326 592634
rect 231562 592398 231646 592634
rect 231882 592398 267326 592634
rect 267562 592398 267646 592634
rect 267882 592398 303326 592634
rect 303562 592398 303646 592634
rect 303882 592398 339326 592634
rect 339562 592398 339646 592634
rect 339882 592398 375326 592634
rect 375562 592398 375646 592634
rect 375882 592398 411326 592634
rect 411562 592398 411646 592634
rect 411882 592398 447326 592634
rect 447562 592398 447646 592634
rect 447882 592398 483326 592634
rect 483562 592398 483646 592634
rect 483882 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 592650 592634
rect -8726 592366 592650 592398
rect -8726 588454 592650 588486
rect -8726 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 82826 588454
rect 83062 588218 83146 588454
rect 83382 588218 118826 588454
rect 119062 588218 119146 588454
rect 119382 588218 154826 588454
rect 155062 588218 155146 588454
rect 155382 588218 190826 588454
rect 191062 588218 191146 588454
rect 191382 588218 226826 588454
rect 227062 588218 227146 588454
rect 227382 588218 262826 588454
rect 263062 588218 263146 588454
rect 263382 588218 298826 588454
rect 299062 588218 299146 588454
rect 299382 588218 334826 588454
rect 335062 588218 335146 588454
rect 335382 588218 370826 588454
rect 371062 588218 371146 588454
rect 371382 588218 406826 588454
rect 407062 588218 407146 588454
rect 407382 588218 442826 588454
rect 443062 588218 443146 588454
rect 443382 588218 478826 588454
rect 479062 588218 479146 588454
rect 479382 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 592650 588454
rect -8726 588134 592650 588218
rect -8726 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 82826 588134
rect 83062 587898 83146 588134
rect 83382 587898 118826 588134
rect 119062 587898 119146 588134
rect 119382 587898 154826 588134
rect 155062 587898 155146 588134
rect 155382 587898 190826 588134
rect 191062 587898 191146 588134
rect 191382 587898 226826 588134
rect 227062 587898 227146 588134
rect 227382 587898 262826 588134
rect 263062 587898 263146 588134
rect 263382 587898 298826 588134
rect 299062 587898 299146 588134
rect 299382 587898 334826 588134
rect 335062 587898 335146 588134
rect 335382 587898 370826 588134
rect 371062 587898 371146 588134
rect 371382 587898 406826 588134
rect 407062 587898 407146 588134
rect 407382 587898 442826 588134
rect 443062 587898 443146 588134
rect 443382 587898 478826 588134
rect 479062 587898 479146 588134
rect 479382 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 592650 588134
rect -8726 587866 592650 587898
rect -8726 583954 592650 583986
rect -8726 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 78326 583954
rect 78562 583718 78646 583954
rect 78882 583718 114326 583954
rect 114562 583718 114646 583954
rect 114882 583718 150326 583954
rect 150562 583718 150646 583954
rect 150882 583718 186326 583954
rect 186562 583718 186646 583954
rect 186882 583718 222326 583954
rect 222562 583718 222646 583954
rect 222882 583718 258326 583954
rect 258562 583718 258646 583954
rect 258882 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 330326 583954
rect 330562 583718 330646 583954
rect 330882 583718 366326 583954
rect 366562 583718 366646 583954
rect 366882 583718 402326 583954
rect 402562 583718 402646 583954
rect 402882 583718 438326 583954
rect 438562 583718 438646 583954
rect 438882 583718 474326 583954
rect 474562 583718 474646 583954
rect 474882 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 592650 583954
rect -8726 583634 592650 583718
rect -8726 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 78326 583634
rect 78562 583398 78646 583634
rect 78882 583398 114326 583634
rect 114562 583398 114646 583634
rect 114882 583398 150326 583634
rect 150562 583398 150646 583634
rect 150882 583398 186326 583634
rect 186562 583398 186646 583634
rect 186882 583398 222326 583634
rect 222562 583398 222646 583634
rect 222882 583398 258326 583634
rect 258562 583398 258646 583634
rect 258882 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 330326 583634
rect 330562 583398 330646 583634
rect 330882 583398 366326 583634
rect 366562 583398 366646 583634
rect 366882 583398 402326 583634
rect 402562 583398 402646 583634
rect 402882 583398 438326 583634
rect 438562 583398 438646 583634
rect 438882 583398 474326 583634
rect 474562 583398 474646 583634
rect 474882 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 592650 583634
rect -8726 583366 592650 583398
rect -8726 579454 592650 579486
rect -8726 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 592650 579454
rect -8726 579134 592650 579218
rect -8726 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 592650 579134
rect -8726 578866 592650 578898
rect -8726 574954 592650 574986
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 69326 574954
rect 69562 574718 69646 574954
rect 69882 574718 105326 574954
rect 105562 574718 105646 574954
rect 105882 574718 141326 574954
rect 141562 574718 141646 574954
rect 141882 574718 177326 574954
rect 177562 574718 177646 574954
rect 177882 574718 213326 574954
rect 213562 574718 213646 574954
rect 213882 574718 249326 574954
rect 249562 574718 249646 574954
rect 249882 574718 285326 574954
rect 285562 574718 285646 574954
rect 285882 574718 321326 574954
rect 321562 574718 321646 574954
rect 321882 574718 357326 574954
rect 357562 574718 357646 574954
rect 357882 574718 393326 574954
rect 393562 574718 393646 574954
rect 393882 574718 429326 574954
rect 429562 574718 429646 574954
rect 429882 574718 465326 574954
rect 465562 574718 465646 574954
rect 465882 574718 501326 574954
rect 501562 574718 501646 574954
rect 501882 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect -8726 574634 592650 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 69326 574634
rect 69562 574398 69646 574634
rect 69882 574398 105326 574634
rect 105562 574398 105646 574634
rect 105882 574398 141326 574634
rect 141562 574398 141646 574634
rect 141882 574398 177326 574634
rect 177562 574398 177646 574634
rect 177882 574398 213326 574634
rect 213562 574398 213646 574634
rect 213882 574398 249326 574634
rect 249562 574398 249646 574634
rect 249882 574398 285326 574634
rect 285562 574398 285646 574634
rect 285882 574398 321326 574634
rect 321562 574398 321646 574634
rect 321882 574398 357326 574634
rect 357562 574398 357646 574634
rect 357882 574398 393326 574634
rect 393562 574398 393646 574634
rect 393882 574398 429326 574634
rect 429562 574398 429646 574634
rect 429882 574398 465326 574634
rect 465562 574398 465646 574634
rect 465882 574398 501326 574634
rect 501562 574398 501646 574634
rect 501882 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect -8726 574366 592650 574398
rect -8726 570454 592650 570486
rect -8726 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 64826 570454
rect 65062 570218 65146 570454
rect 65382 570218 100826 570454
rect 101062 570218 101146 570454
rect 101382 570218 136826 570454
rect 137062 570218 137146 570454
rect 137382 570218 172826 570454
rect 173062 570218 173146 570454
rect 173382 570218 208826 570454
rect 209062 570218 209146 570454
rect 209382 570218 244826 570454
rect 245062 570218 245146 570454
rect 245382 570218 280826 570454
rect 281062 570218 281146 570454
rect 281382 570218 316826 570454
rect 317062 570218 317146 570454
rect 317382 570218 352826 570454
rect 353062 570218 353146 570454
rect 353382 570218 388826 570454
rect 389062 570218 389146 570454
rect 389382 570218 424826 570454
rect 425062 570218 425146 570454
rect 425382 570218 460826 570454
rect 461062 570218 461146 570454
rect 461382 570218 496826 570454
rect 497062 570218 497146 570454
rect 497382 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 592650 570454
rect -8726 570134 592650 570218
rect -8726 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 64826 570134
rect 65062 569898 65146 570134
rect 65382 569898 100826 570134
rect 101062 569898 101146 570134
rect 101382 569898 136826 570134
rect 137062 569898 137146 570134
rect 137382 569898 172826 570134
rect 173062 569898 173146 570134
rect 173382 569898 208826 570134
rect 209062 569898 209146 570134
rect 209382 569898 244826 570134
rect 245062 569898 245146 570134
rect 245382 569898 280826 570134
rect 281062 569898 281146 570134
rect 281382 569898 316826 570134
rect 317062 569898 317146 570134
rect 317382 569898 352826 570134
rect 353062 569898 353146 570134
rect 353382 569898 388826 570134
rect 389062 569898 389146 570134
rect 389382 569898 424826 570134
rect 425062 569898 425146 570134
rect 425382 569898 460826 570134
rect 461062 569898 461146 570134
rect 461382 569898 496826 570134
rect 497062 569898 497146 570134
rect 497382 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 592650 570134
rect -8726 569866 592650 569898
rect -8726 565954 592650 565986
rect -8726 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 60326 565954
rect 60562 565718 60646 565954
rect 60882 565718 96326 565954
rect 96562 565718 96646 565954
rect 96882 565718 132326 565954
rect 132562 565718 132646 565954
rect 132882 565718 168326 565954
rect 168562 565718 168646 565954
rect 168882 565718 204326 565954
rect 204562 565718 204646 565954
rect 204882 565718 240326 565954
rect 240562 565718 240646 565954
rect 240882 565718 276326 565954
rect 276562 565718 276646 565954
rect 276882 565718 312326 565954
rect 312562 565718 312646 565954
rect 312882 565718 348326 565954
rect 348562 565718 348646 565954
rect 348882 565718 384326 565954
rect 384562 565718 384646 565954
rect 384882 565718 420326 565954
rect 420562 565718 420646 565954
rect 420882 565718 456326 565954
rect 456562 565718 456646 565954
rect 456882 565718 492326 565954
rect 492562 565718 492646 565954
rect 492882 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 592650 565954
rect -8726 565634 592650 565718
rect -8726 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 60326 565634
rect 60562 565398 60646 565634
rect 60882 565398 96326 565634
rect 96562 565398 96646 565634
rect 96882 565398 132326 565634
rect 132562 565398 132646 565634
rect 132882 565398 168326 565634
rect 168562 565398 168646 565634
rect 168882 565398 204326 565634
rect 204562 565398 204646 565634
rect 204882 565398 240326 565634
rect 240562 565398 240646 565634
rect 240882 565398 276326 565634
rect 276562 565398 276646 565634
rect 276882 565398 312326 565634
rect 312562 565398 312646 565634
rect 312882 565398 348326 565634
rect 348562 565398 348646 565634
rect 348882 565398 384326 565634
rect 384562 565398 384646 565634
rect 384882 565398 420326 565634
rect 420562 565398 420646 565634
rect 420882 565398 456326 565634
rect 456562 565398 456646 565634
rect 456882 565398 492326 565634
rect 492562 565398 492646 565634
rect 492882 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 592650 565634
rect -8726 565366 592650 565398
rect -8726 561454 592650 561486
rect -8726 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 592650 561454
rect -8726 561134 592650 561218
rect -8726 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 592650 561134
rect -8726 560866 592650 560898
rect -8726 556954 592650 556986
rect -8726 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 51326 556954
rect 51562 556718 51646 556954
rect 51882 556718 87326 556954
rect 87562 556718 87646 556954
rect 87882 556718 123326 556954
rect 123562 556718 123646 556954
rect 123882 556718 159326 556954
rect 159562 556718 159646 556954
rect 159882 556718 195326 556954
rect 195562 556718 195646 556954
rect 195882 556718 231326 556954
rect 231562 556718 231646 556954
rect 231882 556718 267326 556954
rect 267562 556718 267646 556954
rect 267882 556718 303326 556954
rect 303562 556718 303646 556954
rect 303882 556718 339326 556954
rect 339562 556718 339646 556954
rect 339882 556718 375326 556954
rect 375562 556718 375646 556954
rect 375882 556718 411326 556954
rect 411562 556718 411646 556954
rect 411882 556718 447326 556954
rect 447562 556718 447646 556954
rect 447882 556718 483326 556954
rect 483562 556718 483646 556954
rect 483882 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 592650 556954
rect -8726 556634 592650 556718
rect -8726 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 51326 556634
rect 51562 556398 51646 556634
rect 51882 556398 87326 556634
rect 87562 556398 87646 556634
rect 87882 556398 123326 556634
rect 123562 556398 123646 556634
rect 123882 556398 159326 556634
rect 159562 556398 159646 556634
rect 159882 556398 195326 556634
rect 195562 556398 195646 556634
rect 195882 556398 231326 556634
rect 231562 556398 231646 556634
rect 231882 556398 267326 556634
rect 267562 556398 267646 556634
rect 267882 556398 303326 556634
rect 303562 556398 303646 556634
rect 303882 556398 339326 556634
rect 339562 556398 339646 556634
rect 339882 556398 375326 556634
rect 375562 556398 375646 556634
rect 375882 556398 411326 556634
rect 411562 556398 411646 556634
rect 411882 556398 447326 556634
rect 447562 556398 447646 556634
rect 447882 556398 483326 556634
rect 483562 556398 483646 556634
rect 483882 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 592650 556634
rect -8726 556366 592650 556398
rect -8726 552454 592650 552486
rect -8726 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 82826 552454
rect 83062 552218 83146 552454
rect 83382 552218 118826 552454
rect 119062 552218 119146 552454
rect 119382 552218 154826 552454
rect 155062 552218 155146 552454
rect 155382 552218 190826 552454
rect 191062 552218 191146 552454
rect 191382 552218 226826 552454
rect 227062 552218 227146 552454
rect 227382 552218 262826 552454
rect 263062 552218 263146 552454
rect 263382 552218 298826 552454
rect 299062 552218 299146 552454
rect 299382 552218 334826 552454
rect 335062 552218 335146 552454
rect 335382 552218 370826 552454
rect 371062 552218 371146 552454
rect 371382 552218 406826 552454
rect 407062 552218 407146 552454
rect 407382 552218 442826 552454
rect 443062 552218 443146 552454
rect 443382 552218 478826 552454
rect 479062 552218 479146 552454
rect 479382 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 592650 552454
rect -8726 552134 592650 552218
rect -8726 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 82826 552134
rect 83062 551898 83146 552134
rect 83382 551898 118826 552134
rect 119062 551898 119146 552134
rect 119382 551898 154826 552134
rect 155062 551898 155146 552134
rect 155382 551898 190826 552134
rect 191062 551898 191146 552134
rect 191382 551898 226826 552134
rect 227062 551898 227146 552134
rect 227382 551898 262826 552134
rect 263062 551898 263146 552134
rect 263382 551898 298826 552134
rect 299062 551898 299146 552134
rect 299382 551898 334826 552134
rect 335062 551898 335146 552134
rect 335382 551898 370826 552134
rect 371062 551898 371146 552134
rect 371382 551898 406826 552134
rect 407062 551898 407146 552134
rect 407382 551898 442826 552134
rect 443062 551898 443146 552134
rect 443382 551898 478826 552134
rect 479062 551898 479146 552134
rect 479382 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 592650 552134
rect -8726 551866 592650 551898
rect -8726 547954 592650 547986
rect -8726 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 78326 547954
rect 78562 547718 78646 547954
rect 78882 547718 114326 547954
rect 114562 547718 114646 547954
rect 114882 547718 150326 547954
rect 150562 547718 150646 547954
rect 150882 547718 186326 547954
rect 186562 547718 186646 547954
rect 186882 547718 222326 547954
rect 222562 547718 222646 547954
rect 222882 547718 258326 547954
rect 258562 547718 258646 547954
rect 258882 547718 294326 547954
rect 294562 547718 294646 547954
rect 294882 547718 330326 547954
rect 330562 547718 330646 547954
rect 330882 547718 366326 547954
rect 366562 547718 366646 547954
rect 366882 547718 402326 547954
rect 402562 547718 402646 547954
rect 402882 547718 438326 547954
rect 438562 547718 438646 547954
rect 438882 547718 474326 547954
rect 474562 547718 474646 547954
rect 474882 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 592650 547954
rect -8726 547634 592650 547718
rect -8726 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 78326 547634
rect 78562 547398 78646 547634
rect 78882 547398 114326 547634
rect 114562 547398 114646 547634
rect 114882 547398 150326 547634
rect 150562 547398 150646 547634
rect 150882 547398 186326 547634
rect 186562 547398 186646 547634
rect 186882 547398 222326 547634
rect 222562 547398 222646 547634
rect 222882 547398 258326 547634
rect 258562 547398 258646 547634
rect 258882 547398 294326 547634
rect 294562 547398 294646 547634
rect 294882 547398 330326 547634
rect 330562 547398 330646 547634
rect 330882 547398 366326 547634
rect 366562 547398 366646 547634
rect 366882 547398 402326 547634
rect 402562 547398 402646 547634
rect 402882 547398 438326 547634
rect 438562 547398 438646 547634
rect 438882 547398 474326 547634
rect 474562 547398 474646 547634
rect 474882 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 592650 547634
rect -8726 547366 592650 547398
rect -8726 543454 592650 543486
rect -8726 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 592650 543454
rect -8726 543134 592650 543218
rect -8726 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 592650 543134
rect -8726 542866 592650 542898
rect -8726 538954 592650 538986
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 69326 538954
rect 69562 538718 69646 538954
rect 69882 538718 105326 538954
rect 105562 538718 105646 538954
rect 105882 538718 141326 538954
rect 141562 538718 141646 538954
rect 141882 538718 177326 538954
rect 177562 538718 177646 538954
rect 177882 538718 213326 538954
rect 213562 538718 213646 538954
rect 213882 538718 249326 538954
rect 249562 538718 249646 538954
rect 249882 538718 285326 538954
rect 285562 538718 285646 538954
rect 285882 538718 321326 538954
rect 321562 538718 321646 538954
rect 321882 538718 357326 538954
rect 357562 538718 357646 538954
rect 357882 538718 393326 538954
rect 393562 538718 393646 538954
rect 393882 538718 429326 538954
rect 429562 538718 429646 538954
rect 429882 538718 465326 538954
rect 465562 538718 465646 538954
rect 465882 538718 501326 538954
rect 501562 538718 501646 538954
rect 501882 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect -8726 538634 592650 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 69326 538634
rect 69562 538398 69646 538634
rect 69882 538398 105326 538634
rect 105562 538398 105646 538634
rect 105882 538398 141326 538634
rect 141562 538398 141646 538634
rect 141882 538398 177326 538634
rect 177562 538398 177646 538634
rect 177882 538398 213326 538634
rect 213562 538398 213646 538634
rect 213882 538398 249326 538634
rect 249562 538398 249646 538634
rect 249882 538398 285326 538634
rect 285562 538398 285646 538634
rect 285882 538398 321326 538634
rect 321562 538398 321646 538634
rect 321882 538398 357326 538634
rect 357562 538398 357646 538634
rect 357882 538398 393326 538634
rect 393562 538398 393646 538634
rect 393882 538398 429326 538634
rect 429562 538398 429646 538634
rect 429882 538398 465326 538634
rect 465562 538398 465646 538634
rect 465882 538398 501326 538634
rect 501562 538398 501646 538634
rect 501882 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect -8726 538366 592650 538398
rect -8726 534454 592650 534486
rect -8726 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 64826 534454
rect 65062 534218 65146 534454
rect 65382 534218 100826 534454
rect 101062 534218 101146 534454
rect 101382 534218 136826 534454
rect 137062 534218 137146 534454
rect 137382 534218 172826 534454
rect 173062 534218 173146 534454
rect 173382 534218 208826 534454
rect 209062 534218 209146 534454
rect 209382 534218 244826 534454
rect 245062 534218 245146 534454
rect 245382 534218 280826 534454
rect 281062 534218 281146 534454
rect 281382 534218 316826 534454
rect 317062 534218 317146 534454
rect 317382 534218 352826 534454
rect 353062 534218 353146 534454
rect 353382 534218 388826 534454
rect 389062 534218 389146 534454
rect 389382 534218 424826 534454
rect 425062 534218 425146 534454
rect 425382 534218 460826 534454
rect 461062 534218 461146 534454
rect 461382 534218 496826 534454
rect 497062 534218 497146 534454
rect 497382 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 592650 534454
rect -8726 534134 592650 534218
rect -8726 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 64826 534134
rect 65062 533898 65146 534134
rect 65382 533898 100826 534134
rect 101062 533898 101146 534134
rect 101382 533898 136826 534134
rect 137062 533898 137146 534134
rect 137382 533898 172826 534134
rect 173062 533898 173146 534134
rect 173382 533898 208826 534134
rect 209062 533898 209146 534134
rect 209382 533898 244826 534134
rect 245062 533898 245146 534134
rect 245382 533898 280826 534134
rect 281062 533898 281146 534134
rect 281382 533898 316826 534134
rect 317062 533898 317146 534134
rect 317382 533898 352826 534134
rect 353062 533898 353146 534134
rect 353382 533898 388826 534134
rect 389062 533898 389146 534134
rect 389382 533898 424826 534134
rect 425062 533898 425146 534134
rect 425382 533898 460826 534134
rect 461062 533898 461146 534134
rect 461382 533898 496826 534134
rect 497062 533898 497146 534134
rect 497382 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 592650 534134
rect -8726 533866 592650 533898
rect -8726 529954 592650 529986
rect -8726 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 60326 529954
rect 60562 529718 60646 529954
rect 60882 529718 96326 529954
rect 96562 529718 96646 529954
rect 96882 529718 132326 529954
rect 132562 529718 132646 529954
rect 132882 529718 168326 529954
rect 168562 529718 168646 529954
rect 168882 529718 204326 529954
rect 204562 529718 204646 529954
rect 204882 529718 240326 529954
rect 240562 529718 240646 529954
rect 240882 529718 276326 529954
rect 276562 529718 276646 529954
rect 276882 529718 312326 529954
rect 312562 529718 312646 529954
rect 312882 529718 348326 529954
rect 348562 529718 348646 529954
rect 348882 529718 384326 529954
rect 384562 529718 384646 529954
rect 384882 529718 420326 529954
rect 420562 529718 420646 529954
rect 420882 529718 456326 529954
rect 456562 529718 456646 529954
rect 456882 529718 492326 529954
rect 492562 529718 492646 529954
rect 492882 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 592650 529954
rect -8726 529634 592650 529718
rect -8726 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 60326 529634
rect 60562 529398 60646 529634
rect 60882 529398 96326 529634
rect 96562 529398 96646 529634
rect 96882 529398 132326 529634
rect 132562 529398 132646 529634
rect 132882 529398 168326 529634
rect 168562 529398 168646 529634
rect 168882 529398 204326 529634
rect 204562 529398 204646 529634
rect 204882 529398 240326 529634
rect 240562 529398 240646 529634
rect 240882 529398 276326 529634
rect 276562 529398 276646 529634
rect 276882 529398 312326 529634
rect 312562 529398 312646 529634
rect 312882 529398 348326 529634
rect 348562 529398 348646 529634
rect 348882 529398 384326 529634
rect 384562 529398 384646 529634
rect 384882 529398 420326 529634
rect 420562 529398 420646 529634
rect 420882 529398 456326 529634
rect 456562 529398 456646 529634
rect 456882 529398 492326 529634
rect 492562 529398 492646 529634
rect 492882 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 592650 529634
rect -8726 529366 592650 529398
rect -8726 525454 592650 525486
rect -8726 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 592650 525454
rect -8726 525134 592650 525218
rect -8726 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 592650 525134
rect -8726 524866 592650 524898
rect -8726 520954 592650 520986
rect -8726 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 51326 520954
rect 51562 520718 51646 520954
rect 51882 520718 87326 520954
rect 87562 520718 87646 520954
rect 87882 520718 123326 520954
rect 123562 520718 123646 520954
rect 123882 520718 159326 520954
rect 159562 520718 159646 520954
rect 159882 520718 195326 520954
rect 195562 520718 195646 520954
rect 195882 520718 231326 520954
rect 231562 520718 231646 520954
rect 231882 520718 267326 520954
rect 267562 520718 267646 520954
rect 267882 520718 303326 520954
rect 303562 520718 303646 520954
rect 303882 520718 339326 520954
rect 339562 520718 339646 520954
rect 339882 520718 375326 520954
rect 375562 520718 375646 520954
rect 375882 520718 411326 520954
rect 411562 520718 411646 520954
rect 411882 520718 447326 520954
rect 447562 520718 447646 520954
rect 447882 520718 483326 520954
rect 483562 520718 483646 520954
rect 483882 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 592650 520954
rect -8726 520634 592650 520718
rect -8726 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 51326 520634
rect 51562 520398 51646 520634
rect 51882 520398 87326 520634
rect 87562 520398 87646 520634
rect 87882 520398 123326 520634
rect 123562 520398 123646 520634
rect 123882 520398 159326 520634
rect 159562 520398 159646 520634
rect 159882 520398 195326 520634
rect 195562 520398 195646 520634
rect 195882 520398 231326 520634
rect 231562 520398 231646 520634
rect 231882 520398 267326 520634
rect 267562 520398 267646 520634
rect 267882 520398 303326 520634
rect 303562 520398 303646 520634
rect 303882 520398 339326 520634
rect 339562 520398 339646 520634
rect 339882 520398 375326 520634
rect 375562 520398 375646 520634
rect 375882 520398 411326 520634
rect 411562 520398 411646 520634
rect 411882 520398 447326 520634
rect 447562 520398 447646 520634
rect 447882 520398 483326 520634
rect 483562 520398 483646 520634
rect 483882 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 592650 520634
rect -8726 520366 592650 520398
rect -8726 516454 592650 516486
rect -8726 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 82826 516454
rect 83062 516218 83146 516454
rect 83382 516218 118826 516454
rect 119062 516218 119146 516454
rect 119382 516218 154826 516454
rect 155062 516218 155146 516454
rect 155382 516218 190826 516454
rect 191062 516218 191146 516454
rect 191382 516218 226826 516454
rect 227062 516218 227146 516454
rect 227382 516218 262826 516454
rect 263062 516218 263146 516454
rect 263382 516218 298826 516454
rect 299062 516218 299146 516454
rect 299382 516218 334826 516454
rect 335062 516218 335146 516454
rect 335382 516218 370826 516454
rect 371062 516218 371146 516454
rect 371382 516218 406826 516454
rect 407062 516218 407146 516454
rect 407382 516218 442826 516454
rect 443062 516218 443146 516454
rect 443382 516218 478826 516454
rect 479062 516218 479146 516454
rect 479382 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 592650 516454
rect -8726 516134 592650 516218
rect -8726 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 82826 516134
rect 83062 515898 83146 516134
rect 83382 515898 118826 516134
rect 119062 515898 119146 516134
rect 119382 515898 154826 516134
rect 155062 515898 155146 516134
rect 155382 515898 190826 516134
rect 191062 515898 191146 516134
rect 191382 515898 226826 516134
rect 227062 515898 227146 516134
rect 227382 515898 262826 516134
rect 263062 515898 263146 516134
rect 263382 515898 298826 516134
rect 299062 515898 299146 516134
rect 299382 515898 334826 516134
rect 335062 515898 335146 516134
rect 335382 515898 370826 516134
rect 371062 515898 371146 516134
rect 371382 515898 406826 516134
rect 407062 515898 407146 516134
rect 407382 515898 442826 516134
rect 443062 515898 443146 516134
rect 443382 515898 478826 516134
rect 479062 515898 479146 516134
rect 479382 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 592650 516134
rect -8726 515866 592650 515898
rect -8726 511954 592650 511986
rect -8726 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 78326 511954
rect 78562 511718 78646 511954
rect 78882 511718 114326 511954
rect 114562 511718 114646 511954
rect 114882 511718 150326 511954
rect 150562 511718 150646 511954
rect 150882 511718 186326 511954
rect 186562 511718 186646 511954
rect 186882 511718 222326 511954
rect 222562 511718 222646 511954
rect 222882 511718 258326 511954
rect 258562 511718 258646 511954
rect 258882 511718 294326 511954
rect 294562 511718 294646 511954
rect 294882 511718 330326 511954
rect 330562 511718 330646 511954
rect 330882 511718 366326 511954
rect 366562 511718 366646 511954
rect 366882 511718 402326 511954
rect 402562 511718 402646 511954
rect 402882 511718 438326 511954
rect 438562 511718 438646 511954
rect 438882 511718 474326 511954
rect 474562 511718 474646 511954
rect 474882 511718 510326 511954
rect 510562 511718 510646 511954
rect 510882 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 592650 511954
rect -8726 511634 592650 511718
rect -8726 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 78326 511634
rect 78562 511398 78646 511634
rect 78882 511398 114326 511634
rect 114562 511398 114646 511634
rect 114882 511398 150326 511634
rect 150562 511398 150646 511634
rect 150882 511398 186326 511634
rect 186562 511398 186646 511634
rect 186882 511398 222326 511634
rect 222562 511398 222646 511634
rect 222882 511398 258326 511634
rect 258562 511398 258646 511634
rect 258882 511398 294326 511634
rect 294562 511398 294646 511634
rect 294882 511398 330326 511634
rect 330562 511398 330646 511634
rect 330882 511398 366326 511634
rect 366562 511398 366646 511634
rect 366882 511398 402326 511634
rect 402562 511398 402646 511634
rect 402882 511398 438326 511634
rect 438562 511398 438646 511634
rect 438882 511398 474326 511634
rect 474562 511398 474646 511634
rect 474882 511398 510326 511634
rect 510562 511398 510646 511634
rect 510882 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 592650 511634
rect -8726 511366 592650 511398
rect -8726 507454 592650 507486
rect -8726 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 592650 507454
rect -8726 507134 592650 507218
rect -8726 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 592650 507134
rect -8726 506866 592650 506898
rect -8726 502954 592650 502986
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 69326 502954
rect 69562 502718 69646 502954
rect 69882 502718 105326 502954
rect 105562 502718 105646 502954
rect 105882 502718 141326 502954
rect 141562 502718 141646 502954
rect 141882 502718 177326 502954
rect 177562 502718 177646 502954
rect 177882 502718 213326 502954
rect 213562 502718 213646 502954
rect 213882 502718 249326 502954
rect 249562 502718 249646 502954
rect 249882 502718 285326 502954
rect 285562 502718 285646 502954
rect 285882 502718 321326 502954
rect 321562 502718 321646 502954
rect 321882 502718 357326 502954
rect 357562 502718 357646 502954
rect 357882 502718 393326 502954
rect 393562 502718 393646 502954
rect 393882 502718 429326 502954
rect 429562 502718 429646 502954
rect 429882 502718 465326 502954
rect 465562 502718 465646 502954
rect 465882 502718 501326 502954
rect 501562 502718 501646 502954
rect 501882 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect -8726 502634 592650 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 69326 502634
rect 69562 502398 69646 502634
rect 69882 502398 105326 502634
rect 105562 502398 105646 502634
rect 105882 502398 141326 502634
rect 141562 502398 141646 502634
rect 141882 502398 177326 502634
rect 177562 502398 177646 502634
rect 177882 502398 213326 502634
rect 213562 502398 213646 502634
rect 213882 502398 249326 502634
rect 249562 502398 249646 502634
rect 249882 502398 285326 502634
rect 285562 502398 285646 502634
rect 285882 502398 321326 502634
rect 321562 502398 321646 502634
rect 321882 502398 357326 502634
rect 357562 502398 357646 502634
rect 357882 502398 393326 502634
rect 393562 502398 393646 502634
rect 393882 502398 429326 502634
rect 429562 502398 429646 502634
rect 429882 502398 465326 502634
rect 465562 502398 465646 502634
rect 465882 502398 501326 502634
rect 501562 502398 501646 502634
rect 501882 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect -8726 502366 592650 502398
rect -8726 498454 592650 498486
rect -8726 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 64826 498454
rect 65062 498218 65146 498454
rect 65382 498218 100826 498454
rect 101062 498218 101146 498454
rect 101382 498218 136826 498454
rect 137062 498218 137146 498454
rect 137382 498218 172826 498454
rect 173062 498218 173146 498454
rect 173382 498218 208826 498454
rect 209062 498218 209146 498454
rect 209382 498218 244826 498454
rect 245062 498218 245146 498454
rect 245382 498218 280826 498454
rect 281062 498218 281146 498454
rect 281382 498218 316826 498454
rect 317062 498218 317146 498454
rect 317382 498218 352826 498454
rect 353062 498218 353146 498454
rect 353382 498218 388826 498454
rect 389062 498218 389146 498454
rect 389382 498218 424826 498454
rect 425062 498218 425146 498454
rect 425382 498218 460826 498454
rect 461062 498218 461146 498454
rect 461382 498218 496826 498454
rect 497062 498218 497146 498454
rect 497382 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 592650 498454
rect -8726 498134 592650 498218
rect -8726 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 64826 498134
rect 65062 497898 65146 498134
rect 65382 497898 100826 498134
rect 101062 497898 101146 498134
rect 101382 497898 136826 498134
rect 137062 497898 137146 498134
rect 137382 497898 172826 498134
rect 173062 497898 173146 498134
rect 173382 497898 208826 498134
rect 209062 497898 209146 498134
rect 209382 497898 244826 498134
rect 245062 497898 245146 498134
rect 245382 497898 280826 498134
rect 281062 497898 281146 498134
rect 281382 497898 316826 498134
rect 317062 497898 317146 498134
rect 317382 497898 352826 498134
rect 353062 497898 353146 498134
rect 353382 497898 388826 498134
rect 389062 497898 389146 498134
rect 389382 497898 424826 498134
rect 425062 497898 425146 498134
rect 425382 497898 460826 498134
rect 461062 497898 461146 498134
rect 461382 497898 496826 498134
rect 497062 497898 497146 498134
rect 497382 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 592650 498134
rect -8726 497866 592650 497898
rect -8726 493954 592650 493986
rect -8726 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 60326 493954
rect 60562 493718 60646 493954
rect 60882 493718 96326 493954
rect 96562 493718 96646 493954
rect 96882 493718 132326 493954
rect 132562 493718 132646 493954
rect 132882 493718 168326 493954
rect 168562 493718 168646 493954
rect 168882 493718 204326 493954
rect 204562 493718 204646 493954
rect 204882 493718 240326 493954
rect 240562 493718 240646 493954
rect 240882 493718 276326 493954
rect 276562 493718 276646 493954
rect 276882 493718 312326 493954
rect 312562 493718 312646 493954
rect 312882 493718 348326 493954
rect 348562 493718 348646 493954
rect 348882 493718 384326 493954
rect 384562 493718 384646 493954
rect 384882 493718 420326 493954
rect 420562 493718 420646 493954
rect 420882 493718 456326 493954
rect 456562 493718 456646 493954
rect 456882 493718 492326 493954
rect 492562 493718 492646 493954
rect 492882 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 592650 493954
rect -8726 493634 592650 493718
rect -8726 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 60326 493634
rect 60562 493398 60646 493634
rect 60882 493398 96326 493634
rect 96562 493398 96646 493634
rect 96882 493398 132326 493634
rect 132562 493398 132646 493634
rect 132882 493398 168326 493634
rect 168562 493398 168646 493634
rect 168882 493398 204326 493634
rect 204562 493398 204646 493634
rect 204882 493398 240326 493634
rect 240562 493398 240646 493634
rect 240882 493398 276326 493634
rect 276562 493398 276646 493634
rect 276882 493398 312326 493634
rect 312562 493398 312646 493634
rect 312882 493398 348326 493634
rect 348562 493398 348646 493634
rect 348882 493398 384326 493634
rect 384562 493398 384646 493634
rect 384882 493398 420326 493634
rect 420562 493398 420646 493634
rect 420882 493398 456326 493634
rect 456562 493398 456646 493634
rect 456882 493398 492326 493634
rect 492562 493398 492646 493634
rect 492882 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 592650 493634
rect -8726 493366 592650 493398
rect -8726 489454 592650 489486
rect -8726 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 592650 489454
rect -8726 489134 592650 489218
rect -8726 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 592650 489134
rect -8726 488866 592650 488898
rect -8726 484954 592650 484986
rect -8726 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 51326 484954
rect 51562 484718 51646 484954
rect 51882 484718 87326 484954
rect 87562 484718 87646 484954
rect 87882 484718 123326 484954
rect 123562 484718 123646 484954
rect 123882 484718 159326 484954
rect 159562 484718 159646 484954
rect 159882 484718 195326 484954
rect 195562 484718 195646 484954
rect 195882 484718 231326 484954
rect 231562 484718 231646 484954
rect 231882 484718 267326 484954
rect 267562 484718 267646 484954
rect 267882 484718 303326 484954
rect 303562 484718 303646 484954
rect 303882 484718 339326 484954
rect 339562 484718 339646 484954
rect 339882 484718 375326 484954
rect 375562 484718 375646 484954
rect 375882 484718 411326 484954
rect 411562 484718 411646 484954
rect 411882 484718 447326 484954
rect 447562 484718 447646 484954
rect 447882 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 592650 484954
rect -8726 484634 592650 484718
rect -8726 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 51326 484634
rect 51562 484398 51646 484634
rect 51882 484398 87326 484634
rect 87562 484398 87646 484634
rect 87882 484398 123326 484634
rect 123562 484398 123646 484634
rect 123882 484398 159326 484634
rect 159562 484398 159646 484634
rect 159882 484398 195326 484634
rect 195562 484398 195646 484634
rect 195882 484398 231326 484634
rect 231562 484398 231646 484634
rect 231882 484398 267326 484634
rect 267562 484398 267646 484634
rect 267882 484398 303326 484634
rect 303562 484398 303646 484634
rect 303882 484398 339326 484634
rect 339562 484398 339646 484634
rect 339882 484398 375326 484634
rect 375562 484398 375646 484634
rect 375882 484398 411326 484634
rect 411562 484398 411646 484634
rect 411882 484398 447326 484634
rect 447562 484398 447646 484634
rect 447882 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 592650 484634
rect -8726 484366 592650 484398
rect -8726 480454 592650 480486
rect -8726 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 82826 480454
rect 83062 480218 83146 480454
rect 83382 480218 118826 480454
rect 119062 480218 119146 480454
rect 119382 480218 154826 480454
rect 155062 480218 155146 480454
rect 155382 480218 190826 480454
rect 191062 480218 191146 480454
rect 191382 480218 226826 480454
rect 227062 480218 227146 480454
rect 227382 480218 262826 480454
rect 263062 480218 263146 480454
rect 263382 480218 298826 480454
rect 299062 480218 299146 480454
rect 299382 480218 334826 480454
rect 335062 480218 335146 480454
rect 335382 480218 370826 480454
rect 371062 480218 371146 480454
rect 371382 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 442826 480454
rect 443062 480218 443146 480454
rect 443382 480218 478826 480454
rect 479062 480218 479146 480454
rect 479382 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 592650 480454
rect -8726 480134 592650 480218
rect -8726 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 82826 480134
rect 83062 479898 83146 480134
rect 83382 479898 118826 480134
rect 119062 479898 119146 480134
rect 119382 479898 154826 480134
rect 155062 479898 155146 480134
rect 155382 479898 190826 480134
rect 191062 479898 191146 480134
rect 191382 479898 226826 480134
rect 227062 479898 227146 480134
rect 227382 479898 262826 480134
rect 263062 479898 263146 480134
rect 263382 479898 298826 480134
rect 299062 479898 299146 480134
rect 299382 479898 334826 480134
rect 335062 479898 335146 480134
rect 335382 479898 370826 480134
rect 371062 479898 371146 480134
rect 371382 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 442826 480134
rect 443062 479898 443146 480134
rect 443382 479898 478826 480134
rect 479062 479898 479146 480134
rect 479382 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 592650 480134
rect -8726 479866 592650 479898
rect -8726 475954 592650 475986
rect -8726 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 78326 475954
rect 78562 475718 78646 475954
rect 78882 475718 114326 475954
rect 114562 475718 114646 475954
rect 114882 475718 150326 475954
rect 150562 475718 150646 475954
rect 150882 475718 186326 475954
rect 186562 475718 186646 475954
rect 186882 475718 222326 475954
rect 222562 475718 222646 475954
rect 222882 475718 258326 475954
rect 258562 475718 258646 475954
rect 258882 475718 294326 475954
rect 294562 475718 294646 475954
rect 294882 475718 330326 475954
rect 330562 475718 330646 475954
rect 330882 475718 366326 475954
rect 366562 475718 366646 475954
rect 366882 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 438326 475954
rect 438562 475718 438646 475954
rect 438882 475718 474326 475954
rect 474562 475718 474646 475954
rect 474882 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 592650 475954
rect -8726 475634 592650 475718
rect -8726 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 78326 475634
rect 78562 475398 78646 475634
rect 78882 475398 114326 475634
rect 114562 475398 114646 475634
rect 114882 475398 150326 475634
rect 150562 475398 150646 475634
rect 150882 475398 186326 475634
rect 186562 475398 186646 475634
rect 186882 475398 222326 475634
rect 222562 475398 222646 475634
rect 222882 475398 258326 475634
rect 258562 475398 258646 475634
rect 258882 475398 294326 475634
rect 294562 475398 294646 475634
rect 294882 475398 330326 475634
rect 330562 475398 330646 475634
rect 330882 475398 366326 475634
rect 366562 475398 366646 475634
rect 366882 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 438326 475634
rect 438562 475398 438646 475634
rect 438882 475398 474326 475634
rect 474562 475398 474646 475634
rect 474882 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 592650 475634
rect -8726 475366 592650 475398
rect -8726 471454 592650 471486
rect -8726 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 592650 471454
rect -8726 471134 592650 471218
rect -8726 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 592650 471134
rect -8726 470866 592650 470898
rect -8726 466954 592650 466986
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 69326 466954
rect 69562 466718 69646 466954
rect 69882 466718 105326 466954
rect 105562 466718 105646 466954
rect 105882 466718 141326 466954
rect 141562 466718 141646 466954
rect 141882 466718 177326 466954
rect 177562 466718 177646 466954
rect 177882 466718 213326 466954
rect 213562 466718 213646 466954
rect 213882 466718 249326 466954
rect 249562 466718 249646 466954
rect 249882 466718 285326 466954
rect 285562 466718 285646 466954
rect 285882 466718 321326 466954
rect 321562 466718 321646 466954
rect 321882 466718 357326 466954
rect 357562 466718 357646 466954
rect 357882 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 429326 466954
rect 429562 466718 429646 466954
rect 429882 466718 465326 466954
rect 465562 466718 465646 466954
rect 465882 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect -8726 466634 592650 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 69326 466634
rect 69562 466398 69646 466634
rect 69882 466398 105326 466634
rect 105562 466398 105646 466634
rect 105882 466398 141326 466634
rect 141562 466398 141646 466634
rect 141882 466398 177326 466634
rect 177562 466398 177646 466634
rect 177882 466398 213326 466634
rect 213562 466398 213646 466634
rect 213882 466398 249326 466634
rect 249562 466398 249646 466634
rect 249882 466398 285326 466634
rect 285562 466398 285646 466634
rect 285882 466398 321326 466634
rect 321562 466398 321646 466634
rect 321882 466398 357326 466634
rect 357562 466398 357646 466634
rect 357882 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 429326 466634
rect 429562 466398 429646 466634
rect 429882 466398 465326 466634
rect 465562 466398 465646 466634
rect 465882 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect -8726 466366 592650 466398
rect -8726 462454 592650 462486
rect -8726 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 64826 462454
rect 65062 462218 65146 462454
rect 65382 462218 100826 462454
rect 101062 462218 101146 462454
rect 101382 462218 136826 462454
rect 137062 462218 137146 462454
rect 137382 462218 172826 462454
rect 173062 462218 173146 462454
rect 173382 462218 208826 462454
rect 209062 462218 209146 462454
rect 209382 462218 244826 462454
rect 245062 462218 245146 462454
rect 245382 462218 280826 462454
rect 281062 462218 281146 462454
rect 281382 462218 316826 462454
rect 317062 462218 317146 462454
rect 317382 462218 352826 462454
rect 353062 462218 353146 462454
rect 353382 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 424826 462454
rect 425062 462218 425146 462454
rect 425382 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 592650 462454
rect -8726 462134 592650 462218
rect -8726 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 64826 462134
rect 65062 461898 65146 462134
rect 65382 461898 100826 462134
rect 101062 461898 101146 462134
rect 101382 461898 136826 462134
rect 137062 461898 137146 462134
rect 137382 461898 172826 462134
rect 173062 461898 173146 462134
rect 173382 461898 208826 462134
rect 209062 461898 209146 462134
rect 209382 461898 244826 462134
rect 245062 461898 245146 462134
rect 245382 461898 280826 462134
rect 281062 461898 281146 462134
rect 281382 461898 316826 462134
rect 317062 461898 317146 462134
rect 317382 461898 352826 462134
rect 353062 461898 353146 462134
rect 353382 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 424826 462134
rect 425062 461898 425146 462134
rect 425382 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 592650 462134
rect -8726 461866 592650 461898
rect -8726 457954 592650 457986
rect -8726 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 60326 457954
rect 60562 457718 60646 457954
rect 60882 457718 96326 457954
rect 96562 457718 96646 457954
rect 96882 457718 132326 457954
rect 132562 457718 132646 457954
rect 132882 457718 168326 457954
rect 168562 457718 168646 457954
rect 168882 457718 204326 457954
rect 204562 457718 204646 457954
rect 204882 457718 240326 457954
rect 240562 457718 240646 457954
rect 240882 457718 276326 457954
rect 276562 457718 276646 457954
rect 276882 457718 312326 457954
rect 312562 457718 312646 457954
rect 312882 457718 348326 457954
rect 348562 457718 348646 457954
rect 348882 457718 384326 457954
rect 384562 457718 384646 457954
rect 384882 457718 420326 457954
rect 420562 457718 420646 457954
rect 420882 457718 456326 457954
rect 456562 457718 456646 457954
rect 456882 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 592650 457954
rect -8726 457634 592650 457718
rect -8726 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 60326 457634
rect 60562 457398 60646 457634
rect 60882 457398 96326 457634
rect 96562 457398 96646 457634
rect 96882 457398 132326 457634
rect 132562 457398 132646 457634
rect 132882 457398 168326 457634
rect 168562 457398 168646 457634
rect 168882 457398 204326 457634
rect 204562 457398 204646 457634
rect 204882 457398 240326 457634
rect 240562 457398 240646 457634
rect 240882 457398 276326 457634
rect 276562 457398 276646 457634
rect 276882 457398 312326 457634
rect 312562 457398 312646 457634
rect 312882 457398 348326 457634
rect 348562 457398 348646 457634
rect 348882 457398 384326 457634
rect 384562 457398 384646 457634
rect 384882 457398 420326 457634
rect 420562 457398 420646 457634
rect 420882 457398 456326 457634
rect 456562 457398 456646 457634
rect 456882 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 592650 457634
rect -8726 457366 592650 457398
rect -8726 453454 592650 453486
rect -8726 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 592650 453454
rect -8726 453134 592650 453218
rect -8726 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 592650 453134
rect -8726 452866 592650 452898
rect -8726 448954 592650 448986
rect -8726 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 51326 448954
rect 51562 448718 51646 448954
rect 51882 448718 87326 448954
rect 87562 448718 87646 448954
rect 87882 448718 123326 448954
rect 123562 448718 123646 448954
rect 123882 448718 159326 448954
rect 159562 448718 159646 448954
rect 159882 448718 195326 448954
rect 195562 448718 195646 448954
rect 195882 448718 231326 448954
rect 231562 448718 231646 448954
rect 231882 448718 267326 448954
rect 267562 448718 267646 448954
rect 267882 448718 303326 448954
rect 303562 448718 303646 448954
rect 303882 448718 339326 448954
rect 339562 448718 339646 448954
rect 339882 448718 375326 448954
rect 375562 448718 375646 448954
rect 375882 448718 411326 448954
rect 411562 448718 411646 448954
rect 411882 448718 447326 448954
rect 447562 448718 447646 448954
rect 447882 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 592650 448954
rect -8726 448634 592650 448718
rect -8726 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 51326 448634
rect 51562 448398 51646 448634
rect 51882 448398 87326 448634
rect 87562 448398 87646 448634
rect 87882 448398 123326 448634
rect 123562 448398 123646 448634
rect 123882 448398 159326 448634
rect 159562 448398 159646 448634
rect 159882 448398 195326 448634
rect 195562 448398 195646 448634
rect 195882 448398 231326 448634
rect 231562 448398 231646 448634
rect 231882 448398 267326 448634
rect 267562 448398 267646 448634
rect 267882 448398 303326 448634
rect 303562 448398 303646 448634
rect 303882 448398 339326 448634
rect 339562 448398 339646 448634
rect 339882 448398 375326 448634
rect 375562 448398 375646 448634
rect 375882 448398 411326 448634
rect 411562 448398 411646 448634
rect 411882 448398 447326 448634
rect 447562 448398 447646 448634
rect 447882 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 592650 448634
rect -8726 448366 592650 448398
rect -8726 444454 592650 444486
rect -8726 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 82826 444454
rect 83062 444218 83146 444454
rect 83382 444218 118826 444454
rect 119062 444218 119146 444454
rect 119382 444218 154826 444454
rect 155062 444218 155146 444454
rect 155382 444218 190826 444454
rect 191062 444218 191146 444454
rect 191382 444218 226826 444454
rect 227062 444218 227146 444454
rect 227382 444218 262826 444454
rect 263062 444218 263146 444454
rect 263382 444218 298826 444454
rect 299062 444218 299146 444454
rect 299382 444218 334826 444454
rect 335062 444218 335146 444454
rect 335382 444218 370826 444454
rect 371062 444218 371146 444454
rect 371382 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 592650 444454
rect -8726 444134 592650 444218
rect -8726 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 82826 444134
rect 83062 443898 83146 444134
rect 83382 443898 118826 444134
rect 119062 443898 119146 444134
rect 119382 443898 154826 444134
rect 155062 443898 155146 444134
rect 155382 443898 190826 444134
rect 191062 443898 191146 444134
rect 191382 443898 226826 444134
rect 227062 443898 227146 444134
rect 227382 443898 262826 444134
rect 263062 443898 263146 444134
rect 263382 443898 298826 444134
rect 299062 443898 299146 444134
rect 299382 443898 334826 444134
rect 335062 443898 335146 444134
rect 335382 443898 370826 444134
rect 371062 443898 371146 444134
rect 371382 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 592650 444134
rect -8726 443866 592650 443898
rect -8726 439954 592650 439986
rect -8726 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 78326 439954
rect 78562 439718 78646 439954
rect 78882 439718 114326 439954
rect 114562 439718 114646 439954
rect 114882 439718 150326 439954
rect 150562 439718 150646 439954
rect 150882 439718 186326 439954
rect 186562 439718 186646 439954
rect 186882 439718 222326 439954
rect 222562 439718 222646 439954
rect 222882 439718 258326 439954
rect 258562 439718 258646 439954
rect 258882 439718 294326 439954
rect 294562 439718 294646 439954
rect 294882 439718 330326 439954
rect 330562 439718 330646 439954
rect 330882 439718 366326 439954
rect 366562 439718 366646 439954
rect 366882 439718 402326 439954
rect 402562 439718 402646 439954
rect 402882 439718 438326 439954
rect 438562 439718 438646 439954
rect 438882 439718 474326 439954
rect 474562 439718 474646 439954
rect 474882 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 592650 439954
rect -8726 439634 592650 439718
rect -8726 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 78326 439634
rect 78562 439398 78646 439634
rect 78882 439398 114326 439634
rect 114562 439398 114646 439634
rect 114882 439398 150326 439634
rect 150562 439398 150646 439634
rect 150882 439398 186326 439634
rect 186562 439398 186646 439634
rect 186882 439398 222326 439634
rect 222562 439398 222646 439634
rect 222882 439398 258326 439634
rect 258562 439398 258646 439634
rect 258882 439398 294326 439634
rect 294562 439398 294646 439634
rect 294882 439398 330326 439634
rect 330562 439398 330646 439634
rect 330882 439398 366326 439634
rect 366562 439398 366646 439634
rect 366882 439398 402326 439634
rect 402562 439398 402646 439634
rect 402882 439398 438326 439634
rect 438562 439398 438646 439634
rect 438882 439398 474326 439634
rect 474562 439398 474646 439634
rect 474882 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 592650 439634
rect -8726 439366 592650 439398
rect -8726 435454 592650 435486
rect -8726 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 592650 435454
rect -8726 435134 592650 435218
rect -8726 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 592650 435134
rect -8726 434866 592650 434898
rect -8726 430954 592650 430986
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 69326 430954
rect 69562 430718 69646 430954
rect 69882 430718 105326 430954
rect 105562 430718 105646 430954
rect 105882 430718 141326 430954
rect 141562 430718 141646 430954
rect 141882 430718 177326 430954
rect 177562 430718 177646 430954
rect 177882 430718 213326 430954
rect 213562 430718 213646 430954
rect 213882 430718 249326 430954
rect 249562 430718 249646 430954
rect 249882 430718 285326 430954
rect 285562 430718 285646 430954
rect 285882 430718 321326 430954
rect 321562 430718 321646 430954
rect 321882 430718 357326 430954
rect 357562 430718 357646 430954
rect 357882 430718 393326 430954
rect 393562 430718 393646 430954
rect 393882 430718 429326 430954
rect 429562 430718 429646 430954
rect 429882 430718 465326 430954
rect 465562 430718 465646 430954
rect 465882 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect -8726 430634 592650 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 69326 430634
rect 69562 430398 69646 430634
rect 69882 430398 105326 430634
rect 105562 430398 105646 430634
rect 105882 430398 141326 430634
rect 141562 430398 141646 430634
rect 141882 430398 177326 430634
rect 177562 430398 177646 430634
rect 177882 430398 213326 430634
rect 213562 430398 213646 430634
rect 213882 430398 249326 430634
rect 249562 430398 249646 430634
rect 249882 430398 285326 430634
rect 285562 430398 285646 430634
rect 285882 430398 321326 430634
rect 321562 430398 321646 430634
rect 321882 430398 357326 430634
rect 357562 430398 357646 430634
rect 357882 430398 393326 430634
rect 393562 430398 393646 430634
rect 393882 430398 429326 430634
rect 429562 430398 429646 430634
rect 429882 430398 465326 430634
rect 465562 430398 465646 430634
rect 465882 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect -8726 430366 592650 430398
rect -8726 426454 592650 426486
rect -8726 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 64826 426454
rect 65062 426218 65146 426454
rect 65382 426218 100826 426454
rect 101062 426218 101146 426454
rect 101382 426218 136826 426454
rect 137062 426218 137146 426454
rect 137382 426218 172826 426454
rect 173062 426218 173146 426454
rect 173382 426218 208826 426454
rect 209062 426218 209146 426454
rect 209382 426218 244826 426454
rect 245062 426218 245146 426454
rect 245382 426218 280826 426454
rect 281062 426218 281146 426454
rect 281382 426218 316826 426454
rect 317062 426218 317146 426454
rect 317382 426218 352826 426454
rect 353062 426218 353146 426454
rect 353382 426218 388826 426454
rect 389062 426218 389146 426454
rect 389382 426218 424826 426454
rect 425062 426218 425146 426454
rect 425382 426218 460826 426454
rect 461062 426218 461146 426454
rect 461382 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 592650 426454
rect -8726 426134 592650 426218
rect -8726 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 64826 426134
rect 65062 425898 65146 426134
rect 65382 425898 100826 426134
rect 101062 425898 101146 426134
rect 101382 425898 136826 426134
rect 137062 425898 137146 426134
rect 137382 425898 172826 426134
rect 173062 425898 173146 426134
rect 173382 425898 208826 426134
rect 209062 425898 209146 426134
rect 209382 425898 244826 426134
rect 245062 425898 245146 426134
rect 245382 425898 280826 426134
rect 281062 425898 281146 426134
rect 281382 425898 316826 426134
rect 317062 425898 317146 426134
rect 317382 425898 352826 426134
rect 353062 425898 353146 426134
rect 353382 425898 388826 426134
rect 389062 425898 389146 426134
rect 389382 425898 424826 426134
rect 425062 425898 425146 426134
rect 425382 425898 460826 426134
rect 461062 425898 461146 426134
rect 461382 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 592650 426134
rect -8726 425866 592650 425898
rect -8726 421954 592650 421986
rect -8726 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 60326 421954
rect 60562 421718 60646 421954
rect 60882 421718 96326 421954
rect 96562 421718 96646 421954
rect 96882 421718 132326 421954
rect 132562 421718 132646 421954
rect 132882 421718 168326 421954
rect 168562 421718 168646 421954
rect 168882 421718 204326 421954
rect 204562 421718 204646 421954
rect 204882 421718 240326 421954
rect 240562 421718 240646 421954
rect 240882 421718 276326 421954
rect 276562 421718 276646 421954
rect 276882 421718 312326 421954
rect 312562 421718 312646 421954
rect 312882 421718 348326 421954
rect 348562 421718 348646 421954
rect 348882 421718 384326 421954
rect 384562 421718 384646 421954
rect 384882 421718 420326 421954
rect 420562 421718 420646 421954
rect 420882 421718 456326 421954
rect 456562 421718 456646 421954
rect 456882 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 592650 421954
rect -8726 421634 592650 421718
rect -8726 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 60326 421634
rect 60562 421398 60646 421634
rect 60882 421398 96326 421634
rect 96562 421398 96646 421634
rect 96882 421398 132326 421634
rect 132562 421398 132646 421634
rect 132882 421398 168326 421634
rect 168562 421398 168646 421634
rect 168882 421398 204326 421634
rect 204562 421398 204646 421634
rect 204882 421398 240326 421634
rect 240562 421398 240646 421634
rect 240882 421398 276326 421634
rect 276562 421398 276646 421634
rect 276882 421398 312326 421634
rect 312562 421398 312646 421634
rect 312882 421398 348326 421634
rect 348562 421398 348646 421634
rect 348882 421398 384326 421634
rect 384562 421398 384646 421634
rect 384882 421398 420326 421634
rect 420562 421398 420646 421634
rect 420882 421398 456326 421634
rect 456562 421398 456646 421634
rect 456882 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 592650 421634
rect -8726 421366 592650 421398
rect -8726 417454 592650 417486
rect -8726 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 592650 417454
rect -8726 417134 592650 417218
rect -8726 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 592650 417134
rect -8726 416866 592650 416898
rect -8726 412954 592650 412986
rect -8726 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 51326 412954
rect 51562 412718 51646 412954
rect 51882 412718 87326 412954
rect 87562 412718 87646 412954
rect 87882 412718 123326 412954
rect 123562 412718 123646 412954
rect 123882 412718 159326 412954
rect 159562 412718 159646 412954
rect 159882 412718 195326 412954
rect 195562 412718 195646 412954
rect 195882 412718 231326 412954
rect 231562 412718 231646 412954
rect 231882 412718 267326 412954
rect 267562 412718 267646 412954
rect 267882 412718 303326 412954
rect 303562 412718 303646 412954
rect 303882 412718 339326 412954
rect 339562 412718 339646 412954
rect 339882 412718 375326 412954
rect 375562 412718 375646 412954
rect 375882 412718 411326 412954
rect 411562 412718 411646 412954
rect 411882 412718 447326 412954
rect 447562 412718 447646 412954
rect 447882 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 592650 412954
rect -8726 412634 592650 412718
rect -8726 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 51326 412634
rect 51562 412398 51646 412634
rect 51882 412398 87326 412634
rect 87562 412398 87646 412634
rect 87882 412398 123326 412634
rect 123562 412398 123646 412634
rect 123882 412398 159326 412634
rect 159562 412398 159646 412634
rect 159882 412398 195326 412634
rect 195562 412398 195646 412634
rect 195882 412398 231326 412634
rect 231562 412398 231646 412634
rect 231882 412398 267326 412634
rect 267562 412398 267646 412634
rect 267882 412398 303326 412634
rect 303562 412398 303646 412634
rect 303882 412398 339326 412634
rect 339562 412398 339646 412634
rect 339882 412398 375326 412634
rect 375562 412398 375646 412634
rect 375882 412398 411326 412634
rect 411562 412398 411646 412634
rect 411882 412398 447326 412634
rect 447562 412398 447646 412634
rect 447882 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 592650 412634
rect -8726 412366 592650 412398
rect -8726 408454 592650 408486
rect -8726 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 82826 408454
rect 83062 408218 83146 408454
rect 83382 408218 118826 408454
rect 119062 408218 119146 408454
rect 119382 408218 154826 408454
rect 155062 408218 155146 408454
rect 155382 408218 190826 408454
rect 191062 408218 191146 408454
rect 191382 408218 226826 408454
rect 227062 408218 227146 408454
rect 227382 408218 262826 408454
rect 263062 408218 263146 408454
rect 263382 408218 298826 408454
rect 299062 408218 299146 408454
rect 299382 408218 334826 408454
rect 335062 408218 335146 408454
rect 335382 408218 370826 408454
rect 371062 408218 371146 408454
rect 371382 408218 406826 408454
rect 407062 408218 407146 408454
rect 407382 408218 442826 408454
rect 443062 408218 443146 408454
rect 443382 408218 478826 408454
rect 479062 408218 479146 408454
rect 479382 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 592650 408454
rect -8726 408134 592650 408218
rect -8726 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 82826 408134
rect 83062 407898 83146 408134
rect 83382 407898 118826 408134
rect 119062 407898 119146 408134
rect 119382 407898 154826 408134
rect 155062 407898 155146 408134
rect 155382 407898 190826 408134
rect 191062 407898 191146 408134
rect 191382 407898 226826 408134
rect 227062 407898 227146 408134
rect 227382 407898 262826 408134
rect 263062 407898 263146 408134
rect 263382 407898 298826 408134
rect 299062 407898 299146 408134
rect 299382 407898 334826 408134
rect 335062 407898 335146 408134
rect 335382 407898 370826 408134
rect 371062 407898 371146 408134
rect 371382 407898 406826 408134
rect 407062 407898 407146 408134
rect 407382 407898 442826 408134
rect 443062 407898 443146 408134
rect 443382 407898 478826 408134
rect 479062 407898 479146 408134
rect 479382 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 592650 408134
rect -8726 407866 592650 407898
rect -8726 403954 592650 403986
rect -8726 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 78326 403954
rect 78562 403718 78646 403954
rect 78882 403718 114326 403954
rect 114562 403718 114646 403954
rect 114882 403718 150326 403954
rect 150562 403718 150646 403954
rect 150882 403718 186326 403954
rect 186562 403718 186646 403954
rect 186882 403718 222326 403954
rect 222562 403718 222646 403954
rect 222882 403718 258326 403954
rect 258562 403718 258646 403954
rect 258882 403718 294326 403954
rect 294562 403718 294646 403954
rect 294882 403718 330326 403954
rect 330562 403718 330646 403954
rect 330882 403718 366326 403954
rect 366562 403718 366646 403954
rect 366882 403718 402326 403954
rect 402562 403718 402646 403954
rect 402882 403718 438326 403954
rect 438562 403718 438646 403954
rect 438882 403718 474326 403954
rect 474562 403718 474646 403954
rect 474882 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 592650 403954
rect -8726 403634 592650 403718
rect -8726 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 78326 403634
rect 78562 403398 78646 403634
rect 78882 403398 114326 403634
rect 114562 403398 114646 403634
rect 114882 403398 150326 403634
rect 150562 403398 150646 403634
rect 150882 403398 186326 403634
rect 186562 403398 186646 403634
rect 186882 403398 222326 403634
rect 222562 403398 222646 403634
rect 222882 403398 258326 403634
rect 258562 403398 258646 403634
rect 258882 403398 294326 403634
rect 294562 403398 294646 403634
rect 294882 403398 330326 403634
rect 330562 403398 330646 403634
rect 330882 403398 366326 403634
rect 366562 403398 366646 403634
rect 366882 403398 402326 403634
rect 402562 403398 402646 403634
rect 402882 403398 438326 403634
rect 438562 403398 438646 403634
rect 438882 403398 474326 403634
rect 474562 403398 474646 403634
rect 474882 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 592650 403634
rect -8726 403366 592650 403398
rect -8726 399454 592650 399486
rect -8726 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 592650 399454
rect -8726 399134 592650 399218
rect -8726 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 592650 399134
rect -8726 398866 592650 398898
rect -8726 394954 592650 394986
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 69326 394954
rect 69562 394718 69646 394954
rect 69882 394718 105326 394954
rect 105562 394718 105646 394954
rect 105882 394718 141326 394954
rect 141562 394718 141646 394954
rect 141882 394718 177326 394954
rect 177562 394718 177646 394954
rect 177882 394718 213326 394954
rect 213562 394718 213646 394954
rect 213882 394718 249326 394954
rect 249562 394718 249646 394954
rect 249882 394718 285326 394954
rect 285562 394718 285646 394954
rect 285882 394718 321326 394954
rect 321562 394718 321646 394954
rect 321882 394718 357326 394954
rect 357562 394718 357646 394954
rect 357882 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect -8726 394634 592650 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 69326 394634
rect 69562 394398 69646 394634
rect 69882 394398 105326 394634
rect 105562 394398 105646 394634
rect 105882 394398 141326 394634
rect 141562 394398 141646 394634
rect 141882 394398 177326 394634
rect 177562 394398 177646 394634
rect 177882 394398 213326 394634
rect 213562 394398 213646 394634
rect 213882 394398 249326 394634
rect 249562 394398 249646 394634
rect 249882 394398 285326 394634
rect 285562 394398 285646 394634
rect 285882 394398 321326 394634
rect 321562 394398 321646 394634
rect 321882 394398 357326 394634
rect 357562 394398 357646 394634
rect 357882 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect -8726 394366 592650 394398
rect -8726 390454 592650 390486
rect -8726 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 64826 390454
rect 65062 390218 65146 390454
rect 65382 390218 100826 390454
rect 101062 390218 101146 390454
rect 101382 390218 136826 390454
rect 137062 390218 137146 390454
rect 137382 390218 172826 390454
rect 173062 390218 173146 390454
rect 173382 390218 208826 390454
rect 209062 390218 209146 390454
rect 209382 390218 244826 390454
rect 245062 390218 245146 390454
rect 245382 390218 280826 390454
rect 281062 390218 281146 390454
rect 281382 390218 316826 390454
rect 317062 390218 317146 390454
rect 317382 390218 352826 390454
rect 353062 390218 353146 390454
rect 353382 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 592650 390454
rect -8726 390134 592650 390218
rect -8726 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 64826 390134
rect 65062 389898 65146 390134
rect 65382 389898 100826 390134
rect 101062 389898 101146 390134
rect 101382 389898 136826 390134
rect 137062 389898 137146 390134
rect 137382 389898 172826 390134
rect 173062 389898 173146 390134
rect 173382 389898 208826 390134
rect 209062 389898 209146 390134
rect 209382 389898 244826 390134
rect 245062 389898 245146 390134
rect 245382 389898 280826 390134
rect 281062 389898 281146 390134
rect 281382 389898 316826 390134
rect 317062 389898 317146 390134
rect 317382 389898 352826 390134
rect 353062 389898 353146 390134
rect 353382 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 592650 390134
rect -8726 389866 592650 389898
rect -8726 385954 592650 385986
rect -8726 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 60326 385954
rect 60562 385718 60646 385954
rect 60882 385718 96326 385954
rect 96562 385718 96646 385954
rect 96882 385718 132326 385954
rect 132562 385718 132646 385954
rect 132882 385718 168326 385954
rect 168562 385718 168646 385954
rect 168882 385718 204326 385954
rect 204562 385718 204646 385954
rect 204882 385718 240326 385954
rect 240562 385718 240646 385954
rect 240882 385718 276326 385954
rect 276562 385718 276646 385954
rect 276882 385718 312326 385954
rect 312562 385718 312646 385954
rect 312882 385718 348326 385954
rect 348562 385718 348646 385954
rect 348882 385718 384326 385954
rect 384562 385718 384646 385954
rect 384882 385718 420326 385954
rect 420562 385718 420646 385954
rect 420882 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 592650 385954
rect -8726 385634 592650 385718
rect -8726 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 60326 385634
rect 60562 385398 60646 385634
rect 60882 385398 96326 385634
rect 96562 385398 96646 385634
rect 96882 385398 132326 385634
rect 132562 385398 132646 385634
rect 132882 385398 168326 385634
rect 168562 385398 168646 385634
rect 168882 385398 204326 385634
rect 204562 385398 204646 385634
rect 204882 385398 240326 385634
rect 240562 385398 240646 385634
rect 240882 385398 276326 385634
rect 276562 385398 276646 385634
rect 276882 385398 312326 385634
rect 312562 385398 312646 385634
rect 312882 385398 348326 385634
rect 348562 385398 348646 385634
rect 348882 385398 384326 385634
rect 384562 385398 384646 385634
rect 384882 385398 420326 385634
rect 420562 385398 420646 385634
rect 420882 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 592650 385634
rect -8726 385366 592650 385398
rect -8726 381454 592650 381486
rect -8726 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 592650 381454
rect -8726 381134 592650 381218
rect -8726 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 592650 381134
rect -8726 380866 592650 380898
rect -8726 376954 592650 376986
rect -8726 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 51326 376954
rect 51562 376718 51646 376954
rect 51882 376718 87326 376954
rect 87562 376718 87646 376954
rect 87882 376718 123326 376954
rect 123562 376718 123646 376954
rect 123882 376718 159326 376954
rect 159562 376718 159646 376954
rect 159882 376718 195326 376954
rect 195562 376718 195646 376954
rect 195882 376718 231326 376954
rect 231562 376718 231646 376954
rect 231882 376718 267326 376954
rect 267562 376718 267646 376954
rect 267882 376718 303326 376954
rect 303562 376718 303646 376954
rect 303882 376718 339326 376954
rect 339562 376718 339646 376954
rect 339882 376718 375326 376954
rect 375562 376718 375646 376954
rect 375882 376718 411326 376954
rect 411562 376718 411646 376954
rect 411882 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 592650 376954
rect -8726 376634 592650 376718
rect -8726 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 51326 376634
rect 51562 376398 51646 376634
rect 51882 376398 87326 376634
rect 87562 376398 87646 376634
rect 87882 376398 123326 376634
rect 123562 376398 123646 376634
rect 123882 376398 159326 376634
rect 159562 376398 159646 376634
rect 159882 376398 195326 376634
rect 195562 376398 195646 376634
rect 195882 376398 231326 376634
rect 231562 376398 231646 376634
rect 231882 376398 267326 376634
rect 267562 376398 267646 376634
rect 267882 376398 303326 376634
rect 303562 376398 303646 376634
rect 303882 376398 339326 376634
rect 339562 376398 339646 376634
rect 339882 376398 375326 376634
rect 375562 376398 375646 376634
rect 375882 376398 411326 376634
rect 411562 376398 411646 376634
rect 411882 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 592650 376634
rect -8726 376366 592650 376398
rect -8726 372454 592650 372486
rect -8726 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 82826 372454
rect 83062 372218 83146 372454
rect 83382 372218 118826 372454
rect 119062 372218 119146 372454
rect 119382 372218 154826 372454
rect 155062 372218 155146 372454
rect 155382 372218 190826 372454
rect 191062 372218 191146 372454
rect 191382 372218 226826 372454
rect 227062 372218 227146 372454
rect 227382 372218 262826 372454
rect 263062 372218 263146 372454
rect 263382 372218 298826 372454
rect 299062 372218 299146 372454
rect 299382 372218 334826 372454
rect 335062 372218 335146 372454
rect 335382 372218 370826 372454
rect 371062 372218 371146 372454
rect 371382 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 592650 372454
rect -8726 372134 592650 372218
rect -8726 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 82826 372134
rect 83062 371898 83146 372134
rect 83382 371898 118826 372134
rect 119062 371898 119146 372134
rect 119382 371898 154826 372134
rect 155062 371898 155146 372134
rect 155382 371898 190826 372134
rect 191062 371898 191146 372134
rect 191382 371898 226826 372134
rect 227062 371898 227146 372134
rect 227382 371898 262826 372134
rect 263062 371898 263146 372134
rect 263382 371898 298826 372134
rect 299062 371898 299146 372134
rect 299382 371898 334826 372134
rect 335062 371898 335146 372134
rect 335382 371898 370826 372134
rect 371062 371898 371146 372134
rect 371382 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 592650 372134
rect -8726 371866 592650 371898
rect -8726 367954 592650 367986
rect -8726 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 78326 367954
rect 78562 367718 78646 367954
rect 78882 367718 114326 367954
rect 114562 367718 114646 367954
rect 114882 367718 150326 367954
rect 150562 367718 150646 367954
rect 150882 367718 186326 367954
rect 186562 367718 186646 367954
rect 186882 367718 222326 367954
rect 222562 367718 222646 367954
rect 222882 367718 258326 367954
rect 258562 367718 258646 367954
rect 258882 367718 294326 367954
rect 294562 367718 294646 367954
rect 294882 367718 330326 367954
rect 330562 367718 330646 367954
rect 330882 367718 366326 367954
rect 366562 367718 366646 367954
rect 366882 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 592650 367954
rect -8726 367634 592650 367718
rect -8726 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 78326 367634
rect 78562 367398 78646 367634
rect 78882 367398 114326 367634
rect 114562 367398 114646 367634
rect 114882 367398 150326 367634
rect 150562 367398 150646 367634
rect 150882 367398 186326 367634
rect 186562 367398 186646 367634
rect 186882 367398 222326 367634
rect 222562 367398 222646 367634
rect 222882 367398 258326 367634
rect 258562 367398 258646 367634
rect 258882 367398 294326 367634
rect 294562 367398 294646 367634
rect 294882 367398 330326 367634
rect 330562 367398 330646 367634
rect 330882 367398 366326 367634
rect 366562 367398 366646 367634
rect 366882 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 592650 367634
rect -8726 367366 592650 367398
rect -8726 363454 592650 363486
rect -8726 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 592650 363454
rect -8726 363134 592650 363218
rect -8726 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 592650 363134
rect -8726 362866 592650 362898
rect -8726 358954 592650 358986
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 69326 358954
rect 69562 358718 69646 358954
rect 69882 358718 105326 358954
rect 105562 358718 105646 358954
rect 105882 358718 141326 358954
rect 141562 358718 141646 358954
rect 141882 358718 177326 358954
rect 177562 358718 177646 358954
rect 177882 358718 213326 358954
rect 213562 358718 213646 358954
rect 213882 358718 249326 358954
rect 249562 358718 249646 358954
rect 249882 358718 285326 358954
rect 285562 358718 285646 358954
rect 285882 358718 321326 358954
rect 321562 358718 321646 358954
rect 321882 358718 357326 358954
rect 357562 358718 357646 358954
rect 357882 358718 393326 358954
rect 393562 358718 393646 358954
rect 393882 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect -8726 358634 592650 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 69326 358634
rect 69562 358398 69646 358634
rect 69882 358398 105326 358634
rect 105562 358398 105646 358634
rect 105882 358398 141326 358634
rect 141562 358398 141646 358634
rect 141882 358398 177326 358634
rect 177562 358398 177646 358634
rect 177882 358398 213326 358634
rect 213562 358398 213646 358634
rect 213882 358398 249326 358634
rect 249562 358398 249646 358634
rect 249882 358398 285326 358634
rect 285562 358398 285646 358634
rect 285882 358398 321326 358634
rect 321562 358398 321646 358634
rect 321882 358398 357326 358634
rect 357562 358398 357646 358634
rect 357882 358398 393326 358634
rect 393562 358398 393646 358634
rect 393882 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect -8726 358366 592650 358398
rect -8726 354454 592650 354486
rect -8726 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 64826 354454
rect 65062 354218 65146 354454
rect 65382 354218 100826 354454
rect 101062 354218 101146 354454
rect 101382 354218 136826 354454
rect 137062 354218 137146 354454
rect 137382 354218 172826 354454
rect 173062 354218 173146 354454
rect 173382 354218 208826 354454
rect 209062 354218 209146 354454
rect 209382 354218 244826 354454
rect 245062 354218 245146 354454
rect 245382 354218 280826 354454
rect 281062 354218 281146 354454
rect 281382 354218 316826 354454
rect 317062 354218 317146 354454
rect 317382 354218 352826 354454
rect 353062 354218 353146 354454
rect 353382 354218 388826 354454
rect 389062 354218 389146 354454
rect 389382 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 592650 354454
rect -8726 354134 592650 354218
rect -8726 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 64826 354134
rect 65062 353898 65146 354134
rect 65382 353898 100826 354134
rect 101062 353898 101146 354134
rect 101382 353898 136826 354134
rect 137062 353898 137146 354134
rect 137382 353898 172826 354134
rect 173062 353898 173146 354134
rect 173382 353898 208826 354134
rect 209062 353898 209146 354134
rect 209382 353898 244826 354134
rect 245062 353898 245146 354134
rect 245382 353898 280826 354134
rect 281062 353898 281146 354134
rect 281382 353898 316826 354134
rect 317062 353898 317146 354134
rect 317382 353898 352826 354134
rect 353062 353898 353146 354134
rect 353382 353898 388826 354134
rect 389062 353898 389146 354134
rect 389382 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 592650 354134
rect -8726 353866 592650 353898
rect -8726 349954 592650 349986
rect -8726 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 60326 349954
rect 60562 349718 60646 349954
rect 60882 349718 96326 349954
rect 96562 349718 96646 349954
rect 96882 349718 132326 349954
rect 132562 349718 132646 349954
rect 132882 349718 168326 349954
rect 168562 349718 168646 349954
rect 168882 349718 204326 349954
rect 204562 349718 204646 349954
rect 204882 349718 240326 349954
rect 240562 349718 240646 349954
rect 240882 349718 276326 349954
rect 276562 349718 276646 349954
rect 276882 349718 312326 349954
rect 312562 349718 312646 349954
rect 312882 349718 348326 349954
rect 348562 349718 348646 349954
rect 348882 349718 384326 349954
rect 384562 349718 384646 349954
rect 384882 349718 420326 349954
rect 420562 349718 420646 349954
rect 420882 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 592650 349954
rect -8726 349634 592650 349718
rect -8726 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 60326 349634
rect 60562 349398 60646 349634
rect 60882 349398 96326 349634
rect 96562 349398 96646 349634
rect 96882 349398 132326 349634
rect 132562 349398 132646 349634
rect 132882 349398 168326 349634
rect 168562 349398 168646 349634
rect 168882 349398 204326 349634
rect 204562 349398 204646 349634
rect 204882 349398 240326 349634
rect 240562 349398 240646 349634
rect 240882 349398 276326 349634
rect 276562 349398 276646 349634
rect 276882 349398 312326 349634
rect 312562 349398 312646 349634
rect 312882 349398 348326 349634
rect 348562 349398 348646 349634
rect 348882 349398 384326 349634
rect 384562 349398 384646 349634
rect 384882 349398 420326 349634
rect 420562 349398 420646 349634
rect 420882 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 592650 349634
rect -8726 349366 592650 349398
rect -8726 345454 592650 345486
rect -8726 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 592650 345454
rect -8726 345134 592650 345218
rect -8726 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 592650 345134
rect -8726 344866 592650 344898
rect -8726 340954 592650 340986
rect -8726 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 51326 340954
rect 51562 340718 51646 340954
rect 51882 340718 87326 340954
rect 87562 340718 87646 340954
rect 87882 340718 123326 340954
rect 123562 340718 123646 340954
rect 123882 340718 159326 340954
rect 159562 340718 159646 340954
rect 159882 340718 195326 340954
rect 195562 340718 195646 340954
rect 195882 340718 231326 340954
rect 231562 340718 231646 340954
rect 231882 340718 267326 340954
rect 267562 340718 267646 340954
rect 267882 340718 303326 340954
rect 303562 340718 303646 340954
rect 303882 340718 339326 340954
rect 339562 340718 339646 340954
rect 339882 340718 375326 340954
rect 375562 340718 375646 340954
rect 375882 340718 411326 340954
rect 411562 340718 411646 340954
rect 411882 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 592650 340954
rect -8726 340634 592650 340718
rect -8726 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 51326 340634
rect 51562 340398 51646 340634
rect 51882 340398 87326 340634
rect 87562 340398 87646 340634
rect 87882 340398 123326 340634
rect 123562 340398 123646 340634
rect 123882 340398 159326 340634
rect 159562 340398 159646 340634
rect 159882 340398 195326 340634
rect 195562 340398 195646 340634
rect 195882 340398 231326 340634
rect 231562 340398 231646 340634
rect 231882 340398 267326 340634
rect 267562 340398 267646 340634
rect 267882 340398 303326 340634
rect 303562 340398 303646 340634
rect 303882 340398 339326 340634
rect 339562 340398 339646 340634
rect 339882 340398 375326 340634
rect 375562 340398 375646 340634
rect 375882 340398 411326 340634
rect 411562 340398 411646 340634
rect 411882 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 592650 340634
rect -8726 340366 592650 340398
rect -8726 336454 592650 336486
rect -8726 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 82826 336454
rect 83062 336218 83146 336454
rect 83382 336218 118826 336454
rect 119062 336218 119146 336454
rect 119382 336218 154826 336454
rect 155062 336218 155146 336454
rect 155382 336218 190826 336454
rect 191062 336218 191146 336454
rect 191382 336218 226826 336454
rect 227062 336218 227146 336454
rect 227382 336218 262826 336454
rect 263062 336218 263146 336454
rect 263382 336218 298826 336454
rect 299062 336218 299146 336454
rect 299382 336218 334826 336454
rect 335062 336218 335146 336454
rect 335382 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 592650 336454
rect -8726 336134 592650 336218
rect -8726 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 82826 336134
rect 83062 335898 83146 336134
rect 83382 335898 118826 336134
rect 119062 335898 119146 336134
rect 119382 335898 154826 336134
rect 155062 335898 155146 336134
rect 155382 335898 190826 336134
rect 191062 335898 191146 336134
rect 191382 335898 226826 336134
rect 227062 335898 227146 336134
rect 227382 335898 262826 336134
rect 263062 335898 263146 336134
rect 263382 335898 298826 336134
rect 299062 335898 299146 336134
rect 299382 335898 334826 336134
rect 335062 335898 335146 336134
rect 335382 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 592650 336134
rect -8726 335866 592650 335898
rect -8726 331954 592650 331986
rect -8726 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 78326 331954
rect 78562 331718 78646 331954
rect 78882 331718 114326 331954
rect 114562 331718 114646 331954
rect 114882 331718 150326 331954
rect 150562 331718 150646 331954
rect 150882 331718 186326 331954
rect 186562 331718 186646 331954
rect 186882 331718 222326 331954
rect 222562 331718 222646 331954
rect 222882 331718 258326 331954
rect 258562 331718 258646 331954
rect 258882 331718 294326 331954
rect 294562 331718 294646 331954
rect 294882 331718 330326 331954
rect 330562 331718 330646 331954
rect 330882 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 592650 331954
rect -8726 331634 592650 331718
rect -8726 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 78326 331634
rect 78562 331398 78646 331634
rect 78882 331398 114326 331634
rect 114562 331398 114646 331634
rect 114882 331398 150326 331634
rect 150562 331398 150646 331634
rect 150882 331398 186326 331634
rect 186562 331398 186646 331634
rect 186882 331398 222326 331634
rect 222562 331398 222646 331634
rect 222882 331398 258326 331634
rect 258562 331398 258646 331634
rect 258882 331398 294326 331634
rect 294562 331398 294646 331634
rect 294882 331398 330326 331634
rect 330562 331398 330646 331634
rect 330882 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 592650 331634
rect -8726 331366 592650 331398
rect -8726 327454 592650 327486
rect -8726 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 592650 327454
rect -8726 327134 592650 327218
rect -8726 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 592650 327134
rect -8726 326866 592650 326898
rect -8726 322954 592650 322986
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 69326 322954
rect 69562 322718 69646 322954
rect 69882 322718 105326 322954
rect 105562 322718 105646 322954
rect 105882 322718 141326 322954
rect 141562 322718 141646 322954
rect 141882 322718 177326 322954
rect 177562 322718 177646 322954
rect 177882 322718 213326 322954
rect 213562 322718 213646 322954
rect 213882 322718 249326 322954
rect 249562 322718 249646 322954
rect 249882 322718 285326 322954
rect 285562 322718 285646 322954
rect 285882 322718 321326 322954
rect 321562 322718 321646 322954
rect 321882 322718 357326 322954
rect 357562 322718 357646 322954
rect 357882 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect -8726 322634 592650 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 69326 322634
rect 69562 322398 69646 322634
rect 69882 322398 105326 322634
rect 105562 322398 105646 322634
rect 105882 322398 141326 322634
rect 141562 322398 141646 322634
rect 141882 322398 177326 322634
rect 177562 322398 177646 322634
rect 177882 322398 213326 322634
rect 213562 322398 213646 322634
rect 213882 322398 249326 322634
rect 249562 322398 249646 322634
rect 249882 322398 285326 322634
rect 285562 322398 285646 322634
rect 285882 322398 321326 322634
rect 321562 322398 321646 322634
rect 321882 322398 357326 322634
rect 357562 322398 357646 322634
rect 357882 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect -8726 322366 592650 322398
rect -8726 318454 592650 318486
rect -8726 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 64826 318454
rect 65062 318218 65146 318454
rect 65382 318218 100826 318454
rect 101062 318218 101146 318454
rect 101382 318218 136826 318454
rect 137062 318218 137146 318454
rect 137382 318218 172826 318454
rect 173062 318218 173146 318454
rect 173382 318218 208826 318454
rect 209062 318218 209146 318454
rect 209382 318218 244826 318454
rect 245062 318218 245146 318454
rect 245382 318218 280826 318454
rect 281062 318218 281146 318454
rect 281382 318218 316826 318454
rect 317062 318218 317146 318454
rect 317382 318218 352826 318454
rect 353062 318218 353146 318454
rect 353382 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 591102 318454
rect 591338 318218 591422 318454
rect 591658 318218 592650 318454
rect -8726 318134 592650 318218
rect -8726 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 64826 318134
rect 65062 317898 65146 318134
rect 65382 317898 100826 318134
rect 101062 317898 101146 318134
rect 101382 317898 136826 318134
rect 137062 317898 137146 318134
rect 137382 317898 172826 318134
rect 173062 317898 173146 318134
rect 173382 317898 208826 318134
rect 209062 317898 209146 318134
rect 209382 317898 244826 318134
rect 245062 317898 245146 318134
rect 245382 317898 280826 318134
rect 281062 317898 281146 318134
rect 281382 317898 316826 318134
rect 317062 317898 317146 318134
rect 317382 317898 352826 318134
rect 353062 317898 353146 318134
rect 353382 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 591102 318134
rect 591338 317898 591422 318134
rect 591658 317898 592650 318134
rect -8726 317866 592650 317898
rect -8726 313954 592650 313986
rect -8726 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 60326 313954
rect 60562 313718 60646 313954
rect 60882 313718 96326 313954
rect 96562 313718 96646 313954
rect 96882 313718 132326 313954
rect 132562 313718 132646 313954
rect 132882 313718 168326 313954
rect 168562 313718 168646 313954
rect 168882 313718 204326 313954
rect 204562 313718 204646 313954
rect 204882 313718 240326 313954
rect 240562 313718 240646 313954
rect 240882 313718 276326 313954
rect 276562 313718 276646 313954
rect 276882 313718 312326 313954
rect 312562 313718 312646 313954
rect 312882 313718 348326 313954
rect 348562 313718 348646 313954
rect 348882 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 420326 313954
rect 420562 313718 420646 313954
rect 420882 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 592650 313954
rect -8726 313634 592650 313718
rect -8726 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 60326 313634
rect 60562 313398 60646 313634
rect 60882 313398 96326 313634
rect 96562 313398 96646 313634
rect 96882 313398 132326 313634
rect 132562 313398 132646 313634
rect 132882 313398 168326 313634
rect 168562 313398 168646 313634
rect 168882 313398 204326 313634
rect 204562 313398 204646 313634
rect 204882 313398 240326 313634
rect 240562 313398 240646 313634
rect 240882 313398 276326 313634
rect 276562 313398 276646 313634
rect 276882 313398 312326 313634
rect 312562 313398 312646 313634
rect 312882 313398 348326 313634
rect 348562 313398 348646 313634
rect 348882 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 420326 313634
rect 420562 313398 420646 313634
rect 420882 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 592650 313634
rect -8726 313366 592650 313398
rect -8726 309454 592650 309486
rect -8726 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 592650 309454
rect -8726 309134 592650 309218
rect -8726 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 592650 309134
rect -8726 308866 592650 308898
rect -8726 304954 592650 304986
rect -8726 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 51326 304954
rect 51562 304718 51646 304954
rect 51882 304718 87326 304954
rect 87562 304718 87646 304954
rect 87882 304718 123326 304954
rect 123562 304718 123646 304954
rect 123882 304718 159326 304954
rect 159562 304718 159646 304954
rect 159882 304718 195326 304954
rect 195562 304718 195646 304954
rect 195882 304718 231326 304954
rect 231562 304718 231646 304954
rect 231882 304718 267326 304954
rect 267562 304718 267646 304954
rect 267882 304718 303326 304954
rect 303562 304718 303646 304954
rect 303882 304718 339326 304954
rect 339562 304718 339646 304954
rect 339882 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 411326 304954
rect 411562 304718 411646 304954
rect 411882 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 592650 304954
rect -8726 304634 592650 304718
rect -8726 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 51326 304634
rect 51562 304398 51646 304634
rect 51882 304398 87326 304634
rect 87562 304398 87646 304634
rect 87882 304398 123326 304634
rect 123562 304398 123646 304634
rect 123882 304398 159326 304634
rect 159562 304398 159646 304634
rect 159882 304398 195326 304634
rect 195562 304398 195646 304634
rect 195882 304398 231326 304634
rect 231562 304398 231646 304634
rect 231882 304398 267326 304634
rect 267562 304398 267646 304634
rect 267882 304398 303326 304634
rect 303562 304398 303646 304634
rect 303882 304398 339326 304634
rect 339562 304398 339646 304634
rect 339882 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 411326 304634
rect 411562 304398 411646 304634
rect 411882 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 592650 304634
rect -8726 304366 592650 304398
rect -8726 300454 592650 300486
rect -8726 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 82826 300454
rect 83062 300218 83146 300454
rect 83382 300218 118826 300454
rect 119062 300218 119146 300454
rect 119382 300218 154826 300454
rect 155062 300218 155146 300454
rect 155382 300218 190826 300454
rect 191062 300218 191146 300454
rect 191382 300218 226826 300454
rect 227062 300218 227146 300454
rect 227382 300218 262826 300454
rect 263062 300218 263146 300454
rect 263382 300218 298826 300454
rect 299062 300218 299146 300454
rect 299382 300218 334826 300454
rect 335062 300218 335146 300454
rect 335382 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 592650 300454
rect -8726 300134 592650 300218
rect -8726 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 82826 300134
rect 83062 299898 83146 300134
rect 83382 299898 118826 300134
rect 119062 299898 119146 300134
rect 119382 299898 154826 300134
rect 155062 299898 155146 300134
rect 155382 299898 190826 300134
rect 191062 299898 191146 300134
rect 191382 299898 226826 300134
rect 227062 299898 227146 300134
rect 227382 299898 262826 300134
rect 263062 299898 263146 300134
rect 263382 299898 298826 300134
rect 299062 299898 299146 300134
rect 299382 299898 334826 300134
rect 335062 299898 335146 300134
rect 335382 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 592650 300134
rect -8726 299866 592650 299898
rect -8726 295954 592650 295986
rect -8726 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 78326 295954
rect 78562 295718 78646 295954
rect 78882 295718 114326 295954
rect 114562 295718 114646 295954
rect 114882 295718 150326 295954
rect 150562 295718 150646 295954
rect 150882 295718 186326 295954
rect 186562 295718 186646 295954
rect 186882 295718 222326 295954
rect 222562 295718 222646 295954
rect 222882 295718 258326 295954
rect 258562 295718 258646 295954
rect 258882 295718 294326 295954
rect 294562 295718 294646 295954
rect 294882 295718 330326 295954
rect 330562 295718 330646 295954
rect 330882 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 438326 295954
rect 438562 295718 438646 295954
rect 438882 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 592650 295954
rect -8726 295634 592650 295718
rect -8726 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 78326 295634
rect 78562 295398 78646 295634
rect 78882 295398 114326 295634
rect 114562 295398 114646 295634
rect 114882 295398 150326 295634
rect 150562 295398 150646 295634
rect 150882 295398 186326 295634
rect 186562 295398 186646 295634
rect 186882 295398 222326 295634
rect 222562 295398 222646 295634
rect 222882 295398 258326 295634
rect 258562 295398 258646 295634
rect 258882 295398 294326 295634
rect 294562 295398 294646 295634
rect 294882 295398 330326 295634
rect 330562 295398 330646 295634
rect 330882 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 438326 295634
rect 438562 295398 438646 295634
rect 438882 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 592650 295634
rect -8726 295366 592650 295398
rect -8726 291454 592650 291486
rect -8726 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 592650 291454
rect -8726 291134 592650 291218
rect -8726 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 592650 291134
rect -8726 290866 592650 290898
rect -8726 286954 592650 286986
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 69326 286954
rect 69562 286718 69646 286954
rect 69882 286718 105326 286954
rect 105562 286718 105646 286954
rect 105882 286718 141326 286954
rect 141562 286718 141646 286954
rect 141882 286718 177326 286954
rect 177562 286718 177646 286954
rect 177882 286718 213326 286954
rect 213562 286718 213646 286954
rect 213882 286718 249326 286954
rect 249562 286718 249646 286954
rect 249882 286718 285326 286954
rect 285562 286718 285646 286954
rect 285882 286718 321326 286954
rect 321562 286718 321646 286954
rect 321882 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 393326 286954
rect 393562 286718 393646 286954
rect 393882 286718 429326 286954
rect 429562 286718 429646 286954
rect 429882 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect -8726 286634 592650 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 69326 286634
rect 69562 286398 69646 286634
rect 69882 286398 105326 286634
rect 105562 286398 105646 286634
rect 105882 286398 141326 286634
rect 141562 286398 141646 286634
rect 141882 286398 177326 286634
rect 177562 286398 177646 286634
rect 177882 286398 213326 286634
rect 213562 286398 213646 286634
rect 213882 286398 249326 286634
rect 249562 286398 249646 286634
rect 249882 286398 285326 286634
rect 285562 286398 285646 286634
rect 285882 286398 321326 286634
rect 321562 286398 321646 286634
rect 321882 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 393326 286634
rect 393562 286398 393646 286634
rect 393882 286398 429326 286634
rect 429562 286398 429646 286634
rect 429882 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect -8726 286366 592650 286398
rect -8726 282454 592650 282486
rect -8726 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 64826 282454
rect 65062 282218 65146 282454
rect 65382 282218 100826 282454
rect 101062 282218 101146 282454
rect 101382 282218 136826 282454
rect 137062 282218 137146 282454
rect 137382 282218 172826 282454
rect 173062 282218 173146 282454
rect 173382 282218 208826 282454
rect 209062 282218 209146 282454
rect 209382 282218 244826 282454
rect 245062 282218 245146 282454
rect 245382 282218 280826 282454
rect 281062 282218 281146 282454
rect 281382 282218 316826 282454
rect 317062 282218 317146 282454
rect 317382 282218 352826 282454
rect 353062 282218 353146 282454
rect 353382 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 592650 282454
rect -8726 282134 592650 282218
rect -8726 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 64826 282134
rect 65062 281898 65146 282134
rect 65382 281898 100826 282134
rect 101062 281898 101146 282134
rect 101382 281898 136826 282134
rect 137062 281898 137146 282134
rect 137382 281898 172826 282134
rect 173062 281898 173146 282134
rect 173382 281898 208826 282134
rect 209062 281898 209146 282134
rect 209382 281898 244826 282134
rect 245062 281898 245146 282134
rect 245382 281898 280826 282134
rect 281062 281898 281146 282134
rect 281382 281898 316826 282134
rect 317062 281898 317146 282134
rect 317382 281898 352826 282134
rect 353062 281898 353146 282134
rect 353382 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 592650 282134
rect -8726 281866 592650 281898
rect -8726 277954 592650 277986
rect -8726 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 96326 277954
rect 96562 277718 96646 277954
rect 96882 277718 132326 277954
rect 132562 277718 132646 277954
rect 132882 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 204326 277954
rect 204562 277718 204646 277954
rect 204882 277718 240326 277954
rect 240562 277718 240646 277954
rect 240882 277718 276326 277954
rect 276562 277718 276646 277954
rect 276882 277718 312326 277954
rect 312562 277718 312646 277954
rect 312882 277718 348326 277954
rect 348562 277718 348646 277954
rect 348882 277718 384326 277954
rect 384562 277718 384646 277954
rect 384882 277718 420326 277954
rect 420562 277718 420646 277954
rect 420882 277718 456326 277954
rect 456562 277718 456646 277954
rect 456882 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 592650 277954
rect -8726 277634 592650 277718
rect -8726 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 96326 277634
rect 96562 277398 96646 277634
rect 96882 277398 132326 277634
rect 132562 277398 132646 277634
rect 132882 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 204326 277634
rect 204562 277398 204646 277634
rect 204882 277398 240326 277634
rect 240562 277398 240646 277634
rect 240882 277398 276326 277634
rect 276562 277398 276646 277634
rect 276882 277398 312326 277634
rect 312562 277398 312646 277634
rect 312882 277398 348326 277634
rect 348562 277398 348646 277634
rect 348882 277398 384326 277634
rect 384562 277398 384646 277634
rect 384882 277398 420326 277634
rect 420562 277398 420646 277634
rect 420882 277398 456326 277634
rect 456562 277398 456646 277634
rect 456882 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 592650 277634
rect -8726 277366 592650 277398
rect -8726 273454 592650 273486
rect -8726 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 592650 273454
rect -8726 273134 592650 273218
rect -8726 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 592650 273134
rect -8726 272866 592650 272898
rect -8726 268954 592650 268986
rect -8726 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 87326 268954
rect 87562 268718 87646 268954
rect 87882 268718 123326 268954
rect 123562 268718 123646 268954
rect 123882 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 195326 268954
rect 195562 268718 195646 268954
rect 195882 268718 231326 268954
rect 231562 268718 231646 268954
rect 231882 268718 267326 268954
rect 267562 268718 267646 268954
rect 267882 268718 303326 268954
rect 303562 268718 303646 268954
rect 303882 268718 339326 268954
rect 339562 268718 339646 268954
rect 339882 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 411326 268954
rect 411562 268718 411646 268954
rect 411882 268718 447326 268954
rect 447562 268718 447646 268954
rect 447882 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 592650 268954
rect -8726 268634 592650 268718
rect -8726 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 87326 268634
rect 87562 268398 87646 268634
rect 87882 268398 123326 268634
rect 123562 268398 123646 268634
rect 123882 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 195326 268634
rect 195562 268398 195646 268634
rect 195882 268398 231326 268634
rect 231562 268398 231646 268634
rect 231882 268398 267326 268634
rect 267562 268398 267646 268634
rect 267882 268398 303326 268634
rect 303562 268398 303646 268634
rect 303882 268398 339326 268634
rect 339562 268398 339646 268634
rect 339882 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 411326 268634
rect 411562 268398 411646 268634
rect 411882 268398 447326 268634
rect 447562 268398 447646 268634
rect 447882 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 592650 268634
rect -8726 268366 592650 268398
rect -8726 264454 592650 264486
rect -8726 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 82826 264454
rect 83062 264218 83146 264454
rect 83382 264218 118826 264454
rect 119062 264218 119146 264454
rect 119382 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 190826 264454
rect 191062 264218 191146 264454
rect 191382 264218 226826 264454
rect 227062 264218 227146 264454
rect 227382 264218 262826 264454
rect 263062 264218 263146 264454
rect 263382 264218 298826 264454
rect 299062 264218 299146 264454
rect 299382 264218 334826 264454
rect 335062 264218 335146 264454
rect 335382 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 406826 264454
rect 407062 264218 407146 264454
rect 407382 264218 442826 264454
rect 443062 264218 443146 264454
rect 443382 264218 478826 264454
rect 479062 264218 479146 264454
rect 479382 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 592650 264454
rect -8726 264134 592650 264218
rect -8726 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 82826 264134
rect 83062 263898 83146 264134
rect 83382 263898 118826 264134
rect 119062 263898 119146 264134
rect 119382 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 190826 264134
rect 191062 263898 191146 264134
rect 191382 263898 226826 264134
rect 227062 263898 227146 264134
rect 227382 263898 262826 264134
rect 263062 263898 263146 264134
rect 263382 263898 298826 264134
rect 299062 263898 299146 264134
rect 299382 263898 334826 264134
rect 335062 263898 335146 264134
rect 335382 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 406826 264134
rect 407062 263898 407146 264134
rect 407382 263898 442826 264134
rect 443062 263898 443146 264134
rect 443382 263898 478826 264134
rect 479062 263898 479146 264134
rect 479382 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 592650 264134
rect -8726 263866 592650 263898
rect -8726 259954 592650 259986
rect -8726 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 78326 259954
rect 78562 259718 78646 259954
rect 78882 259718 114326 259954
rect 114562 259718 114646 259954
rect 114882 259718 222326 259954
rect 222562 259718 222646 259954
rect 222882 259718 258326 259954
rect 258562 259718 258646 259954
rect 258882 259718 294326 259954
rect 294562 259718 294646 259954
rect 294882 259718 330326 259954
rect 330562 259718 330646 259954
rect 330882 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 402326 259954
rect 402562 259718 402646 259954
rect 402882 259718 438326 259954
rect 438562 259718 438646 259954
rect 438882 259718 474326 259954
rect 474562 259718 474646 259954
rect 474882 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 592650 259954
rect -8726 259634 592650 259718
rect -8726 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 78326 259634
rect 78562 259398 78646 259634
rect 78882 259398 114326 259634
rect 114562 259398 114646 259634
rect 114882 259398 222326 259634
rect 222562 259398 222646 259634
rect 222882 259398 258326 259634
rect 258562 259398 258646 259634
rect 258882 259398 294326 259634
rect 294562 259398 294646 259634
rect 294882 259398 330326 259634
rect 330562 259398 330646 259634
rect 330882 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 402326 259634
rect 402562 259398 402646 259634
rect 402882 259398 438326 259634
rect 438562 259398 438646 259634
rect 438882 259398 474326 259634
rect 474562 259398 474646 259634
rect 474882 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 592650 259634
rect -8726 259366 592650 259398
rect -8726 255454 592650 255486
rect -8726 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 124250 255454
rect 124486 255218 154970 255454
rect 155206 255218 185690 255454
rect 185926 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 592650 255454
rect -8726 255134 592650 255218
rect -8726 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 124250 255134
rect 124486 254898 154970 255134
rect 155206 254898 185690 255134
rect 185926 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 592650 255134
rect -8726 254866 592650 254898
rect -8726 250954 592650 250986
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 69326 250954
rect 69562 250718 69646 250954
rect 69882 250718 105326 250954
rect 105562 250718 105646 250954
rect 105882 250718 213326 250954
rect 213562 250718 213646 250954
rect 213882 250718 249326 250954
rect 249562 250718 249646 250954
rect 249882 250718 285326 250954
rect 285562 250718 285646 250954
rect 285882 250718 321326 250954
rect 321562 250718 321646 250954
rect 321882 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 393326 250954
rect 393562 250718 393646 250954
rect 393882 250718 429326 250954
rect 429562 250718 429646 250954
rect 429882 250718 465326 250954
rect 465562 250718 465646 250954
rect 465882 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect -8726 250634 592650 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 69326 250634
rect 69562 250398 69646 250634
rect 69882 250398 105326 250634
rect 105562 250398 105646 250634
rect 105882 250398 213326 250634
rect 213562 250398 213646 250634
rect 213882 250398 249326 250634
rect 249562 250398 249646 250634
rect 249882 250398 285326 250634
rect 285562 250398 285646 250634
rect 285882 250398 321326 250634
rect 321562 250398 321646 250634
rect 321882 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 393326 250634
rect 393562 250398 393646 250634
rect 393882 250398 429326 250634
rect 429562 250398 429646 250634
rect 429882 250398 465326 250634
rect 465562 250398 465646 250634
rect 465882 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect -8726 250366 592650 250398
rect -8726 246454 592650 246486
rect -8726 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246218 64826 246454
rect 65062 246218 65146 246454
rect 65382 246218 100826 246454
rect 101062 246218 101146 246454
rect 101382 246218 208826 246454
rect 209062 246218 209146 246454
rect 209382 246218 244826 246454
rect 245062 246218 245146 246454
rect 245382 246218 280826 246454
rect 281062 246218 281146 246454
rect 281382 246218 316826 246454
rect 317062 246218 317146 246454
rect 317382 246218 352826 246454
rect 353062 246218 353146 246454
rect 353382 246218 388826 246454
rect 389062 246218 389146 246454
rect 389382 246218 424826 246454
rect 425062 246218 425146 246454
rect 425382 246218 460826 246454
rect 461062 246218 461146 246454
rect 461382 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 592650 246454
rect -8726 246134 592650 246218
rect -8726 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 245898 64826 246134
rect 65062 245898 65146 246134
rect 65382 245898 100826 246134
rect 101062 245898 101146 246134
rect 101382 245898 208826 246134
rect 209062 245898 209146 246134
rect 209382 245898 244826 246134
rect 245062 245898 245146 246134
rect 245382 245898 280826 246134
rect 281062 245898 281146 246134
rect 281382 245898 316826 246134
rect 317062 245898 317146 246134
rect 317382 245898 352826 246134
rect 353062 245898 353146 246134
rect 353382 245898 388826 246134
rect 389062 245898 389146 246134
rect 389382 245898 424826 246134
rect 425062 245898 425146 246134
rect 425382 245898 460826 246134
rect 461062 245898 461146 246134
rect 461382 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 592650 246134
rect -8726 245866 592650 245898
rect -8726 241954 592650 241986
rect -8726 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241718 60326 241954
rect 60562 241718 60646 241954
rect 60882 241718 96326 241954
rect 96562 241718 96646 241954
rect 96882 241718 204326 241954
rect 204562 241718 204646 241954
rect 204882 241718 240326 241954
rect 240562 241718 240646 241954
rect 240882 241718 276326 241954
rect 276562 241718 276646 241954
rect 276882 241718 312326 241954
rect 312562 241718 312646 241954
rect 312882 241718 348326 241954
rect 348562 241718 348646 241954
rect 348882 241718 384326 241954
rect 384562 241718 384646 241954
rect 384882 241718 420326 241954
rect 420562 241718 420646 241954
rect 420882 241718 456326 241954
rect 456562 241718 456646 241954
rect 456882 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 592650 241954
rect -8726 241634 592650 241718
rect -8726 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241398 60326 241634
rect 60562 241398 60646 241634
rect 60882 241398 96326 241634
rect 96562 241398 96646 241634
rect 96882 241398 204326 241634
rect 204562 241398 204646 241634
rect 204882 241398 240326 241634
rect 240562 241398 240646 241634
rect 240882 241398 276326 241634
rect 276562 241398 276646 241634
rect 276882 241398 312326 241634
rect 312562 241398 312646 241634
rect 312882 241398 348326 241634
rect 348562 241398 348646 241634
rect 348882 241398 384326 241634
rect 384562 241398 384646 241634
rect 384882 241398 420326 241634
rect 420562 241398 420646 241634
rect 420882 241398 456326 241634
rect 456562 241398 456646 241634
rect 456882 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 592650 241634
rect -8726 241366 592650 241398
rect -8726 237454 592650 237486
rect -8726 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 592650 237454
rect -8726 237134 592650 237218
rect -8726 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 592650 237134
rect -8726 236866 592650 236898
rect -8726 232954 592650 232986
rect -8726 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 51326 232954
rect 51562 232718 51646 232954
rect 51882 232718 87326 232954
rect 87562 232718 87646 232954
rect 87882 232718 195326 232954
rect 195562 232718 195646 232954
rect 195882 232718 231326 232954
rect 231562 232718 231646 232954
rect 231882 232718 267326 232954
rect 267562 232718 267646 232954
rect 267882 232718 303326 232954
rect 303562 232718 303646 232954
rect 303882 232718 339326 232954
rect 339562 232718 339646 232954
rect 339882 232718 375326 232954
rect 375562 232718 375646 232954
rect 375882 232718 411326 232954
rect 411562 232718 411646 232954
rect 411882 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 592650 232954
rect -8726 232634 592650 232718
rect -8726 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 51326 232634
rect 51562 232398 51646 232634
rect 51882 232398 87326 232634
rect 87562 232398 87646 232634
rect 87882 232398 195326 232634
rect 195562 232398 195646 232634
rect 195882 232398 231326 232634
rect 231562 232398 231646 232634
rect 231882 232398 267326 232634
rect 267562 232398 267646 232634
rect 267882 232398 303326 232634
rect 303562 232398 303646 232634
rect 303882 232398 339326 232634
rect 339562 232398 339646 232634
rect 339882 232398 375326 232634
rect 375562 232398 375646 232634
rect 375882 232398 411326 232634
rect 411562 232398 411646 232634
rect 411882 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 592650 232634
rect -8726 232366 592650 232398
rect -8726 228454 592650 228486
rect -8726 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 46826 228454
rect 47062 228218 47146 228454
rect 47382 228218 82826 228454
rect 83062 228218 83146 228454
rect 83382 228218 226826 228454
rect 227062 228218 227146 228454
rect 227382 228218 262826 228454
rect 263062 228218 263146 228454
rect 263382 228218 298826 228454
rect 299062 228218 299146 228454
rect 299382 228218 334826 228454
rect 335062 228218 335146 228454
rect 335382 228218 370826 228454
rect 371062 228218 371146 228454
rect 371382 228218 406826 228454
rect 407062 228218 407146 228454
rect 407382 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 592650 228454
rect -8726 228134 592650 228218
rect -8726 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 46826 228134
rect 47062 227898 47146 228134
rect 47382 227898 82826 228134
rect 83062 227898 83146 228134
rect 83382 227898 226826 228134
rect 227062 227898 227146 228134
rect 227382 227898 262826 228134
rect 263062 227898 263146 228134
rect 263382 227898 298826 228134
rect 299062 227898 299146 228134
rect 299382 227898 334826 228134
rect 335062 227898 335146 228134
rect 335382 227898 370826 228134
rect 371062 227898 371146 228134
rect 371382 227898 406826 228134
rect 407062 227898 407146 228134
rect 407382 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 592650 228134
rect -8726 227866 592650 227898
rect -8726 223954 592650 223986
rect -8726 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 78326 223954
rect 78562 223718 78646 223954
rect 78882 223718 114326 223954
rect 114562 223718 114646 223954
rect 114882 223718 139610 223954
rect 139846 223718 170330 223954
rect 170566 223718 222326 223954
rect 222562 223718 222646 223954
rect 222882 223718 258326 223954
rect 258562 223718 258646 223954
rect 258882 223718 294326 223954
rect 294562 223718 294646 223954
rect 294882 223718 330326 223954
rect 330562 223718 330646 223954
rect 330882 223718 366326 223954
rect 366562 223718 366646 223954
rect 366882 223718 402326 223954
rect 402562 223718 402646 223954
rect 402882 223718 438326 223954
rect 438562 223718 438646 223954
rect 438882 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 592650 223954
rect -8726 223634 592650 223718
rect -8726 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 78326 223634
rect 78562 223398 78646 223634
rect 78882 223398 114326 223634
rect 114562 223398 114646 223634
rect 114882 223398 139610 223634
rect 139846 223398 170330 223634
rect 170566 223398 222326 223634
rect 222562 223398 222646 223634
rect 222882 223398 258326 223634
rect 258562 223398 258646 223634
rect 258882 223398 294326 223634
rect 294562 223398 294646 223634
rect 294882 223398 330326 223634
rect 330562 223398 330646 223634
rect 330882 223398 366326 223634
rect 366562 223398 366646 223634
rect 366882 223398 402326 223634
rect 402562 223398 402646 223634
rect 402882 223398 438326 223634
rect 438562 223398 438646 223634
rect 438882 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 592650 223634
rect -8726 223366 592650 223398
rect -8726 219454 592650 219486
rect -8726 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 124250 219454
rect 124486 219218 154970 219454
rect 155206 219218 185690 219454
rect 185926 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 592650 219454
rect -8726 219134 592650 219218
rect -8726 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 124250 219134
rect 124486 218898 154970 219134
rect 155206 218898 185690 219134
rect 185926 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 592650 219134
rect -8726 218866 592650 218898
rect -8726 214954 592650 214986
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 69326 214954
rect 69562 214718 69646 214954
rect 69882 214718 105326 214954
rect 105562 214718 105646 214954
rect 105882 214718 213326 214954
rect 213562 214718 213646 214954
rect 213882 214718 249326 214954
rect 249562 214718 249646 214954
rect 249882 214718 285326 214954
rect 285562 214718 285646 214954
rect 285882 214718 321326 214954
rect 321562 214718 321646 214954
rect 321882 214718 357326 214954
rect 357562 214718 357646 214954
rect 357882 214718 393326 214954
rect 393562 214718 393646 214954
rect 393882 214718 429326 214954
rect 429562 214718 429646 214954
rect 429882 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect -8726 214634 592650 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 69326 214634
rect 69562 214398 69646 214634
rect 69882 214398 105326 214634
rect 105562 214398 105646 214634
rect 105882 214398 213326 214634
rect 213562 214398 213646 214634
rect 213882 214398 249326 214634
rect 249562 214398 249646 214634
rect 249882 214398 285326 214634
rect 285562 214398 285646 214634
rect 285882 214398 321326 214634
rect 321562 214398 321646 214634
rect 321882 214398 357326 214634
rect 357562 214398 357646 214634
rect 357882 214398 393326 214634
rect 393562 214398 393646 214634
rect 393882 214398 429326 214634
rect 429562 214398 429646 214634
rect 429882 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect -8726 214366 592650 214398
rect -8726 210454 592650 210486
rect -8726 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 64826 210454
rect 65062 210218 65146 210454
rect 65382 210218 100826 210454
rect 101062 210218 101146 210454
rect 101382 210218 208826 210454
rect 209062 210218 209146 210454
rect 209382 210218 244826 210454
rect 245062 210218 245146 210454
rect 245382 210218 280826 210454
rect 281062 210218 281146 210454
rect 281382 210218 316826 210454
rect 317062 210218 317146 210454
rect 317382 210218 352826 210454
rect 353062 210218 353146 210454
rect 353382 210218 388826 210454
rect 389062 210218 389146 210454
rect 389382 210218 424826 210454
rect 425062 210218 425146 210454
rect 425382 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 592650 210454
rect -8726 210134 592650 210218
rect -8726 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 64826 210134
rect 65062 209898 65146 210134
rect 65382 209898 100826 210134
rect 101062 209898 101146 210134
rect 101382 209898 208826 210134
rect 209062 209898 209146 210134
rect 209382 209898 244826 210134
rect 245062 209898 245146 210134
rect 245382 209898 280826 210134
rect 281062 209898 281146 210134
rect 281382 209898 316826 210134
rect 317062 209898 317146 210134
rect 317382 209898 352826 210134
rect 353062 209898 353146 210134
rect 353382 209898 388826 210134
rect 389062 209898 389146 210134
rect 389382 209898 424826 210134
rect 425062 209898 425146 210134
rect 425382 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 592650 210134
rect -8726 209866 592650 209898
rect -8726 205954 592650 205986
rect -8726 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 60326 205954
rect 60562 205718 60646 205954
rect 60882 205718 96326 205954
rect 96562 205718 96646 205954
rect 96882 205718 204326 205954
rect 204562 205718 204646 205954
rect 204882 205718 240326 205954
rect 240562 205718 240646 205954
rect 240882 205718 276326 205954
rect 276562 205718 276646 205954
rect 276882 205718 312326 205954
rect 312562 205718 312646 205954
rect 312882 205718 348326 205954
rect 348562 205718 348646 205954
rect 348882 205718 384326 205954
rect 384562 205718 384646 205954
rect 384882 205718 420326 205954
rect 420562 205718 420646 205954
rect 420882 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 592650 205954
rect -8726 205634 592650 205718
rect -8726 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 60326 205634
rect 60562 205398 60646 205634
rect 60882 205398 96326 205634
rect 96562 205398 96646 205634
rect 96882 205398 204326 205634
rect 204562 205398 204646 205634
rect 204882 205398 240326 205634
rect 240562 205398 240646 205634
rect 240882 205398 276326 205634
rect 276562 205398 276646 205634
rect 276882 205398 312326 205634
rect 312562 205398 312646 205634
rect 312882 205398 348326 205634
rect 348562 205398 348646 205634
rect 348882 205398 384326 205634
rect 384562 205398 384646 205634
rect 384882 205398 420326 205634
rect 420562 205398 420646 205634
rect 420882 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 592650 205634
rect -8726 205366 592650 205398
rect -8726 201454 592650 201486
rect -8726 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 592650 201454
rect -8726 201134 592650 201218
rect -8726 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 592650 201134
rect -8726 200866 592650 200898
rect -8726 196954 592650 196986
rect -8726 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 123326 196954
rect 123562 196718 123646 196954
rect 123882 196718 159326 196954
rect 159562 196718 159646 196954
rect 159882 196718 195326 196954
rect 195562 196718 195646 196954
rect 195882 196718 231326 196954
rect 231562 196718 231646 196954
rect 231882 196718 267326 196954
rect 267562 196718 267646 196954
rect 267882 196718 303326 196954
rect 303562 196718 303646 196954
rect 303882 196718 339326 196954
rect 339562 196718 339646 196954
rect 339882 196718 375326 196954
rect 375562 196718 375646 196954
rect 375882 196718 411326 196954
rect 411562 196718 411646 196954
rect 411882 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 592650 196954
rect -8726 196634 592650 196718
rect -8726 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 123326 196634
rect 123562 196398 123646 196634
rect 123882 196398 159326 196634
rect 159562 196398 159646 196634
rect 159882 196398 195326 196634
rect 195562 196398 195646 196634
rect 195882 196398 231326 196634
rect 231562 196398 231646 196634
rect 231882 196398 267326 196634
rect 267562 196398 267646 196634
rect 267882 196398 303326 196634
rect 303562 196398 303646 196634
rect 303882 196398 339326 196634
rect 339562 196398 339646 196634
rect 339882 196398 375326 196634
rect 375562 196398 375646 196634
rect 375882 196398 411326 196634
rect 411562 196398 411646 196634
rect 411882 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 592650 196634
rect -8726 196366 592650 196398
rect -8726 192454 592650 192486
rect -8726 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 82826 192454
rect 83062 192218 83146 192454
rect 83382 192218 118826 192454
rect 119062 192218 119146 192454
rect 119382 192218 154826 192454
rect 155062 192218 155146 192454
rect 155382 192218 190826 192454
rect 191062 192218 191146 192454
rect 191382 192218 226826 192454
rect 227062 192218 227146 192454
rect 227382 192218 262826 192454
rect 263062 192218 263146 192454
rect 263382 192218 298826 192454
rect 299062 192218 299146 192454
rect 299382 192218 334826 192454
rect 335062 192218 335146 192454
rect 335382 192218 370826 192454
rect 371062 192218 371146 192454
rect 371382 192218 406826 192454
rect 407062 192218 407146 192454
rect 407382 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 592650 192454
rect -8726 192134 592650 192218
rect -8726 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 82826 192134
rect 83062 191898 83146 192134
rect 83382 191898 118826 192134
rect 119062 191898 119146 192134
rect 119382 191898 154826 192134
rect 155062 191898 155146 192134
rect 155382 191898 190826 192134
rect 191062 191898 191146 192134
rect 191382 191898 226826 192134
rect 227062 191898 227146 192134
rect 227382 191898 262826 192134
rect 263062 191898 263146 192134
rect 263382 191898 298826 192134
rect 299062 191898 299146 192134
rect 299382 191898 334826 192134
rect 335062 191898 335146 192134
rect 335382 191898 370826 192134
rect 371062 191898 371146 192134
rect 371382 191898 406826 192134
rect 407062 191898 407146 192134
rect 407382 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 592650 192134
rect -8726 191866 592650 191898
rect -8726 187954 592650 187986
rect -8726 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 78326 187954
rect 78562 187718 78646 187954
rect 78882 187718 114326 187954
rect 114562 187718 114646 187954
rect 114882 187718 150326 187954
rect 150562 187718 150646 187954
rect 150882 187718 186326 187954
rect 186562 187718 186646 187954
rect 186882 187718 222326 187954
rect 222562 187718 222646 187954
rect 222882 187718 258326 187954
rect 258562 187718 258646 187954
rect 258882 187718 294326 187954
rect 294562 187718 294646 187954
rect 294882 187718 330326 187954
rect 330562 187718 330646 187954
rect 330882 187718 366326 187954
rect 366562 187718 366646 187954
rect 366882 187718 402326 187954
rect 402562 187718 402646 187954
rect 402882 187718 438326 187954
rect 438562 187718 438646 187954
rect 438882 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 592650 187954
rect -8726 187634 592650 187718
rect -8726 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 78326 187634
rect 78562 187398 78646 187634
rect 78882 187398 114326 187634
rect 114562 187398 114646 187634
rect 114882 187398 150326 187634
rect 150562 187398 150646 187634
rect 150882 187398 186326 187634
rect 186562 187398 186646 187634
rect 186882 187398 222326 187634
rect 222562 187398 222646 187634
rect 222882 187398 258326 187634
rect 258562 187398 258646 187634
rect 258882 187398 294326 187634
rect 294562 187398 294646 187634
rect 294882 187398 330326 187634
rect 330562 187398 330646 187634
rect 330882 187398 366326 187634
rect 366562 187398 366646 187634
rect 366882 187398 402326 187634
rect 402562 187398 402646 187634
rect 402882 187398 438326 187634
rect 438562 187398 438646 187634
rect 438882 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 592650 187634
rect -8726 187366 592650 187398
rect -8726 183454 592650 183486
rect -8726 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 592650 183454
rect -8726 183134 592650 183218
rect -8726 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 592650 183134
rect -8726 182866 592650 182898
rect -8726 178954 592650 178986
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 69326 178954
rect 69562 178718 69646 178954
rect 69882 178718 105326 178954
rect 105562 178718 105646 178954
rect 105882 178718 141326 178954
rect 141562 178718 141646 178954
rect 141882 178718 177326 178954
rect 177562 178718 177646 178954
rect 177882 178718 213326 178954
rect 213562 178718 213646 178954
rect 213882 178718 249326 178954
rect 249562 178718 249646 178954
rect 249882 178718 285326 178954
rect 285562 178718 285646 178954
rect 285882 178718 321326 178954
rect 321562 178718 321646 178954
rect 321882 178718 357326 178954
rect 357562 178718 357646 178954
rect 357882 178718 393326 178954
rect 393562 178718 393646 178954
rect 393882 178718 429326 178954
rect 429562 178718 429646 178954
rect 429882 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect -8726 178634 592650 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 69326 178634
rect 69562 178398 69646 178634
rect 69882 178398 105326 178634
rect 105562 178398 105646 178634
rect 105882 178398 141326 178634
rect 141562 178398 141646 178634
rect 141882 178398 177326 178634
rect 177562 178398 177646 178634
rect 177882 178398 213326 178634
rect 213562 178398 213646 178634
rect 213882 178398 249326 178634
rect 249562 178398 249646 178634
rect 249882 178398 285326 178634
rect 285562 178398 285646 178634
rect 285882 178398 321326 178634
rect 321562 178398 321646 178634
rect 321882 178398 357326 178634
rect 357562 178398 357646 178634
rect 357882 178398 393326 178634
rect 393562 178398 393646 178634
rect 393882 178398 429326 178634
rect 429562 178398 429646 178634
rect 429882 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect -8726 178366 592650 178398
rect -8726 174454 592650 174486
rect -8726 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 64826 174454
rect 65062 174218 65146 174454
rect 65382 174218 100826 174454
rect 101062 174218 101146 174454
rect 101382 174218 208826 174454
rect 209062 174218 209146 174454
rect 209382 174218 244826 174454
rect 245062 174218 245146 174454
rect 245382 174218 280826 174454
rect 281062 174218 281146 174454
rect 281382 174218 316826 174454
rect 317062 174218 317146 174454
rect 317382 174218 352826 174454
rect 353062 174218 353146 174454
rect 353382 174218 388826 174454
rect 389062 174218 389146 174454
rect 389382 174218 424826 174454
rect 425062 174218 425146 174454
rect 425382 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 592650 174454
rect -8726 174134 592650 174218
rect -8726 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 64826 174134
rect 65062 173898 65146 174134
rect 65382 173898 100826 174134
rect 101062 173898 101146 174134
rect 101382 173898 208826 174134
rect 209062 173898 209146 174134
rect 209382 173898 244826 174134
rect 245062 173898 245146 174134
rect 245382 173898 280826 174134
rect 281062 173898 281146 174134
rect 281382 173898 316826 174134
rect 317062 173898 317146 174134
rect 317382 173898 352826 174134
rect 353062 173898 353146 174134
rect 353382 173898 388826 174134
rect 389062 173898 389146 174134
rect 389382 173898 424826 174134
rect 425062 173898 425146 174134
rect 425382 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 592650 174134
rect -8726 173866 592650 173898
rect -8726 169954 592650 169986
rect -8726 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 60326 169954
rect 60562 169718 60646 169954
rect 60882 169718 96326 169954
rect 96562 169718 96646 169954
rect 96882 169718 204326 169954
rect 204562 169718 204646 169954
rect 204882 169718 240326 169954
rect 240562 169718 240646 169954
rect 240882 169718 276326 169954
rect 276562 169718 276646 169954
rect 276882 169718 312326 169954
rect 312562 169718 312646 169954
rect 312882 169718 348326 169954
rect 348562 169718 348646 169954
rect 348882 169718 384326 169954
rect 384562 169718 384646 169954
rect 384882 169718 420326 169954
rect 420562 169718 420646 169954
rect 420882 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 592650 169954
rect -8726 169634 592650 169718
rect -8726 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 60326 169634
rect 60562 169398 60646 169634
rect 60882 169398 96326 169634
rect 96562 169398 96646 169634
rect 96882 169398 204326 169634
rect 204562 169398 204646 169634
rect 204882 169398 240326 169634
rect 240562 169398 240646 169634
rect 240882 169398 276326 169634
rect 276562 169398 276646 169634
rect 276882 169398 312326 169634
rect 312562 169398 312646 169634
rect 312882 169398 348326 169634
rect 348562 169398 348646 169634
rect 348882 169398 384326 169634
rect 384562 169398 384646 169634
rect 384882 169398 420326 169634
rect 420562 169398 420646 169634
rect 420882 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 592650 169634
rect -8726 169366 592650 169398
rect -8726 165454 592650 165486
rect -8726 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 592650 165454
rect -8726 165134 592650 165218
rect -8726 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 592650 165134
rect -8726 164866 592650 164898
rect -8726 160954 592650 160986
rect -8726 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 87326 160954
rect 87562 160718 87646 160954
rect 87882 160718 123326 160954
rect 123562 160718 123646 160954
rect 123882 160718 159326 160954
rect 159562 160718 159646 160954
rect 159882 160718 195326 160954
rect 195562 160718 195646 160954
rect 195882 160718 231326 160954
rect 231562 160718 231646 160954
rect 231882 160718 267326 160954
rect 267562 160718 267646 160954
rect 267882 160718 303326 160954
rect 303562 160718 303646 160954
rect 303882 160718 339326 160954
rect 339562 160718 339646 160954
rect 339882 160718 375326 160954
rect 375562 160718 375646 160954
rect 375882 160718 411326 160954
rect 411562 160718 411646 160954
rect 411882 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 592650 160954
rect -8726 160634 592650 160718
rect -8726 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 87326 160634
rect 87562 160398 87646 160634
rect 87882 160398 123326 160634
rect 123562 160398 123646 160634
rect 123882 160398 159326 160634
rect 159562 160398 159646 160634
rect 159882 160398 195326 160634
rect 195562 160398 195646 160634
rect 195882 160398 231326 160634
rect 231562 160398 231646 160634
rect 231882 160398 267326 160634
rect 267562 160398 267646 160634
rect 267882 160398 303326 160634
rect 303562 160398 303646 160634
rect 303882 160398 339326 160634
rect 339562 160398 339646 160634
rect 339882 160398 375326 160634
rect 375562 160398 375646 160634
rect 375882 160398 411326 160634
rect 411562 160398 411646 160634
rect 411882 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 592650 160634
rect -8726 160366 592650 160398
rect -8726 156454 592650 156486
rect -8726 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 82826 156454
rect 83062 156218 83146 156454
rect 83382 156218 118826 156454
rect 119062 156218 119146 156454
rect 119382 156218 154826 156454
rect 155062 156218 155146 156454
rect 155382 156218 190826 156454
rect 191062 156218 191146 156454
rect 191382 156218 226826 156454
rect 227062 156218 227146 156454
rect 227382 156218 262826 156454
rect 263062 156218 263146 156454
rect 263382 156218 298826 156454
rect 299062 156218 299146 156454
rect 299382 156218 334826 156454
rect 335062 156218 335146 156454
rect 335382 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 592650 156454
rect -8726 156134 592650 156218
rect -8726 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 82826 156134
rect 83062 155898 83146 156134
rect 83382 155898 118826 156134
rect 119062 155898 119146 156134
rect 119382 155898 154826 156134
rect 155062 155898 155146 156134
rect 155382 155898 190826 156134
rect 191062 155898 191146 156134
rect 191382 155898 226826 156134
rect 227062 155898 227146 156134
rect 227382 155898 262826 156134
rect 263062 155898 263146 156134
rect 263382 155898 298826 156134
rect 299062 155898 299146 156134
rect 299382 155898 334826 156134
rect 335062 155898 335146 156134
rect 335382 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 592650 156134
rect -8726 155866 592650 155898
rect -8726 151954 592650 151986
rect -8726 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 78326 151954
rect 78562 151718 78646 151954
rect 78882 151718 114326 151954
rect 114562 151718 114646 151954
rect 114882 151718 150326 151954
rect 150562 151718 150646 151954
rect 150882 151718 186326 151954
rect 186562 151718 186646 151954
rect 186882 151718 222326 151954
rect 222562 151718 222646 151954
rect 222882 151718 258326 151954
rect 258562 151718 258646 151954
rect 258882 151718 294326 151954
rect 294562 151718 294646 151954
rect 294882 151718 330326 151954
rect 330562 151718 330646 151954
rect 330882 151718 366326 151954
rect 366562 151718 366646 151954
rect 366882 151718 402326 151954
rect 402562 151718 402646 151954
rect 402882 151718 438326 151954
rect 438562 151718 438646 151954
rect 438882 151718 474326 151954
rect 474562 151718 474646 151954
rect 474882 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 592650 151954
rect -8726 151634 592650 151718
rect -8726 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 78326 151634
rect 78562 151398 78646 151634
rect 78882 151398 114326 151634
rect 114562 151398 114646 151634
rect 114882 151398 150326 151634
rect 150562 151398 150646 151634
rect 150882 151398 186326 151634
rect 186562 151398 186646 151634
rect 186882 151398 222326 151634
rect 222562 151398 222646 151634
rect 222882 151398 258326 151634
rect 258562 151398 258646 151634
rect 258882 151398 294326 151634
rect 294562 151398 294646 151634
rect 294882 151398 330326 151634
rect 330562 151398 330646 151634
rect 330882 151398 366326 151634
rect 366562 151398 366646 151634
rect 366882 151398 402326 151634
rect 402562 151398 402646 151634
rect 402882 151398 438326 151634
rect 438562 151398 438646 151634
rect 438882 151398 474326 151634
rect 474562 151398 474646 151634
rect 474882 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 592650 151634
rect -8726 151366 592650 151398
rect -8726 147454 592650 147486
rect -8726 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 592650 147454
rect -8726 147134 592650 147218
rect -8726 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 592650 147134
rect -8726 146866 592650 146898
rect -8726 142954 592650 142986
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 69326 142954
rect 69562 142718 69646 142954
rect 69882 142718 105326 142954
rect 105562 142718 105646 142954
rect 105882 142718 141326 142954
rect 141562 142718 141646 142954
rect 141882 142718 177326 142954
rect 177562 142718 177646 142954
rect 177882 142718 213326 142954
rect 213562 142718 213646 142954
rect 213882 142718 249326 142954
rect 249562 142718 249646 142954
rect 249882 142718 285326 142954
rect 285562 142718 285646 142954
rect 285882 142718 321326 142954
rect 321562 142718 321646 142954
rect 321882 142718 357326 142954
rect 357562 142718 357646 142954
rect 357882 142718 393326 142954
rect 393562 142718 393646 142954
rect 393882 142718 429326 142954
rect 429562 142718 429646 142954
rect 429882 142718 465326 142954
rect 465562 142718 465646 142954
rect 465882 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect -8726 142634 592650 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 69326 142634
rect 69562 142398 69646 142634
rect 69882 142398 105326 142634
rect 105562 142398 105646 142634
rect 105882 142398 141326 142634
rect 141562 142398 141646 142634
rect 141882 142398 177326 142634
rect 177562 142398 177646 142634
rect 177882 142398 213326 142634
rect 213562 142398 213646 142634
rect 213882 142398 249326 142634
rect 249562 142398 249646 142634
rect 249882 142398 285326 142634
rect 285562 142398 285646 142634
rect 285882 142398 321326 142634
rect 321562 142398 321646 142634
rect 321882 142398 357326 142634
rect 357562 142398 357646 142634
rect 357882 142398 393326 142634
rect 393562 142398 393646 142634
rect 393882 142398 429326 142634
rect 429562 142398 429646 142634
rect 429882 142398 465326 142634
rect 465562 142398 465646 142634
rect 465882 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect -8726 142366 592650 142398
rect -8726 138454 592650 138486
rect -8726 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 64826 138454
rect 65062 138218 65146 138454
rect 65382 138218 100826 138454
rect 101062 138218 101146 138454
rect 101382 138218 208826 138454
rect 209062 138218 209146 138454
rect 209382 138218 244826 138454
rect 245062 138218 245146 138454
rect 245382 138218 280826 138454
rect 281062 138218 281146 138454
rect 281382 138218 316826 138454
rect 317062 138218 317146 138454
rect 317382 138218 352826 138454
rect 353062 138218 353146 138454
rect 353382 138218 388826 138454
rect 389062 138218 389146 138454
rect 389382 138218 424826 138454
rect 425062 138218 425146 138454
rect 425382 138218 460826 138454
rect 461062 138218 461146 138454
rect 461382 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 592650 138454
rect -8726 138134 592650 138218
rect -8726 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 64826 138134
rect 65062 137898 65146 138134
rect 65382 137898 100826 138134
rect 101062 137898 101146 138134
rect 101382 137898 208826 138134
rect 209062 137898 209146 138134
rect 209382 137898 244826 138134
rect 245062 137898 245146 138134
rect 245382 137898 280826 138134
rect 281062 137898 281146 138134
rect 281382 137898 316826 138134
rect 317062 137898 317146 138134
rect 317382 137898 352826 138134
rect 353062 137898 353146 138134
rect 353382 137898 388826 138134
rect 389062 137898 389146 138134
rect 389382 137898 424826 138134
rect 425062 137898 425146 138134
rect 425382 137898 460826 138134
rect 461062 137898 461146 138134
rect 461382 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 592650 138134
rect -8726 137866 592650 137898
rect -8726 133954 592650 133986
rect -8726 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 60326 133954
rect 60562 133718 60646 133954
rect 60882 133718 96326 133954
rect 96562 133718 96646 133954
rect 96882 133718 204326 133954
rect 204562 133718 204646 133954
rect 204882 133718 240326 133954
rect 240562 133718 240646 133954
rect 240882 133718 276326 133954
rect 276562 133718 276646 133954
rect 276882 133718 312326 133954
rect 312562 133718 312646 133954
rect 312882 133718 348326 133954
rect 348562 133718 348646 133954
rect 348882 133718 384326 133954
rect 384562 133718 384646 133954
rect 384882 133718 420326 133954
rect 420562 133718 420646 133954
rect 420882 133718 456326 133954
rect 456562 133718 456646 133954
rect 456882 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 592650 133954
rect -8726 133634 592650 133718
rect -8726 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 60326 133634
rect 60562 133398 60646 133634
rect 60882 133398 96326 133634
rect 96562 133398 96646 133634
rect 96882 133398 204326 133634
rect 204562 133398 204646 133634
rect 204882 133398 240326 133634
rect 240562 133398 240646 133634
rect 240882 133398 276326 133634
rect 276562 133398 276646 133634
rect 276882 133398 312326 133634
rect 312562 133398 312646 133634
rect 312882 133398 348326 133634
rect 348562 133398 348646 133634
rect 348882 133398 384326 133634
rect 384562 133398 384646 133634
rect 384882 133398 420326 133634
rect 420562 133398 420646 133634
rect 420882 133398 456326 133634
rect 456562 133398 456646 133634
rect 456882 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 592650 133634
rect -8726 133366 592650 133398
rect -8726 129454 592650 129486
rect -8726 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 592650 129454
rect -8726 129134 592650 129218
rect -8726 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 592650 129134
rect -8726 128866 592650 128898
rect -8726 124954 592650 124986
rect -8726 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 87326 124954
rect 87562 124718 87646 124954
rect 87882 124718 195326 124954
rect 195562 124718 195646 124954
rect 195882 124718 231326 124954
rect 231562 124718 231646 124954
rect 231882 124718 267326 124954
rect 267562 124718 267646 124954
rect 267882 124718 303326 124954
rect 303562 124718 303646 124954
rect 303882 124718 339326 124954
rect 339562 124718 339646 124954
rect 339882 124718 375326 124954
rect 375562 124718 375646 124954
rect 375882 124718 411326 124954
rect 411562 124718 411646 124954
rect 411882 124718 447326 124954
rect 447562 124718 447646 124954
rect 447882 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 592650 124954
rect -8726 124634 592650 124718
rect -8726 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 87326 124634
rect 87562 124398 87646 124634
rect 87882 124398 195326 124634
rect 195562 124398 195646 124634
rect 195882 124398 231326 124634
rect 231562 124398 231646 124634
rect 231882 124398 267326 124634
rect 267562 124398 267646 124634
rect 267882 124398 303326 124634
rect 303562 124398 303646 124634
rect 303882 124398 339326 124634
rect 339562 124398 339646 124634
rect 339882 124398 375326 124634
rect 375562 124398 375646 124634
rect 375882 124398 411326 124634
rect 411562 124398 411646 124634
rect 411882 124398 447326 124634
rect 447562 124398 447646 124634
rect 447882 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 592650 124634
rect -8726 124366 592650 124398
rect -8726 120454 592650 120486
rect -8726 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 82826 120454
rect 83062 120218 83146 120454
rect 83382 120218 226826 120454
rect 227062 120218 227146 120454
rect 227382 120218 262826 120454
rect 263062 120218 263146 120454
rect 263382 120218 298826 120454
rect 299062 120218 299146 120454
rect 299382 120218 334826 120454
rect 335062 120218 335146 120454
rect 335382 120218 370826 120454
rect 371062 120218 371146 120454
rect 371382 120218 406826 120454
rect 407062 120218 407146 120454
rect 407382 120218 442826 120454
rect 443062 120218 443146 120454
rect 443382 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 592650 120454
rect -8726 120134 592650 120218
rect -8726 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 82826 120134
rect 83062 119898 83146 120134
rect 83382 119898 226826 120134
rect 227062 119898 227146 120134
rect 227382 119898 262826 120134
rect 263062 119898 263146 120134
rect 263382 119898 298826 120134
rect 299062 119898 299146 120134
rect 299382 119898 334826 120134
rect 335062 119898 335146 120134
rect 335382 119898 370826 120134
rect 371062 119898 371146 120134
rect 371382 119898 406826 120134
rect 407062 119898 407146 120134
rect 407382 119898 442826 120134
rect 443062 119898 443146 120134
rect 443382 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 592650 120134
rect -8726 119866 592650 119898
rect -8726 115954 592650 115986
rect -8726 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 78326 115954
rect 78562 115718 78646 115954
rect 78882 115718 114326 115954
rect 114562 115718 114646 115954
rect 114882 115718 139610 115954
rect 139846 115718 170330 115954
rect 170566 115718 222326 115954
rect 222562 115718 222646 115954
rect 222882 115718 258326 115954
rect 258562 115718 258646 115954
rect 258882 115718 294326 115954
rect 294562 115718 294646 115954
rect 294882 115718 330326 115954
rect 330562 115718 330646 115954
rect 330882 115718 366326 115954
rect 366562 115718 366646 115954
rect 366882 115718 402326 115954
rect 402562 115718 402646 115954
rect 402882 115718 438326 115954
rect 438562 115718 438646 115954
rect 438882 115718 474326 115954
rect 474562 115718 474646 115954
rect 474882 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 592650 115954
rect -8726 115634 592650 115718
rect -8726 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 78326 115634
rect 78562 115398 78646 115634
rect 78882 115398 114326 115634
rect 114562 115398 114646 115634
rect 114882 115398 139610 115634
rect 139846 115398 170330 115634
rect 170566 115398 222326 115634
rect 222562 115398 222646 115634
rect 222882 115398 258326 115634
rect 258562 115398 258646 115634
rect 258882 115398 294326 115634
rect 294562 115398 294646 115634
rect 294882 115398 330326 115634
rect 330562 115398 330646 115634
rect 330882 115398 366326 115634
rect 366562 115398 366646 115634
rect 366882 115398 402326 115634
rect 402562 115398 402646 115634
rect 402882 115398 438326 115634
rect 438562 115398 438646 115634
rect 438882 115398 474326 115634
rect 474562 115398 474646 115634
rect 474882 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 592650 115634
rect -8726 115366 592650 115398
rect -8726 111454 592650 111486
rect -8726 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 124250 111454
rect 124486 111218 154970 111454
rect 155206 111218 185690 111454
rect 185926 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 592650 111454
rect -8726 111134 592650 111218
rect -8726 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 124250 111134
rect 124486 110898 154970 111134
rect 155206 110898 185690 111134
rect 185926 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 592650 111134
rect -8726 110866 592650 110898
rect -8726 106954 592650 106986
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 69326 106954
rect 69562 106718 69646 106954
rect 69882 106718 105326 106954
rect 105562 106718 105646 106954
rect 105882 106718 213326 106954
rect 213562 106718 213646 106954
rect 213882 106718 249326 106954
rect 249562 106718 249646 106954
rect 249882 106718 285326 106954
rect 285562 106718 285646 106954
rect 285882 106718 321326 106954
rect 321562 106718 321646 106954
rect 321882 106718 357326 106954
rect 357562 106718 357646 106954
rect 357882 106718 393326 106954
rect 393562 106718 393646 106954
rect 393882 106718 429326 106954
rect 429562 106718 429646 106954
rect 429882 106718 465326 106954
rect 465562 106718 465646 106954
rect 465882 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect -8726 106634 592650 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 69326 106634
rect 69562 106398 69646 106634
rect 69882 106398 105326 106634
rect 105562 106398 105646 106634
rect 105882 106398 213326 106634
rect 213562 106398 213646 106634
rect 213882 106398 249326 106634
rect 249562 106398 249646 106634
rect 249882 106398 285326 106634
rect 285562 106398 285646 106634
rect 285882 106398 321326 106634
rect 321562 106398 321646 106634
rect 321882 106398 357326 106634
rect 357562 106398 357646 106634
rect 357882 106398 393326 106634
rect 393562 106398 393646 106634
rect 393882 106398 429326 106634
rect 429562 106398 429646 106634
rect 429882 106398 465326 106634
rect 465562 106398 465646 106634
rect 465882 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect -8726 106366 592650 106398
rect -8726 102454 592650 102486
rect -8726 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 64826 102454
rect 65062 102218 65146 102454
rect 65382 102218 100826 102454
rect 101062 102218 101146 102454
rect 101382 102218 208826 102454
rect 209062 102218 209146 102454
rect 209382 102218 244826 102454
rect 245062 102218 245146 102454
rect 245382 102218 280826 102454
rect 281062 102218 281146 102454
rect 281382 102218 316826 102454
rect 317062 102218 317146 102454
rect 317382 102218 352826 102454
rect 353062 102218 353146 102454
rect 353382 102218 388826 102454
rect 389062 102218 389146 102454
rect 389382 102218 424826 102454
rect 425062 102218 425146 102454
rect 425382 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 592650 102454
rect -8726 102134 592650 102218
rect -8726 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 64826 102134
rect 65062 101898 65146 102134
rect 65382 101898 100826 102134
rect 101062 101898 101146 102134
rect 101382 101898 208826 102134
rect 209062 101898 209146 102134
rect 209382 101898 244826 102134
rect 245062 101898 245146 102134
rect 245382 101898 280826 102134
rect 281062 101898 281146 102134
rect 281382 101898 316826 102134
rect 317062 101898 317146 102134
rect 317382 101898 352826 102134
rect 353062 101898 353146 102134
rect 353382 101898 388826 102134
rect 389062 101898 389146 102134
rect 389382 101898 424826 102134
rect 425062 101898 425146 102134
rect 425382 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 592650 102134
rect -8726 101866 592650 101898
rect -8726 97954 592650 97986
rect -8726 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 60326 97954
rect 60562 97718 60646 97954
rect 60882 97718 96326 97954
rect 96562 97718 96646 97954
rect 96882 97718 204326 97954
rect 204562 97718 204646 97954
rect 204882 97718 240326 97954
rect 240562 97718 240646 97954
rect 240882 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 312326 97954
rect 312562 97718 312646 97954
rect 312882 97718 348326 97954
rect 348562 97718 348646 97954
rect 348882 97718 384326 97954
rect 384562 97718 384646 97954
rect 384882 97718 420326 97954
rect 420562 97718 420646 97954
rect 420882 97718 456326 97954
rect 456562 97718 456646 97954
rect 456882 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 592650 97954
rect -8726 97634 592650 97718
rect -8726 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 60326 97634
rect 60562 97398 60646 97634
rect 60882 97398 96326 97634
rect 96562 97398 96646 97634
rect 96882 97398 204326 97634
rect 204562 97398 204646 97634
rect 204882 97398 240326 97634
rect 240562 97398 240646 97634
rect 240882 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 312326 97634
rect 312562 97398 312646 97634
rect 312882 97398 348326 97634
rect 348562 97398 348646 97634
rect 348882 97398 384326 97634
rect 384562 97398 384646 97634
rect 384882 97398 420326 97634
rect 420562 97398 420646 97634
rect 420882 97398 456326 97634
rect 456562 97398 456646 97634
rect 456882 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 592650 97634
rect -8726 97366 592650 97398
rect -8726 93454 592650 93486
rect -8726 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 592650 93454
rect -8726 93134 592650 93218
rect -8726 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 592650 93134
rect -8726 92866 592650 92898
rect -8726 88954 592650 88986
rect -8726 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 87326 88954
rect 87562 88718 87646 88954
rect 87882 88718 195326 88954
rect 195562 88718 195646 88954
rect 195882 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 303326 88954
rect 303562 88718 303646 88954
rect 303882 88718 339326 88954
rect 339562 88718 339646 88954
rect 339882 88718 375326 88954
rect 375562 88718 375646 88954
rect 375882 88718 411326 88954
rect 411562 88718 411646 88954
rect 411882 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 592650 88954
rect -8726 88634 592650 88718
rect -8726 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 87326 88634
rect 87562 88398 87646 88634
rect 87882 88398 195326 88634
rect 195562 88398 195646 88634
rect 195882 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 303326 88634
rect 303562 88398 303646 88634
rect 303882 88398 339326 88634
rect 339562 88398 339646 88634
rect 339882 88398 375326 88634
rect 375562 88398 375646 88634
rect 375882 88398 411326 88634
rect 411562 88398 411646 88634
rect 411882 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 592650 88634
rect -8726 88366 592650 88398
rect -8726 84454 592650 84486
rect -8726 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 82826 84454
rect 83062 84218 83146 84454
rect 83382 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 298826 84454
rect 299062 84218 299146 84454
rect 299382 84218 334826 84454
rect 335062 84218 335146 84454
rect 335382 84218 370826 84454
rect 371062 84218 371146 84454
rect 371382 84218 406826 84454
rect 407062 84218 407146 84454
rect 407382 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 592650 84454
rect -8726 84134 592650 84218
rect -8726 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 82826 84134
rect 83062 83898 83146 84134
rect 83382 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 298826 84134
rect 299062 83898 299146 84134
rect 299382 83898 334826 84134
rect 335062 83898 335146 84134
rect 335382 83898 370826 84134
rect 371062 83898 371146 84134
rect 371382 83898 406826 84134
rect 407062 83898 407146 84134
rect 407382 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 592650 84134
rect -8726 83866 592650 83898
rect -8726 79954 592650 79986
rect -8726 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 78326 79954
rect 78562 79718 78646 79954
rect 78882 79718 114326 79954
rect 114562 79718 114646 79954
rect 114882 79718 222326 79954
rect 222562 79718 222646 79954
rect 222882 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 330326 79954
rect 330562 79718 330646 79954
rect 330882 79718 366326 79954
rect 366562 79718 366646 79954
rect 366882 79718 402326 79954
rect 402562 79718 402646 79954
rect 402882 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 592650 79954
rect -8726 79634 592650 79718
rect -8726 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 78326 79634
rect 78562 79398 78646 79634
rect 78882 79398 114326 79634
rect 114562 79398 114646 79634
rect 114882 79398 222326 79634
rect 222562 79398 222646 79634
rect 222882 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 330326 79634
rect 330562 79398 330646 79634
rect 330882 79398 366326 79634
rect 366562 79398 366646 79634
rect 366882 79398 402326 79634
rect 402562 79398 402646 79634
rect 402882 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 592650 79634
rect -8726 79366 592650 79398
rect -8726 75454 592650 75486
rect -8726 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 592650 75454
rect -8726 75134 592650 75218
rect -8726 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 592650 75134
rect -8726 74866 592650 74898
rect -8726 70954 592650 70986
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 69326 70954
rect 69562 70718 69646 70954
rect 69882 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 213326 70954
rect 213562 70718 213646 70954
rect 213882 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 321326 70954
rect 321562 70718 321646 70954
rect 321882 70718 357326 70954
rect 357562 70718 357646 70954
rect 357882 70718 393326 70954
rect 393562 70718 393646 70954
rect 393882 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect -8726 70634 592650 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 69326 70634
rect 69562 70398 69646 70634
rect 69882 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 213326 70634
rect 213562 70398 213646 70634
rect 213882 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 321326 70634
rect 321562 70398 321646 70634
rect 321882 70398 357326 70634
rect 357562 70398 357646 70634
rect 357882 70398 393326 70634
rect 393562 70398 393646 70634
rect 393882 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect -8726 70366 592650 70398
rect -8726 66454 592650 66486
rect -8726 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 64826 66454
rect 65062 66218 65146 66454
rect 65382 66218 100826 66454
rect 101062 66218 101146 66454
rect 101382 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 316826 66454
rect 317062 66218 317146 66454
rect 317382 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 592650 66454
rect -8726 66134 592650 66218
rect -8726 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 64826 66134
rect 65062 65898 65146 66134
rect 65382 65898 100826 66134
rect 101062 65898 101146 66134
rect 101382 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 316826 66134
rect 317062 65898 317146 66134
rect 317382 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 592650 66134
rect -8726 65866 592650 65898
rect -8726 61954 592650 61986
rect -8726 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 60326 61954
rect 60562 61718 60646 61954
rect 60882 61718 96326 61954
rect 96562 61718 96646 61954
rect 96882 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 312326 61954
rect 312562 61718 312646 61954
rect 312882 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 592650 61954
rect -8726 61634 592650 61718
rect -8726 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 60326 61634
rect 60562 61398 60646 61634
rect 60882 61398 96326 61634
rect 96562 61398 96646 61634
rect 96882 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 312326 61634
rect 312562 61398 312646 61634
rect 312882 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 592650 61634
rect -8726 61366 592650 61398
rect -8726 57454 592650 57486
rect -8726 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 592650 57454
rect -8726 57134 592650 57218
rect -8726 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 592650 57134
rect -8726 56866 592650 56898
rect -8726 52954 592650 52986
rect -8726 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 592650 52954
rect -8726 52634 592650 52718
rect -8726 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 592650 52634
rect -8726 52366 592650 52398
rect -8726 48454 592650 48486
rect -8726 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 592650 48454
rect -8726 48134 592650 48218
rect -8726 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 592650 48134
rect -8726 47866 592650 47898
rect -8726 43954 592650 43986
rect -8726 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 592650 43954
rect -8726 43634 592650 43718
rect -8726 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 592650 43634
rect -8726 43366 592650 43398
rect -8726 39454 592650 39486
rect -8726 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 592650 39454
rect -8726 39134 592650 39218
rect -8726 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 592650 39134
rect -8726 38866 592650 38898
rect -8726 34954 592650 34986
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect -8726 34634 592650 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect -8726 34366 592650 34398
rect -8726 30454 592650 30486
rect -8726 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 592650 30454
rect -8726 30134 592650 30218
rect -8726 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 592650 30134
rect -8726 29866 592650 29898
rect -8726 25954 592650 25986
rect -8726 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 592650 25954
rect -8726 25634 592650 25718
rect -8726 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 592650 25634
rect -8726 25366 592650 25398
rect -8726 21454 592650 21486
rect -8726 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 592650 21454
rect -8726 21134 592650 21218
rect -8726 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 592650 21134
rect -8726 20866 592650 20898
rect -8726 16954 592650 16986
rect -8726 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 592650 16954
rect -8726 16634 592650 16718
rect -8726 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 592650 16634
rect -8726 16366 592650 16398
rect -8726 12454 592650 12486
rect -8726 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 592650 12454
rect -8726 12134 592650 12218
rect -8726 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 592650 12134
rect -8726 11866 592650 11898
rect -8726 7954 592650 7986
rect -8726 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 592650 7954
rect -8726 7634 592650 7718
rect -8726 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 592650 7634
rect -8726 7366 592650 7398
rect -8726 3454 592650 3486
rect -8726 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 592650 3454
rect -8726 3134 592650 3218
rect -8726 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 592650 3134
rect -8726 2866 592650 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 19826 -4186
rect 20062 -4422 20146 -4186
rect 20382 -4422 55826 -4186
rect 56062 -4422 56146 -4186
rect 56382 -4422 91826 -4186
rect 92062 -4422 92146 -4186
rect 92382 -4422 127826 -4186
rect 128062 -4422 128146 -4186
rect 128382 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 19826 -4506
rect 20062 -4742 20146 -4506
rect 20382 -4742 55826 -4506
rect 56062 -4742 56146 -4506
rect 56382 -4742 91826 -4506
rect 92062 -4742 92146 -4506
rect 92382 -4742 127826 -4506
rect 128062 -4742 128146 -4506
rect 128382 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 24326 -5146
rect 24562 -5382 24646 -5146
rect 24882 -5382 60326 -5146
rect 60562 -5382 60646 -5146
rect 60882 -5382 96326 -5146
rect 96562 -5382 96646 -5146
rect 96882 -5382 132326 -5146
rect 132562 -5382 132646 -5146
rect 132882 -5382 168326 -5146
rect 168562 -5382 168646 -5146
rect 168882 -5382 204326 -5146
rect 204562 -5382 204646 -5146
rect 204882 -5382 240326 -5146
rect 240562 -5382 240646 -5146
rect 240882 -5382 276326 -5146
rect 276562 -5382 276646 -5146
rect 276882 -5382 312326 -5146
rect 312562 -5382 312646 -5146
rect 312882 -5382 348326 -5146
rect 348562 -5382 348646 -5146
rect 348882 -5382 384326 -5146
rect 384562 -5382 384646 -5146
rect 384882 -5382 420326 -5146
rect 420562 -5382 420646 -5146
rect 420882 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 24326 -5466
rect 24562 -5702 24646 -5466
rect 24882 -5702 60326 -5466
rect 60562 -5702 60646 -5466
rect 60882 -5702 96326 -5466
rect 96562 -5702 96646 -5466
rect 96882 -5702 132326 -5466
rect 132562 -5702 132646 -5466
rect 132882 -5702 168326 -5466
rect 168562 -5702 168646 -5466
rect 168882 -5702 204326 -5466
rect 204562 -5702 204646 -5466
rect 204882 -5702 240326 -5466
rect 240562 -5702 240646 -5466
rect 240882 -5702 276326 -5466
rect 276562 -5702 276646 -5466
rect 276882 -5702 312326 -5466
rect 312562 -5702 312646 -5466
rect 312882 -5702 348326 -5466
rect 348562 -5702 348646 -5466
rect 348882 -5702 384326 -5466
rect 384562 -5702 384646 -5466
rect 384882 -5702 420326 -5466
rect 420562 -5702 420646 -5466
rect 420882 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 28826 -6106
rect 29062 -6342 29146 -6106
rect 29382 -6342 64826 -6106
rect 65062 -6342 65146 -6106
rect 65382 -6342 100826 -6106
rect 101062 -6342 101146 -6106
rect 101382 -6342 136826 -6106
rect 137062 -6342 137146 -6106
rect 137382 -6342 172826 -6106
rect 173062 -6342 173146 -6106
rect 173382 -6342 208826 -6106
rect 209062 -6342 209146 -6106
rect 209382 -6342 244826 -6106
rect 245062 -6342 245146 -6106
rect 245382 -6342 280826 -6106
rect 281062 -6342 281146 -6106
rect 281382 -6342 316826 -6106
rect 317062 -6342 317146 -6106
rect 317382 -6342 352826 -6106
rect 353062 -6342 353146 -6106
rect 353382 -6342 388826 -6106
rect 389062 -6342 389146 -6106
rect 389382 -6342 424826 -6106
rect 425062 -6342 425146 -6106
rect 425382 -6342 460826 -6106
rect 461062 -6342 461146 -6106
rect 461382 -6342 496826 -6106
rect 497062 -6342 497146 -6106
rect 497382 -6342 532826 -6106
rect 533062 -6342 533146 -6106
rect 533382 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 28826 -6426
rect 29062 -6662 29146 -6426
rect 29382 -6662 64826 -6426
rect 65062 -6662 65146 -6426
rect 65382 -6662 100826 -6426
rect 101062 -6662 101146 -6426
rect 101382 -6662 136826 -6426
rect 137062 -6662 137146 -6426
rect 137382 -6662 172826 -6426
rect 173062 -6662 173146 -6426
rect 173382 -6662 208826 -6426
rect 209062 -6662 209146 -6426
rect 209382 -6662 244826 -6426
rect 245062 -6662 245146 -6426
rect 245382 -6662 280826 -6426
rect 281062 -6662 281146 -6426
rect 281382 -6662 316826 -6426
rect 317062 -6662 317146 -6426
rect 317382 -6662 352826 -6426
rect 353062 -6662 353146 -6426
rect 353382 -6662 388826 -6426
rect 389062 -6662 389146 -6426
rect 389382 -6662 424826 -6426
rect 425062 -6662 425146 -6426
rect 425382 -6662 460826 -6426
rect 461062 -6662 461146 -6426
rect 461382 -6662 496826 -6426
rect 497062 -6662 497146 -6426
rect 497382 -6662 532826 -6426
rect 533062 -6662 533146 -6426
rect 533382 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 33326 -7066
rect 33562 -7302 33646 -7066
rect 33882 -7302 69326 -7066
rect 69562 -7302 69646 -7066
rect 69882 -7302 105326 -7066
rect 105562 -7302 105646 -7066
rect 105882 -7302 141326 -7066
rect 141562 -7302 141646 -7066
rect 141882 -7302 177326 -7066
rect 177562 -7302 177646 -7066
rect 177882 -7302 213326 -7066
rect 213562 -7302 213646 -7066
rect 213882 -7302 249326 -7066
rect 249562 -7302 249646 -7066
rect 249882 -7302 285326 -7066
rect 285562 -7302 285646 -7066
rect 285882 -7302 321326 -7066
rect 321562 -7302 321646 -7066
rect 321882 -7302 357326 -7066
rect 357562 -7302 357646 -7066
rect 357882 -7302 393326 -7066
rect 393562 -7302 393646 -7066
rect 393882 -7302 429326 -7066
rect 429562 -7302 429646 -7066
rect 429882 -7302 465326 -7066
rect 465562 -7302 465646 -7066
rect 465882 -7302 501326 -7066
rect 501562 -7302 501646 -7066
rect 501882 -7302 537326 -7066
rect 537562 -7302 537646 -7066
rect 537882 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 33326 -7386
rect 33562 -7622 33646 -7386
rect 33882 -7622 69326 -7386
rect 69562 -7622 69646 -7386
rect 69882 -7622 105326 -7386
rect 105562 -7622 105646 -7386
rect 105882 -7622 141326 -7386
rect 141562 -7622 141646 -7386
rect 141882 -7622 177326 -7386
rect 177562 -7622 177646 -7386
rect 177882 -7622 213326 -7386
rect 213562 -7622 213646 -7386
rect 213882 -7622 249326 -7386
rect 249562 -7622 249646 -7386
rect 249882 -7622 285326 -7386
rect 285562 -7622 285646 -7386
rect 285882 -7622 321326 -7386
rect 321562 -7622 321646 -7386
rect 321882 -7622 357326 -7386
rect 357562 -7622 357646 -7386
rect 357882 -7622 393326 -7386
rect 393562 -7622 393646 -7386
rect 393882 -7622 429326 -7386
rect 429562 -7622 429646 -7386
rect 429882 -7622 465326 -7386
rect 465562 -7622 465646 -7386
rect 465882 -7622 501326 -7386
rect 501562 -7622 501646 -7386
rect 501882 -7622 537326 -7386
rect 537562 -7622 537646 -7386
rect 537882 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use pixel_macro  pixel_macro0
timestamp 0
transform 1 0 120000 0 1 200000
box 1066 0 68854 60000
use rlbp_macro  rlbp_macro0
timestamp 0
transform 1 0 120000 0 1 80000
box 1066 0 68854 60000
<< labels >>
flabel metal3 s 583520 285276 584960 285516 0 FreeSans 960 0 0 0 analog_io[0]
port 0 nsew signal bidirectional
flabel metal2 s 446098 703520 446210 704960 0 FreeSans 448 90 0 0 analog_io[10]
port 1 nsew signal bidirectional
flabel metal2 s 381146 703520 381258 704960 0 FreeSans 448 90 0 0 analog_io[11]
port 2 nsew signal bidirectional
flabel metal2 s 316286 703520 316398 704960 0 FreeSans 448 90 0 0 analog_io[12]
port 3 nsew signal bidirectional
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 448 90 0 0 analog_io[13]
port 4 nsew signal bidirectional
flabel metal2 s 186474 703520 186586 704960 0 FreeSans 448 90 0 0 analog_io[14]
port 5 nsew signal bidirectional
flabel metal2 s 121614 703520 121726 704960 0 FreeSans 448 90 0 0 analog_io[15]
port 6 nsew signal bidirectional
flabel metal2 s 56754 703520 56866 704960 0 FreeSans 448 90 0 0 analog_io[16]
port 7 nsew signal bidirectional
flabel metal3 s -960 697220 480 697460 0 FreeSans 960 0 0 0 analog_io[17]
port 8 nsew signal bidirectional
flabel metal3 s -960 644996 480 645236 0 FreeSans 960 0 0 0 analog_io[18]
port 9 nsew signal bidirectional
flabel metal3 s -960 592908 480 593148 0 FreeSans 960 0 0 0 analog_io[19]
port 10 nsew signal bidirectional
flabel metal3 s 583520 338452 584960 338692 0 FreeSans 960 0 0 0 analog_io[1]
port 11 nsew signal bidirectional
flabel metal3 s -960 540684 480 540924 0 FreeSans 960 0 0 0 analog_io[20]
port 12 nsew signal bidirectional
flabel metal3 s -960 488596 480 488836 0 FreeSans 960 0 0 0 analog_io[21]
port 13 nsew signal bidirectional
flabel metal3 s -960 436508 480 436748 0 FreeSans 960 0 0 0 analog_io[22]
port 14 nsew signal bidirectional
flabel metal3 s -960 384284 480 384524 0 FreeSans 960 0 0 0 analog_io[23]
port 15 nsew signal bidirectional
flabel metal3 s -960 332196 480 332436 0 FreeSans 960 0 0 0 analog_io[24]
port 16 nsew signal bidirectional
flabel metal3 s -960 279972 480 280212 0 FreeSans 960 0 0 0 analog_io[25]
port 17 nsew signal bidirectional
flabel metal3 s -960 227884 480 228124 0 FreeSans 960 0 0 0 analog_io[26]
port 18 nsew signal bidirectional
flabel metal3 s -960 175796 480 176036 0 FreeSans 960 0 0 0 analog_io[27]
port 19 nsew signal bidirectional
flabel metal3 s -960 123572 480 123812 0 FreeSans 960 0 0 0 analog_io[28]
port 20 nsew signal bidirectional
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 960 0 0 0 analog_io[2]
port 21 nsew signal bidirectional
flabel metal3 s 583520 444668 584960 444908 0 FreeSans 960 0 0 0 analog_io[3]
port 22 nsew signal bidirectional
flabel metal3 s 583520 497844 584960 498084 0 FreeSans 960 0 0 0 analog_io[4]
port 23 nsew signal bidirectional
flabel metal3 s 583520 551020 584960 551260 0 FreeSans 960 0 0 0 analog_io[5]
port 24 nsew signal bidirectional
flabel metal3 s 583520 604060 584960 604300 0 FreeSans 960 0 0 0 analog_io[6]
port 25 nsew signal bidirectional
flabel metal3 s 583520 657236 584960 657476 0 FreeSans 960 0 0 0 analog_io[7]
port 26 nsew signal bidirectional
flabel metal2 s 575818 703520 575930 704960 0 FreeSans 448 90 0 0 analog_io[8]
port 27 nsew signal bidirectional
flabel metal2 s 510958 703520 511070 704960 0 FreeSans 448 90 0 0 analog_io[9]
port 28 nsew signal bidirectional
flabel metal3 s 583520 6476 584960 6716 0 FreeSans 960 0 0 0 io_in[0]
port 29 nsew signal input
flabel metal3 s 583520 457996 584960 458236 0 FreeSans 960 0 0 0 io_in[10]
port 30 nsew signal input
flabel metal3 s 583520 511172 584960 511412 0 FreeSans 960 0 0 0 io_in[11]
port 31 nsew signal input
flabel metal3 s 583520 564212 584960 564452 0 FreeSans 960 0 0 0 io_in[12]
port 32 nsew signal input
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 960 0 0 0 io_in[13]
port 33 nsew signal input
flabel metal3 s 583520 670564 584960 670804 0 FreeSans 960 0 0 0 io_in[14]
port 34 nsew signal input
flabel metal2 s 559626 703520 559738 704960 0 FreeSans 448 90 0 0 io_in[15]
port 35 nsew signal input
flabel metal2 s 494766 703520 494878 704960 0 FreeSans 448 90 0 0 io_in[16]
port 36 nsew signal input
flabel metal2 s 429814 703520 429926 704960 0 FreeSans 448 90 0 0 io_in[17]
port 37 nsew signal input
flabel metal2 s 364954 703520 365066 704960 0 FreeSans 448 90 0 0 io_in[18]
port 38 nsew signal input
flabel metal2 s 300094 703520 300206 704960 0 FreeSans 448 90 0 0 io_in[19]
port 39 nsew signal input
flabel metal3 s 583520 46188 584960 46428 0 FreeSans 960 0 0 0 io_in[1]
port 40 nsew signal input
flabel metal2 s 235142 703520 235254 704960 0 FreeSans 448 90 0 0 io_in[20]
port 41 nsew signal input
flabel metal2 s 170282 703520 170394 704960 0 FreeSans 448 90 0 0 io_in[21]
port 42 nsew signal input
flabel metal2 s 105422 703520 105534 704960 0 FreeSans 448 90 0 0 io_in[22]
port 43 nsew signal input
flabel metal2 s 40470 703520 40582 704960 0 FreeSans 448 90 0 0 io_in[23]
port 44 nsew signal input
flabel metal3 s -960 684164 480 684404 0 FreeSans 960 0 0 0 io_in[24]
port 45 nsew signal input
flabel metal3 s -960 631940 480 632180 0 FreeSans 960 0 0 0 io_in[25]
port 46 nsew signal input
flabel metal3 s -960 579852 480 580092 0 FreeSans 960 0 0 0 io_in[26]
port 47 nsew signal input
flabel metal3 s -960 527764 480 528004 0 FreeSans 960 0 0 0 io_in[27]
port 48 nsew signal input
flabel metal3 s -960 475540 480 475780 0 FreeSans 960 0 0 0 io_in[28]
port 49 nsew signal input
flabel metal3 s -960 423452 480 423692 0 FreeSans 960 0 0 0 io_in[29]
port 50 nsew signal input
flabel metal3 s 583520 86036 584960 86276 0 FreeSans 960 0 0 0 io_in[2]
port 51 nsew signal input
flabel metal3 s -960 371228 480 371468 0 FreeSans 960 0 0 0 io_in[30]
port 52 nsew signal input
flabel metal3 s -960 319140 480 319380 0 FreeSans 960 0 0 0 io_in[31]
port 53 nsew signal input
flabel metal3 s -960 267052 480 267292 0 FreeSans 960 0 0 0 io_in[32]
port 54 nsew signal input
flabel metal3 s -960 214828 480 215068 0 FreeSans 960 0 0 0 io_in[33]
port 55 nsew signal input
flabel metal3 s -960 162740 480 162980 0 FreeSans 960 0 0 0 io_in[34]
port 56 nsew signal input
flabel metal3 s -960 110516 480 110756 0 FreeSans 960 0 0 0 io_in[35]
port 57 nsew signal input
flabel metal3 s -960 71484 480 71724 0 FreeSans 960 0 0 0 io_in[36]
port 58 nsew signal input
flabel metal3 s -960 32316 480 32556 0 FreeSans 960 0 0 0 io_in[37]
port 59 nsew signal input
flabel metal3 s 583520 125884 584960 126124 0 FreeSans 960 0 0 0 io_in[3]
port 60 nsew signal input
flabel metal3 s 583520 165732 584960 165972 0 FreeSans 960 0 0 0 io_in[4]
port 61 nsew signal input
flabel metal3 s 583520 205580 584960 205820 0 FreeSans 960 0 0 0 io_in[5]
port 62 nsew signal input
flabel metal3 s 583520 245428 584960 245668 0 FreeSans 960 0 0 0 io_in[6]
port 63 nsew signal input
flabel metal3 s 583520 298604 584960 298844 0 FreeSans 960 0 0 0 io_in[7]
port 64 nsew signal input
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 960 0 0 0 io_in[8]
port 65 nsew signal input
flabel metal3 s 583520 404820 584960 405060 0 FreeSans 960 0 0 0 io_in[9]
port 66 nsew signal input
flabel metal3 s 583520 32996 584960 33236 0 FreeSans 960 0 0 0 io_oeb[0]
port 67 nsew signal tristate
flabel metal3 s 583520 484516 584960 484756 0 FreeSans 960 0 0 0 io_oeb[10]
port 68 nsew signal tristate
flabel metal3 s 583520 537692 584960 537932 0 FreeSans 960 0 0 0 io_oeb[11]
port 69 nsew signal tristate
flabel metal3 s 583520 590868 584960 591108 0 FreeSans 960 0 0 0 io_oeb[12]
port 70 nsew signal tristate
flabel metal3 s 583520 643908 584960 644148 0 FreeSans 960 0 0 0 io_oeb[13]
port 71 nsew signal tristate
flabel metal3 s 583520 697084 584960 697324 0 FreeSans 960 0 0 0 io_oeb[14]
port 72 nsew signal tristate
flabel metal2 s 527150 703520 527262 704960 0 FreeSans 448 90 0 0 io_oeb[15]
port 73 nsew signal tristate
flabel metal2 s 462290 703520 462402 704960 0 FreeSans 448 90 0 0 io_oeb[16]
port 74 nsew signal tristate
flabel metal2 s 397430 703520 397542 704960 0 FreeSans 448 90 0 0 io_oeb[17]
port 75 nsew signal tristate
flabel metal2 s 332478 703520 332590 704960 0 FreeSans 448 90 0 0 io_oeb[18]
port 76 nsew signal tristate
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 448 90 0 0 io_oeb[19]
port 77 nsew signal tristate
flabel metal3 s 583520 72844 584960 73084 0 FreeSans 960 0 0 0 io_oeb[1]
port 78 nsew signal tristate
flabel metal2 s 202758 703520 202870 704960 0 FreeSans 448 90 0 0 io_oeb[20]
port 79 nsew signal tristate
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 448 90 0 0 io_oeb[21]
port 80 nsew signal tristate
flabel metal2 s 72946 703520 73058 704960 0 FreeSans 448 90 0 0 io_oeb[22]
port 81 nsew signal tristate
flabel metal2 s 8086 703520 8198 704960 0 FreeSans 448 90 0 0 io_oeb[23]
port 82 nsew signal tristate
flabel metal3 s -960 658052 480 658292 0 FreeSans 960 0 0 0 io_oeb[24]
port 83 nsew signal tristate
flabel metal3 s -960 605964 480 606204 0 FreeSans 960 0 0 0 io_oeb[25]
port 84 nsew signal tristate
flabel metal3 s -960 553740 480 553980 0 FreeSans 960 0 0 0 io_oeb[26]
port 85 nsew signal tristate
flabel metal3 s -960 501652 480 501892 0 FreeSans 960 0 0 0 io_oeb[27]
port 86 nsew signal tristate
flabel metal3 s -960 449428 480 449668 0 FreeSans 960 0 0 0 io_oeb[28]
port 87 nsew signal tristate
flabel metal3 s -960 397340 480 397580 0 FreeSans 960 0 0 0 io_oeb[29]
port 88 nsew signal tristate
flabel metal3 s 583520 112692 584960 112932 0 FreeSans 960 0 0 0 io_oeb[2]
port 89 nsew signal tristate
flabel metal3 s -960 345252 480 345492 0 FreeSans 960 0 0 0 io_oeb[30]
port 90 nsew signal tristate
flabel metal3 s -960 293028 480 293268 0 FreeSans 960 0 0 0 io_oeb[31]
port 91 nsew signal tristate
flabel metal3 s -960 240940 480 241180 0 FreeSans 960 0 0 0 io_oeb[32]
port 92 nsew signal tristate
flabel metal3 s -960 188716 480 188956 0 FreeSans 960 0 0 0 io_oeb[33]
port 93 nsew signal tristate
flabel metal3 s -960 136628 480 136868 0 FreeSans 960 0 0 0 io_oeb[34]
port 94 nsew signal tristate
flabel metal3 s -960 84540 480 84780 0 FreeSans 960 0 0 0 io_oeb[35]
port 95 nsew signal tristate
flabel metal3 s -960 45372 480 45612 0 FreeSans 960 0 0 0 io_oeb[36]
port 96 nsew signal tristate
flabel metal3 s -960 6340 480 6580 0 FreeSans 960 0 0 0 io_oeb[37]
port 97 nsew signal tristate
flabel metal3 s 583520 152540 584960 152780 0 FreeSans 960 0 0 0 io_oeb[3]
port 98 nsew signal tristate
flabel metal3 s 583520 192388 584960 192628 0 FreeSans 960 0 0 0 io_oeb[4]
port 99 nsew signal tristate
flabel metal3 s 583520 232236 584960 232476 0 FreeSans 960 0 0 0 io_oeb[5]
port 100 nsew signal tristate
flabel metal3 s 583520 272084 584960 272324 0 FreeSans 960 0 0 0 io_oeb[6]
port 101 nsew signal tristate
flabel metal3 s 583520 325124 584960 325364 0 FreeSans 960 0 0 0 io_oeb[7]
port 102 nsew signal tristate
flabel metal3 s 583520 378300 584960 378540 0 FreeSans 960 0 0 0 io_oeb[8]
port 103 nsew signal tristate
flabel metal3 s 583520 431476 584960 431716 0 FreeSans 960 0 0 0 io_oeb[9]
port 104 nsew signal tristate
flabel metal3 s 583520 19668 584960 19908 0 FreeSans 960 0 0 0 io_out[0]
port 105 nsew signal tristate
flabel metal3 s 583520 471324 584960 471564 0 FreeSans 960 0 0 0 io_out[10]
port 106 nsew signal tristate
flabel metal3 s 583520 524364 584960 524604 0 FreeSans 960 0 0 0 io_out[11]
port 107 nsew signal tristate
flabel metal3 s 583520 577540 584960 577780 0 FreeSans 960 0 0 0 io_out[12]
port 108 nsew signal tristate
flabel metal3 s 583520 630716 584960 630956 0 FreeSans 960 0 0 0 io_out[13]
port 109 nsew signal tristate
flabel metal3 s 583520 683756 584960 683996 0 FreeSans 960 0 0 0 io_out[14]
port 110 nsew signal tristate
flabel metal2 s 543434 703520 543546 704960 0 FreeSans 448 90 0 0 io_out[15]
port 111 nsew signal tristate
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 448 90 0 0 io_out[16]
port 112 nsew signal tristate
flabel metal2 s 413622 703520 413734 704960 0 FreeSans 448 90 0 0 io_out[17]
port 113 nsew signal tristate
flabel metal2 s 348762 703520 348874 704960 0 FreeSans 448 90 0 0 io_out[18]
port 114 nsew signal tristate
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 448 90 0 0 io_out[19]
port 115 nsew signal tristate
flabel metal3 s 583520 59516 584960 59756 0 FreeSans 960 0 0 0 io_out[1]
port 116 nsew signal tristate
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 448 90 0 0 io_out[20]
port 117 nsew signal tristate
flabel metal2 s 154090 703520 154202 704960 0 FreeSans 448 90 0 0 io_out[21]
port 118 nsew signal tristate
flabel metal2 s 89138 703520 89250 704960 0 FreeSans 448 90 0 0 io_out[22]
port 119 nsew signal tristate
flabel metal2 s 24278 703520 24390 704960 0 FreeSans 448 90 0 0 io_out[23]
port 120 nsew signal tristate
flabel metal3 s -960 671108 480 671348 0 FreeSans 960 0 0 0 io_out[24]
port 121 nsew signal tristate
flabel metal3 s -960 619020 480 619260 0 FreeSans 960 0 0 0 io_out[25]
port 122 nsew signal tristate
flabel metal3 s -960 566796 480 567036 0 FreeSans 960 0 0 0 io_out[26]
port 123 nsew signal tristate
flabel metal3 s -960 514708 480 514948 0 FreeSans 960 0 0 0 io_out[27]
port 124 nsew signal tristate
flabel metal3 s -960 462484 480 462724 0 FreeSans 960 0 0 0 io_out[28]
port 125 nsew signal tristate
flabel metal3 s -960 410396 480 410636 0 FreeSans 960 0 0 0 io_out[29]
port 126 nsew signal tristate
flabel metal3 s 583520 99364 584960 99604 0 FreeSans 960 0 0 0 io_out[2]
port 127 nsew signal tristate
flabel metal3 s -960 358308 480 358548 0 FreeSans 960 0 0 0 io_out[30]
port 128 nsew signal tristate
flabel metal3 s -960 306084 480 306324 0 FreeSans 960 0 0 0 io_out[31]
port 129 nsew signal tristate
flabel metal3 s -960 253996 480 254236 0 FreeSans 960 0 0 0 io_out[32]
port 130 nsew signal tristate
flabel metal3 s -960 201772 480 202012 0 FreeSans 960 0 0 0 io_out[33]
port 131 nsew signal tristate
flabel metal3 s -960 149684 480 149924 0 FreeSans 960 0 0 0 io_out[34]
port 132 nsew signal tristate
flabel metal3 s -960 97460 480 97700 0 FreeSans 960 0 0 0 io_out[35]
port 133 nsew signal tristate
flabel metal3 s -960 58428 480 58668 0 FreeSans 960 0 0 0 io_out[36]
port 134 nsew signal tristate
flabel metal3 s -960 19260 480 19500 0 FreeSans 960 0 0 0 io_out[37]
port 135 nsew signal tristate
flabel metal3 s 583520 139212 584960 139452 0 FreeSans 960 0 0 0 io_out[3]
port 136 nsew signal tristate
flabel metal3 s 583520 179060 584960 179300 0 FreeSans 960 0 0 0 io_out[4]
port 137 nsew signal tristate
flabel metal3 s 583520 218908 584960 219148 0 FreeSans 960 0 0 0 io_out[5]
port 138 nsew signal tristate
flabel metal3 s 583520 258756 584960 258996 0 FreeSans 960 0 0 0 io_out[6]
port 139 nsew signal tristate
flabel metal3 s 583520 311932 584960 312172 0 FreeSans 960 0 0 0 io_out[7]
port 140 nsew signal tristate
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 960 0 0 0 io_out[8]
port 141 nsew signal tristate
flabel metal3 s 583520 418148 584960 418388 0 FreeSans 960 0 0 0 io_out[9]
port 142 nsew signal tristate
flabel metal2 s 125846 -960 125958 480 0 FreeSans 448 90 0 0 la_data_in[0]
port 143 nsew signal input
flabel metal2 s 480506 -960 480618 480 0 FreeSans 448 90 0 0 la_data_in[100]
port 144 nsew signal input
flabel metal2 s 484002 -960 484114 480 0 FreeSans 448 90 0 0 la_data_in[101]
port 145 nsew signal input
flabel metal2 s 487590 -960 487702 480 0 FreeSans 448 90 0 0 la_data_in[102]
port 146 nsew signal input
flabel metal2 s 491086 -960 491198 480 0 FreeSans 448 90 0 0 la_data_in[103]
port 147 nsew signal input
flabel metal2 s 494674 -960 494786 480 0 FreeSans 448 90 0 0 la_data_in[104]
port 148 nsew signal input
flabel metal2 s 498170 -960 498282 480 0 FreeSans 448 90 0 0 la_data_in[105]
port 149 nsew signal input
flabel metal2 s 501758 -960 501870 480 0 FreeSans 448 90 0 0 la_data_in[106]
port 150 nsew signal input
flabel metal2 s 505346 -960 505458 480 0 FreeSans 448 90 0 0 la_data_in[107]
port 151 nsew signal input
flabel metal2 s 508842 -960 508954 480 0 FreeSans 448 90 0 0 la_data_in[108]
port 152 nsew signal input
flabel metal2 s 512430 -960 512542 480 0 FreeSans 448 90 0 0 la_data_in[109]
port 153 nsew signal input
flabel metal2 s 161266 -960 161378 480 0 FreeSans 448 90 0 0 la_data_in[10]
port 154 nsew signal input
flabel metal2 s 515926 -960 516038 480 0 FreeSans 448 90 0 0 la_data_in[110]
port 155 nsew signal input
flabel metal2 s 519514 -960 519626 480 0 FreeSans 448 90 0 0 la_data_in[111]
port 156 nsew signal input
flabel metal2 s 523010 -960 523122 480 0 FreeSans 448 90 0 0 la_data_in[112]
port 157 nsew signal input
flabel metal2 s 526598 -960 526710 480 0 FreeSans 448 90 0 0 la_data_in[113]
port 158 nsew signal input
flabel metal2 s 530094 -960 530206 480 0 FreeSans 448 90 0 0 la_data_in[114]
port 159 nsew signal input
flabel metal2 s 533682 -960 533794 480 0 FreeSans 448 90 0 0 la_data_in[115]
port 160 nsew signal input
flabel metal2 s 537178 -960 537290 480 0 FreeSans 448 90 0 0 la_data_in[116]
port 161 nsew signal input
flabel metal2 s 540766 -960 540878 480 0 FreeSans 448 90 0 0 la_data_in[117]
port 162 nsew signal input
flabel metal2 s 544354 -960 544466 480 0 FreeSans 448 90 0 0 la_data_in[118]
port 163 nsew signal input
flabel metal2 s 547850 -960 547962 480 0 FreeSans 448 90 0 0 la_data_in[119]
port 164 nsew signal input
flabel metal2 s 164854 -960 164966 480 0 FreeSans 448 90 0 0 la_data_in[11]
port 165 nsew signal input
flabel metal2 s 551438 -960 551550 480 0 FreeSans 448 90 0 0 la_data_in[120]
port 166 nsew signal input
flabel metal2 s 554934 -960 555046 480 0 FreeSans 448 90 0 0 la_data_in[121]
port 167 nsew signal input
flabel metal2 s 558522 -960 558634 480 0 FreeSans 448 90 0 0 la_data_in[122]
port 168 nsew signal input
flabel metal2 s 562018 -960 562130 480 0 FreeSans 448 90 0 0 la_data_in[123]
port 169 nsew signal input
flabel metal2 s 565606 -960 565718 480 0 FreeSans 448 90 0 0 la_data_in[124]
port 170 nsew signal input
flabel metal2 s 569102 -960 569214 480 0 FreeSans 448 90 0 0 la_data_in[125]
port 171 nsew signal input
flabel metal2 s 572690 -960 572802 480 0 FreeSans 448 90 0 0 la_data_in[126]
port 172 nsew signal input
flabel metal2 s 576278 -960 576390 480 0 FreeSans 448 90 0 0 la_data_in[127]
port 173 nsew signal input
flabel metal2 s 168350 -960 168462 480 0 FreeSans 448 90 0 0 la_data_in[12]
port 174 nsew signal input
flabel metal2 s 171938 -960 172050 480 0 FreeSans 448 90 0 0 la_data_in[13]
port 175 nsew signal input
flabel metal2 s 175434 -960 175546 480 0 FreeSans 448 90 0 0 la_data_in[14]
port 176 nsew signal input
flabel metal2 s 179022 -960 179134 480 0 FreeSans 448 90 0 0 la_data_in[15]
port 177 nsew signal input
flabel metal2 s 182518 -960 182630 480 0 FreeSans 448 90 0 0 la_data_in[16]
port 178 nsew signal input
flabel metal2 s 186106 -960 186218 480 0 FreeSans 448 90 0 0 la_data_in[17]
port 179 nsew signal input
flabel metal2 s 189694 -960 189806 480 0 FreeSans 448 90 0 0 la_data_in[18]
port 180 nsew signal input
flabel metal2 s 193190 -960 193302 480 0 FreeSans 448 90 0 0 la_data_in[19]
port 181 nsew signal input
flabel metal2 s 129342 -960 129454 480 0 FreeSans 448 90 0 0 la_data_in[1]
port 182 nsew signal input
flabel metal2 s 196778 -960 196890 480 0 FreeSans 448 90 0 0 la_data_in[20]
port 183 nsew signal input
flabel metal2 s 200274 -960 200386 480 0 FreeSans 448 90 0 0 la_data_in[21]
port 184 nsew signal input
flabel metal2 s 203862 -960 203974 480 0 FreeSans 448 90 0 0 la_data_in[22]
port 185 nsew signal input
flabel metal2 s 207358 -960 207470 480 0 FreeSans 448 90 0 0 la_data_in[23]
port 186 nsew signal input
flabel metal2 s 210946 -960 211058 480 0 FreeSans 448 90 0 0 la_data_in[24]
port 187 nsew signal input
flabel metal2 s 214442 -960 214554 480 0 FreeSans 448 90 0 0 la_data_in[25]
port 188 nsew signal input
flabel metal2 s 218030 -960 218142 480 0 FreeSans 448 90 0 0 la_data_in[26]
port 189 nsew signal input
flabel metal2 s 221526 -960 221638 480 0 FreeSans 448 90 0 0 la_data_in[27]
port 190 nsew signal input
flabel metal2 s 225114 -960 225226 480 0 FreeSans 448 90 0 0 la_data_in[28]
port 191 nsew signal input
flabel metal2 s 228702 -960 228814 480 0 FreeSans 448 90 0 0 la_data_in[29]
port 192 nsew signal input
flabel metal2 s 132930 -960 133042 480 0 FreeSans 448 90 0 0 la_data_in[2]
port 193 nsew signal input
flabel metal2 s 232198 -960 232310 480 0 FreeSans 448 90 0 0 la_data_in[30]
port 194 nsew signal input
flabel metal2 s 235786 -960 235898 480 0 FreeSans 448 90 0 0 la_data_in[31]
port 195 nsew signal input
flabel metal2 s 239282 -960 239394 480 0 FreeSans 448 90 0 0 la_data_in[32]
port 196 nsew signal input
flabel metal2 s 242870 -960 242982 480 0 FreeSans 448 90 0 0 la_data_in[33]
port 197 nsew signal input
flabel metal2 s 246366 -960 246478 480 0 FreeSans 448 90 0 0 la_data_in[34]
port 198 nsew signal input
flabel metal2 s 249954 -960 250066 480 0 FreeSans 448 90 0 0 la_data_in[35]
port 199 nsew signal input
flabel metal2 s 253450 -960 253562 480 0 FreeSans 448 90 0 0 la_data_in[36]
port 200 nsew signal input
flabel metal2 s 257038 -960 257150 480 0 FreeSans 448 90 0 0 la_data_in[37]
port 201 nsew signal input
flabel metal2 s 260626 -960 260738 480 0 FreeSans 448 90 0 0 la_data_in[38]
port 202 nsew signal input
flabel metal2 s 264122 -960 264234 480 0 FreeSans 448 90 0 0 la_data_in[39]
port 203 nsew signal input
flabel metal2 s 136426 -960 136538 480 0 FreeSans 448 90 0 0 la_data_in[3]
port 204 nsew signal input
flabel metal2 s 267710 -960 267822 480 0 FreeSans 448 90 0 0 la_data_in[40]
port 205 nsew signal input
flabel metal2 s 271206 -960 271318 480 0 FreeSans 448 90 0 0 la_data_in[41]
port 206 nsew signal input
flabel metal2 s 274794 -960 274906 480 0 FreeSans 448 90 0 0 la_data_in[42]
port 207 nsew signal input
flabel metal2 s 278290 -960 278402 480 0 FreeSans 448 90 0 0 la_data_in[43]
port 208 nsew signal input
flabel metal2 s 281878 -960 281990 480 0 FreeSans 448 90 0 0 la_data_in[44]
port 209 nsew signal input
flabel metal2 s 285374 -960 285486 480 0 FreeSans 448 90 0 0 la_data_in[45]
port 210 nsew signal input
flabel metal2 s 288962 -960 289074 480 0 FreeSans 448 90 0 0 la_data_in[46]
port 211 nsew signal input
flabel metal2 s 292550 -960 292662 480 0 FreeSans 448 90 0 0 la_data_in[47]
port 212 nsew signal input
flabel metal2 s 296046 -960 296158 480 0 FreeSans 448 90 0 0 la_data_in[48]
port 213 nsew signal input
flabel metal2 s 299634 -960 299746 480 0 FreeSans 448 90 0 0 la_data_in[49]
port 214 nsew signal input
flabel metal2 s 140014 -960 140126 480 0 FreeSans 448 90 0 0 la_data_in[4]
port 215 nsew signal input
flabel metal2 s 303130 -960 303242 480 0 FreeSans 448 90 0 0 la_data_in[50]
port 216 nsew signal input
flabel metal2 s 306718 -960 306830 480 0 FreeSans 448 90 0 0 la_data_in[51]
port 217 nsew signal input
flabel metal2 s 310214 -960 310326 480 0 FreeSans 448 90 0 0 la_data_in[52]
port 218 nsew signal input
flabel metal2 s 313802 -960 313914 480 0 FreeSans 448 90 0 0 la_data_in[53]
port 219 nsew signal input
flabel metal2 s 317298 -960 317410 480 0 FreeSans 448 90 0 0 la_data_in[54]
port 220 nsew signal input
flabel metal2 s 320886 -960 320998 480 0 FreeSans 448 90 0 0 la_data_in[55]
port 221 nsew signal input
flabel metal2 s 324382 -960 324494 480 0 FreeSans 448 90 0 0 la_data_in[56]
port 222 nsew signal input
flabel metal2 s 327970 -960 328082 480 0 FreeSans 448 90 0 0 la_data_in[57]
port 223 nsew signal input
flabel metal2 s 331558 -960 331670 480 0 FreeSans 448 90 0 0 la_data_in[58]
port 224 nsew signal input
flabel metal2 s 335054 -960 335166 480 0 FreeSans 448 90 0 0 la_data_in[59]
port 225 nsew signal input
flabel metal2 s 143510 -960 143622 480 0 FreeSans 448 90 0 0 la_data_in[5]
port 226 nsew signal input
flabel metal2 s 338642 -960 338754 480 0 FreeSans 448 90 0 0 la_data_in[60]
port 227 nsew signal input
flabel metal2 s 342138 -960 342250 480 0 FreeSans 448 90 0 0 la_data_in[61]
port 228 nsew signal input
flabel metal2 s 345726 -960 345838 480 0 FreeSans 448 90 0 0 la_data_in[62]
port 229 nsew signal input
flabel metal2 s 349222 -960 349334 480 0 FreeSans 448 90 0 0 la_data_in[63]
port 230 nsew signal input
flabel metal2 s 352810 -960 352922 480 0 FreeSans 448 90 0 0 la_data_in[64]
port 231 nsew signal input
flabel metal2 s 356306 -960 356418 480 0 FreeSans 448 90 0 0 la_data_in[65]
port 232 nsew signal input
flabel metal2 s 359894 -960 360006 480 0 FreeSans 448 90 0 0 la_data_in[66]
port 233 nsew signal input
flabel metal2 s 363482 -960 363594 480 0 FreeSans 448 90 0 0 la_data_in[67]
port 234 nsew signal input
flabel metal2 s 366978 -960 367090 480 0 FreeSans 448 90 0 0 la_data_in[68]
port 235 nsew signal input
flabel metal2 s 370566 -960 370678 480 0 FreeSans 448 90 0 0 la_data_in[69]
port 236 nsew signal input
flabel metal2 s 147098 -960 147210 480 0 FreeSans 448 90 0 0 la_data_in[6]
port 237 nsew signal input
flabel metal2 s 374062 -960 374174 480 0 FreeSans 448 90 0 0 la_data_in[70]
port 238 nsew signal input
flabel metal2 s 377650 -960 377762 480 0 FreeSans 448 90 0 0 la_data_in[71]
port 239 nsew signal input
flabel metal2 s 381146 -960 381258 480 0 FreeSans 448 90 0 0 la_data_in[72]
port 240 nsew signal input
flabel metal2 s 384734 -960 384846 480 0 FreeSans 448 90 0 0 la_data_in[73]
port 241 nsew signal input
flabel metal2 s 388230 -960 388342 480 0 FreeSans 448 90 0 0 la_data_in[74]
port 242 nsew signal input
flabel metal2 s 391818 -960 391930 480 0 FreeSans 448 90 0 0 la_data_in[75]
port 243 nsew signal input
flabel metal2 s 395314 -960 395426 480 0 FreeSans 448 90 0 0 la_data_in[76]
port 244 nsew signal input
flabel metal2 s 398902 -960 399014 480 0 FreeSans 448 90 0 0 la_data_in[77]
port 245 nsew signal input
flabel metal2 s 402490 -960 402602 480 0 FreeSans 448 90 0 0 la_data_in[78]
port 246 nsew signal input
flabel metal2 s 405986 -960 406098 480 0 FreeSans 448 90 0 0 la_data_in[79]
port 247 nsew signal input
flabel metal2 s 150594 -960 150706 480 0 FreeSans 448 90 0 0 la_data_in[7]
port 248 nsew signal input
flabel metal2 s 409574 -960 409686 480 0 FreeSans 448 90 0 0 la_data_in[80]
port 249 nsew signal input
flabel metal2 s 413070 -960 413182 480 0 FreeSans 448 90 0 0 la_data_in[81]
port 250 nsew signal input
flabel metal2 s 416658 -960 416770 480 0 FreeSans 448 90 0 0 la_data_in[82]
port 251 nsew signal input
flabel metal2 s 420154 -960 420266 480 0 FreeSans 448 90 0 0 la_data_in[83]
port 252 nsew signal input
flabel metal2 s 423742 -960 423854 480 0 FreeSans 448 90 0 0 la_data_in[84]
port 253 nsew signal input
flabel metal2 s 427238 -960 427350 480 0 FreeSans 448 90 0 0 la_data_in[85]
port 254 nsew signal input
flabel metal2 s 430826 -960 430938 480 0 FreeSans 448 90 0 0 la_data_in[86]
port 255 nsew signal input
flabel metal2 s 434414 -960 434526 480 0 FreeSans 448 90 0 0 la_data_in[87]
port 256 nsew signal input
flabel metal2 s 437910 -960 438022 480 0 FreeSans 448 90 0 0 la_data_in[88]
port 257 nsew signal input
flabel metal2 s 441498 -960 441610 480 0 FreeSans 448 90 0 0 la_data_in[89]
port 258 nsew signal input
flabel metal2 s 154182 -960 154294 480 0 FreeSans 448 90 0 0 la_data_in[8]
port 259 nsew signal input
flabel metal2 s 444994 -960 445106 480 0 FreeSans 448 90 0 0 la_data_in[90]
port 260 nsew signal input
flabel metal2 s 448582 -960 448694 480 0 FreeSans 448 90 0 0 la_data_in[91]
port 261 nsew signal input
flabel metal2 s 452078 -960 452190 480 0 FreeSans 448 90 0 0 la_data_in[92]
port 262 nsew signal input
flabel metal2 s 455666 -960 455778 480 0 FreeSans 448 90 0 0 la_data_in[93]
port 263 nsew signal input
flabel metal2 s 459162 -960 459274 480 0 FreeSans 448 90 0 0 la_data_in[94]
port 264 nsew signal input
flabel metal2 s 462750 -960 462862 480 0 FreeSans 448 90 0 0 la_data_in[95]
port 265 nsew signal input
flabel metal2 s 466246 -960 466358 480 0 FreeSans 448 90 0 0 la_data_in[96]
port 266 nsew signal input
flabel metal2 s 469834 -960 469946 480 0 FreeSans 448 90 0 0 la_data_in[97]
port 267 nsew signal input
flabel metal2 s 473422 -960 473534 480 0 FreeSans 448 90 0 0 la_data_in[98]
port 268 nsew signal input
flabel metal2 s 476918 -960 477030 480 0 FreeSans 448 90 0 0 la_data_in[99]
port 269 nsew signal input
flabel metal2 s 157770 -960 157882 480 0 FreeSans 448 90 0 0 la_data_in[9]
port 270 nsew signal input
flabel metal2 s 126950 -960 127062 480 0 FreeSans 448 90 0 0 la_data_out[0]
port 271 nsew signal tristate
flabel metal2 s 481702 -960 481814 480 0 FreeSans 448 90 0 0 la_data_out[100]
port 272 nsew signal tristate
flabel metal2 s 485198 -960 485310 480 0 FreeSans 448 90 0 0 la_data_out[101]
port 273 nsew signal tristate
flabel metal2 s 488786 -960 488898 480 0 FreeSans 448 90 0 0 la_data_out[102]
port 274 nsew signal tristate
flabel metal2 s 492282 -960 492394 480 0 FreeSans 448 90 0 0 la_data_out[103]
port 275 nsew signal tristate
flabel metal2 s 495870 -960 495982 480 0 FreeSans 448 90 0 0 la_data_out[104]
port 276 nsew signal tristate
flabel metal2 s 499366 -960 499478 480 0 FreeSans 448 90 0 0 la_data_out[105]
port 277 nsew signal tristate
flabel metal2 s 502954 -960 503066 480 0 FreeSans 448 90 0 0 la_data_out[106]
port 278 nsew signal tristate
flabel metal2 s 506450 -960 506562 480 0 FreeSans 448 90 0 0 la_data_out[107]
port 279 nsew signal tristate
flabel metal2 s 510038 -960 510150 480 0 FreeSans 448 90 0 0 la_data_out[108]
port 280 nsew signal tristate
flabel metal2 s 513534 -960 513646 480 0 FreeSans 448 90 0 0 la_data_out[109]
port 281 nsew signal tristate
flabel metal2 s 162462 -960 162574 480 0 FreeSans 448 90 0 0 la_data_out[10]
port 282 nsew signal tristate
flabel metal2 s 517122 -960 517234 480 0 FreeSans 448 90 0 0 la_data_out[110]
port 283 nsew signal tristate
flabel metal2 s 520710 -960 520822 480 0 FreeSans 448 90 0 0 la_data_out[111]
port 284 nsew signal tristate
flabel metal2 s 524206 -960 524318 480 0 FreeSans 448 90 0 0 la_data_out[112]
port 285 nsew signal tristate
flabel metal2 s 527794 -960 527906 480 0 FreeSans 448 90 0 0 la_data_out[113]
port 286 nsew signal tristate
flabel metal2 s 531290 -960 531402 480 0 FreeSans 448 90 0 0 la_data_out[114]
port 287 nsew signal tristate
flabel metal2 s 534878 -960 534990 480 0 FreeSans 448 90 0 0 la_data_out[115]
port 288 nsew signal tristate
flabel metal2 s 538374 -960 538486 480 0 FreeSans 448 90 0 0 la_data_out[116]
port 289 nsew signal tristate
flabel metal2 s 541962 -960 542074 480 0 FreeSans 448 90 0 0 la_data_out[117]
port 290 nsew signal tristate
flabel metal2 s 545458 -960 545570 480 0 FreeSans 448 90 0 0 la_data_out[118]
port 291 nsew signal tristate
flabel metal2 s 549046 -960 549158 480 0 FreeSans 448 90 0 0 la_data_out[119]
port 292 nsew signal tristate
flabel metal2 s 166050 -960 166162 480 0 FreeSans 448 90 0 0 la_data_out[11]
port 293 nsew signal tristate
flabel metal2 s 552634 -960 552746 480 0 FreeSans 448 90 0 0 la_data_out[120]
port 294 nsew signal tristate
flabel metal2 s 556130 -960 556242 480 0 FreeSans 448 90 0 0 la_data_out[121]
port 295 nsew signal tristate
flabel metal2 s 559718 -960 559830 480 0 FreeSans 448 90 0 0 la_data_out[122]
port 296 nsew signal tristate
flabel metal2 s 563214 -960 563326 480 0 FreeSans 448 90 0 0 la_data_out[123]
port 297 nsew signal tristate
flabel metal2 s 566802 -960 566914 480 0 FreeSans 448 90 0 0 la_data_out[124]
port 298 nsew signal tristate
flabel metal2 s 570298 -960 570410 480 0 FreeSans 448 90 0 0 la_data_out[125]
port 299 nsew signal tristate
flabel metal2 s 573886 -960 573998 480 0 FreeSans 448 90 0 0 la_data_out[126]
port 300 nsew signal tristate
flabel metal2 s 577382 -960 577494 480 0 FreeSans 448 90 0 0 la_data_out[127]
port 301 nsew signal tristate
flabel metal2 s 169546 -960 169658 480 0 FreeSans 448 90 0 0 la_data_out[12]
port 302 nsew signal tristate
flabel metal2 s 173134 -960 173246 480 0 FreeSans 448 90 0 0 la_data_out[13]
port 303 nsew signal tristate
flabel metal2 s 176630 -960 176742 480 0 FreeSans 448 90 0 0 la_data_out[14]
port 304 nsew signal tristate
flabel metal2 s 180218 -960 180330 480 0 FreeSans 448 90 0 0 la_data_out[15]
port 305 nsew signal tristate
flabel metal2 s 183714 -960 183826 480 0 FreeSans 448 90 0 0 la_data_out[16]
port 306 nsew signal tristate
flabel metal2 s 187302 -960 187414 480 0 FreeSans 448 90 0 0 la_data_out[17]
port 307 nsew signal tristate
flabel metal2 s 190798 -960 190910 480 0 FreeSans 448 90 0 0 la_data_out[18]
port 308 nsew signal tristate
flabel metal2 s 194386 -960 194498 480 0 FreeSans 448 90 0 0 la_data_out[19]
port 309 nsew signal tristate
flabel metal2 s 130538 -960 130650 480 0 FreeSans 448 90 0 0 la_data_out[1]
port 310 nsew signal tristate
flabel metal2 s 197882 -960 197994 480 0 FreeSans 448 90 0 0 la_data_out[20]
port 311 nsew signal tristate
flabel metal2 s 201470 -960 201582 480 0 FreeSans 448 90 0 0 la_data_out[21]
port 312 nsew signal tristate
flabel metal2 s 205058 -960 205170 480 0 FreeSans 448 90 0 0 la_data_out[22]
port 313 nsew signal tristate
flabel metal2 s 208554 -960 208666 480 0 FreeSans 448 90 0 0 la_data_out[23]
port 314 nsew signal tristate
flabel metal2 s 212142 -960 212254 480 0 FreeSans 448 90 0 0 la_data_out[24]
port 315 nsew signal tristate
flabel metal2 s 215638 -960 215750 480 0 FreeSans 448 90 0 0 la_data_out[25]
port 316 nsew signal tristate
flabel metal2 s 219226 -960 219338 480 0 FreeSans 448 90 0 0 la_data_out[26]
port 317 nsew signal tristate
flabel metal2 s 222722 -960 222834 480 0 FreeSans 448 90 0 0 la_data_out[27]
port 318 nsew signal tristate
flabel metal2 s 226310 -960 226422 480 0 FreeSans 448 90 0 0 la_data_out[28]
port 319 nsew signal tristate
flabel metal2 s 229806 -960 229918 480 0 FreeSans 448 90 0 0 la_data_out[29]
port 320 nsew signal tristate
flabel metal2 s 134126 -960 134238 480 0 FreeSans 448 90 0 0 la_data_out[2]
port 321 nsew signal tristate
flabel metal2 s 233394 -960 233506 480 0 FreeSans 448 90 0 0 la_data_out[30]
port 322 nsew signal tristate
flabel metal2 s 236982 -960 237094 480 0 FreeSans 448 90 0 0 la_data_out[31]
port 323 nsew signal tristate
flabel metal2 s 240478 -960 240590 480 0 FreeSans 448 90 0 0 la_data_out[32]
port 324 nsew signal tristate
flabel metal2 s 244066 -960 244178 480 0 FreeSans 448 90 0 0 la_data_out[33]
port 325 nsew signal tristate
flabel metal2 s 247562 -960 247674 480 0 FreeSans 448 90 0 0 la_data_out[34]
port 326 nsew signal tristate
flabel metal2 s 251150 -960 251262 480 0 FreeSans 448 90 0 0 la_data_out[35]
port 327 nsew signal tristate
flabel metal2 s 254646 -960 254758 480 0 FreeSans 448 90 0 0 la_data_out[36]
port 328 nsew signal tristate
flabel metal2 s 258234 -960 258346 480 0 FreeSans 448 90 0 0 la_data_out[37]
port 329 nsew signal tristate
flabel metal2 s 261730 -960 261842 480 0 FreeSans 448 90 0 0 la_data_out[38]
port 330 nsew signal tristate
flabel metal2 s 265318 -960 265430 480 0 FreeSans 448 90 0 0 la_data_out[39]
port 331 nsew signal tristate
flabel metal2 s 137622 -960 137734 480 0 FreeSans 448 90 0 0 la_data_out[3]
port 332 nsew signal tristate
flabel metal2 s 268814 -960 268926 480 0 FreeSans 448 90 0 0 la_data_out[40]
port 333 nsew signal tristate
flabel metal2 s 272402 -960 272514 480 0 FreeSans 448 90 0 0 la_data_out[41]
port 334 nsew signal tristate
flabel metal2 s 275990 -960 276102 480 0 FreeSans 448 90 0 0 la_data_out[42]
port 335 nsew signal tristate
flabel metal2 s 279486 -960 279598 480 0 FreeSans 448 90 0 0 la_data_out[43]
port 336 nsew signal tristate
flabel metal2 s 283074 -960 283186 480 0 FreeSans 448 90 0 0 la_data_out[44]
port 337 nsew signal tristate
flabel metal2 s 286570 -960 286682 480 0 FreeSans 448 90 0 0 la_data_out[45]
port 338 nsew signal tristate
flabel metal2 s 290158 -960 290270 480 0 FreeSans 448 90 0 0 la_data_out[46]
port 339 nsew signal tristate
flabel metal2 s 293654 -960 293766 480 0 FreeSans 448 90 0 0 la_data_out[47]
port 340 nsew signal tristate
flabel metal2 s 297242 -960 297354 480 0 FreeSans 448 90 0 0 la_data_out[48]
port 341 nsew signal tristate
flabel metal2 s 300738 -960 300850 480 0 FreeSans 448 90 0 0 la_data_out[49]
port 342 nsew signal tristate
flabel metal2 s 141210 -960 141322 480 0 FreeSans 448 90 0 0 la_data_out[4]
port 343 nsew signal tristate
flabel metal2 s 304326 -960 304438 480 0 FreeSans 448 90 0 0 la_data_out[50]
port 344 nsew signal tristate
flabel metal2 s 307914 -960 308026 480 0 FreeSans 448 90 0 0 la_data_out[51]
port 345 nsew signal tristate
flabel metal2 s 311410 -960 311522 480 0 FreeSans 448 90 0 0 la_data_out[52]
port 346 nsew signal tristate
flabel metal2 s 314998 -960 315110 480 0 FreeSans 448 90 0 0 la_data_out[53]
port 347 nsew signal tristate
flabel metal2 s 318494 -960 318606 480 0 FreeSans 448 90 0 0 la_data_out[54]
port 348 nsew signal tristate
flabel metal2 s 322082 -960 322194 480 0 FreeSans 448 90 0 0 la_data_out[55]
port 349 nsew signal tristate
flabel metal2 s 325578 -960 325690 480 0 FreeSans 448 90 0 0 la_data_out[56]
port 350 nsew signal tristate
flabel metal2 s 329166 -960 329278 480 0 FreeSans 448 90 0 0 la_data_out[57]
port 351 nsew signal tristate
flabel metal2 s 332662 -960 332774 480 0 FreeSans 448 90 0 0 la_data_out[58]
port 352 nsew signal tristate
flabel metal2 s 336250 -960 336362 480 0 FreeSans 448 90 0 0 la_data_out[59]
port 353 nsew signal tristate
flabel metal2 s 144706 -960 144818 480 0 FreeSans 448 90 0 0 la_data_out[5]
port 354 nsew signal tristate
flabel metal2 s 339838 -960 339950 480 0 FreeSans 448 90 0 0 la_data_out[60]
port 355 nsew signal tristate
flabel metal2 s 343334 -960 343446 480 0 FreeSans 448 90 0 0 la_data_out[61]
port 356 nsew signal tristate
flabel metal2 s 346922 -960 347034 480 0 FreeSans 448 90 0 0 la_data_out[62]
port 357 nsew signal tristate
flabel metal2 s 350418 -960 350530 480 0 FreeSans 448 90 0 0 la_data_out[63]
port 358 nsew signal tristate
flabel metal2 s 354006 -960 354118 480 0 FreeSans 448 90 0 0 la_data_out[64]
port 359 nsew signal tristate
flabel metal2 s 357502 -960 357614 480 0 FreeSans 448 90 0 0 la_data_out[65]
port 360 nsew signal tristate
flabel metal2 s 361090 -960 361202 480 0 FreeSans 448 90 0 0 la_data_out[66]
port 361 nsew signal tristate
flabel metal2 s 364586 -960 364698 480 0 FreeSans 448 90 0 0 la_data_out[67]
port 362 nsew signal tristate
flabel metal2 s 368174 -960 368286 480 0 FreeSans 448 90 0 0 la_data_out[68]
port 363 nsew signal tristate
flabel metal2 s 371670 -960 371782 480 0 FreeSans 448 90 0 0 la_data_out[69]
port 364 nsew signal tristate
flabel metal2 s 148294 -960 148406 480 0 FreeSans 448 90 0 0 la_data_out[6]
port 365 nsew signal tristate
flabel metal2 s 375258 -960 375370 480 0 FreeSans 448 90 0 0 la_data_out[70]
port 366 nsew signal tristate
flabel metal2 s 378846 -960 378958 480 0 FreeSans 448 90 0 0 la_data_out[71]
port 367 nsew signal tristate
flabel metal2 s 382342 -960 382454 480 0 FreeSans 448 90 0 0 la_data_out[72]
port 368 nsew signal tristate
flabel metal2 s 385930 -960 386042 480 0 FreeSans 448 90 0 0 la_data_out[73]
port 369 nsew signal tristate
flabel metal2 s 389426 -960 389538 480 0 FreeSans 448 90 0 0 la_data_out[74]
port 370 nsew signal tristate
flabel metal2 s 393014 -960 393126 480 0 FreeSans 448 90 0 0 la_data_out[75]
port 371 nsew signal tristate
flabel metal2 s 396510 -960 396622 480 0 FreeSans 448 90 0 0 la_data_out[76]
port 372 nsew signal tristate
flabel metal2 s 400098 -960 400210 480 0 FreeSans 448 90 0 0 la_data_out[77]
port 373 nsew signal tristate
flabel metal2 s 403594 -960 403706 480 0 FreeSans 448 90 0 0 la_data_out[78]
port 374 nsew signal tristate
flabel metal2 s 407182 -960 407294 480 0 FreeSans 448 90 0 0 la_data_out[79]
port 375 nsew signal tristate
flabel metal2 s 151790 -960 151902 480 0 FreeSans 448 90 0 0 la_data_out[7]
port 376 nsew signal tristate
flabel metal2 s 410770 -960 410882 480 0 FreeSans 448 90 0 0 la_data_out[80]
port 377 nsew signal tristate
flabel metal2 s 414266 -960 414378 480 0 FreeSans 448 90 0 0 la_data_out[81]
port 378 nsew signal tristate
flabel metal2 s 417854 -960 417966 480 0 FreeSans 448 90 0 0 la_data_out[82]
port 379 nsew signal tristate
flabel metal2 s 421350 -960 421462 480 0 FreeSans 448 90 0 0 la_data_out[83]
port 380 nsew signal tristate
flabel metal2 s 424938 -960 425050 480 0 FreeSans 448 90 0 0 la_data_out[84]
port 381 nsew signal tristate
flabel metal2 s 428434 -960 428546 480 0 FreeSans 448 90 0 0 la_data_out[85]
port 382 nsew signal tristate
flabel metal2 s 432022 -960 432134 480 0 FreeSans 448 90 0 0 la_data_out[86]
port 383 nsew signal tristate
flabel metal2 s 435518 -960 435630 480 0 FreeSans 448 90 0 0 la_data_out[87]
port 384 nsew signal tristate
flabel metal2 s 439106 -960 439218 480 0 FreeSans 448 90 0 0 la_data_out[88]
port 385 nsew signal tristate
flabel metal2 s 442602 -960 442714 480 0 FreeSans 448 90 0 0 la_data_out[89]
port 386 nsew signal tristate
flabel metal2 s 155378 -960 155490 480 0 FreeSans 448 90 0 0 la_data_out[8]
port 387 nsew signal tristate
flabel metal2 s 446190 -960 446302 480 0 FreeSans 448 90 0 0 la_data_out[90]
port 388 nsew signal tristate
flabel metal2 s 449778 -960 449890 480 0 FreeSans 448 90 0 0 la_data_out[91]
port 389 nsew signal tristate
flabel metal2 s 453274 -960 453386 480 0 FreeSans 448 90 0 0 la_data_out[92]
port 390 nsew signal tristate
flabel metal2 s 456862 -960 456974 480 0 FreeSans 448 90 0 0 la_data_out[93]
port 391 nsew signal tristate
flabel metal2 s 460358 -960 460470 480 0 FreeSans 448 90 0 0 la_data_out[94]
port 392 nsew signal tristate
flabel metal2 s 463946 -960 464058 480 0 FreeSans 448 90 0 0 la_data_out[95]
port 393 nsew signal tristate
flabel metal2 s 467442 -960 467554 480 0 FreeSans 448 90 0 0 la_data_out[96]
port 394 nsew signal tristate
flabel metal2 s 471030 -960 471142 480 0 FreeSans 448 90 0 0 la_data_out[97]
port 395 nsew signal tristate
flabel metal2 s 474526 -960 474638 480 0 FreeSans 448 90 0 0 la_data_out[98]
port 396 nsew signal tristate
flabel metal2 s 478114 -960 478226 480 0 FreeSans 448 90 0 0 la_data_out[99]
port 397 nsew signal tristate
flabel metal2 s 158874 -960 158986 480 0 FreeSans 448 90 0 0 la_data_out[9]
port 398 nsew signal tristate
flabel metal2 s 128146 -960 128258 480 0 FreeSans 448 90 0 0 la_oenb[0]
port 399 nsew signal input
flabel metal2 s 482806 -960 482918 480 0 FreeSans 448 90 0 0 la_oenb[100]
port 400 nsew signal input
flabel metal2 s 486394 -960 486506 480 0 FreeSans 448 90 0 0 la_oenb[101]
port 401 nsew signal input
flabel metal2 s 489890 -960 490002 480 0 FreeSans 448 90 0 0 la_oenb[102]
port 402 nsew signal input
flabel metal2 s 493478 -960 493590 480 0 FreeSans 448 90 0 0 la_oenb[103]
port 403 nsew signal input
flabel metal2 s 497066 -960 497178 480 0 FreeSans 448 90 0 0 la_oenb[104]
port 404 nsew signal input
flabel metal2 s 500562 -960 500674 480 0 FreeSans 448 90 0 0 la_oenb[105]
port 405 nsew signal input
flabel metal2 s 504150 -960 504262 480 0 FreeSans 448 90 0 0 la_oenb[106]
port 406 nsew signal input
flabel metal2 s 507646 -960 507758 480 0 FreeSans 448 90 0 0 la_oenb[107]
port 407 nsew signal input
flabel metal2 s 511234 -960 511346 480 0 FreeSans 448 90 0 0 la_oenb[108]
port 408 nsew signal input
flabel metal2 s 514730 -960 514842 480 0 FreeSans 448 90 0 0 la_oenb[109]
port 409 nsew signal input
flabel metal2 s 163658 -960 163770 480 0 FreeSans 448 90 0 0 la_oenb[10]
port 410 nsew signal input
flabel metal2 s 518318 -960 518430 480 0 FreeSans 448 90 0 0 la_oenb[110]
port 411 nsew signal input
flabel metal2 s 521814 -960 521926 480 0 FreeSans 448 90 0 0 la_oenb[111]
port 412 nsew signal input
flabel metal2 s 525402 -960 525514 480 0 FreeSans 448 90 0 0 la_oenb[112]
port 413 nsew signal input
flabel metal2 s 528990 -960 529102 480 0 FreeSans 448 90 0 0 la_oenb[113]
port 414 nsew signal input
flabel metal2 s 532486 -960 532598 480 0 FreeSans 448 90 0 0 la_oenb[114]
port 415 nsew signal input
flabel metal2 s 536074 -960 536186 480 0 FreeSans 448 90 0 0 la_oenb[115]
port 416 nsew signal input
flabel metal2 s 539570 -960 539682 480 0 FreeSans 448 90 0 0 la_oenb[116]
port 417 nsew signal input
flabel metal2 s 543158 -960 543270 480 0 FreeSans 448 90 0 0 la_oenb[117]
port 418 nsew signal input
flabel metal2 s 546654 -960 546766 480 0 FreeSans 448 90 0 0 la_oenb[118]
port 419 nsew signal input
flabel metal2 s 550242 -960 550354 480 0 FreeSans 448 90 0 0 la_oenb[119]
port 420 nsew signal input
flabel metal2 s 167154 -960 167266 480 0 FreeSans 448 90 0 0 la_oenb[11]
port 421 nsew signal input
flabel metal2 s 553738 -960 553850 480 0 FreeSans 448 90 0 0 la_oenb[120]
port 422 nsew signal input
flabel metal2 s 557326 -960 557438 480 0 FreeSans 448 90 0 0 la_oenb[121]
port 423 nsew signal input
flabel metal2 s 560822 -960 560934 480 0 FreeSans 448 90 0 0 la_oenb[122]
port 424 nsew signal input
flabel metal2 s 564410 -960 564522 480 0 FreeSans 448 90 0 0 la_oenb[123]
port 425 nsew signal input
flabel metal2 s 567998 -960 568110 480 0 FreeSans 448 90 0 0 la_oenb[124]
port 426 nsew signal input
flabel metal2 s 571494 -960 571606 480 0 FreeSans 448 90 0 0 la_oenb[125]
port 427 nsew signal input
flabel metal2 s 575082 -960 575194 480 0 FreeSans 448 90 0 0 la_oenb[126]
port 428 nsew signal input
flabel metal2 s 578578 -960 578690 480 0 FreeSans 448 90 0 0 la_oenb[127]
port 429 nsew signal input
flabel metal2 s 170742 -960 170854 480 0 FreeSans 448 90 0 0 la_oenb[12]
port 430 nsew signal input
flabel metal2 s 174238 -960 174350 480 0 FreeSans 448 90 0 0 la_oenb[13]
port 431 nsew signal input
flabel metal2 s 177826 -960 177938 480 0 FreeSans 448 90 0 0 la_oenb[14]
port 432 nsew signal input
flabel metal2 s 181414 -960 181526 480 0 FreeSans 448 90 0 0 la_oenb[15]
port 433 nsew signal input
flabel metal2 s 184910 -960 185022 480 0 FreeSans 448 90 0 0 la_oenb[16]
port 434 nsew signal input
flabel metal2 s 188498 -960 188610 480 0 FreeSans 448 90 0 0 la_oenb[17]
port 435 nsew signal input
flabel metal2 s 191994 -960 192106 480 0 FreeSans 448 90 0 0 la_oenb[18]
port 436 nsew signal input
flabel metal2 s 195582 -960 195694 480 0 FreeSans 448 90 0 0 la_oenb[19]
port 437 nsew signal input
flabel metal2 s 131734 -960 131846 480 0 FreeSans 448 90 0 0 la_oenb[1]
port 438 nsew signal input
flabel metal2 s 199078 -960 199190 480 0 FreeSans 448 90 0 0 la_oenb[20]
port 439 nsew signal input
flabel metal2 s 202666 -960 202778 480 0 FreeSans 448 90 0 0 la_oenb[21]
port 440 nsew signal input
flabel metal2 s 206162 -960 206274 480 0 FreeSans 448 90 0 0 la_oenb[22]
port 441 nsew signal input
flabel metal2 s 209750 -960 209862 480 0 FreeSans 448 90 0 0 la_oenb[23]
port 442 nsew signal input
flabel metal2 s 213338 -960 213450 480 0 FreeSans 448 90 0 0 la_oenb[24]
port 443 nsew signal input
flabel metal2 s 216834 -960 216946 480 0 FreeSans 448 90 0 0 la_oenb[25]
port 444 nsew signal input
flabel metal2 s 220422 -960 220534 480 0 FreeSans 448 90 0 0 la_oenb[26]
port 445 nsew signal input
flabel metal2 s 223918 -960 224030 480 0 FreeSans 448 90 0 0 la_oenb[27]
port 446 nsew signal input
flabel metal2 s 227506 -960 227618 480 0 FreeSans 448 90 0 0 la_oenb[28]
port 447 nsew signal input
flabel metal2 s 231002 -960 231114 480 0 FreeSans 448 90 0 0 la_oenb[29]
port 448 nsew signal input
flabel metal2 s 135230 -960 135342 480 0 FreeSans 448 90 0 0 la_oenb[2]
port 449 nsew signal input
flabel metal2 s 234590 -960 234702 480 0 FreeSans 448 90 0 0 la_oenb[30]
port 450 nsew signal input
flabel metal2 s 238086 -960 238198 480 0 FreeSans 448 90 0 0 la_oenb[31]
port 451 nsew signal input
flabel metal2 s 241674 -960 241786 480 0 FreeSans 448 90 0 0 la_oenb[32]
port 452 nsew signal input
flabel metal2 s 245170 -960 245282 480 0 FreeSans 448 90 0 0 la_oenb[33]
port 453 nsew signal input
flabel metal2 s 248758 -960 248870 480 0 FreeSans 448 90 0 0 la_oenb[34]
port 454 nsew signal input
flabel metal2 s 252346 -960 252458 480 0 FreeSans 448 90 0 0 la_oenb[35]
port 455 nsew signal input
flabel metal2 s 255842 -960 255954 480 0 FreeSans 448 90 0 0 la_oenb[36]
port 456 nsew signal input
flabel metal2 s 259430 -960 259542 480 0 FreeSans 448 90 0 0 la_oenb[37]
port 457 nsew signal input
flabel metal2 s 262926 -960 263038 480 0 FreeSans 448 90 0 0 la_oenb[38]
port 458 nsew signal input
flabel metal2 s 266514 -960 266626 480 0 FreeSans 448 90 0 0 la_oenb[39]
port 459 nsew signal input
flabel metal2 s 138818 -960 138930 480 0 FreeSans 448 90 0 0 la_oenb[3]
port 460 nsew signal input
flabel metal2 s 270010 -960 270122 480 0 FreeSans 448 90 0 0 la_oenb[40]
port 461 nsew signal input
flabel metal2 s 273598 -960 273710 480 0 FreeSans 448 90 0 0 la_oenb[41]
port 462 nsew signal input
flabel metal2 s 277094 -960 277206 480 0 FreeSans 448 90 0 0 la_oenb[42]
port 463 nsew signal input
flabel metal2 s 280682 -960 280794 480 0 FreeSans 448 90 0 0 la_oenb[43]
port 464 nsew signal input
flabel metal2 s 284270 -960 284382 480 0 FreeSans 448 90 0 0 la_oenb[44]
port 465 nsew signal input
flabel metal2 s 287766 -960 287878 480 0 FreeSans 448 90 0 0 la_oenb[45]
port 466 nsew signal input
flabel metal2 s 291354 -960 291466 480 0 FreeSans 448 90 0 0 la_oenb[46]
port 467 nsew signal input
flabel metal2 s 294850 -960 294962 480 0 FreeSans 448 90 0 0 la_oenb[47]
port 468 nsew signal input
flabel metal2 s 298438 -960 298550 480 0 FreeSans 448 90 0 0 la_oenb[48]
port 469 nsew signal input
flabel metal2 s 301934 -960 302046 480 0 FreeSans 448 90 0 0 la_oenb[49]
port 470 nsew signal input
flabel metal2 s 142406 -960 142518 480 0 FreeSans 448 90 0 0 la_oenb[4]
port 471 nsew signal input
flabel metal2 s 305522 -960 305634 480 0 FreeSans 448 90 0 0 la_oenb[50]
port 472 nsew signal input
flabel metal2 s 309018 -960 309130 480 0 FreeSans 448 90 0 0 la_oenb[51]
port 473 nsew signal input
flabel metal2 s 312606 -960 312718 480 0 FreeSans 448 90 0 0 la_oenb[52]
port 474 nsew signal input
flabel metal2 s 316194 -960 316306 480 0 FreeSans 448 90 0 0 la_oenb[53]
port 475 nsew signal input
flabel metal2 s 319690 -960 319802 480 0 FreeSans 448 90 0 0 la_oenb[54]
port 476 nsew signal input
flabel metal2 s 323278 -960 323390 480 0 FreeSans 448 90 0 0 la_oenb[55]
port 477 nsew signal input
flabel metal2 s 326774 -960 326886 480 0 FreeSans 448 90 0 0 la_oenb[56]
port 478 nsew signal input
flabel metal2 s 330362 -960 330474 480 0 FreeSans 448 90 0 0 la_oenb[57]
port 479 nsew signal input
flabel metal2 s 333858 -960 333970 480 0 FreeSans 448 90 0 0 la_oenb[58]
port 480 nsew signal input
flabel metal2 s 337446 -960 337558 480 0 FreeSans 448 90 0 0 la_oenb[59]
port 481 nsew signal input
flabel metal2 s 145902 -960 146014 480 0 FreeSans 448 90 0 0 la_oenb[5]
port 482 nsew signal input
flabel metal2 s 340942 -960 341054 480 0 FreeSans 448 90 0 0 la_oenb[60]
port 483 nsew signal input
flabel metal2 s 344530 -960 344642 480 0 FreeSans 448 90 0 0 la_oenb[61]
port 484 nsew signal input
flabel metal2 s 348026 -960 348138 480 0 FreeSans 448 90 0 0 la_oenb[62]
port 485 nsew signal input
flabel metal2 s 351614 -960 351726 480 0 FreeSans 448 90 0 0 la_oenb[63]
port 486 nsew signal input
flabel metal2 s 355202 -960 355314 480 0 FreeSans 448 90 0 0 la_oenb[64]
port 487 nsew signal input
flabel metal2 s 358698 -960 358810 480 0 FreeSans 448 90 0 0 la_oenb[65]
port 488 nsew signal input
flabel metal2 s 362286 -960 362398 480 0 FreeSans 448 90 0 0 la_oenb[66]
port 489 nsew signal input
flabel metal2 s 365782 -960 365894 480 0 FreeSans 448 90 0 0 la_oenb[67]
port 490 nsew signal input
flabel metal2 s 369370 -960 369482 480 0 FreeSans 448 90 0 0 la_oenb[68]
port 491 nsew signal input
flabel metal2 s 372866 -960 372978 480 0 FreeSans 448 90 0 0 la_oenb[69]
port 492 nsew signal input
flabel metal2 s 149490 -960 149602 480 0 FreeSans 448 90 0 0 la_oenb[6]
port 493 nsew signal input
flabel metal2 s 376454 -960 376566 480 0 FreeSans 448 90 0 0 la_oenb[70]
port 494 nsew signal input
flabel metal2 s 379950 -960 380062 480 0 FreeSans 448 90 0 0 la_oenb[71]
port 495 nsew signal input
flabel metal2 s 383538 -960 383650 480 0 FreeSans 448 90 0 0 la_oenb[72]
port 496 nsew signal input
flabel metal2 s 387126 -960 387238 480 0 FreeSans 448 90 0 0 la_oenb[73]
port 497 nsew signal input
flabel metal2 s 390622 -960 390734 480 0 FreeSans 448 90 0 0 la_oenb[74]
port 498 nsew signal input
flabel metal2 s 394210 -960 394322 480 0 FreeSans 448 90 0 0 la_oenb[75]
port 499 nsew signal input
flabel metal2 s 397706 -960 397818 480 0 FreeSans 448 90 0 0 la_oenb[76]
port 500 nsew signal input
flabel metal2 s 401294 -960 401406 480 0 FreeSans 448 90 0 0 la_oenb[77]
port 501 nsew signal input
flabel metal2 s 404790 -960 404902 480 0 FreeSans 448 90 0 0 la_oenb[78]
port 502 nsew signal input
flabel metal2 s 408378 -960 408490 480 0 FreeSans 448 90 0 0 la_oenb[79]
port 503 nsew signal input
flabel metal2 s 152986 -960 153098 480 0 FreeSans 448 90 0 0 la_oenb[7]
port 504 nsew signal input
flabel metal2 s 411874 -960 411986 480 0 FreeSans 448 90 0 0 la_oenb[80]
port 505 nsew signal input
flabel metal2 s 415462 -960 415574 480 0 FreeSans 448 90 0 0 la_oenb[81]
port 506 nsew signal input
flabel metal2 s 418958 -960 419070 480 0 FreeSans 448 90 0 0 la_oenb[82]
port 507 nsew signal input
flabel metal2 s 422546 -960 422658 480 0 FreeSans 448 90 0 0 la_oenb[83]
port 508 nsew signal input
flabel metal2 s 426134 -960 426246 480 0 FreeSans 448 90 0 0 la_oenb[84]
port 509 nsew signal input
flabel metal2 s 429630 -960 429742 480 0 FreeSans 448 90 0 0 la_oenb[85]
port 510 nsew signal input
flabel metal2 s 433218 -960 433330 480 0 FreeSans 448 90 0 0 la_oenb[86]
port 511 nsew signal input
flabel metal2 s 436714 -960 436826 480 0 FreeSans 448 90 0 0 la_oenb[87]
port 512 nsew signal input
flabel metal2 s 440302 -960 440414 480 0 FreeSans 448 90 0 0 la_oenb[88]
port 513 nsew signal input
flabel metal2 s 443798 -960 443910 480 0 FreeSans 448 90 0 0 la_oenb[89]
port 514 nsew signal input
flabel metal2 s 156574 -960 156686 480 0 FreeSans 448 90 0 0 la_oenb[8]
port 515 nsew signal input
flabel metal2 s 447386 -960 447498 480 0 FreeSans 448 90 0 0 la_oenb[90]
port 516 nsew signal input
flabel metal2 s 450882 -960 450994 480 0 FreeSans 448 90 0 0 la_oenb[91]
port 517 nsew signal input
flabel metal2 s 454470 -960 454582 480 0 FreeSans 448 90 0 0 la_oenb[92]
port 518 nsew signal input
flabel metal2 s 458058 -960 458170 480 0 FreeSans 448 90 0 0 la_oenb[93]
port 519 nsew signal input
flabel metal2 s 461554 -960 461666 480 0 FreeSans 448 90 0 0 la_oenb[94]
port 520 nsew signal input
flabel metal2 s 465142 -960 465254 480 0 FreeSans 448 90 0 0 la_oenb[95]
port 521 nsew signal input
flabel metal2 s 468638 -960 468750 480 0 FreeSans 448 90 0 0 la_oenb[96]
port 522 nsew signal input
flabel metal2 s 472226 -960 472338 480 0 FreeSans 448 90 0 0 la_oenb[97]
port 523 nsew signal input
flabel metal2 s 475722 -960 475834 480 0 FreeSans 448 90 0 0 la_oenb[98]
port 524 nsew signal input
flabel metal2 s 479310 -960 479422 480 0 FreeSans 448 90 0 0 la_oenb[99]
port 525 nsew signal input
flabel metal2 s 160070 -960 160182 480 0 FreeSans 448 90 0 0 la_oenb[9]
port 526 nsew signal input
flabel metal2 s 579774 -960 579886 480 0 FreeSans 448 90 0 0 user_clock2
port 527 nsew signal input
flabel metal2 s 580970 -960 581082 480 0 FreeSans 448 90 0 0 user_irq[0]
port 528 nsew signal tristate
flabel metal2 s 582166 -960 582278 480 0 FreeSans 448 90 0 0 user_irq[1]
port 529 nsew signal tristate
flabel metal2 s 583362 -960 583474 480 0 FreeSans 448 90 0 0 user_irq[2]
port 530 nsew signal tristate
flabel metal4 s -2006 -934 -1386 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 -934 585930 -314 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 704250 585930 704870 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 585310 -934 585930 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 1794 -7654 2414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 37794 -7654 38414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 -7654 74414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 -7654 110414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 -7654 146414 78000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 142000 146414 198000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 262000 146414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 -7654 182414 78000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 142000 182414 198000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 262000 182414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 -7654 218414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 -7654 254414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 -7654 290414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 -7654 326414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 -7654 362414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 -7654 398414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 -7654 434414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 -7654 470414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 -7654 506414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 541794 -7654 542414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 577794 -7654 578414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 2866 592650 3486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 38866 592650 39486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 74866 592650 75486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 110866 592650 111486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 146866 592650 147486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 182866 592650 183486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 218866 592650 219486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 254866 592650 255486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 290866 592650 291486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 326866 592650 327486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 362866 592650 363486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 398866 592650 399486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 434866 592650 435486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 470866 592650 471486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 506866 592650 507486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 542866 592650 543486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 578866 592650 579486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 614866 592650 615486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 650866 592650 651486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 686866 592650 687486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s -3926 -2854 -3306 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 -2854 587850 -2234 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 706170 587850 706790 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 587230 -2854 587850 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 10794 -7654 11414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 46794 -7654 47414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 82794 -7654 83414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 -7654 119414 78000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 142000 119414 198000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 262000 119414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 154794 -7654 155414 78000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 154794 142000 155414 198000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 154794 262000 155414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 190794 -7654 191414 78000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 190794 142000 191414 198000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 190794 262000 191414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 226794 -7654 227414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 262794 -7654 263414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 298794 -7654 299414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 334794 -7654 335414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 370794 -7654 371414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 406794 -7654 407414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 442794 -7654 443414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 478794 -7654 479414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 514794 -7654 515414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 550794 -7654 551414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 11866 592650 12486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 47866 592650 48486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 83866 592650 84486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 119866 592650 120486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 155866 592650 156486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 191866 592650 192486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 227866 592650 228486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 263866 592650 264486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 299866 592650 300486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 335866 592650 336486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 371866 592650 372486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 407866 592650 408486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 443866 592650 444486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 479866 592650 480486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 515866 592650 516486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 551866 592650 552486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 587866 592650 588486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 623866 592650 624486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 659866 592650 660486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 695866 592650 696486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s -5846 -4774 -5226 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 -4774 589770 -4154 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 708090 589770 708710 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 589150 -4774 589770 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 19794 -7654 20414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 55794 -7654 56414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 91794 -7654 92414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 127794 -7654 128414 78000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 127794 262000 128414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 163794 -7654 164414 78000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 163794 262000 164414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 199794 -7654 200414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 235794 -7654 236414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 271794 -7654 272414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 307794 -7654 308414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 343794 -7654 344414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 379794 -7654 380414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 415794 -7654 416414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 451794 -7654 452414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 487794 -7654 488414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 523794 -7654 524414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 559794 -7654 560414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 20866 592650 21486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 56866 592650 57486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 92866 592650 93486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 128866 592650 129486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 164866 592650 165486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 200866 592650 201486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 236866 592650 237486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 272866 592650 273486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 308866 592650 309486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 344866 592650 345486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 380866 592650 381486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 416866 592650 417486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 452866 592650 453486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 488866 592650 489486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 524866 592650 525486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 560866 592650 561486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 596866 592650 597486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 632866 592650 633486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 668866 592650 669486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s -7766 -6694 -7146 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 -6694 591690 -6074 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 710010 591690 710630 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 591070 -6694 591690 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 28794 -7654 29414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 64794 -7654 65414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 100794 -7654 101414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 136794 -7654 137414 78000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 136794 262000 137414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 172794 -7654 173414 78000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 172794 262000 173414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 208794 -7654 209414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 244794 -7654 245414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 280794 -7654 281414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 316794 -7654 317414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 352794 -7654 353414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 388794 -7654 389414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 424794 -7654 425414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 460794 -7654 461414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 496794 -7654 497414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 532794 -7654 533414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 568794 -7654 569414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 29866 592650 30486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 65866 592650 66486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 101866 592650 102486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 137866 592650 138486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 173866 592650 174486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 209866 592650 210486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 245866 592650 246486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 281866 592650 282486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 317866 592650 318486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 353866 592650 354486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 389866 592650 390486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 425866 592650 426486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 461866 592650 462486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 497866 592650 498486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 533866 592650 534486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 569866 592650 570486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 605866 592650 606486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 641866 592650 642486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 677866 592650 678486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s -6806 -5734 -6186 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 -5734 590730 -5114 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 709050 590730 709670 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 590110 -5734 590730 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 24294 -7654 24914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 60294 -7654 60914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 96294 -7654 96914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 132294 -7654 132914 78000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 132294 262000 132914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 168294 -7654 168914 78000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 168294 262000 168914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 204294 -7654 204914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 240294 -7654 240914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 276294 -7654 276914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 312294 -7654 312914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 348294 -7654 348914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 384294 -7654 384914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 420294 -7654 420914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 456294 -7654 456914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 492294 -7654 492914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 528294 -7654 528914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 564294 -7654 564914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 25366 592650 25986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 61366 592650 61986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 97366 592650 97986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 133366 592650 133986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 169366 592650 169986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 205366 592650 205986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 241366 592650 241986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 277366 592650 277986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 313366 592650 313986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 349366 592650 349986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 385366 592650 385986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 421366 592650 421986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 457366 592650 457986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 493366 592650 493986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 529366 592650 529986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 565366 592650 565986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 601366 592650 601986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 637366 592650 637986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 673366 592650 673986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s -8726 -7654 -8106 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 -7654 592650 -7034 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 710970 592650 711590 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 592030 -7654 592650 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 33294 -7654 33914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 69294 -7654 69914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 105294 -7654 105914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 141294 -7654 141914 78000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 141294 142000 141914 198000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 141294 262000 141914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 177294 -7654 177914 78000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 177294 142000 177914 198000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 177294 262000 177914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 213294 -7654 213914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 249294 -7654 249914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 285294 -7654 285914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 321294 -7654 321914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 357294 -7654 357914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 393294 -7654 393914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 429294 -7654 429914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 465294 -7654 465914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 501294 -7654 501914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 537294 -7654 537914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 573294 -7654 573914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 34366 592650 34986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 70366 592650 70986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 106366 592650 106986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 142366 592650 142986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 178366 592650 178986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 214366 592650 214986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 250366 592650 250986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 286366 592650 286986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 322366 592650 322986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 358366 592650 358986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 394366 592650 394986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 430366 592650 430986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 466366 592650 466986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 502366 592650 502986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 538366 592650 538986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 574366 592650 574986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 610366 592650 610986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 646366 592650 646986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 682366 592650 682986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s -2966 -1894 -2346 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 -1894 586890 -1274 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 705210 586890 705830 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 586270 -1894 586890 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 6294 -7654 6914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 42294 -7654 42914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 78294 -7654 78914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 114294 -7654 114914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 150294 -7654 150914 78000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 150294 142000 150914 198000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 150294 262000 150914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 186294 -7654 186914 78000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 186294 142000 186914 198000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 186294 262000 186914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 222294 -7654 222914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 258294 -7654 258914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 294294 -7654 294914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 330294 -7654 330914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 366294 -7654 366914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 402294 -7654 402914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 438294 -7654 438914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 474294 -7654 474914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 510294 -7654 510914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 546294 -7654 546914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 582294 -7654 582914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 7366 592650 7986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 43366 592650 43986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 79366 592650 79986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 115366 592650 115986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 151366 592650 151986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 187366 592650 187986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 223366 592650 223986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 259366 592650 259986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 295366 592650 295986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 331366 592650 331986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 367366 592650 367986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 403366 592650 403986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 439366 592650 439986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 475366 592650 475986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 511366 592650 511986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 547366 592650 547986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 583366 592650 583986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 619366 592650 619986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 655366 592650 655986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 691366 592650 691986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s -4886 -3814 -4266 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 -3814 588810 -3194 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 707130 588810 707750 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 588190 -3814 588810 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 15294 -7654 15914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 51294 -7654 51914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 87294 -7654 87914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 -7654 123914 78000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 142000 123914 198000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 262000 123914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 159294 -7654 159914 78000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 159294 142000 159914 198000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 159294 262000 159914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 195294 -7654 195914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 231294 -7654 231914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 267294 -7654 267914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 303294 -7654 303914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 339294 -7654 339914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 375294 -7654 375914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 411294 -7654 411914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 447294 -7654 447914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 483294 -7654 483914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 519294 -7654 519914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 555294 -7654 555914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 16366 592650 16986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 52366 592650 52986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 88366 592650 88986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 124366 592650 124986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 160366 592650 160986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 196366 592650 196986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 232366 592650 232986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 268366 592650 268986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 304366 592650 304986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 340366 592650 340986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 376366 592650 376986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 412366 592650 412986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 448366 592650 448986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 484366 592650 484986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 520366 592650 520986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 556366 592650 556986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 592366 592650 592986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 628366 592650 628986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 664366 592650 664986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 700366 592650 700986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal2 s 542 -960 654 480 0 FreeSans 448 90 0 0 wb_clk_i
port 539 nsew signal input
flabel metal2 s 1646 -960 1758 480 0 FreeSans 448 90 0 0 wb_rst_i
port 540 nsew signal input
flabel metal2 s 2842 -960 2954 480 0 FreeSans 448 90 0 0 wbs_ack_o
port 541 nsew signal tristate
flabel metal2 s 7626 -960 7738 480 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 542 nsew signal input
flabel metal2 s 47830 -960 47942 480 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 543 nsew signal input
flabel metal2 s 51326 -960 51438 480 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 544 nsew signal input
flabel metal2 s 54914 -960 55026 480 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 545 nsew signal input
flabel metal2 s 58410 -960 58522 480 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 546 nsew signal input
flabel metal2 s 61998 -960 62110 480 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 547 nsew signal input
flabel metal2 s 65494 -960 65606 480 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 548 nsew signal input
flabel metal2 s 69082 -960 69194 480 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 549 nsew signal input
flabel metal2 s 72578 -960 72690 480 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 550 nsew signal input
flabel metal2 s 76166 -960 76278 480 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 551 nsew signal input
flabel metal2 s 79662 -960 79774 480 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 552 nsew signal input
flabel metal2 s 12318 -960 12430 480 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 553 nsew signal input
flabel metal2 s 83250 -960 83362 480 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 554 nsew signal input
flabel metal2 s 86838 -960 86950 480 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 555 nsew signal input
flabel metal2 s 90334 -960 90446 480 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 556 nsew signal input
flabel metal2 s 93922 -960 94034 480 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 557 nsew signal input
flabel metal2 s 97418 -960 97530 480 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 558 nsew signal input
flabel metal2 s 101006 -960 101118 480 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 559 nsew signal input
flabel metal2 s 104502 -960 104614 480 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 560 nsew signal input
flabel metal2 s 108090 -960 108202 480 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 561 nsew signal input
flabel metal2 s 111586 -960 111698 480 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 562 nsew signal input
flabel metal2 s 115174 -960 115286 480 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 563 nsew signal input
flabel metal2 s 17010 -960 17122 480 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 564 nsew signal input
flabel metal2 s 118762 -960 118874 480 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 565 nsew signal input
flabel metal2 s 122258 -960 122370 480 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 566 nsew signal input
flabel metal2 s 21794 -960 21906 480 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 567 nsew signal input
flabel metal2 s 26486 -960 26598 480 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 568 nsew signal input
flabel metal2 s 30074 -960 30186 480 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 569 nsew signal input
flabel metal2 s 33570 -960 33682 480 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 570 nsew signal input
flabel metal2 s 37158 -960 37270 480 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 571 nsew signal input
flabel metal2 s 40654 -960 40766 480 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 572 nsew signal input
flabel metal2 s 44242 -960 44354 480 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 573 nsew signal input
flabel metal2 s 4038 -960 4150 480 0 FreeSans 448 90 0 0 wbs_cyc_i
port 574 nsew signal input
flabel metal2 s 8730 -960 8842 480 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 575 nsew signal input
flabel metal2 s 48934 -960 49046 480 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 576 nsew signal input
flabel metal2 s 52522 -960 52634 480 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 577 nsew signal input
flabel metal2 s 56018 -960 56130 480 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 578 nsew signal input
flabel metal2 s 59606 -960 59718 480 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 579 nsew signal input
flabel metal2 s 63194 -960 63306 480 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 580 nsew signal input
flabel metal2 s 66690 -960 66802 480 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 581 nsew signal input
flabel metal2 s 70278 -960 70390 480 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 582 nsew signal input
flabel metal2 s 73774 -960 73886 480 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 583 nsew signal input
flabel metal2 s 77362 -960 77474 480 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 584 nsew signal input
flabel metal2 s 80858 -960 80970 480 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 585 nsew signal input
flabel metal2 s 13514 -960 13626 480 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 586 nsew signal input
flabel metal2 s 84446 -960 84558 480 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 587 nsew signal input
flabel metal2 s 87942 -960 88054 480 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 588 nsew signal input
flabel metal2 s 91530 -960 91642 480 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 589 nsew signal input
flabel metal2 s 95118 -960 95230 480 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 590 nsew signal input
flabel metal2 s 98614 -960 98726 480 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 591 nsew signal input
flabel metal2 s 102202 -960 102314 480 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 592 nsew signal input
flabel metal2 s 105698 -960 105810 480 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 593 nsew signal input
flabel metal2 s 109286 -960 109398 480 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 594 nsew signal input
flabel metal2 s 112782 -960 112894 480 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 595 nsew signal input
flabel metal2 s 116370 -960 116482 480 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 596 nsew signal input
flabel metal2 s 18206 -960 18318 480 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 597 nsew signal input
flabel metal2 s 119866 -960 119978 480 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 598 nsew signal input
flabel metal2 s 123454 -960 123566 480 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 599 nsew signal input
flabel metal2 s 22990 -960 23102 480 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 600 nsew signal input
flabel metal2 s 27682 -960 27794 480 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 601 nsew signal input
flabel metal2 s 31270 -960 31382 480 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 602 nsew signal input
flabel metal2 s 34766 -960 34878 480 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 603 nsew signal input
flabel metal2 s 38354 -960 38466 480 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 604 nsew signal input
flabel metal2 s 41850 -960 41962 480 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 605 nsew signal input
flabel metal2 s 45438 -960 45550 480 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 606 nsew signal input
flabel metal2 s 9926 -960 10038 480 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 607 nsew signal tristate
flabel metal2 s 50130 -960 50242 480 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 608 nsew signal tristate
flabel metal2 s 53718 -960 53830 480 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 609 nsew signal tristate
flabel metal2 s 57214 -960 57326 480 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 610 nsew signal tristate
flabel metal2 s 60802 -960 60914 480 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 611 nsew signal tristate
flabel metal2 s 64298 -960 64410 480 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 612 nsew signal tristate
flabel metal2 s 67886 -960 67998 480 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 613 nsew signal tristate
flabel metal2 s 71474 -960 71586 480 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 614 nsew signal tristate
flabel metal2 s 74970 -960 75082 480 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 615 nsew signal tristate
flabel metal2 s 78558 -960 78670 480 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 616 nsew signal tristate
flabel metal2 s 82054 -960 82166 480 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 617 nsew signal tristate
flabel metal2 s 14710 -960 14822 480 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 618 nsew signal tristate
flabel metal2 s 85642 -960 85754 480 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 619 nsew signal tristate
flabel metal2 s 89138 -960 89250 480 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 620 nsew signal tristate
flabel metal2 s 92726 -960 92838 480 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 621 nsew signal tristate
flabel metal2 s 96222 -960 96334 480 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 622 nsew signal tristate
flabel metal2 s 99810 -960 99922 480 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 623 nsew signal tristate
flabel metal2 s 103306 -960 103418 480 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 624 nsew signal tristate
flabel metal2 s 106894 -960 107006 480 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 625 nsew signal tristate
flabel metal2 s 110482 -960 110594 480 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 626 nsew signal tristate
flabel metal2 s 113978 -960 114090 480 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 627 nsew signal tristate
flabel metal2 s 117566 -960 117678 480 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 628 nsew signal tristate
flabel metal2 s 19402 -960 19514 480 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 629 nsew signal tristate
flabel metal2 s 121062 -960 121174 480 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 630 nsew signal tristate
flabel metal2 s 124650 -960 124762 480 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 631 nsew signal tristate
flabel metal2 s 24186 -960 24298 480 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 632 nsew signal tristate
flabel metal2 s 28878 -960 28990 480 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 633 nsew signal tristate
flabel metal2 s 32374 -960 32486 480 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 634 nsew signal tristate
flabel metal2 s 35962 -960 36074 480 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 635 nsew signal tristate
flabel metal2 s 39550 -960 39662 480 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 636 nsew signal tristate
flabel metal2 s 43046 -960 43158 480 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 637 nsew signal tristate
flabel metal2 s 46634 -960 46746 480 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 638 nsew signal tristate
flabel metal2 s 11122 -960 11234 480 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 639 nsew signal input
flabel metal2 s 15906 -960 16018 480 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 640 nsew signal input
flabel metal2 s 20598 -960 20710 480 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 641 nsew signal input
flabel metal2 s 25290 -960 25402 480 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 642 nsew signal input
flabel metal2 s 5234 -960 5346 480 0 FreeSans 448 90 0 0 wbs_stb_i
port 643 nsew signal input
flabel metal2 s 6430 -960 6542 480 0 FreeSans 448 90 0 0 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
