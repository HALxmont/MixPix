VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO APS
  CLASS BLOCK ;
  FOREIGN APS ;
  ORIGIN -150.000 13.000 ;
  SIZE 126.500 BY 84.000 ;
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 246.500 67.000 270.500 71.000 ;
        RECT 246.500 63.000 270.470 67.000 ;
    END
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 150.000 33.500 251.500 35.000 ;
        RECT 150.000 1.500 151.500 33.500 ;
        RECT 250.000 1.500 251.500 33.500 ;
        RECT 150.000 0.000 251.500 1.500 ;
        RECT 212.000 -3.500 214.960 0.000 ;
        RECT 215.000 -3.500 217.960 0.000 ;
        RECT 218.000 -2.600 220.960 0.000 ;
        RECT 221.000 -2.600 235.570 0.000 ;
        RECT 218.000 -2.900 235.570 -2.600 ;
        RECT 218.000 -3.500 220.960 -2.900 ;
        RECT 221.000 -3.500 235.570 -2.900 ;
      LAYER li1 ;
        RECT 258.500 38.000 262.500 47.500 ;
        RECT 150.500 34.000 266.000 38.000 ;
        RECT 150.500 1.000 151.000 34.000 ;
        RECT 250.500 1.000 251.000 34.000 ;
        RECT 150.500 0.500 251.000 1.000 ;
        RECT 212.500 0.110 235.500 0.500 ;
        RECT 212.180 0.000 235.500 0.110 ;
        RECT 212.180 -0.060 214.780 0.000 ;
        RECT 212.180 -3.150 212.350 -0.060 ;
        RECT 214.040 -2.470 214.210 -0.430 ;
        RECT 214.610 -3.150 214.780 -0.060 ;
        RECT 212.180 -3.320 214.780 -3.150 ;
        RECT 215.180 -0.060 217.780 0.000 ;
        RECT 215.180 -3.150 215.350 -0.060 ;
        RECT 215.750 -2.470 215.920 -0.430 ;
        RECT 217.610 -3.150 217.780 -0.060 ;
        RECT 215.180 -3.320 217.780 -3.150 ;
        RECT 218.180 -0.060 220.780 0.000 ;
        RECT 218.180 -3.150 218.350 -0.060 ;
        RECT 220.100 -0.430 220.780 -0.060 ;
        RECT 220.040 -2.300 220.780 -0.430 ;
        RECT 220.040 -2.470 220.210 -2.300 ;
        RECT 220.610 -3.150 220.780 -2.300 ;
        RECT 218.180 -3.320 220.780 -3.150 ;
        RECT 221.180 -0.060 235.390 0.000 ;
        RECT 221.180 -3.150 221.350 -0.060 ;
        RECT 221.700 -0.900 222.000 -0.060 ;
        RECT 224.300 -0.900 224.600 -0.060 ;
        RECT 226.800 -0.900 227.100 -0.060 ;
        RECT 229.400 -0.900 229.700 -0.060 ;
        RECT 232.000 -0.900 232.300 -0.060 ;
        RECT 234.600 -0.900 234.900 -0.060 ;
        RECT 221.750 -2.470 221.920 -0.900 ;
        RECT 224.330 -2.470 224.500 -0.900 ;
        RECT 226.910 -2.470 227.080 -0.900 ;
        RECT 229.490 -2.470 229.660 -0.900 ;
        RECT 232.070 -2.470 232.240 -0.900 ;
        RECT 234.650 -2.470 234.820 -0.900 ;
        RECT 235.220 -3.150 235.390 -0.060 ;
        RECT 221.180 -3.320 235.390 -3.150 ;
      LAYER mcon ;
        RECT 258.500 43.500 262.500 47.500 ;
        RECT 214.040 -2.390 214.210 -0.510 ;
        RECT 215.750 -2.390 215.920 -0.510 ;
        RECT 220.040 -2.390 220.210 -0.510 ;
        RECT 221.750 -2.390 221.920 -0.510 ;
        RECT 224.330 -2.390 224.500 -0.510 ;
        RECT 226.910 -2.390 227.080 -0.510 ;
        RECT 229.490 -2.390 229.660 -0.510 ;
        RECT 232.070 -2.390 232.240 -0.510 ;
        RECT 234.650 -2.390 234.820 -0.510 ;
      LAYER met1 ;
        RECT 258.470 47.530 262.530 47.560 ;
        RECT 258.440 43.470 262.560 47.530 ;
        RECT 250.250 0.750 250.750 43.030 ;
        RECT 214.000 0.250 250.750 0.750 ;
        RECT 214.000 -1.750 214.500 0.250 ;
        RECT 214.010 -2.450 214.240 -1.750 ;
        RECT 215.500 -2.250 216.000 0.250 ;
        RECT 215.720 -2.450 215.950 -2.250 ;
        RECT 220.010 -2.450 220.240 -0.450 ;
        RECT 221.720 -2.450 221.950 -0.450 ;
        RECT 224.300 -2.450 224.530 -0.450 ;
        RECT 226.880 -2.450 227.110 -0.450 ;
        RECT 229.460 -2.450 229.690 -0.450 ;
        RECT 232.040 -2.450 232.270 -0.450 ;
        RECT 234.620 -2.450 234.850 -0.450 ;
      LAYER via ;
        RECT 258.470 43.530 262.530 47.530 ;
        RECT 250.250 42.500 250.750 43.000 ;
      LAYER met2 ;
        RECT 250.250 43.000 250.750 43.045 ;
        RECT 258.000 43.000 263.000 48.000 ;
        RECT 250.220 42.500 250.780 43.000 ;
        RECT 250.250 42.455 250.750 42.500 ;
      LAYER via2 ;
        RECT 258.470 43.530 262.530 47.530 ;
        RECT 250.250 42.500 250.750 43.000 ;
      LAYER met3 ;
        RECT 250.225 42.475 250.775 43.055 ;
        RECT 258.000 43.000 263.000 48.000 ;
      LAYER via3 ;
        RECT 258.445 43.505 262.555 47.555 ;
        RECT 250.225 42.525 250.775 43.025 ;
      LAYER met4 ;
        RECT 258.440 47.530 262.560 47.560 ;
        RECT 258.440 47.500 275.500 47.530 ;
        RECT 246.500 43.500 276.500 47.500 ;
        RECT 250.250 43.030 250.750 43.500 ;
        RECT 250.220 42.520 250.780 43.030 ;
    END
  END VSS
  PIN RST
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.000000 ;
    PORT
      LAYER li1 ;
        RECT 212.980 -2.810 213.980 -2.640 ;
      LAYER mcon ;
        RECT 213.060 -2.810 213.900 -2.640 ;
      LAYER met1 ;
        RECT 213.250 -2.610 213.750 -2.500 ;
        RECT 213.000 -2.840 213.960 -2.610 ;
        RECT 213.250 -4.000 213.750 -2.840 ;
        RECT 205.000 -4.500 213.750 -4.000 ;
        RECT 205.000 -5.200 205.500 -4.500 ;
        RECT 204.950 -5.800 205.550 -5.200 ;
      LAYER via ;
        RECT 205.000 -5.750 205.500 -5.250 ;
      LAYER met2 ;
        RECT 204.800 -6.000 205.800 -5.150 ;
        RECT 203.000 -13.000 207.500 -6.000 ;
    END
  END RST
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.160000 ;
    PORT
      LAYER li1 ;
        RECT 217.040 -2.470 217.210 -0.430 ;
        RECT 218.750 -2.470 218.920 -0.430 ;
      LAYER mcon ;
        RECT 217.040 -2.390 217.210 -0.510 ;
        RECT 218.750 -2.390 218.920 -0.510 ;
      LAYER met1 ;
        RECT 217.010 -1.000 217.240 -0.450 ;
        RECT 218.720 -1.000 218.950 -0.450 ;
        RECT 217.000 -2.000 218.950 -1.000 ;
        RECT 217.010 -2.450 217.240 -2.000 ;
        RECT 217.700 -5.430 218.300 -2.000 ;
        RECT 218.720 -2.450 218.950 -2.000 ;
      LAYER via ;
        RECT 217.700 -5.400 218.300 -4.800 ;
      LAYER met2 ;
        RECT 217.670 -5.400 218.330 -4.800 ;
        RECT 217.700 -6.000 218.300 -5.400 ;
        RECT 216.000 -13.000 220.500 -6.000 ;
    END
  END OUT
  PIN IP
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.000000 ;
    ANTENNADIFFAREA 2.900000 ;
    PORT
      LAYER li1 ;
        RECT 223.040 -2.470 223.210 -0.430 ;
        RECT 225.620 -2.470 225.790 -0.430 ;
        RECT 228.200 -2.470 228.370 -0.430 ;
        RECT 230.780 -2.470 230.950 -0.430 ;
        RECT 233.360 -2.470 233.530 -0.430 ;
        RECT 218.980 -2.810 219.980 -2.640 ;
      LAYER mcon ;
        RECT 223.040 -2.390 223.210 -0.510 ;
        RECT 225.620 -2.390 225.790 -0.510 ;
        RECT 228.200 -2.390 228.370 -0.510 ;
        RECT 230.780 -2.390 230.950 -0.510 ;
        RECT 233.360 -2.390 233.530 -0.510 ;
        RECT 219.060 -2.810 219.900 -2.640 ;
      LAYER met1 ;
        RECT 223.010 -2.200 223.240 -0.450 ;
        RECT 225.590 -2.200 225.820 -0.450 ;
        RECT 228.170 -2.200 228.400 -0.450 ;
        RECT 230.750 -2.200 230.980 -0.450 ;
        RECT 233.330 -2.200 233.560 -0.450 ;
        RECT 223.000 -2.600 223.300 -2.200 ;
        RECT 225.590 -2.450 225.900 -2.200 ;
        RECT 225.600 -2.600 225.900 -2.450 ;
        RECT 228.100 -2.600 228.400 -2.200 ;
        RECT 230.700 -2.600 231.000 -2.200 ;
        RECT 233.300 -2.600 233.600 -2.200 ;
        RECT 218.900 -2.900 234.800 -2.600 ;
        RECT 227.200 -5.530 227.800 -2.900 ;
      LAYER via ;
        RECT 227.200 -5.500 227.800 -4.900 ;
      LAYER met2 ;
        RECT 227.170 -5.500 227.830 -4.900 ;
        RECT 227.200 -6.000 227.800 -5.500 ;
        RECT 226.000 -13.000 230.500 -6.000 ;
    END
  END IP
  OBS
      LAYER nwell ;
        RECT 151.500 30.500 250.000 33.500 ;
        RECT 151.500 4.500 154.500 30.500 ;
        RECT 185.500 25.000 215.500 27.500 ;
        RECT 185.500 10.000 188.000 25.000 ;
        RECT 199.300 17.300 200.700 18.700 ;
        RECT 213.000 10.000 215.500 25.000 ;
        RECT 185.500 7.500 215.500 10.000 ;
        RECT 247.000 4.500 250.000 30.500 ;
        RECT 151.500 1.500 250.000 4.500 ;
      LAYER li1 ;
        RECT 152.500 2.500 153.500 32.500 ;
        RECT 196.500 31.500 203.500 32.500 ;
        RECT 186.500 14.500 187.500 21.500 ;
        RECT 199.500 17.500 200.500 18.500 ;
        RECT 199.750 6.150 200.250 17.500 ;
        RECT 213.500 14.500 214.500 21.500 ;
        RECT 199.750 5.650 205.400 6.150 ;
        RECT 196.500 2.500 203.500 3.500 ;
        RECT 204.900 1.500 205.400 5.650 ;
        RECT 248.000 2.500 249.000 32.500 ;
        RECT 212.750 -2.470 212.920 -0.430 ;
        RECT 215.980 -2.810 216.980 -2.640 ;
        RECT 221.980 -2.810 222.980 -2.640 ;
        RECT 223.270 -2.810 224.270 -2.640 ;
        RECT 224.560 -2.810 225.560 -2.640 ;
        RECT 225.850 -2.810 226.850 -2.640 ;
        RECT 227.140 -2.810 228.140 -2.640 ;
        RECT 228.430 -2.810 229.430 -2.640 ;
        RECT 229.720 -2.810 230.720 -2.640 ;
        RECT 231.010 -2.810 232.010 -2.640 ;
        RECT 232.300 -2.810 233.300 -2.640 ;
        RECT 233.590 -2.810 234.590 -2.640 ;
      LAYER mcon ;
        RECT 212.750 -2.390 212.920 -0.510 ;
        RECT 216.060 -2.810 216.900 -2.640 ;
      LAYER met1 ;
        RECT 154.500 4.500 247.000 30.500 ;
      LAYER met1 ;
        RECT 204.840 1.470 205.460 2.030 ;
        RECT 204.900 -0.750 205.400 1.470 ;
        RECT 212.720 -0.750 212.950 -0.450 ;
        RECT 204.900 -1.250 213.000 -0.750 ;
        RECT 210.500 -2.780 211.000 -1.250 ;
        RECT 212.720 -2.450 212.950 -1.250 ;
        RECT 216.250 -2.610 216.750 -2.500 ;
        RECT 216.000 -2.840 216.960 -2.610 ;
        RECT 215.250 -4.000 215.750 -3.970 ;
        RECT 216.250 -4.000 216.750 -2.840 ;
        RECT 215.250 -4.500 216.750 -4.000 ;
        RECT 215.250 -4.530 215.750 -4.500 ;
      LAYER via ;
        RECT 210.500 -2.750 211.000 -2.250 ;
      LAYER met2 ;
        RECT 150.500 0.500 250.500 34.500 ;
      LAYER met2 ;
        RECT 210.470 -2.750 211.030 -2.250 ;
        RECT 210.500 -4.000 211.000 -2.750 ;
        RECT 210.500 -4.500 215.780 -4.000 ;
  END
END APS
END LIBRARY

