magic
tech sky130B
magscale 1 2
timestamp 1668033436
<< viali >>
rect 22109 57545 22143 57579
rect 30849 57545 30883 57579
rect 40049 57545 40083 57579
rect 48329 57545 48363 57579
rect 57069 57545 57103 57579
rect 65809 57545 65843 57579
rect 47593 57477 47627 57511
rect 4445 57409 4479 57443
rect 13185 57409 13219 57443
rect 21925 57409 21959 57443
rect 30665 57409 30699 57443
rect 39865 57409 39899 57443
rect 48145 57409 48179 57443
rect 56885 57409 56919 57443
rect 65073 57409 65107 57443
rect 65625 57409 65659 57443
rect 67649 57409 67683 57443
rect 30113 57205 30147 57239
rect 39221 57205 39255 57239
rect 56333 57205 56367 57239
rect 21741 56661 21775 56695
rect 67649 56117 67683 56151
rect 68109 54621 68143 54655
rect 68109 53533 68143 53567
rect 67649 51765 67683 51799
rect 68109 50269 68143 50303
rect 67649 48569 67683 48603
rect 67649 47413 67683 47447
rect 68109 45917 68143 45951
rect 67649 44149 67683 44183
rect 68109 42653 68143 42687
rect 68109 41565 68143 41599
rect 67649 39797 67683 39831
rect 68109 38301 68143 38335
rect 67649 36601 67683 36635
rect 67649 35445 67683 35479
rect 68109 33949 68143 33983
rect 67649 32181 67683 32215
rect 68109 30685 68143 30719
rect 7205 30209 7239 30243
rect 8033 30209 8067 30243
rect 6929 30141 6963 30175
rect 27169 29801 27203 29835
rect 7303 29597 7337 29631
rect 7481 29597 7515 29631
rect 26157 29597 26191 29631
rect 26433 29597 26467 29631
rect 68109 29597 68143 29631
rect 7389 29461 7423 29495
rect 5089 29121 5123 29155
rect 6745 29121 6779 29155
rect 7849 29121 7883 29155
rect 19349 29121 19383 29155
rect 24501 29121 24535 29155
rect 4813 29053 4847 29087
rect 6561 29053 6595 29087
rect 19441 29053 19475 29087
rect 5825 28985 5859 29019
rect 7757 28985 7791 29019
rect 8309 28985 8343 29019
rect 18981 28985 19015 29019
rect 6929 28917 6963 28951
rect 9229 28917 9263 28951
rect 24409 28917 24443 28951
rect 6745 28713 6779 28747
rect 8309 28713 8343 28747
rect 16957 28713 16991 28747
rect 17785 28713 17819 28747
rect 18245 28713 18279 28747
rect 19717 28713 19751 28747
rect 23857 28713 23891 28747
rect 6101 28645 6135 28679
rect 4813 28577 4847 28611
rect 9321 28577 9355 28611
rect 16773 28577 16807 28611
rect 17969 28577 18003 28611
rect 21741 28577 21775 28611
rect 25789 28577 25823 28611
rect 4537 28509 4571 28543
rect 5457 28509 5491 28543
rect 5641 28509 5675 28543
rect 6285 28509 6319 28543
rect 6929 28509 6963 28543
rect 7941 28509 7975 28543
rect 8125 28509 8159 28543
rect 9597 28509 9631 28543
rect 9686 28509 9720 28543
rect 9781 28509 9815 28543
rect 9977 28509 10011 28543
rect 15577 28509 15611 28543
rect 16681 28509 16715 28543
rect 18061 28509 18095 28543
rect 19901 28509 19935 28543
rect 19993 28509 20027 28543
rect 20637 28509 20671 28543
rect 20821 28509 20855 28543
rect 21097 28509 21131 28543
rect 22017 28509 22051 28543
rect 23213 28509 23247 28543
rect 23305 28509 23339 28543
rect 23732 28509 23766 28543
rect 25053 28509 25087 28543
rect 25145 28509 25179 28543
rect 26065 28509 26099 28543
rect 5549 28441 5583 28475
rect 8401 28441 8435 28475
rect 15393 28441 15427 28475
rect 17785 28441 17819 28475
rect 19717 28441 19751 28475
rect 3801 28373 3835 28407
rect 7757 28373 7791 28407
rect 15761 28373 15795 28407
rect 20177 28373 20211 28407
rect 21281 28373 21315 28407
rect 22753 28373 22787 28407
rect 23673 28373 23707 28407
rect 25329 28373 25363 28407
rect 26801 28373 26835 28407
rect 7389 28169 7423 28203
rect 9137 28169 9171 28203
rect 9505 28169 9539 28203
rect 11621 28169 11655 28203
rect 20545 28169 20579 28203
rect 23949 28169 23983 28203
rect 25789 28169 25823 28203
rect 14013 28101 14047 28135
rect 15301 28101 15335 28135
rect 7573 28033 7607 28067
rect 7849 28033 7883 28067
rect 8033 28033 8067 28067
rect 9413 28033 9447 28067
rect 11529 28033 11563 28067
rect 11713 28033 11747 28067
rect 13829 28033 13863 28067
rect 15117 28033 15151 28067
rect 18153 28033 18187 28067
rect 18337 28033 18371 28067
rect 19349 28033 19383 28067
rect 19533 28033 19567 28067
rect 20177 28033 20211 28067
rect 23489 28033 23523 28067
rect 23673 28033 23707 28067
rect 23765 28033 23799 28067
rect 24409 28033 24443 28067
rect 24593 28033 24627 28067
rect 25605 28033 25639 28067
rect 19717 27965 19751 27999
rect 20269 27965 20303 27999
rect 9137 27897 9171 27931
rect 9229 27829 9263 27863
rect 9321 27829 9355 27863
rect 10609 27829 10643 27863
rect 13645 27829 13679 27863
rect 14933 27829 14967 27863
rect 17417 27829 17451 27863
rect 17969 27829 18003 27863
rect 20361 27829 20395 27863
rect 23765 27829 23799 27863
rect 24593 27829 24627 27863
rect 67649 27829 67683 27863
rect 4426 27625 4460 27659
rect 8401 27625 8435 27659
rect 10241 27625 10275 27659
rect 10885 27625 10919 27659
rect 25973 27625 26007 27659
rect 27457 27625 27491 27659
rect 2421 27557 2455 27591
rect 5917 27557 5951 27591
rect 9873 27557 9907 27591
rect 1961 27489 1995 27523
rect 9965 27489 9999 27523
rect 10057 27489 10091 27523
rect 10885 27489 10919 27523
rect 10977 27489 11011 27523
rect 21097 27489 21131 27523
rect 2053 27421 2087 27455
rect 2881 27421 2915 27455
rect 4169 27421 4203 27455
rect 7757 27421 7791 27455
rect 7905 27421 7939 27455
rect 8033 27421 8067 27455
rect 8263 27421 8297 27455
rect 9781 27421 9815 27455
rect 11069 27421 11103 27455
rect 11805 27421 11839 27455
rect 14381 27421 14415 27455
rect 14565 27421 14599 27455
rect 14657 27421 14691 27455
rect 14749 27421 14783 27455
rect 15485 27421 15519 27455
rect 17785 27421 17819 27455
rect 17877 27421 17911 27455
rect 17969 27421 18003 27455
rect 18153 27421 18187 27455
rect 19901 27421 19935 27455
rect 20085 27421 20119 27455
rect 20177 27421 20211 27455
rect 20269 27421 20303 27455
rect 27721 27421 27755 27455
rect 8125 27353 8159 27387
rect 10701 27353 10735 27387
rect 12072 27353 12106 27387
rect 15025 27353 15059 27387
rect 15730 27353 15764 27387
rect 20545 27353 20579 27387
rect 21342 27353 21376 27387
rect 7205 27285 7239 27319
rect 8953 27285 8987 27319
rect 9689 27285 9723 27319
rect 13185 27285 13219 27319
rect 16865 27285 16899 27319
rect 17509 27285 17543 27319
rect 19441 27285 19475 27319
rect 22477 27285 22511 27319
rect 2053 27081 2087 27115
rect 5273 27081 5307 27115
rect 8769 27081 8803 27115
rect 11529 27081 11563 27115
rect 13461 27081 13495 27115
rect 20913 27081 20947 27115
rect 25789 27081 25823 27115
rect 27077 27081 27111 27115
rect 6653 27013 6687 27047
rect 14657 27013 14691 27047
rect 17938 27013 17972 27047
rect 20453 27013 20487 27047
rect 23314 27013 23348 27047
rect 24317 27013 24351 27047
rect 1685 26945 1719 26979
rect 2513 26945 2547 26979
rect 3321 26945 3355 26979
rect 5365 26945 5399 26979
rect 9229 26945 9263 26979
rect 9413 26945 9447 26979
rect 11805 26945 11839 26979
rect 13691 26945 13725 26979
rect 13829 26945 13863 26979
rect 13921 26945 13955 26979
rect 14105 26945 14139 26979
rect 17693 26945 17727 26979
rect 19809 26945 19843 26979
rect 19993 26945 20027 26979
rect 20085 26945 20119 26979
rect 20177 26945 20211 26979
rect 21097 26945 21131 26979
rect 21281 26945 21315 26979
rect 26985 26945 27019 26979
rect 27629 26945 27663 26979
rect 1777 26877 1811 26911
rect 3065 26877 3099 26911
rect 6377 26877 6411 26911
rect 11529 26877 11563 26911
rect 12265 26877 12299 26911
rect 13001 26877 13035 26911
rect 23581 26877 23615 26911
rect 24041 26877 24075 26911
rect 8125 26809 8159 26843
rect 9597 26809 9631 26843
rect 4445 26741 4479 26775
rect 9321 26741 9355 26775
rect 10333 26741 10367 26775
rect 10885 26741 10919 26775
rect 11713 26741 11747 26775
rect 19073 26741 19107 26775
rect 22201 26741 22235 26775
rect 7113 26537 7147 26571
rect 9505 26537 9539 26571
rect 13369 26537 13403 26571
rect 21097 26537 21131 26571
rect 25237 26537 25271 26571
rect 36829 26537 36863 26571
rect 12909 26469 12943 26503
rect 17141 26469 17175 26503
rect 11989 26401 12023 26435
rect 14657 26401 14691 26435
rect 7021 26333 7055 26367
rect 9413 26333 9447 26367
rect 10793 26333 10827 26367
rect 10977 26333 11011 26367
rect 11069 26333 11103 26367
rect 11161 26333 11195 26367
rect 13093 26333 13127 26367
rect 13185 26333 13219 26367
rect 14933 26333 14967 26367
rect 15761 26333 15795 26367
rect 21281 26333 21315 26367
rect 25329 26333 25363 26367
rect 25789 26333 25823 26367
rect 32229 26333 32263 26367
rect 32505 26333 32539 26367
rect 33977 26333 34011 26367
rect 34989 26333 35023 26367
rect 35173 26333 35207 26367
rect 35817 26333 35851 26367
rect 36093 26333 36127 26367
rect 68109 26333 68143 26367
rect 5549 26265 5583 26299
rect 7757 26265 7791 26299
rect 13369 26265 13403 26299
rect 16006 26265 16040 26299
rect 19717 26265 19751 26299
rect 10057 26197 10091 26231
rect 11437 26197 11471 26231
rect 33241 26197 33275 26231
rect 34069 26197 34103 26231
rect 35357 26197 35391 26231
rect 3157 25993 3191 26027
rect 7757 25993 7791 26027
rect 19257 25993 19291 26027
rect 34805 25993 34839 26027
rect 2697 25925 2731 25959
rect 11774 25925 11808 25959
rect 33333 25925 33367 25959
rect 2329 25857 2363 25891
rect 2513 25857 2547 25891
rect 3387 25857 3421 25891
rect 3506 25857 3540 25891
rect 3617 25857 3651 25891
rect 3801 25857 3835 25891
rect 6644 25857 6678 25891
rect 8677 25857 8711 25891
rect 8933 25857 8967 25891
rect 11529 25857 11563 25891
rect 15229 25857 15263 25891
rect 15485 25857 15519 25891
rect 16681 25857 16715 25891
rect 17877 25857 17911 25891
rect 18133 25857 18167 25891
rect 20177 25857 20211 25891
rect 22946 25857 22980 25891
rect 23673 25857 23707 25891
rect 23857 25857 23891 25891
rect 25309 25857 25343 25891
rect 35357 25857 35391 25891
rect 6377 25789 6411 25823
rect 19901 25789 19935 25823
rect 23213 25789 23247 25823
rect 25053 25789 25087 25823
rect 33057 25789 33091 25823
rect 4353 25721 4387 25755
rect 10057 25653 10091 25687
rect 12909 25653 12943 25687
rect 14105 25653 14139 25687
rect 16037 25653 16071 25687
rect 16865 25653 16899 25687
rect 21833 25653 21867 25687
rect 24041 25653 24075 25687
rect 24593 25653 24627 25687
rect 26433 25653 26467 25687
rect 35541 25653 35575 25687
rect 6561 25449 6595 25483
rect 8401 25449 8435 25483
rect 16221 25449 16255 25483
rect 17785 25449 17819 25483
rect 25145 25449 25179 25483
rect 35541 25449 35575 25483
rect 26525 25381 26559 25415
rect 33425 25381 33459 25415
rect 2881 25313 2915 25347
rect 12909 25313 12943 25347
rect 13185 25313 13219 25347
rect 21005 25313 21039 25347
rect 23857 25313 23891 25347
rect 32137 25313 32171 25347
rect 33517 25313 33551 25347
rect 3893 25245 3927 25279
rect 6837 25245 6871 25279
rect 6929 25245 6963 25279
rect 7021 25242 7055 25276
rect 7205 25245 7239 25279
rect 7757 25245 7791 25279
rect 7941 25245 7975 25279
rect 8033 25245 8067 25279
rect 8125 25245 8159 25279
rect 9781 25245 9815 25279
rect 10701 25245 10735 25279
rect 10977 25245 11011 25279
rect 14841 25245 14875 25279
rect 15117 25245 15151 25279
rect 15577 25245 15611 25279
rect 15761 25245 15795 25279
rect 15853 25245 15887 25279
rect 15945 25245 15979 25279
rect 17141 25245 17175 25279
rect 17325 25245 17359 25279
rect 17417 25245 17451 25279
rect 17509 25245 17543 25279
rect 20729 25245 20763 25279
rect 21741 25245 21775 25279
rect 24501 25245 24535 25279
rect 24685 25245 24719 25279
rect 24777 25245 24811 25279
rect 24869 25245 24903 25279
rect 27905 25245 27939 25279
rect 31033 25245 31067 25279
rect 31861 25245 31895 25279
rect 33977 25245 34011 25279
rect 34161 25245 34195 25279
rect 35357 25245 35391 25279
rect 36461 25245 36495 25279
rect 4160 25177 4194 25211
rect 23489 25177 23523 25211
rect 23673 25177 23707 25211
rect 27638 25177 27672 25211
rect 33057 25177 33091 25211
rect 36737 25177 36771 25211
rect 5273 25109 5307 25143
rect 6009 25109 6043 25143
rect 9551 25109 9585 25143
rect 18337 25109 18371 25143
rect 21557 25109 21591 25143
rect 22569 25109 22603 25143
rect 34069 25109 34103 25143
rect 38209 25109 38243 25143
rect 7021 24905 7055 24939
rect 8217 24905 8251 24939
rect 17325 24905 17359 24939
rect 34253 24905 34287 24939
rect 36093 24905 36127 24939
rect 2421 24837 2455 24871
rect 11897 24837 11931 24871
rect 16957 24837 16991 24871
rect 2605 24769 2639 24803
rect 3249 24769 3283 24803
rect 3412 24769 3446 24803
rect 3512 24775 3546 24809
rect 3617 24769 3651 24803
rect 7205 24769 7239 24803
rect 7389 24769 7423 24803
rect 8401 24769 8435 24803
rect 8585 24769 8619 24803
rect 11713 24769 11747 24803
rect 13645 24769 13679 24803
rect 14381 24769 14415 24803
rect 14565 24769 14599 24803
rect 15209 24769 15243 24803
rect 15393 24769 15427 24803
rect 15485 24769 15519 24803
rect 15577 24769 15611 24803
rect 17141 24769 17175 24803
rect 18337 24769 18371 24803
rect 18593 24769 18627 24803
rect 20177 24769 20211 24803
rect 20361 24769 20395 24803
rect 20453 24769 20487 24803
rect 20545 24769 20579 24803
rect 21833 24769 21867 24803
rect 22017 24769 22051 24803
rect 22109 24769 22143 24803
rect 22201 24769 22235 24803
rect 23765 24769 23799 24803
rect 24317 24769 24351 24803
rect 24501 24769 24535 24803
rect 24593 24769 24627 24803
rect 24685 24769 24719 24803
rect 28621 24769 28655 24803
rect 32413 24769 32447 24803
rect 32597 24769 32631 24803
rect 33241 24769 33275 24803
rect 33609 24769 33643 24803
rect 34161 24769 34195 24803
rect 34437 24769 34471 24803
rect 34621 24769 34655 24803
rect 35357 24769 35391 24803
rect 37657 24769 37691 24803
rect 37749 24769 37783 24803
rect 43177 24769 43211 24803
rect 2789 24701 2823 24735
rect 3893 24701 3927 24735
rect 13921 24701 13955 24735
rect 14749 24701 14783 24735
rect 15853 24701 15887 24735
rect 20821 24701 20855 24735
rect 23673 24701 23707 24735
rect 24961 24701 24995 24735
rect 28365 24701 28399 24735
rect 35081 24701 35115 24735
rect 39037 24701 39071 24735
rect 39313 24701 39347 24735
rect 42901 24701 42935 24735
rect 4353 24633 4387 24667
rect 5825 24633 5859 24667
rect 11529 24633 11563 24667
rect 32413 24633 32447 24667
rect 67649 24633 67683 24667
rect 6561 24565 6595 24599
rect 9137 24565 9171 24599
rect 19717 24565 19751 24599
rect 22477 24565 22511 24599
rect 23397 24565 23431 24599
rect 23765 24565 23799 24599
rect 29745 24565 29779 24599
rect 33057 24565 33091 24599
rect 33517 24565 33551 24599
rect 40785 24565 40819 24599
rect 43913 24565 43947 24599
rect 6653 24361 6687 24395
rect 8033 24361 8067 24395
rect 13093 24361 13127 24395
rect 15485 24361 15519 24395
rect 16037 24361 16071 24395
rect 17969 24361 18003 24395
rect 19901 24361 19935 24395
rect 20453 24361 20487 24395
rect 21649 24361 21683 24395
rect 24501 24361 24535 24395
rect 32781 24361 32815 24395
rect 35357 24361 35391 24395
rect 39957 24361 39991 24395
rect 41797 24361 41831 24395
rect 43269 24361 43303 24395
rect 35265 24293 35299 24327
rect 5273 24225 5307 24259
rect 11713 24225 11747 24259
rect 16865 24225 16899 24259
rect 34897 24225 34931 24259
rect 7297 24157 7331 24191
rect 7481 24157 7515 24191
rect 8125 24157 8159 24191
rect 8953 24157 8987 24191
rect 9137 24157 9171 24191
rect 9781 24157 9815 24191
rect 14105 24157 14139 24191
rect 16497 24157 16531 24191
rect 17325 24157 17359 24191
rect 17509 24157 17543 24191
rect 17601 24157 17635 24191
rect 17693 24157 17727 24191
rect 19809 24157 19843 24191
rect 19993 24157 20027 24191
rect 21281 24157 21315 24191
rect 23222 24157 23256 24191
rect 23489 24157 23523 24191
rect 24961 24157 24995 24191
rect 26801 24157 26835 24191
rect 29837 24157 29871 24191
rect 32689 24157 32723 24191
rect 32781 24157 32815 24191
rect 38669 24157 38703 24191
rect 39865 24157 39899 24191
rect 41153 24157 41187 24191
rect 42533 24157 42567 24191
rect 42809 24157 42843 24191
rect 43269 24157 43303 24191
rect 5540 24089 5574 24123
rect 10026 24089 10060 24123
rect 11958 24089 11992 24123
rect 14350 24089 14384 24123
rect 16681 24089 16715 24123
rect 21465 24089 21499 24123
rect 25206 24089 25240 24123
rect 27068 24089 27102 24123
rect 30104 24089 30138 24123
rect 32505 24089 32539 24123
rect 33241 24089 33275 24123
rect 38402 24089 38436 24123
rect 3157 24021 3191 24055
rect 4721 24021 4755 24055
rect 7481 24021 7515 24055
rect 8953 24021 8987 24055
rect 11161 24021 11195 24055
rect 18429 24021 18463 24055
rect 22109 24021 22143 24055
rect 26341 24021 26375 24055
rect 28181 24021 28215 24055
rect 31217 24021 31251 24055
rect 37289 24021 37323 24055
rect 41245 24021 41279 24055
rect 4353 23817 4387 23851
rect 5549 23817 5583 23851
rect 9413 23817 9447 23851
rect 10701 23817 10735 23851
rect 13461 23817 13495 23851
rect 17877 23817 17911 23851
rect 22385 23817 22419 23851
rect 24869 23817 24903 23851
rect 30297 23817 30331 23851
rect 37933 23817 37967 23851
rect 42625 23817 42659 23851
rect 1869 23749 1903 23783
rect 3218 23749 3252 23783
rect 21925 23749 21959 23783
rect 23397 23749 23431 23783
rect 23765 23749 23799 23783
rect 2145 23681 2179 23715
rect 2237 23681 2271 23715
rect 2329 23681 2363 23715
rect 2513 23681 2547 23715
rect 4905 23681 4939 23715
rect 5089 23681 5123 23715
rect 5184 23681 5218 23715
rect 5273 23681 5307 23715
rect 7895 23681 7929 23715
rect 8033 23681 8067 23715
rect 8125 23681 8159 23715
rect 8309 23681 8343 23715
rect 8769 23681 8803 23715
rect 8953 23681 8987 23715
rect 9064 23681 9098 23715
rect 9183 23681 9217 23715
rect 10793 23681 10827 23715
rect 13645 23681 13679 23715
rect 13829 23681 13863 23715
rect 16681 23681 16715 23715
rect 16865 23681 16899 23715
rect 16957 23681 16991 23715
rect 17049 23681 17083 23715
rect 18797 23681 18831 23715
rect 19441 23681 19475 23715
rect 19625 23681 19659 23715
rect 19717 23681 19751 23715
rect 19809 23681 19843 23715
rect 22201 23681 22235 23715
rect 23581 23681 23615 23715
rect 24225 23681 24259 23715
rect 24409 23681 24443 23715
rect 24501 23681 24535 23715
rect 24639 23681 24673 23715
rect 25329 23681 25363 23715
rect 29653 23681 29687 23715
rect 29837 23681 29871 23715
rect 29929 23681 29963 23715
rect 30021 23681 30055 23715
rect 34069 23681 34103 23715
rect 34253 23681 34287 23715
rect 36277 23681 36311 23715
rect 36461 23681 36495 23715
rect 37289 23681 37323 23715
rect 37452 23681 37486 23715
rect 37568 23681 37602 23715
rect 37657 23681 37691 23715
rect 41705 23681 41739 23715
rect 42441 23681 42475 23715
rect 42625 23681 42659 23715
rect 2973 23613 3007 23647
rect 12725 23613 12759 23647
rect 15393 23613 15427 23647
rect 15669 23613 15703 23647
rect 22109 23613 22143 23647
rect 36645 23613 36679 23647
rect 7665 23477 7699 23511
rect 9965 23477 9999 23511
rect 14381 23477 14415 23511
rect 17325 23477 17359 23511
rect 18889 23477 18923 23511
rect 20085 23477 20119 23511
rect 21925 23477 21959 23511
rect 27997 23477 28031 23511
rect 29193 23477 29227 23511
rect 33425 23477 33459 23511
rect 33885 23477 33919 23511
rect 41797 23477 41831 23511
rect 67649 23477 67683 23511
rect 2145 23273 2179 23307
rect 5181 23273 5215 23307
rect 5641 23273 5675 23307
rect 11805 23273 11839 23307
rect 13553 23273 13587 23307
rect 16589 23273 16623 23307
rect 21373 23273 21407 23307
rect 23121 23273 23155 23307
rect 26985 23273 27019 23307
rect 29929 23273 29963 23307
rect 36277 23273 36311 23307
rect 37657 23273 37691 23307
rect 41613 23273 41647 23307
rect 31493 23205 31527 23239
rect 42625 23205 42659 23239
rect 6285 23137 6319 23171
rect 8953 23137 8987 23171
rect 9229 23137 9263 23171
rect 19993 23137 20027 23171
rect 22385 23137 22419 23171
rect 32873 23137 32907 23171
rect 34897 23137 34931 23171
rect 40141 23137 40175 23171
rect 2329 23069 2363 23103
rect 4813 23069 4847 23103
rect 6552 23069 6586 23103
rect 11345 23069 11379 23103
rect 12081 23069 12115 23103
rect 12170 23069 12204 23103
rect 12270 23069 12304 23103
rect 12449 23069 12483 23103
rect 12909 23069 12943 23103
rect 13093 23069 13127 23103
rect 13188 23066 13222 23100
rect 13323 23069 13357 23103
rect 14473 23069 14507 23103
rect 15301 23069 15335 23103
rect 17325 23069 17359 23103
rect 20249 23069 20283 23103
rect 22661 23069 22695 23103
rect 24869 23069 24903 23103
rect 26525 23069 26559 23103
rect 27261 23069 27295 23103
rect 27350 23066 27384 23100
rect 27445 23066 27479 23100
rect 27629 23069 27663 23103
rect 29745 23069 29779 23103
rect 33793 23069 33827 23103
rect 33885 23069 33919 23103
rect 33977 23069 34011 23103
rect 34161 23069 34195 23103
rect 39865 23069 39899 23103
rect 43361 23069 43395 23103
rect 43637 23069 43671 23103
rect 2513 23001 2547 23035
rect 4997 23001 5031 23035
rect 16221 23001 16255 23035
rect 16405 23001 16439 23035
rect 17592 23001 17626 23035
rect 23305 23001 23339 23035
rect 23489 23001 23523 23035
rect 25053 23001 25087 23035
rect 28089 23001 28123 23035
rect 28917 23001 28951 23035
rect 29561 23001 29595 23035
rect 30389 23001 30423 23035
rect 30573 23001 30607 23035
rect 32628 23001 32662 23035
rect 33517 23001 33551 23035
rect 35142 23001 35176 23035
rect 36737 23001 36771 23035
rect 36921 23001 36955 23035
rect 3065 22933 3099 22967
rect 7665 22933 7699 22967
rect 8401 22933 8435 22967
rect 18705 22933 18739 22967
rect 30757 22933 30791 22967
rect 37105 22933 37139 22967
rect 3157 22729 3191 22763
rect 12173 22729 12207 22763
rect 14105 22729 14139 22763
rect 17785 22729 17819 22763
rect 27353 22729 27387 22763
rect 28365 22729 28399 22763
rect 34805 22729 34839 22763
rect 37657 22729 37691 22763
rect 40141 22729 40175 22763
rect 41797 22729 41831 22763
rect 2237 22661 2271 22695
rect 8861 22661 8895 22695
rect 12357 22661 12391 22695
rect 14473 22661 14507 22695
rect 15301 22661 15335 22695
rect 16129 22661 16163 22695
rect 17417 22661 17451 22695
rect 22753 22661 22787 22695
rect 23857 22661 23891 22695
rect 23949 22661 23983 22695
rect 26065 22661 26099 22695
rect 27169 22661 27203 22695
rect 36185 22661 36219 22695
rect 2421 22593 2455 22627
rect 5457 22593 5491 22627
rect 5549 22593 5583 22627
rect 5641 22593 5675 22627
rect 5825 22593 5859 22627
rect 7665 22593 7699 22627
rect 8125 22593 8159 22627
rect 10721 22593 10755 22627
rect 10977 22593 11011 22627
rect 12541 22593 12575 22627
rect 14289 22593 14323 22627
rect 15117 22593 15151 22627
rect 15761 22593 15795 22627
rect 15945 22593 15979 22627
rect 17141 22593 17175 22627
rect 17234 22593 17268 22627
rect 17509 22593 17543 22627
rect 17647 22593 17681 22627
rect 19717 22593 19751 22627
rect 19993 22593 20027 22627
rect 22656 22593 22690 22627
rect 22845 22593 22879 22627
rect 23028 22593 23062 22627
rect 23121 22593 23155 22627
rect 23719 22593 23753 22627
rect 24132 22593 24166 22627
rect 24225 22593 24259 22627
rect 24961 22593 24995 22627
rect 25053 22593 25087 22627
rect 25145 22593 25179 22627
rect 25329 22593 25363 22627
rect 25973 22593 26007 22627
rect 26157 22593 26191 22627
rect 26341 22593 26375 22627
rect 26985 22593 27019 22627
rect 28621 22593 28655 22627
rect 28733 22593 28767 22627
rect 28825 22593 28859 22627
rect 29009 22593 29043 22627
rect 29837 22593 29871 22627
rect 30021 22593 30055 22627
rect 30113 22593 30147 22627
rect 30251 22593 30285 22627
rect 33517 22593 33551 22627
rect 33701 22593 33735 22627
rect 34161 22593 34195 22627
rect 34324 22593 34358 22627
rect 34437 22593 34471 22627
rect 34575 22593 34609 22627
rect 35449 22593 35483 22627
rect 38770 22593 38804 22627
rect 39037 22593 39071 22627
rect 40049 22593 40083 22627
rect 41705 22593 41739 22627
rect 41889 22593 41923 22627
rect 42625 22593 42659 22627
rect 42809 22593 42843 22627
rect 6377 22525 6411 22559
rect 33333 22525 33367 22559
rect 24777 22457 24811 22491
rect 25789 22457 25823 22491
rect 2605 22389 2639 22423
rect 3709 22389 3743 22423
rect 5181 22389 5215 22423
rect 9597 22389 9631 22423
rect 14933 22389 14967 22423
rect 22477 22389 22511 22423
rect 23581 22389 23615 22423
rect 27905 22389 27939 22423
rect 30481 22389 30515 22423
rect 42441 22389 42475 22423
rect 6009 22185 6043 22219
rect 10885 22185 10919 22219
rect 18061 22185 18095 22219
rect 35817 22185 35851 22219
rect 25697 22117 25731 22151
rect 68109 22117 68143 22151
rect 4169 22049 4203 22083
rect 8953 22049 8987 22083
rect 17877 22049 17911 22083
rect 27721 22049 27755 22083
rect 29561 22049 29595 22083
rect 34069 22049 34103 22083
rect 35909 22049 35943 22083
rect 37841 22049 37875 22083
rect 39865 22049 39899 22083
rect 2421 21981 2455 22015
rect 2584 21981 2618 22015
rect 2684 21981 2718 22015
rect 2835 21981 2869 22015
rect 4436 21981 4470 22015
rect 6193 21981 6227 22015
rect 7389 21981 7423 22015
rect 9229 21981 9263 22015
rect 10241 21981 10275 22015
rect 10425 21981 10459 22015
rect 10517 21981 10551 22015
rect 10609 21981 10643 22015
rect 12541 21981 12575 22015
rect 12704 21981 12738 22015
rect 12817 21981 12851 22015
rect 12909 21981 12943 22015
rect 14105 21981 14139 22015
rect 16221 21981 16255 22015
rect 16313 21981 16347 22015
rect 16405 21981 16439 22015
rect 16589 21981 16623 22015
rect 17785 21981 17819 22015
rect 19436 21981 19470 22015
rect 19533 21981 19567 22015
rect 19808 21981 19842 22015
rect 19901 21981 19935 22015
rect 21833 21981 21867 22015
rect 21925 21981 21959 22015
rect 22201 21981 22235 22015
rect 22845 21981 22879 22015
rect 23029 21981 23063 22015
rect 23213 21981 23247 22015
rect 25881 21981 25915 22015
rect 25973 21981 26007 22015
rect 26249 21981 26283 22015
rect 27997 21981 28031 22015
rect 29929 21981 29963 22015
rect 30481 21981 30515 22015
rect 32146 21981 32180 22015
rect 32413 21981 32447 22015
rect 36001 21981 36035 22015
rect 37197 21981 37231 22015
rect 37381 21981 37415 22015
rect 37473 21981 37507 22015
rect 37611 21981 37645 22015
rect 38301 21981 38335 22015
rect 42073 21981 42107 22015
rect 6377 21913 6411 21947
rect 7573 21913 7607 21947
rect 8033 21913 8067 21947
rect 8217 21913 8251 21947
rect 8401 21913 8435 21947
rect 12081 21913 12115 21947
rect 13185 21913 13219 21947
rect 14350 21913 14384 21947
rect 18061 21913 18095 21947
rect 19625 21913 19659 21947
rect 22017 21913 22051 21947
rect 23121 21913 23155 21947
rect 26065 21913 26099 21947
rect 29745 21913 29779 21947
rect 35725 21913 35759 21947
rect 36645 21913 36679 21947
rect 40110 21913 40144 21947
rect 3065 21845 3099 21879
rect 5549 21845 5583 21879
rect 7205 21845 7239 21879
rect 15485 21845 15519 21879
rect 15945 21845 15979 21879
rect 17601 21845 17635 21879
rect 19257 21845 19291 21879
rect 21649 21845 21683 21879
rect 23397 21845 23431 21879
rect 24501 21845 24535 21879
rect 31033 21845 31067 21879
rect 35265 21845 35299 21879
rect 36185 21845 36219 21879
rect 41245 21845 41279 21879
rect 42257 21845 42291 21879
rect 17049 21641 17083 21675
rect 17877 21641 17911 21675
rect 20913 21641 20947 21675
rect 34713 21641 34747 21675
rect 38209 21641 38243 21675
rect 41705 21641 41739 21675
rect 43085 21641 43119 21675
rect 8585 21573 8619 21607
rect 12725 21573 12759 21607
rect 15669 21573 15703 21607
rect 18521 21573 18555 21607
rect 20085 21573 20119 21607
rect 24409 21573 24443 21607
rect 27261 21573 27295 21607
rect 29285 21573 29319 21607
rect 30450 21573 30484 21607
rect 33578 21573 33612 21607
rect 2881 21505 2915 21539
rect 3148 21505 3182 21539
rect 6644 21505 6678 21539
rect 8217 21505 8251 21539
rect 8401 21505 8435 21539
rect 9045 21505 9079 21539
rect 9229 21505 9263 21539
rect 9321 21505 9355 21539
rect 9413 21505 9447 21539
rect 11759 21505 11793 21539
rect 11910 21508 11944 21542
rect 12010 21505 12044 21539
rect 12173 21505 12207 21539
rect 15577 21505 15611 21539
rect 15761 21505 15795 21539
rect 16681 21505 16715 21539
rect 16873 21505 16907 21539
rect 17877 21505 17911 21539
rect 18061 21505 18095 21539
rect 19947 21505 19981 21539
rect 20177 21505 20211 21539
rect 20360 21505 20394 21539
rect 20453 21505 20487 21539
rect 20913 21505 20947 21539
rect 21097 21505 21131 21539
rect 22845 21505 22879 21539
rect 24179 21505 24213 21539
rect 24317 21505 24351 21539
rect 24592 21505 24626 21539
rect 24685 21505 24719 21539
rect 27721 21505 27755 21539
rect 27997 21505 28031 21539
rect 28641 21505 28675 21539
rect 28825 21508 28859 21542
rect 28917 21505 28951 21539
rect 29055 21505 29089 21539
rect 30205 21505 30239 21539
rect 33333 21505 33367 21539
rect 35449 21505 35483 21539
rect 37565 21505 37599 21539
rect 37749 21505 37783 21539
rect 37841 21505 37875 21539
rect 37933 21505 37967 21539
rect 41245 21505 41279 21539
rect 41521 21505 41555 21539
rect 42441 21505 42475 21539
rect 42625 21505 42659 21539
rect 42901 21505 42935 21539
rect 6377 21437 6411 21471
rect 22569 21437 22603 21471
rect 25145 21437 25179 21471
rect 27813 21437 27847 21471
rect 35173 21437 35207 21471
rect 41429 21437 41463 21471
rect 4261 21301 4295 21335
rect 7757 21301 7791 21335
rect 9689 21301 9723 21335
rect 10241 21301 10275 21335
rect 11529 21301 11563 21335
rect 19809 21301 19843 21335
rect 22109 21301 22143 21335
rect 24041 21301 24075 21335
rect 27813 21301 27847 21335
rect 28181 21301 28215 21335
rect 31585 21301 31619 21335
rect 32505 21301 32539 21335
rect 36645 21301 36679 21335
rect 38669 21301 38703 21335
rect 41521 21301 41555 21335
rect 2615 21097 2649 21131
rect 6837 21097 6871 21131
rect 7941 21097 7975 21131
rect 8401 21097 8435 21131
rect 16681 21097 16715 21131
rect 17693 21097 17727 21131
rect 21465 21097 21499 21131
rect 27721 21097 27755 21131
rect 28273 21097 28307 21131
rect 28917 21097 28951 21131
rect 30113 21097 30147 21131
rect 30573 21097 30607 21131
rect 31033 21097 31067 21131
rect 35725 21097 35759 21131
rect 37565 21097 37599 21131
rect 38301 21097 38335 21131
rect 38669 21097 38703 21131
rect 3249 21029 3283 21063
rect 24409 21029 24443 21063
rect 36185 21029 36219 21063
rect 22661 20961 22695 20995
rect 22937 20961 22971 20995
rect 30757 20961 30791 20995
rect 35817 20961 35851 20995
rect 38393 20961 38427 20995
rect 41797 20961 41831 20995
rect 1593 20893 1627 20927
rect 1869 20893 1903 20927
rect 7093 20893 7127 20927
rect 7205 20893 7239 20927
rect 7302 20893 7336 20927
rect 7481 20893 7515 20927
rect 8125 20893 8159 20927
rect 8217 20893 8251 20927
rect 9597 20893 9631 20927
rect 9853 20893 9887 20927
rect 11621 20893 11655 20927
rect 11877 20893 11911 20927
rect 14105 20893 14139 20927
rect 14381 20893 14415 20927
rect 14473 20893 14507 20927
rect 15301 20893 15335 20927
rect 15568 20893 15602 20927
rect 17877 20893 17911 20927
rect 17969 20893 18003 20927
rect 18153 20893 18187 20927
rect 18245 20893 18279 20927
rect 19436 20893 19470 20927
rect 19533 20893 19567 20927
rect 19808 20893 19842 20927
rect 19901 20893 19935 20927
rect 21649 20893 21683 20927
rect 21741 20893 21775 20927
rect 22017 20893 22051 20927
rect 24547 20893 24581 20927
rect 24961 20893 24995 20927
rect 26341 20893 26375 20927
rect 28181 20893 28215 20927
rect 28365 20893 28399 20927
rect 29009 20893 29043 20927
rect 29561 20893 29595 20927
rect 29653 20893 29687 20927
rect 29837 20893 29871 20927
rect 29929 20893 29963 20927
rect 30849 20893 30883 20927
rect 32229 20893 32263 20927
rect 32413 20893 32447 20927
rect 33333 20893 33367 20927
rect 33609 20893 33643 20927
rect 34713 20893 34747 20927
rect 36001 20893 36035 20927
rect 37381 20893 37415 20927
rect 38301 20893 38335 20927
rect 41521 20893 41555 20927
rect 41613 20893 41647 20927
rect 41889 20893 41923 20927
rect 8401 20825 8435 20859
rect 13461 20825 13495 20859
rect 14289 20825 14323 20859
rect 19625 20825 19659 20859
rect 21833 20825 21867 20859
rect 24685 20825 24719 20859
rect 24777 20825 24811 20859
rect 25421 20825 25455 20859
rect 25605 20825 25639 20859
rect 26586 20825 26620 20859
rect 30573 20825 30607 20859
rect 35725 20825 35759 20859
rect 37197 20825 37231 20859
rect 39129 20825 39163 20859
rect 40785 20825 40819 20859
rect 5641 20757 5675 20791
rect 6377 20757 6411 20791
rect 9045 20757 9079 20791
rect 10977 20757 11011 20791
rect 13001 20757 13035 20791
rect 14657 20757 14691 20791
rect 17141 20757 17175 20791
rect 19257 20757 19291 20791
rect 20729 20757 20763 20791
rect 25789 20757 25823 20791
rect 31677 20757 31711 20791
rect 32597 20757 32631 20791
rect 34897 20757 34931 20791
rect 36645 20757 36679 20791
rect 41337 20757 41371 20791
rect 7481 20553 7515 20587
rect 12173 20553 12207 20587
rect 15301 20553 15335 20587
rect 17785 20553 17819 20587
rect 22017 20553 22051 20587
rect 24593 20553 24627 20587
rect 32965 20553 32999 20587
rect 36461 20553 36495 20587
rect 38025 20553 38059 20587
rect 41245 20553 41279 20587
rect 42901 20553 42935 20587
rect 5457 20485 5491 20519
rect 7941 20485 7975 20519
rect 12357 20485 12391 20519
rect 12541 20485 12575 20519
rect 14105 20485 14139 20519
rect 16681 20485 16715 20519
rect 20361 20485 20395 20519
rect 22201 20485 22235 20519
rect 27261 20485 27295 20519
rect 34345 20485 34379 20519
rect 37565 20485 37599 20519
rect 1961 20417 1995 20451
rect 5549 20417 5583 20451
rect 6561 20417 6595 20451
rect 10149 20417 10183 20451
rect 14289 20417 14323 20451
rect 15485 20417 15519 20451
rect 15761 20417 15795 20451
rect 16865 20417 16899 20451
rect 17693 20417 17727 20451
rect 20177 20417 20211 20451
rect 20269 20417 20303 20451
rect 20545 20417 20579 20451
rect 21833 20417 21867 20451
rect 21925 20417 21959 20451
rect 22109 20417 22143 20451
rect 22293 20417 22327 20451
rect 23169 20417 23203 20451
rect 23305 20417 23339 20451
rect 23397 20417 23431 20451
rect 23580 20417 23614 20451
rect 23673 20417 23707 20451
rect 24409 20417 24443 20451
rect 27445 20417 27479 20451
rect 28273 20417 28307 20451
rect 31493 20417 31527 20451
rect 32321 20417 32355 20451
rect 32500 20417 32534 20451
rect 32597 20417 32631 20451
rect 32709 20417 32743 20451
rect 33517 20417 33551 20451
rect 34529 20417 34563 20451
rect 35081 20417 35115 20451
rect 35337 20417 35371 20451
rect 37841 20417 37875 20451
rect 39109 20417 39143 20451
rect 41613 20417 41647 20451
rect 42441 20417 42475 20451
rect 42717 20417 42751 20451
rect 1685 20349 1719 20383
rect 4629 20349 4663 20383
rect 4905 20349 4939 20383
rect 8677 20349 8711 20383
rect 9873 20349 9907 20383
rect 15669 20349 15703 20383
rect 18337 20349 18371 20383
rect 25329 20349 25363 20383
rect 29009 20349 29043 20383
rect 37657 20349 37691 20383
rect 38853 20349 38887 20383
rect 40693 20349 40727 20383
rect 41705 20349 41739 20383
rect 41889 20349 41923 20383
rect 42533 20349 42567 20383
rect 2697 20281 2731 20315
rect 19993 20281 20027 20315
rect 33701 20281 33735 20315
rect 3157 20213 3191 20247
rect 6377 20213 6411 20247
rect 14473 20213 14507 20247
rect 15485 20213 15519 20247
rect 21189 20213 21223 20247
rect 23029 20213 23063 20247
rect 25559 20213 25593 20247
rect 27629 20213 27663 20247
rect 30941 20213 30975 20247
rect 34161 20213 34195 20247
rect 37749 20213 37783 20247
rect 40233 20213 40267 20247
rect 42441 20213 42475 20247
rect 67649 20213 67683 20247
rect 8125 20009 8159 20043
rect 8401 20009 8435 20043
rect 22569 20009 22603 20043
rect 24685 20009 24719 20043
rect 26157 20009 26191 20043
rect 26801 20009 26835 20043
rect 30205 20009 30239 20043
rect 32137 20009 32171 20043
rect 34161 20009 34195 20043
rect 37933 20009 37967 20043
rect 40141 20009 40175 20043
rect 40601 20009 40635 20043
rect 42165 20009 42199 20043
rect 8033 19873 8067 19907
rect 19533 19873 19567 19907
rect 20545 19873 20579 19907
rect 23029 19873 23063 19907
rect 30573 19873 30607 19907
rect 31769 19873 31803 19907
rect 36277 19873 36311 19907
rect 40233 19873 40267 19907
rect 41061 19873 41095 19907
rect 2329 19805 2363 19839
rect 4997 19805 5031 19839
rect 7113 19805 7147 19839
rect 7205 19805 7239 19839
rect 7297 19805 7331 19839
rect 7481 19805 7515 19839
rect 8217 19805 8251 19839
rect 8953 19805 8987 19839
rect 9116 19802 9150 19836
rect 9229 19805 9263 19839
rect 9321 19805 9355 19839
rect 11437 19805 11471 19839
rect 15853 19805 15887 19839
rect 16129 19805 16163 19839
rect 16221 19805 16255 19839
rect 17141 19805 17175 19839
rect 17417 19805 17451 19839
rect 17509 19805 17543 19839
rect 18153 19805 18187 19839
rect 18429 19805 18463 19839
rect 18521 19805 18555 19839
rect 19257 19805 19291 19839
rect 20821 19805 20855 19839
rect 22201 19805 22235 19839
rect 22385 19805 22419 19839
rect 23305 19805 23339 19839
rect 25513 19805 25547 19839
rect 25697 19805 25731 19839
rect 25789 19805 25823 19839
rect 25881 19805 25915 19839
rect 26617 19805 26651 19839
rect 27721 19805 27755 19839
rect 27905 19805 27939 19839
rect 27997 19805 28031 19839
rect 28089 19805 28123 19839
rect 30481 19805 30515 19839
rect 30665 19805 30699 19839
rect 30941 19805 30975 19839
rect 31953 19805 31987 19839
rect 32597 19805 32631 19839
rect 32781 19805 32815 19839
rect 33517 19805 33551 19839
rect 33701 19805 33735 19839
rect 33793 19805 33827 19839
rect 33885 19805 33919 19839
rect 37289 19805 37323 19839
rect 37452 19805 37486 19839
rect 37565 19805 37599 19839
rect 37703 19805 37737 19839
rect 38393 19805 38427 19839
rect 40141 19805 40175 19839
rect 40417 19805 40451 19839
rect 5264 19737 5298 19771
rect 6837 19737 6871 19771
rect 7941 19737 7975 19771
rect 9597 19737 9631 19771
rect 11170 19737 11204 19771
rect 13553 19737 13587 19771
rect 14473 19737 14507 19771
rect 15301 19737 15335 19771
rect 16037 19737 16071 19771
rect 17325 19737 17359 19771
rect 18337 19737 18371 19771
rect 24961 19737 24995 19771
rect 28825 19737 28859 19771
rect 35449 19737 35483 19771
rect 38945 19737 38979 19771
rect 41613 19737 41647 19771
rect 2145 19669 2179 19703
rect 6377 19669 6411 19703
rect 10057 19669 10091 19703
rect 16405 19669 16439 19703
rect 17693 19669 17727 19703
rect 18705 19669 18739 19703
rect 28365 19669 28399 19703
rect 30849 19669 30883 19703
rect 32781 19669 32815 19703
rect 34897 19669 34931 19703
rect 2237 19465 2271 19499
rect 8769 19465 8803 19499
rect 13553 19465 13587 19499
rect 15485 19465 15519 19499
rect 16681 19465 16715 19499
rect 18245 19465 18279 19499
rect 24777 19465 24811 19499
rect 29745 19465 29779 19499
rect 37289 19465 37323 19499
rect 6377 19397 6411 19431
rect 8401 19397 8435 19431
rect 28632 19397 28666 19431
rect 36185 19397 36219 19431
rect 37657 19397 37691 19431
rect 38117 19397 38151 19431
rect 38945 19397 38979 19431
rect 39497 19397 39531 19431
rect 2421 19329 2455 19363
rect 6561 19329 6595 19363
rect 8585 19329 8619 19363
rect 12173 19329 12207 19363
rect 12440 19329 12474 19363
rect 15669 19329 15703 19363
rect 16865 19329 16899 19363
rect 17509 19329 17543 19363
rect 17693 19329 17727 19363
rect 20453 19329 20487 19363
rect 22109 19329 22143 19363
rect 23489 19329 23523 19363
rect 24593 19329 24627 19363
rect 24777 19329 24811 19363
rect 25513 19329 25547 19363
rect 25697 19329 25731 19363
rect 25789 19329 25823 19363
rect 25927 19329 25961 19363
rect 28365 19329 28399 19363
rect 31033 19329 31067 19363
rect 31125 19329 31159 19363
rect 32597 19329 32631 19363
rect 33701 19329 33735 19363
rect 34989 19329 35023 19363
rect 36277 19329 36311 19363
rect 37473 19329 37507 19363
rect 38301 19329 38335 19363
rect 40049 19329 40083 19363
rect 40785 19329 40819 19363
rect 2605 19261 2639 19295
rect 6745 19261 6779 19295
rect 9781 19261 9815 19295
rect 14749 19261 14783 19295
rect 15025 19261 15059 19295
rect 17049 19261 17083 19295
rect 18889 19261 18923 19295
rect 19165 19261 19199 19295
rect 20177 19261 20211 19295
rect 21833 19261 21867 19295
rect 23213 19261 23247 19295
rect 33425 19261 33459 19295
rect 34713 19261 34747 19295
rect 40693 19261 40727 19295
rect 41613 19261 41647 19295
rect 27077 19193 27111 19227
rect 7297 19125 7331 19159
rect 7849 19125 7883 19159
rect 17601 19125 17635 19159
rect 26157 19125 26191 19159
rect 27629 19125 27663 19159
rect 32689 19125 32723 19159
rect 38485 19125 38519 19159
rect 41061 19125 41095 19159
rect 7297 18921 7331 18955
rect 14105 18921 14139 18955
rect 15577 18921 15611 18955
rect 24777 18921 24811 18955
rect 25605 18921 25639 18955
rect 30297 18921 30331 18955
rect 39313 18921 39347 18955
rect 40233 18921 40267 18955
rect 19349 18853 19383 18887
rect 22753 18853 22787 18887
rect 23857 18853 23891 18887
rect 41797 18853 41831 18887
rect 1501 18785 1535 18819
rect 10333 18785 10367 18819
rect 18613 18785 18647 18819
rect 20545 18785 20579 18819
rect 30021 18785 30055 18819
rect 34161 18785 34195 18819
rect 41337 18785 41371 18819
rect 1777 18717 1811 18751
rect 5089 18717 5123 18751
rect 5641 18717 5675 18751
rect 13553 18717 13587 18751
rect 14335 18717 14369 18751
rect 14473 18717 14507 18751
rect 14565 18717 14599 18751
rect 14749 18717 14783 18751
rect 15209 18717 15243 18751
rect 15393 18717 15427 18751
rect 16037 18717 16071 18751
rect 19533 18717 19567 18751
rect 20821 18717 20855 18751
rect 21557 18717 21591 18751
rect 21925 18717 21959 18751
rect 22477 18717 22511 18751
rect 25237 18717 25271 18751
rect 26341 18717 26375 18751
rect 26608 18717 26642 18751
rect 29929 18717 29963 18751
rect 33149 18717 33183 18751
rect 33793 18717 33827 18751
rect 34713 18717 34747 18751
rect 34897 18717 34931 18751
rect 34989 18717 35023 18751
rect 35081 18717 35115 18751
rect 36829 18717 36863 18751
rect 37013 18717 37047 18751
rect 37105 18717 37139 18751
rect 37197 18717 37231 18751
rect 37933 18717 37967 18751
rect 41429 18717 41463 18751
rect 68109 18717 68143 18751
rect 10578 18649 10612 18683
rect 18346 18649 18380 18683
rect 21649 18649 21683 18683
rect 21741 18649 21775 18683
rect 25421 18649 25455 18683
rect 32882 18649 32916 18683
rect 33977 18649 34011 18683
rect 36001 18649 36035 18683
rect 36185 18649 36219 18683
rect 37473 18649 37507 18683
rect 38178 18649 38212 18683
rect 2513 18581 2547 18615
rect 4997 18581 5031 18615
rect 11713 18581 11747 18615
rect 16221 18581 16255 18615
rect 16773 18581 16807 18615
rect 17233 18581 17267 18615
rect 21373 18581 21407 18615
rect 27721 18581 27755 18615
rect 31769 18581 31803 18615
rect 35357 18581 35391 18615
rect 36369 18581 36403 18615
rect 2881 18377 2915 18411
rect 10333 18377 10367 18411
rect 10885 18377 10919 18411
rect 17601 18377 17635 18411
rect 18337 18377 18371 18411
rect 32137 18377 32171 18411
rect 36185 18377 36219 18411
rect 40417 18377 40451 18411
rect 14657 18309 14691 18343
rect 19441 18309 19475 18343
rect 20146 18309 20180 18343
rect 23704 18309 23738 18343
rect 24409 18309 24443 18343
rect 25605 18309 25639 18343
rect 27629 18309 27663 18343
rect 28816 18309 28850 18343
rect 35072 18309 35106 18343
rect 38117 18309 38151 18343
rect 39282 18309 39316 18343
rect 2421 18241 2455 18275
rect 6745 18241 6779 18275
rect 6837 18241 6871 18275
rect 6929 18241 6963 18275
rect 7113 18241 7147 18275
rect 8024 18241 8058 18275
rect 9689 18241 9723 18275
rect 9873 18241 9907 18275
rect 9965 18241 9999 18275
rect 10057 18241 10091 18275
rect 14841 18241 14875 18275
rect 15025 18241 15059 18275
rect 15715 18241 15749 18275
rect 15853 18241 15887 18275
rect 15950 18241 15984 18275
rect 16129 18241 16163 18275
rect 16957 18241 16991 18275
rect 17120 18241 17154 18275
rect 17233 18241 17267 18275
rect 17325 18241 17359 18275
rect 18797 18241 18831 18275
rect 18981 18241 19015 18275
rect 19073 18241 19107 18275
rect 19211 18241 19245 18275
rect 19901 18241 19935 18275
rect 21833 18241 21867 18275
rect 24685 18241 24719 18275
rect 24777 18241 24811 18275
rect 24869 18241 24903 18275
rect 25053 18241 25087 18275
rect 25789 18241 25823 18275
rect 27905 18241 27939 18275
rect 32689 18241 32723 18275
rect 34805 18241 34839 18275
rect 37473 18241 37507 18275
rect 37657 18241 37691 18275
rect 37749 18241 37783 18275
rect 37841 18241 37875 18275
rect 39037 18241 39071 18275
rect 4353 18173 4387 18207
rect 4629 18173 4663 18207
rect 7757 18173 7791 18207
rect 23949 18173 23983 18207
rect 27721 18173 27755 18207
rect 28549 18173 28583 18207
rect 34345 18173 34379 18207
rect 22017 18105 22051 18139
rect 33425 18105 33459 18139
rect 2329 18037 2363 18071
rect 6469 18037 6503 18071
rect 9137 18037 9171 18071
rect 14105 18037 14139 18071
rect 15485 18037 15519 18071
rect 21281 18037 21315 18071
rect 22569 18037 22603 18071
rect 25973 18037 26007 18071
rect 27721 18037 27755 18071
rect 28089 18037 28123 18071
rect 29929 18037 29963 18071
rect 32873 18037 32907 18071
rect 36645 18037 36679 18071
rect 1961 17833 1995 17867
rect 8033 17833 8067 17867
rect 10333 17833 10367 17867
rect 14105 17833 14139 17867
rect 19625 17833 19659 17867
rect 21465 17833 21499 17867
rect 22845 17833 22879 17867
rect 23765 17833 23799 17867
rect 24777 17833 24811 17867
rect 27997 17833 28031 17867
rect 32689 17833 32723 17867
rect 17785 17765 17819 17799
rect 21005 17765 21039 17799
rect 31401 17765 31435 17799
rect 12173 17697 12207 17731
rect 16221 17697 16255 17731
rect 26617 17697 26651 17731
rect 1961 17629 1995 17663
rect 2145 17629 2179 17663
rect 6386 17629 6420 17663
rect 6653 17629 6687 17663
rect 7389 17629 7423 17663
rect 7573 17629 7607 17663
rect 7665 17629 7699 17663
rect 7757 17629 7791 17663
rect 9321 17629 9355 17663
rect 9965 17629 9999 17663
rect 10149 17629 10183 17663
rect 15229 17629 15263 17663
rect 15485 17629 15519 17663
rect 15945 17629 15979 17663
rect 19441 17629 19475 17663
rect 21649 17629 21683 17663
rect 21741 17629 21775 17663
rect 24409 17629 24443 17663
rect 25519 17629 25553 17663
rect 25697 17629 25731 17663
rect 25789 17629 25823 17663
rect 25881 17629 25915 17663
rect 31309 17629 31343 17663
rect 31493 17629 31527 17663
rect 32945 17629 32979 17663
rect 33057 17629 33091 17663
rect 33170 17626 33204 17660
rect 33333 17629 33367 17663
rect 36829 17629 36863 17663
rect 38485 17629 38519 17663
rect 68109 17629 68143 17663
rect 8953 17561 8987 17595
rect 9137 17561 9171 17595
rect 11345 17561 11379 17595
rect 11529 17561 11563 17595
rect 12418 17561 12452 17595
rect 18613 17561 18647 17595
rect 19257 17561 19291 17595
rect 24593 17561 24627 17595
rect 26157 17561 26191 17595
rect 26862 17561 26896 17595
rect 37013 17561 37047 17595
rect 37657 17561 37691 17595
rect 37841 17561 37875 17595
rect 5273 17493 5307 17527
rect 11713 17493 11747 17527
rect 13553 17493 13587 17527
rect 17233 17493 17267 17527
rect 20361 17493 20395 17527
rect 22293 17493 22327 17527
rect 32229 17493 32263 17527
rect 34805 17493 34839 17527
rect 36277 17493 36311 17527
rect 37197 17493 37231 17527
rect 38025 17493 38059 17527
rect 1409 17289 1443 17323
rect 1593 17289 1627 17323
rect 5825 17289 5859 17323
rect 12265 17289 12299 17323
rect 21925 17289 21959 17323
rect 29009 17289 29043 17323
rect 40417 17289 40451 17323
rect 5641 17221 5675 17255
rect 10701 17221 10735 17255
rect 23704 17221 23738 17255
rect 24869 17221 24903 17255
rect 37933 17221 37967 17255
rect 39282 17221 39316 17255
rect 1590 17153 1624 17187
rect 2743 17153 2777 17187
rect 2881 17153 2915 17187
rect 2973 17153 3007 17187
rect 3157 17153 3191 17187
rect 3617 17153 3651 17187
rect 3873 17153 3907 17187
rect 5457 17153 5491 17187
rect 7389 17153 7423 17187
rect 8125 17153 8159 17187
rect 8309 17153 8343 17187
rect 8401 17153 8435 17187
rect 8493 17153 8527 17187
rect 9229 17153 9263 17187
rect 10885 17153 10919 17187
rect 11621 17153 11655 17187
rect 11805 17153 11839 17187
rect 11897 17153 11931 17187
rect 11989 17153 12023 17187
rect 12725 17153 12759 17187
rect 15485 17153 15519 17187
rect 15669 17153 15703 17187
rect 15761 17153 15795 17187
rect 15899 17153 15933 17187
rect 16670 17153 16704 17187
rect 16937 17153 16971 17187
rect 19257 17153 19291 17187
rect 19441 17153 19475 17187
rect 19533 17153 19567 17187
rect 19625 17153 19659 17187
rect 21281 17153 21315 17187
rect 22109 17153 22143 17187
rect 23949 17153 23983 17187
rect 25125 17153 25159 17187
rect 25237 17153 25271 17187
rect 25329 17159 25363 17193
rect 25513 17153 25547 17187
rect 28365 17153 28399 17187
rect 28528 17153 28562 17187
rect 28641 17153 28675 17187
rect 28733 17153 28767 17187
rect 30461 17153 30495 17187
rect 33241 17153 33275 17187
rect 35826 17153 35860 17187
rect 36093 17153 36127 17187
rect 37289 17153 37323 17187
rect 37473 17153 37507 17187
rect 37565 17153 37599 17187
rect 37703 17153 37737 17187
rect 39037 17153 39071 17187
rect 2053 17085 2087 17119
rect 2513 17085 2547 17119
rect 7665 17085 7699 17119
rect 16129 17085 16163 17119
rect 27905 17085 27939 17119
rect 30205 17085 30239 17119
rect 32965 17085 32999 17119
rect 18797 17017 18831 17051
rect 21097 17017 21131 17051
rect 1961 16949 1995 16983
rect 4997 16949 5031 16983
rect 8769 16949 8803 16983
rect 18061 16949 18095 16983
rect 19901 16949 19935 16983
rect 20453 16949 20487 16983
rect 22569 16949 22603 16983
rect 26341 16949 26375 16983
rect 31585 16949 31619 16983
rect 34713 16949 34747 16983
rect 36737 16949 36771 16983
rect 2053 16745 2087 16779
rect 2513 16745 2547 16779
rect 4353 16745 4387 16779
rect 7573 16745 7607 16779
rect 15669 16745 15703 16779
rect 25237 16745 25271 16779
rect 26525 16745 26559 16779
rect 28641 16745 28675 16779
rect 29929 16745 29963 16779
rect 32873 16745 32907 16779
rect 35357 16745 35391 16779
rect 35817 16745 35851 16779
rect 36829 16745 36863 16779
rect 3893 16677 3927 16711
rect 8125 16677 8159 16711
rect 16497 16677 16531 16711
rect 22201 16677 22235 16711
rect 2421 16609 2455 16643
rect 5917 16609 5951 16643
rect 8953 16609 8987 16643
rect 12173 16609 12207 16643
rect 20361 16609 20395 16643
rect 23397 16609 23431 16643
rect 26985 16609 27019 16643
rect 27813 16609 27847 16643
rect 33057 16609 33091 16643
rect 34161 16609 34195 16643
rect 2237 16541 2271 16575
rect 4537 16541 4571 16575
rect 5641 16541 5675 16575
rect 7481 16541 7515 16575
rect 7665 16541 7699 16575
rect 9209 16541 9243 16575
rect 11069 16541 11103 16575
rect 11253 16541 11287 16575
rect 11345 16541 11379 16575
rect 11437 16541 11471 16575
rect 19533 16541 19567 16575
rect 19625 16541 19659 16575
rect 19717 16541 19751 16575
rect 19901 16541 19935 16575
rect 20617 16541 20651 16575
rect 24869 16541 24903 16575
rect 25053 16541 25087 16575
rect 25697 16541 25731 16575
rect 30159 16541 30193 16575
rect 30310 16535 30344 16569
rect 30410 16541 30444 16575
rect 30573 16541 30607 16575
rect 31217 16541 31251 16575
rect 32873 16541 32907 16575
rect 34713 16541 34747 16575
rect 34897 16541 34931 16575
rect 34989 16541 35023 16575
rect 35081 16541 35115 16575
rect 37289 16541 37323 16575
rect 37452 16538 37486 16572
rect 37552 16541 37586 16575
rect 37703 16541 37737 16575
rect 2513 16473 2547 16507
rect 4721 16473 4755 16507
rect 11713 16473 11747 16507
rect 12418 16473 12452 16507
rect 15853 16473 15887 16507
rect 16037 16473 16071 16507
rect 22385 16473 22419 16507
rect 28273 16473 28307 16507
rect 28457 16473 28491 16507
rect 31033 16473 31067 16507
rect 33149 16473 33183 16507
rect 33793 16473 33827 16507
rect 33977 16473 34011 16507
rect 7021 16405 7055 16439
rect 10333 16405 10367 16439
rect 13553 16405 13587 16439
rect 19257 16405 19291 16439
rect 21741 16405 21775 16439
rect 25881 16405 25915 16439
rect 31401 16405 31435 16439
rect 32689 16405 32723 16439
rect 37933 16405 37967 16439
rect 9413 16201 9447 16235
rect 10977 16201 11011 16235
rect 18245 16201 18279 16235
rect 19349 16201 19383 16235
rect 20545 16201 20579 16235
rect 22937 16201 22971 16235
rect 23581 16201 23615 16235
rect 40049 16201 40083 16235
rect 10609 16133 10643 16167
rect 10793 16133 10827 16167
rect 14933 16133 14967 16167
rect 17785 16133 17819 16167
rect 18981 16133 19015 16167
rect 19165 16133 19199 16167
rect 25452 16133 25486 16167
rect 28181 16133 28215 16167
rect 38914 16133 38948 16167
rect 2973 16065 3007 16099
rect 3157 16068 3191 16102
rect 3249 16065 3283 16099
rect 3387 16065 3421 16099
rect 4077 16065 4111 16099
rect 5825 16065 5859 16099
rect 6745 16065 6779 16099
rect 6837 16065 6871 16099
rect 7021 16065 7055 16099
rect 7113 16065 7147 16099
rect 9505 16065 9539 16099
rect 11529 16065 11563 16099
rect 14565 16065 14599 16099
rect 14658 16065 14692 16099
rect 14841 16065 14875 16099
rect 15030 16065 15064 16099
rect 17969 16065 18003 16099
rect 18061 16065 18095 16099
rect 21097 16065 21131 16099
rect 22569 16065 22603 16099
rect 23029 16065 23063 16099
rect 23765 16065 23799 16099
rect 25697 16065 25731 16099
rect 26985 16065 27019 16099
rect 28411 16065 28445 16099
rect 28549 16065 28583 16099
rect 28641 16065 28675 16099
rect 28825 16065 28859 16099
rect 30757 16065 30791 16099
rect 33250 16065 33284 16099
rect 33517 16065 33551 16099
rect 35541 16065 35575 16099
rect 35704 16065 35738 16099
rect 35817 16065 35851 16099
rect 35955 16065 35989 16099
rect 37473 16065 37507 16099
rect 37657 16065 37691 16099
rect 38669 16065 38703 16099
rect 11805 15997 11839 16031
rect 21281 15997 21315 16031
rect 26341 15997 26375 16031
rect 31033 15997 31067 16031
rect 34805 15997 34839 16031
rect 35081 15997 35115 16031
rect 22293 15929 22327 15963
rect 22661 15929 22695 15963
rect 3617 15861 3651 15895
rect 5641 15861 5675 15895
rect 6561 15861 6595 15895
rect 15209 15861 15243 15895
rect 18061 15861 18095 15895
rect 22753 15861 22787 15895
rect 24317 15861 24351 15895
rect 27169 15861 27203 15895
rect 29653 15861 29687 15895
rect 32137 15861 32171 15895
rect 36185 15861 36219 15895
rect 37289 15861 37323 15895
rect 67649 15861 67683 15895
rect 1501 15657 1535 15691
rect 2789 15657 2823 15691
rect 7205 15657 7239 15691
rect 11069 15657 11103 15691
rect 11529 15657 11563 15691
rect 11989 15657 12023 15691
rect 14841 15657 14875 15691
rect 18521 15657 18555 15691
rect 19625 15657 19659 15691
rect 24593 15657 24627 15691
rect 28641 15657 28675 15691
rect 32873 15657 32907 15691
rect 36921 15657 36955 15691
rect 9505 15589 9539 15623
rect 23305 15589 23339 15623
rect 25421 15589 25455 15623
rect 34069 15589 34103 15623
rect 7205 15521 7239 15555
rect 7297 15521 7331 15555
rect 30941 15521 30975 15555
rect 31493 15521 31527 15555
rect 34713 15521 34747 15555
rect 1685 15453 1719 15487
rect 1961 15453 1995 15487
rect 2145 15453 2179 15487
rect 2789 15453 2823 15487
rect 2881 15453 2915 15487
rect 3801 15453 3835 15487
rect 4057 15453 4091 15487
rect 6193 15453 6227 15487
rect 6285 15453 6319 15487
rect 6469 15453 6503 15487
rect 6561 15453 6595 15487
rect 7389 15453 7423 15487
rect 7849 15453 7883 15487
rect 8033 15453 8067 15487
rect 8217 15453 8251 15487
rect 8953 15453 8987 15487
rect 9137 15453 9171 15487
rect 9321 15453 9355 15487
rect 10057 15453 10091 15487
rect 10333 15453 10367 15487
rect 10425 15453 10459 15487
rect 11253 15453 11287 15487
rect 11345 15453 11379 15487
rect 11529 15453 11563 15487
rect 12173 15453 12207 15487
rect 12357 15453 12391 15487
rect 12909 15453 12943 15487
rect 13057 15453 13091 15487
rect 13415 15453 13449 15487
rect 14749 15453 14783 15487
rect 14933 15453 14967 15487
rect 15577 15453 15611 15487
rect 15853 15453 15887 15487
rect 16865 15453 16899 15487
rect 17013 15453 17047 15487
rect 17233 15453 17267 15487
rect 17330 15453 17364 15487
rect 19441 15453 19475 15487
rect 24409 15453 24443 15487
rect 25237 15453 25271 15487
rect 27445 15453 27479 15487
rect 29837 15453 29871 15487
rect 29929 15453 29963 15487
rect 30021 15453 30055 15487
rect 30205 15453 30239 15487
rect 31769 15453 31803 15487
rect 33149 15453 33183 15487
rect 33241 15453 33275 15487
rect 33333 15453 33367 15487
rect 33517 15453 33551 15487
rect 34897 15453 34931 15487
rect 35541 15453 35575 15487
rect 35808 15453 35842 15487
rect 39313 15453 39347 15487
rect 3065 15385 3099 15419
rect 6009 15385 6043 15419
rect 7021 15385 7055 15419
rect 8125 15385 8159 15419
rect 9229 15385 9263 15419
rect 10241 15385 10275 15419
rect 13185 15385 13219 15419
rect 13277 15385 13311 15419
rect 17141 15385 17175 15419
rect 18613 15385 18647 15419
rect 19257 15385 19291 15419
rect 20913 15385 20947 15419
rect 22017 15385 22051 15419
rect 27200 15385 27234 15419
rect 28273 15385 28307 15419
rect 28457 15385 28491 15419
rect 35081 15385 35115 15419
rect 39046 15385 39080 15419
rect 2605 15317 2639 15351
rect 5181 15317 5215 15351
rect 8401 15317 8435 15351
rect 10609 15317 10643 15351
rect 13553 15317 13587 15351
rect 14289 15317 14323 15351
rect 17509 15317 17543 15351
rect 21557 15317 21591 15351
rect 26065 15317 26099 15351
rect 29561 15317 29595 15351
rect 37933 15317 37967 15351
rect 3341 15113 3375 15147
rect 4905 15113 4939 15147
rect 8217 15113 8251 15147
rect 9505 15113 9539 15147
rect 11805 15113 11839 15147
rect 20269 15113 20303 15147
rect 21833 15113 21867 15147
rect 22845 15113 22879 15147
rect 27997 15113 28031 15147
rect 29653 15113 29687 15147
rect 30665 15113 30699 15147
rect 31401 15113 31435 15147
rect 33885 15113 33919 15147
rect 36645 15113 36679 15147
rect 37933 15113 37967 15147
rect 40509 15113 40543 15147
rect 12817 15045 12851 15079
rect 14381 15045 14415 15079
rect 15853 15045 15887 15079
rect 17601 15045 17635 15079
rect 17693 15045 17727 15079
rect 18429 15045 18463 15079
rect 19156 15045 19190 15079
rect 22201 15045 22235 15079
rect 25237 15045 25271 15079
rect 27261 15045 27295 15079
rect 29285 15045 29319 15079
rect 33517 15045 33551 15079
rect 33701 15045 33735 15079
rect 2973 14977 3007 15011
rect 3157 14977 3191 15011
rect 5089 14977 5123 15011
rect 5365 14977 5399 15011
rect 8401 14977 8435 15011
rect 9413 14977 9447 15011
rect 9597 14977 9631 15011
rect 11805 14977 11839 15011
rect 11989 14977 12023 15011
rect 12541 14977 12575 15011
rect 12689 14977 12723 15011
rect 12909 14977 12943 15011
rect 13006 14977 13040 15011
rect 14013 14977 14047 15011
rect 14105 14977 14139 15011
rect 14289 14977 14323 15011
rect 14473 14977 14507 15011
rect 15577 14977 15611 15011
rect 15761 14977 15795 15011
rect 15945 14977 15979 15011
rect 17509 14977 17543 15011
rect 17877 14977 17911 15011
rect 20729 14977 20763 15011
rect 20913 14977 20947 15011
rect 21005 14977 21039 15011
rect 21097 14977 21131 15011
rect 22017 14977 22051 15011
rect 22109 14977 22143 15011
rect 22385 14977 22419 15011
rect 23969 14977 24003 15011
rect 25053 14977 25087 15011
rect 27813 14977 27847 15011
rect 28457 14977 28491 15011
rect 28641 14977 28675 15011
rect 29469 14977 29503 15011
rect 30297 14977 30331 15011
rect 30481 14977 30515 15011
rect 31217 14977 31251 15011
rect 31401 14977 31435 15011
rect 32137 14977 32171 15011
rect 32321 14977 32355 15011
rect 32432 14977 32466 15011
rect 32551 14977 32585 15011
rect 34897 14977 34931 15011
rect 37289 14977 37323 15011
rect 37473 14977 37507 15011
rect 37565 14977 37599 15011
rect 37703 14977 37737 15011
rect 39385 14977 39419 15011
rect 3893 14909 3927 14943
rect 5273 14909 5307 14943
rect 8585 14909 8619 14943
rect 14565 14909 14599 14943
rect 18889 14909 18923 14943
rect 24225 14909 24259 14943
rect 35173 14909 35207 14943
rect 39129 14909 39163 14943
rect 25881 14841 25915 14875
rect 5365 14773 5399 14807
rect 6929 14773 6963 14807
rect 13185 14773 13219 14807
rect 16129 14773 16163 14807
rect 17325 14773 17359 14807
rect 21281 14773 21315 14807
rect 25421 14773 25455 14807
rect 28825 14773 28859 14807
rect 30297 14773 30331 14807
rect 32781 14773 32815 14807
rect 2697 14569 2731 14603
rect 8401 14569 8435 14603
rect 23213 14569 23247 14603
rect 24409 14569 24443 14603
rect 28365 14569 28399 14603
rect 30205 14569 30239 14603
rect 30389 14569 30423 14603
rect 31217 14569 31251 14603
rect 33149 14569 33183 14603
rect 38393 14569 38427 14603
rect 11437 14501 11471 14535
rect 12265 14501 12299 14535
rect 19349 14501 19383 14535
rect 16313 14433 16347 14467
rect 16773 14433 16807 14467
rect 21833 14433 21867 14467
rect 30021 14433 30055 14467
rect 31677 14433 31711 14467
rect 35265 14433 35299 14467
rect 38853 14433 38887 14467
rect 2513 14365 2547 14399
rect 5641 14365 5675 14399
rect 5825 14365 5859 14399
rect 7205 14365 7239 14399
rect 7297 14365 7331 14399
rect 9873 14365 9907 14399
rect 10241 14365 10275 14399
rect 10885 14365 10919 14399
rect 11161 14365 11195 14399
rect 11253 14365 11287 14399
rect 12081 14365 12115 14399
rect 12725 14365 12759 14399
rect 14381 14365 14415 14399
rect 14529 14365 14563 14399
rect 14846 14365 14880 14399
rect 16037 14365 16071 14399
rect 17049 14365 17083 14399
rect 18705 14365 18739 14399
rect 19533 14365 19567 14399
rect 21005 14365 21039 14399
rect 21281 14365 21315 14399
rect 25145 14365 25179 14399
rect 25329 14365 25363 14399
rect 25421 14365 25455 14399
rect 25513 14365 25547 14399
rect 26249 14365 26283 14399
rect 30205 14365 30239 14399
rect 31033 14365 31067 14399
rect 32965 14365 32999 14399
rect 35541 14365 35575 14399
rect 37749 14365 37783 14399
rect 37933 14365 37967 14399
rect 38025 14365 38059 14399
rect 38117 14365 38151 14399
rect 68109 14365 68143 14399
rect 10057 14297 10091 14331
rect 10149 14297 10183 14331
rect 11069 14297 11103 14331
rect 14657 14297 14691 14331
rect 14749 14297 14783 14331
rect 20545 14297 20579 14331
rect 21189 14297 21223 14331
rect 25789 14297 25823 14331
rect 26494 14297 26528 14331
rect 28273 14297 28307 14331
rect 29929 14297 29963 14331
rect 30849 14297 30883 14331
rect 36921 14297 36955 14331
rect 37105 14297 37139 14331
rect 37289 14297 37323 14331
rect 2053 14229 2087 14263
rect 5733 14229 5767 14263
rect 6377 14229 6411 14263
rect 10425 14229 10459 14263
rect 12955 14229 12989 14263
rect 15025 14229 15059 14263
rect 21097 14229 21131 14263
rect 22385 14229 22419 14263
rect 27629 14229 27663 14263
rect 28917 14229 28951 14263
rect 4997 14025 5031 14059
rect 7757 14025 7791 14059
rect 9045 14025 9079 14059
rect 17693 14025 17727 14059
rect 19901 14025 19935 14059
rect 22385 14025 22419 14059
rect 24961 14025 24995 14059
rect 27445 14025 27479 14059
rect 29009 14025 29043 14059
rect 32137 14025 32171 14059
rect 36737 14025 36771 14059
rect 3157 13957 3191 13991
rect 3862 13957 3896 13991
rect 8769 13957 8803 13991
rect 17325 13957 17359 13991
rect 19441 13957 19475 13991
rect 26065 13957 26099 13991
rect 29285 13957 29319 13991
rect 33250 13957 33284 13991
rect 34529 13957 34563 13991
rect 1593 13889 1627 13923
rect 2513 13889 2547 13923
rect 2697 13889 2731 13923
rect 2789 13889 2823 13923
rect 2881 13889 2915 13923
rect 3617 13889 3651 13923
rect 6633 13889 6667 13923
rect 8493 13889 8527 13923
rect 8631 13889 8665 13923
rect 8861 13889 8895 13923
rect 10057 13889 10091 13923
rect 11805 13889 11839 13923
rect 13369 13889 13403 13923
rect 14105 13889 14139 13923
rect 15485 13889 15519 13923
rect 15669 13889 15703 13923
rect 17049 13889 17083 13923
rect 17197 13889 17231 13923
rect 17417 13889 17451 13923
rect 17514 13889 17548 13923
rect 18153 13889 18187 13923
rect 18337 13889 18371 13923
rect 19717 13889 19751 13923
rect 20361 13889 20395 13923
rect 23765 13889 23799 13923
rect 23949 13889 23983 13923
rect 25191 13889 25225 13923
rect 25326 13889 25360 13923
rect 25426 13889 25460 13923
rect 25605 13889 25639 13923
rect 27077 13889 27111 13923
rect 27261 13889 27295 13923
rect 27997 13889 28031 13923
rect 29193 13889 29227 13923
rect 29377 13889 29411 13923
rect 29561 13889 29595 13923
rect 34713 13889 34747 13923
rect 35357 13889 35391 13923
rect 35624 13889 35658 13923
rect 37657 13889 37691 13923
rect 37820 13892 37854 13926
rect 37936 13889 37970 13923
rect 38071 13889 38105 13923
rect 1501 13821 1535 13855
rect 6377 13821 6411 13855
rect 10333 13821 10367 13855
rect 11529 13821 11563 13855
rect 13645 13821 13679 13855
rect 15301 13821 15335 13855
rect 18521 13821 18555 13855
rect 19625 13821 19659 13855
rect 23121 13821 23155 13855
rect 33517 13821 33551 13855
rect 38301 13821 38335 13855
rect 1869 13685 1903 13719
rect 14289 13685 14323 13719
rect 19717 13685 19751 13719
rect 34897 13685 34931 13719
rect 2881 13481 2915 13515
rect 3801 13481 3835 13515
rect 6101 13481 6135 13515
rect 9505 13481 9539 13515
rect 14565 13481 14599 13515
rect 15301 13481 15335 13515
rect 19257 13481 19291 13515
rect 20453 13481 20487 13515
rect 21649 13481 21683 13515
rect 22753 13481 22787 13515
rect 28733 13481 28767 13515
rect 34069 13481 34103 13515
rect 35633 13481 35667 13515
rect 36553 13481 36587 13515
rect 37749 13481 37783 13515
rect 38209 13481 38243 13515
rect 17417 13413 17451 13447
rect 18337 13413 18371 13447
rect 26525 13413 26559 13447
rect 27629 13413 27663 13447
rect 31401 13413 31435 13447
rect 11713 13345 11747 13379
rect 12633 13345 12667 13379
rect 21741 13345 21775 13379
rect 2697 13277 2731 13311
rect 5457 13277 5491 13311
rect 5641 13277 5675 13311
rect 5733 13277 5767 13311
rect 5825 13277 5859 13311
rect 6561 13277 6595 13311
rect 8033 13277 8067 13311
rect 8217 13277 8251 13311
rect 8953 13277 8987 13311
rect 9321 13277 9355 13311
rect 11437 13277 11471 13311
rect 12909 13277 12943 13311
rect 15485 13277 15519 13311
rect 15577 13277 15611 13311
rect 15761 13277 15795 13311
rect 15853 13277 15887 13311
rect 16405 13277 16439 13311
rect 17601 13277 17635 13311
rect 18521 13277 18555 13311
rect 18705 13277 18739 13311
rect 19441 13277 19475 13311
rect 19625 13277 19659 13311
rect 20637 13277 20671 13311
rect 20729 13277 20763 13311
rect 21005 13277 21039 13311
rect 21649 13277 21683 13311
rect 22385 13277 22419 13311
rect 22569 13277 22603 13311
rect 23397 13277 23431 13311
rect 23581 13277 23615 13311
rect 23765 13277 23799 13311
rect 25421 13277 25455 13311
rect 27077 13277 27111 13311
rect 27261 13277 27295 13311
rect 27445 13277 27479 13311
rect 28089 13277 28123 13311
rect 28237 13277 28271 13311
rect 28365 13277 28399 13311
rect 28595 13277 28629 13311
rect 30021 13277 30055 13311
rect 30297 13277 30331 13311
rect 30389 13277 30423 13311
rect 31539 13277 31573 13311
rect 31677 13277 31711 13311
rect 31953 13277 31987 13311
rect 34989 13277 35023 13311
rect 35173 13277 35207 13311
rect 35268 13271 35302 13305
rect 35377 13277 35411 13311
rect 37381 13277 37415 13311
rect 39865 13277 39899 13311
rect 40121 13277 40155 13311
rect 2513 13209 2547 13243
rect 9137 13209 9171 13243
rect 9229 13209 9263 13243
rect 14657 13209 14691 13243
rect 16589 13209 16623 13243
rect 20821 13209 20855 13243
rect 21925 13209 21959 13243
rect 23489 13209 23523 13243
rect 25237 13209 25271 13243
rect 26341 13209 26375 13243
rect 27353 13209 27387 13243
rect 28457 13209 28491 13243
rect 30205 13209 30239 13243
rect 31769 13209 31803 13243
rect 37565 13209 37599 13243
rect 7849 13141 7883 13175
rect 21465 13141 21499 13175
rect 23213 13141 23247 13175
rect 24685 13141 24719 13175
rect 25605 13141 25639 13175
rect 30573 13141 30607 13175
rect 41245 13141 41279 13175
rect 10885 12937 10919 12971
rect 11713 12937 11747 12971
rect 15669 12937 15703 12971
rect 18429 12937 18463 12971
rect 18981 12937 19015 12971
rect 20545 12937 20579 12971
rect 21833 12937 21867 12971
rect 22001 12937 22035 12971
rect 36507 12937 36541 12971
rect 37933 12937 37967 12971
rect 41337 12937 41371 12971
rect 2513 12869 2547 12903
rect 7573 12869 7607 12903
rect 9965 12869 9999 12903
rect 11621 12869 11655 12903
rect 22201 12869 22235 12903
rect 23397 12869 23431 12903
rect 23489 12869 23523 12903
rect 26985 12869 27019 12903
rect 30941 12869 30975 12903
rect 31033 12869 31067 12903
rect 33701 12869 33735 12903
rect 1685 12801 1719 12835
rect 2329 12801 2363 12835
rect 3065 12801 3099 12835
rect 3321 12801 3355 12835
rect 7757 12801 7791 12835
rect 9689 12801 9723 12835
rect 9873 12801 9907 12835
rect 10057 12801 10091 12835
rect 10793 12801 10827 12835
rect 12541 12801 12575 12835
rect 13093 12801 13127 12835
rect 13360 12801 13394 12835
rect 15853 12801 15887 12835
rect 16129 12801 16163 12835
rect 17049 12801 17083 12835
rect 17305 12801 17339 12835
rect 20177 12801 20211 12835
rect 20361 12801 20395 12835
rect 23305 12801 23339 12835
rect 23673 12801 23707 12835
rect 24409 12801 24443 12835
rect 25697 12801 25731 12835
rect 25786 12807 25820 12841
rect 25881 12801 25915 12835
rect 26065 12801 26099 12835
rect 27261 12801 27295 12835
rect 27997 12801 28031 12835
rect 28273 12801 28307 12835
rect 29285 12801 29319 12835
rect 29561 12801 29595 12835
rect 30665 12801 30699 12835
rect 30758 12801 30792 12835
rect 31130 12801 31164 12835
rect 33333 12801 33367 12835
rect 33517 12801 33551 12835
rect 34161 12801 34195 12835
rect 34345 12801 34379 12835
rect 34437 12801 34471 12835
rect 34529 12801 34563 12835
rect 36737 12801 36771 12835
rect 37473 12801 37507 12835
rect 37749 12801 37783 12835
rect 40601 12801 40635 12835
rect 40785 12801 40819 12835
rect 41245 12801 41279 12835
rect 16037 12733 16071 12767
rect 24133 12733 24167 12767
rect 27077 12733 27111 12767
rect 37565 12733 37599 12767
rect 4445 12665 4479 12699
rect 10241 12665 10275 12699
rect 23121 12665 23155 12699
rect 67649 12665 67683 12699
rect 2145 12597 2179 12631
rect 7389 12597 7423 12631
rect 8309 12597 8343 12631
rect 12357 12597 12391 12631
rect 14473 12597 14507 12631
rect 15025 12597 15059 12631
rect 15945 12597 15979 12631
rect 22017 12597 22051 12631
rect 25421 12597 25455 12631
rect 26985 12597 27019 12631
rect 27445 12597 27479 12631
rect 31309 12597 31343 12631
rect 34805 12597 34839 12631
rect 37473 12597 37507 12631
rect 38393 12597 38427 12631
rect 40693 12597 40727 12631
rect 3157 12393 3191 12427
rect 3801 12393 3835 12427
rect 13277 12393 13311 12427
rect 16497 12393 16531 12427
rect 17785 12393 17819 12427
rect 20913 12393 20947 12427
rect 23765 12393 23799 12427
rect 26525 12393 26559 12427
rect 26985 12393 27019 12427
rect 36093 12393 36127 12427
rect 41245 12393 41279 12427
rect 2053 12325 2087 12359
rect 10425 12325 10459 12359
rect 25421 12325 25455 12359
rect 12357 12257 12391 12291
rect 23029 12257 23063 12291
rect 33057 12257 33091 12291
rect 33793 12257 33827 12291
rect 2513 12189 2547 12223
rect 2697 12189 2731 12223
rect 2789 12189 2823 12223
rect 2881 12189 2915 12223
rect 4353 12189 4387 12223
rect 6469 12189 6503 12223
rect 6561 12189 6595 12223
rect 6653 12189 6687 12223
rect 6837 12189 6871 12223
rect 7297 12189 7331 12223
rect 7481 12189 7515 12223
rect 7573 12189 7607 12223
rect 7665 12189 7699 12223
rect 9873 12189 9907 12223
rect 10057 12189 10091 12223
rect 10241 12189 10275 12223
rect 10885 12189 10919 12223
rect 11713 12189 11747 12223
rect 11897 12189 11931 12223
rect 11989 12189 12023 12223
rect 12081 12189 12115 12223
rect 13001 12189 13035 12223
rect 13093 12189 13127 12223
rect 14657 12189 14691 12223
rect 14933 12189 14967 12223
rect 15393 12189 15427 12223
rect 15485 12189 15519 12223
rect 15669 12189 15703 12223
rect 15761 12189 15795 12223
rect 16681 12189 16715 12223
rect 17601 12189 17635 12223
rect 17693 12189 17727 12223
rect 17877 12189 17911 12223
rect 20545 12189 20579 12223
rect 20729 12189 20763 12223
rect 24409 12189 24443 12223
rect 24593 12189 24627 12223
rect 25605 12189 25639 12223
rect 25697 12189 25731 12223
rect 25973 12189 26007 12223
rect 27721 12189 27755 12223
rect 27813 12189 27847 12223
rect 28089 12189 28123 12223
rect 29653 12189 29687 12223
rect 29929 12189 29963 12223
rect 30021 12189 30055 12223
rect 31309 12189 31343 12223
rect 31677 12189 31711 12223
rect 32321 12189 32355 12223
rect 32597 12189 32631 12223
rect 32781 12189 32815 12223
rect 33149 12189 33183 12223
rect 34713 12189 34747 12223
rect 36645 12189 36679 12223
rect 36829 12189 36863 12223
rect 36921 12189 36955 12223
rect 37013 12189 37047 12223
rect 37841 12189 37875 12223
rect 38025 12189 38059 12223
rect 38117 12189 38151 12223
rect 38209 12189 38243 12223
rect 39865 12189 39899 12223
rect 1869 12121 1903 12155
rect 4620 12121 4654 12155
rect 6193 12121 6227 12155
rect 10149 12121 10183 12155
rect 11069 12121 11103 12155
rect 11253 12121 11287 12155
rect 13277 12121 13311 12155
rect 22109 12121 22143 12155
rect 22845 12121 22879 12155
rect 25789 12121 25823 12155
rect 27905 12121 27939 12155
rect 28641 12121 28675 12155
rect 29837 12121 29871 12155
rect 31493 12121 31527 12155
rect 31585 12121 31619 12155
rect 32413 12121 32447 12155
rect 33977 12121 34011 12155
rect 34958 12121 34992 12155
rect 38485 12121 38519 12155
rect 40110 12121 40144 12155
rect 5733 12053 5767 12087
rect 7941 12053 7975 12087
rect 8953 12053 8987 12087
rect 12817 12053 12851 12087
rect 15945 12053 15979 12087
rect 17417 12053 17451 12087
rect 18337 12053 18371 12087
rect 22201 12053 22235 12087
rect 24409 12053 24443 12087
rect 27537 12053 27571 12087
rect 28733 12053 28767 12087
rect 30205 12053 30239 12087
rect 31861 12053 31895 12087
rect 37289 12053 37323 12087
rect 2237 11849 2271 11883
rect 2697 11849 2731 11883
rect 4169 11849 4203 11883
rect 6745 11849 6779 11883
rect 7205 11849 7239 11883
rect 9137 11849 9171 11883
rect 17877 11849 17911 11883
rect 18797 11849 18831 11883
rect 23305 11849 23339 11883
rect 29101 11849 29135 11883
rect 35265 11849 35299 11883
rect 1777 11781 1811 11815
rect 6561 11781 6595 11815
rect 11713 11781 11747 11815
rect 15025 11781 15059 11815
rect 23581 11781 23615 11815
rect 23673 11781 23707 11815
rect 24409 11781 24443 11815
rect 25145 11781 25179 11815
rect 30113 11781 30147 11815
rect 36461 11781 36495 11815
rect 2053 11713 2087 11747
rect 3065 11713 3099 11747
rect 5641 11713 5675 11747
rect 6377 11713 6411 11747
rect 8024 11713 8058 11747
rect 11529 11713 11563 11747
rect 12909 11713 12943 11747
rect 14197 11713 14231 11747
rect 15761 11713 15795 11747
rect 15945 11713 15979 11747
rect 17049 11713 17083 11747
rect 17233 11713 17267 11747
rect 17417 11713 17451 11747
rect 18705 11713 18739 11747
rect 19073 11713 19107 11747
rect 20361 11713 20395 11747
rect 20545 11713 20579 11747
rect 20637 11713 20671 11747
rect 20729 11713 20763 11747
rect 22201 11713 22235 11747
rect 22385 11713 22419 11747
rect 22569 11713 22603 11747
rect 22845 11713 22879 11747
rect 23489 11713 23523 11747
rect 23857 11713 23891 11747
rect 24593 11713 24627 11747
rect 26249 11713 26283 11747
rect 27353 11713 27387 11747
rect 27537 11713 27571 11747
rect 27629 11713 27663 11747
rect 27721 11713 27755 11747
rect 29883 11713 29917 11747
rect 30024 11713 30058 11747
rect 30241 11713 30275 11747
rect 30389 11713 30423 11747
rect 33425 11713 33459 11747
rect 33609 11713 33643 11747
rect 35081 11713 35115 11747
rect 35725 11713 35759 11747
rect 37289 11713 37323 11747
rect 37565 11713 37599 11747
rect 1961 11645 1995 11679
rect 2973 11645 3007 11679
rect 7757 11645 7791 11679
rect 16957 11645 16991 11679
rect 19165 11645 19199 11679
rect 22017 11645 22051 11679
rect 34529 11645 34563 11679
rect 17141 11577 17175 11611
rect 19441 11577 19475 11611
rect 25697 11577 25731 11611
rect 26433 11577 26467 11611
rect 33517 11577 33551 11611
rect 2053 11509 2087 11543
rect 2881 11509 2915 11543
rect 3525 11509 3559 11543
rect 5825 11509 5859 11543
rect 10977 11509 11011 11543
rect 11897 11509 11931 11543
rect 12449 11509 12483 11543
rect 15577 11509 15611 11543
rect 16681 11509 16715 11543
rect 18981 11509 19015 11543
rect 20913 11509 20947 11543
rect 27997 11509 28031 11543
rect 28457 11509 28491 11543
rect 29745 11509 29779 11543
rect 32873 11509 32907 11543
rect 67649 11509 67683 11543
rect 9229 11305 9263 11339
rect 12817 11305 12851 11339
rect 15025 11305 15059 11339
rect 15117 11305 15151 11339
rect 16589 11305 16623 11339
rect 18337 11305 18371 11339
rect 19717 11305 19751 11339
rect 21097 11305 21131 11339
rect 22385 11305 22419 11339
rect 23765 11305 23799 11339
rect 37105 11305 37139 11339
rect 5181 11237 5215 11271
rect 24409 11237 24443 11271
rect 29837 11237 29871 11271
rect 32873 11237 32907 11271
rect 6469 11169 6503 11203
rect 7481 11169 7515 11203
rect 15209 11169 15243 11203
rect 16681 11169 16715 11203
rect 18429 11169 18463 11203
rect 22017 11169 22051 11203
rect 23121 11169 23155 11203
rect 27629 11169 27663 11203
rect 28181 11169 28215 11203
rect 30573 11169 30607 11203
rect 35909 11169 35943 11203
rect 2237 11101 2271 11135
rect 3801 11101 3835 11135
rect 5825 11101 5859 11135
rect 10609 11101 10643 11135
rect 12173 11101 12207 11135
rect 12357 11101 12391 11135
rect 12449 11101 12483 11135
rect 12587 11101 12621 11135
rect 15301 11101 15335 11135
rect 15485 11101 15519 11135
rect 16773 11101 16807 11135
rect 17049 11101 17083 11135
rect 17969 11101 18003 11135
rect 18153 11101 18187 11135
rect 18245 11101 18279 11135
rect 19901 11101 19935 11135
rect 20085 11101 20119 11135
rect 20729 11101 20763 11135
rect 20913 11101 20947 11135
rect 22201 11101 22235 11135
rect 24593 11101 24627 11135
rect 24777 11101 24811 11135
rect 24961 11101 24995 11135
rect 25789 11101 25823 11135
rect 27353 11101 27387 11135
rect 30297 11101 30331 11135
rect 32229 11101 32263 11135
rect 32322 11101 32356 11135
rect 32505 11101 32539 11135
rect 32735 11101 32769 11135
rect 33333 11101 33367 11135
rect 33517 11101 33551 11135
rect 34161 11101 34195 11135
rect 34989 11101 35023 11135
rect 35081 11101 35115 11135
rect 35173 11101 35207 11135
rect 35357 11101 35391 11135
rect 38945 11101 38979 11135
rect 4068 11033 4102 11067
rect 6009 11033 6043 11067
rect 6653 11033 6687 11067
rect 6837 11033 6871 11067
rect 8309 11033 8343 11067
rect 10342 11033 10376 11067
rect 11345 11033 11379 11067
rect 11529 11033 11563 11067
rect 11713 11033 11747 11067
rect 13369 11033 13403 11067
rect 14749 11033 14783 11067
rect 16313 11033 16347 11067
rect 18705 11033 18739 11067
rect 22937 11033 22971 11067
rect 23673 11033 23707 11067
rect 24685 11033 24719 11067
rect 25973 11033 26007 11067
rect 26157 11033 26191 11067
rect 29009 11033 29043 11067
rect 32597 11033 32631 11067
rect 33425 11033 33459 11067
rect 36093 11033 36127 11067
rect 36277 11033 36311 11067
rect 36737 11033 36771 11067
rect 36921 11033 36955 11067
rect 38678 11033 38712 11067
rect 2697 10965 2731 10999
rect 5641 10965 5675 10999
rect 16957 10965 16991 10999
rect 34713 10965 34747 10999
rect 37565 10965 37599 10999
rect 1409 10761 1443 10795
rect 5181 10761 5215 10795
rect 8493 10761 8527 10795
rect 10241 10761 10275 10795
rect 14565 10761 14599 10795
rect 17233 10761 17267 10795
rect 22385 10761 22419 10795
rect 25329 10761 25363 10795
rect 27445 10761 27479 10795
rect 34069 10761 34103 10795
rect 40417 10761 40451 10795
rect 41337 10761 41371 10795
rect 12541 10693 12575 10727
rect 13430 10693 13464 10727
rect 24216 10693 24250 10727
rect 25789 10693 25823 10727
rect 27077 10693 27111 10727
rect 27261 10693 27295 10727
rect 29101 10693 29135 10727
rect 31125 10693 31159 10727
rect 32413 10693 32447 10727
rect 33701 10693 33735 10727
rect 33885 10693 33919 10727
rect 35734 10693 35768 10727
rect 1777 10625 1811 10659
rect 4721 10625 4755 10659
rect 5411 10625 5445 10659
rect 5549 10625 5583 10659
rect 5641 10625 5675 10659
rect 5825 10625 5859 10659
rect 6653 10625 6687 10659
rect 7113 10625 7147 10659
rect 7380 10625 7414 10659
rect 8953 10625 8987 10659
rect 9137 10625 9171 10659
rect 9597 10625 9631 10659
rect 9781 10625 9815 10659
rect 9873 10625 9907 10659
rect 9965 10625 9999 10659
rect 10793 10625 10827 10659
rect 11897 10625 11931 10659
rect 12081 10625 12115 10659
rect 12173 10625 12207 10659
rect 12265 10625 12299 10659
rect 13185 10625 13219 10659
rect 18429 10625 18463 10659
rect 22201 10625 22235 10659
rect 26065 10625 26099 10659
rect 26157 10625 26191 10659
rect 26249 10625 26283 10659
rect 26433 10625 26467 10659
rect 27905 10625 27939 10659
rect 29004 10625 29038 10659
rect 29193 10625 29227 10659
rect 29376 10625 29410 10659
rect 29469 10625 29503 10659
rect 30205 10625 30239 10659
rect 30389 10625 30423 10659
rect 30989 10625 31023 10659
rect 31217 10625 31251 10659
rect 31400 10625 31434 10659
rect 31493 10625 31527 10659
rect 32321 10625 32355 10659
rect 32505 10625 32539 10659
rect 32689 10625 32723 10659
rect 36001 10625 36035 10659
rect 36461 10625 36495 10659
rect 37749 10625 37783 10659
rect 38025 10625 38059 10659
rect 39037 10625 39071 10659
rect 39293 10625 39327 10659
rect 40877 10625 40911 10659
rect 41153 10625 41187 10659
rect 1869 10557 1903 10591
rect 18153 10557 18187 10591
rect 20453 10557 20487 10591
rect 20729 10557 20763 10591
rect 23949 10557 23983 10591
rect 40969 10557 41003 10591
rect 30849 10489 30883 10523
rect 32137 10489 32171 10523
rect 34621 10489 34655 10523
rect 2513 10421 2547 10455
rect 6469 10421 6503 10455
rect 9045 10421 9079 10455
rect 15209 10421 15243 10455
rect 23213 10421 23247 10455
rect 28089 10421 28123 10455
rect 28825 10421 28859 10455
rect 30297 10421 30331 10455
rect 33241 10421 33275 10455
rect 36645 10421 36679 10455
rect 40877 10421 40911 10455
rect 5181 10217 5215 10251
rect 7481 10217 7515 10251
rect 11897 10217 11931 10251
rect 12265 10217 12299 10251
rect 17141 10217 17175 10251
rect 21281 10217 21315 10251
rect 23489 10217 23523 10251
rect 25605 10217 25639 10251
rect 26341 10217 26375 10251
rect 29009 10217 29043 10251
rect 30113 10217 30147 10251
rect 33701 10217 33735 10251
rect 35633 10217 35667 10251
rect 37749 10217 37783 10251
rect 22753 10149 22787 10183
rect 36553 10149 36587 10183
rect 3801 10081 3835 10115
rect 11437 10081 11471 10115
rect 20085 10081 20119 10115
rect 20729 10081 20763 10115
rect 27353 10081 27387 10115
rect 32045 10081 32079 10115
rect 33333 10081 33367 10115
rect 5917 10013 5951 10047
rect 6009 10013 6043 10047
rect 6101 10013 6135 10047
rect 6285 10013 6319 10047
rect 6837 10013 6871 10047
rect 7711 10013 7745 10047
rect 7846 10013 7880 10047
rect 7941 10013 7975 10047
rect 8125 10013 8159 10047
rect 8953 10013 8987 10047
rect 9137 10013 9171 10047
rect 9965 10013 9999 10047
rect 10149 10013 10183 10047
rect 11161 10013 11195 10047
rect 12081 10013 12115 10047
rect 12265 10013 12299 10047
rect 14105 10013 14139 10047
rect 14197 10013 14231 10047
rect 14381 10013 14415 10047
rect 14473 10013 14507 10047
rect 16221 10013 16255 10047
rect 16313 10013 16347 10047
rect 16497 10013 16531 10047
rect 16589 10013 16623 10047
rect 18153 10013 18187 10047
rect 18429 10013 18463 10047
rect 19993 10013 20027 10047
rect 20269 10013 20303 10047
rect 20637 10013 20671 10047
rect 21465 10013 21499 10047
rect 21557 10013 21591 10047
rect 22385 10013 22419 10047
rect 22569 10013 22603 10047
rect 23305 10013 23339 10047
rect 26525 10013 26559 10047
rect 27169 10013 27203 10047
rect 27813 10013 27847 10047
rect 28457 10013 28491 10047
rect 28641 10013 28675 10047
rect 28825 10013 28859 10047
rect 29561 10013 29595 10047
rect 29745 10013 29779 10047
rect 29929 10013 29963 10047
rect 30665 10013 30699 10047
rect 31309 10013 31343 10047
rect 33517 10013 33551 10047
rect 34713 10013 34747 10047
rect 37105 10013 37139 10047
rect 37289 10013 37323 10047
rect 37381 10013 37415 10047
rect 37473 10013 37507 10047
rect 68109 10013 68143 10047
rect 4068 9945 4102 9979
rect 5641 9945 5675 9979
rect 9321 9945 9355 9979
rect 26985 9945 27019 9979
rect 28733 9945 28767 9979
rect 29837 9945 29871 9979
rect 31125 9945 31159 9979
rect 34897 9945 34931 9979
rect 7021 9877 7055 9911
rect 9781 9877 9815 9911
rect 14657 9877 14691 9911
rect 15209 9877 15243 9911
rect 16037 9877 16071 9911
rect 19993 9877 20027 9911
rect 25145 9877 25179 9911
rect 27997 9877 28031 9911
rect 31493 9877 31527 9911
rect 32275 9877 32309 9911
rect 35081 9877 35115 9911
rect 38209 9877 38243 9911
rect 40693 9877 40727 9911
rect 20545 9673 20579 9707
rect 25605 9673 25639 9707
rect 26433 9673 26467 9707
rect 4997 9605 5031 9639
rect 7757 9605 7791 9639
rect 9137 9605 9171 9639
rect 19349 9605 19383 9639
rect 22569 9605 22603 9639
rect 24492 9605 24526 9639
rect 36737 9605 36771 9639
rect 38301 9605 38335 9639
rect 39190 9605 39224 9639
rect 5457 9537 5491 9571
rect 5641 9537 5675 9571
rect 6929 9537 6963 9571
rect 9597 9537 9631 9571
rect 9781 9537 9815 9571
rect 9965 9537 9999 9571
rect 10609 9537 10643 9571
rect 10793 9537 10827 9571
rect 11529 9537 11563 9571
rect 11692 9537 11726 9571
rect 11792 9543 11826 9577
rect 11943 9537 11977 9571
rect 14289 9537 14323 9571
rect 14749 9537 14783 9571
rect 14933 9537 14967 9571
rect 15301 9537 15335 9571
rect 16865 9537 16899 9571
rect 16957 9537 16991 9571
rect 17141 9537 17175 9571
rect 17233 9537 17267 9571
rect 18521 9537 18555 9571
rect 18705 9537 18739 9571
rect 18797 9537 18831 9571
rect 19533 9537 19567 9571
rect 20729 9537 20763 9571
rect 20821 9537 20855 9571
rect 22201 9537 22235 9571
rect 22385 9537 22419 9571
rect 23397 9537 23431 9571
rect 23581 9537 23615 9571
rect 27629 9537 27663 9571
rect 27905 9537 27939 9571
rect 29101 9537 29135 9571
rect 29285 9537 29319 9571
rect 29377 9537 29411 9571
rect 29469 9537 29503 9571
rect 30757 9537 30791 9571
rect 33057 9537 33091 9571
rect 33885 9537 33919 9571
rect 34069 9537 34103 9571
rect 34161 9537 34195 9571
rect 34253 9537 34287 9571
rect 34989 9537 35023 9571
rect 35173 9537 35207 9571
rect 35265 9537 35299 9571
rect 35357 9537 35391 9571
rect 36369 9537 36403 9571
rect 36553 9537 36587 9571
rect 37657 9537 37691 9571
rect 37841 9537 37875 9571
rect 37936 9540 37970 9574
rect 38071 9537 38105 9571
rect 4445 9469 4479 9503
rect 7205 9469 7239 9503
rect 8401 9469 8435 9503
rect 10977 9469 11011 9503
rect 13461 9469 13495 9503
rect 15019 9469 15053 9503
rect 15117 9469 15151 9503
rect 19717 9469 19751 9503
rect 24225 9469 24259 9503
rect 28641 9469 28675 9503
rect 31033 9469 31067 9503
rect 33333 9469 33367 9503
rect 38945 9469 38979 9503
rect 16681 9401 16715 9435
rect 18245 9401 18279 9435
rect 5825 9333 5859 9367
rect 12173 9333 12207 9367
rect 15485 9333 15519 9367
rect 23765 9333 23799 9367
rect 29745 9333 29779 9367
rect 34529 9333 34563 9367
rect 35633 9333 35667 9367
rect 40325 9333 40359 9367
rect 1961 9129 1995 9163
rect 5181 9129 5215 9163
rect 10333 9129 10367 9163
rect 13277 9129 13311 9163
rect 17233 9129 17267 9163
rect 18061 9129 18095 9163
rect 20085 9129 20119 9163
rect 23305 9129 23339 9163
rect 27077 9129 27111 9163
rect 29561 9129 29595 9163
rect 17877 9061 17911 9095
rect 22661 9061 22695 9095
rect 36645 9061 36679 9095
rect 6745 8993 6779 9027
rect 9781 8993 9815 9027
rect 11897 8993 11931 9027
rect 15945 8993 15979 9027
rect 20453 8993 20487 9027
rect 30757 8993 30791 9027
rect 37841 8993 37875 9027
rect 2329 8925 2363 8959
rect 3801 8925 3835 8959
rect 6469 8925 6503 8959
rect 7757 8925 7791 8959
rect 7941 8925 7975 8959
rect 8033 8925 8067 8959
rect 8125 8925 8159 8959
rect 9505 8925 9539 8959
rect 10241 8925 10275 8959
rect 10425 8925 10459 8959
rect 12164 8925 12198 8959
rect 15678 8925 15712 8959
rect 19441 8925 19475 8959
rect 19625 8925 19659 8959
rect 20269 8925 20303 8959
rect 20545 8925 20579 8959
rect 22569 8925 22603 8959
rect 25697 8925 25731 8959
rect 27537 8925 27571 8959
rect 29745 8925 29779 8959
rect 29929 8925 29963 8959
rect 30481 8925 30515 8959
rect 31769 8925 31803 8959
rect 31953 8925 31987 8959
rect 32045 8925 32079 8959
rect 32137 8925 32171 8959
rect 33241 8925 33275 8959
rect 33333 8925 33367 8959
rect 33425 8925 33459 8959
rect 33609 8925 33643 8959
rect 37197 8925 37231 8959
rect 37381 8925 37415 8959
rect 37473 8925 37507 8959
rect 37565 8925 37599 8959
rect 38301 8925 38335 8959
rect 2145 8857 2179 8891
rect 4068 8857 4102 8891
rect 18052 8857 18086 8891
rect 18429 8857 18463 8891
rect 19257 8857 19291 8891
rect 21189 8857 21223 8891
rect 21925 8857 21959 8891
rect 24593 8857 24627 8891
rect 24777 8857 24811 8891
rect 25942 8857 25976 8891
rect 27804 8857 27838 8891
rect 35173 8857 35207 8891
rect 35909 8857 35943 8891
rect 38485 8857 38519 8891
rect 39129 8857 39163 8891
rect 2881 8789 2915 8823
rect 7297 8789 7331 8823
rect 8401 8789 8435 8823
rect 11161 8789 11195 8823
rect 14565 8789 14599 8823
rect 21833 8789 21867 8823
rect 23857 8789 23891 8823
rect 24409 8789 24443 8823
rect 28917 8789 28951 8823
rect 32413 8789 32447 8823
rect 32965 8789 32999 8823
rect 34069 8789 34103 8823
rect 38669 8789 38703 8823
rect 5181 8585 5215 8619
rect 8125 8585 8159 8619
rect 23397 8585 23431 8619
rect 31493 8585 31527 8619
rect 35081 8585 35115 8619
rect 36737 8585 36771 8619
rect 9014 8517 9048 8551
rect 14657 8517 14691 8551
rect 20085 8517 20119 8551
rect 22284 8517 22318 8551
rect 23857 8517 23891 8551
rect 28549 8517 28583 8551
rect 29929 8517 29963 8551
rect 33250 8517 33284 8551
rect 34713 8517 34747 8551
rect 36369 8517 36403 8551
rect 39098 8517 39132 8551
rect 1961 8449 1995 8483
rect 2053 8449 2087 8483
rect 2166 8449 2200 8483
rect 2329 8449 2363 8483
rect 2789 8449 2823 8483
rect 3045 8449 3079 8483
rect 5411 8449 5445 8483
rect 5549 8449 5583 8483
rect 5641 8449 5675 8483
rect 5825 8449 5859 8483
rect 7757 8449 7791 8483
rect 7941 8449 7975 8483
rect 14473 8449 14507 8483
rect 14749 8449 14783 8483
rect 16937 8449 16971 8483
rect 18797 8449 18831 8483
rect 18981 8449 19015 8483
rect 19073 8449 19107 8483
rect 19165 8449 19199 8483
rect 21005 8449 21039 8483
rect 22017 8449 22051 8483
rect 24133 8449 24167 8483
rect 24225 8449 24259 8483
rect 24317 8449 24351 8483
rect 24501 8449 24535 8483
rect 25145 8449 25179 8483
rect 25329 8449 25363 8483
rect 34161 8449 34195 8483
rect 34897 8449 34931 8483
rect 36553 8449 36587 8483
rect 37381 8449 37415 8483
rect 37560 8455 37594 8489
rect 37657 8449 37691 8483
rect 37795 8449 37829 8483
rect 7021 8381 7055 8415
rect 7297 8381 7331 8415
rect 8769 8381 8803 8415
rect 16681 8381 16715 8415
rect 19901 8381 19935 8415
rect 29285 8381 29319 8415
rect 33517 8381 33551 8415
rect 38853 8381 38887 8415
rect 4169 8313 4203 8347
rect 10149 8313 10183 8347
rect 15393 8313 15427 8347
rect 16129 8313 16163 8347
rect 18061 8313 18095 8347
rect 27813 8313 27847 8347
rect 40233 8313 40267 8347
rect 67649 8313 67683 8347
rect 1685 8245 1719 8279
rect 10701 8245 10735 8279
rect 14289 8245 14323 8279
rect 19441 8245 19475 8279
rect 21189 8245 21223 8279
rect 25513 8245 25547 8279
rect 32137 8245 32171 8279
rect 34069 8245 34103 8279
rect 38025 8245 38059 8279
rect 2789 8041 2823 8075
rect 16681 8041 16715 8075
rect 18705 8041 18739 8075
rect 25697 8041 25731 8075
rect 28641 8041 28675 8075
rect 31033 8041 31067 8075
rect 31677 8041 31711 8075
rect 34161 8041 34195 8075
rect 36001 8041 36035 8075
rect 39313 8041 39347 8075
rect 11161 7973 11195 8007
rect 2237 7905 2271 7939
rect 6837 7905 6871 7939
rect 21649 7905 21683 7939
rect 26157 7905 26191 7939
rect 28549 7905 28583 7939
rect 31585 7905 31619 7939
rect 1869 7837 1903 7871
rect 6561 7837 6595 7871
rect 12541 7837 12575 7871
rect 14565 7837 14599 7871
rect 14654 7837 14688 7871
rect 14749 7837 14783 7871
rect 14933 7837 14967 7871
rect 15577 7837 15611 7871
rect 16037 7837 16071 7871
rect 16221 7837 16255 7871
rect 16313 7837 16347 7871
rect 16451 7837 16485 7871
rect 17141 7837 17175 7871
rect 17417 7837 17451 7871
rect 18245 7837 18279 7871
rect 18521 7837 18555 7871
rect 19809 7837 19843 7871
rect 21925 7837 21959 7871
rect 25053 7837 25087 7871
rect 25237 7837 25271 7871
rect 25329 7837 25363 7871
rect 25421 7837 25455 7871
rect 28641 7837 28675 7871
rect 29653 7837 29687 7871
rect 29909 7837 29943 7871
rect 31769 7837 31803 7871
rect 32781 7837 32815 7871
rect 33048 7837 33082 7871
rect 37381 7837 37415 7871
rect 37933 7837 37967 7871
rect 38189 7837 38223 7871
rect 2053 7769 2087 7803
rect 5733 7769 5767 7803
rect 5917 7769 5951 7803
rect 8953 7769 8987 7803
rect 12274 7769 12308 7803
rect 17601 7769 17635 7803
rect 20054 7769 20088 7803
rect 23857 7769 23891 7803
rect 28365 7769 28399 7803
rect 31493 7769 31527 7803
rect 37114 7769 37148 7803
rect 5549 7701 5583 7735
rect 8309 7701 8343 7735
rect 13553 7701 13587 7735
rect 14289 7701 14323 7735
rect 17233 7701 17267 7735
rect 18337 7701 18371 7735
rect 21189 7701 21223 7735
rect 23213 7701 23247 7735
rect 24501 7701 24535 7735
rect 28825 7701 28859 7735
rect 31953 7701 31987 7735
rect 2421 7497 2455 7531
rect 5549 7497 5583 7531
rect 8677 7497 8711 7531
rect 9781 7497 9815 7531
rect 12265 7497 12299 7531
rect 19993 7497 20027 7531
rect 20453 7497 20487 7531
rect 29285 7497 29319 7531
rect 32873 7497 32907 7531
rect 34713 7497 34747 7531
rect 37381 7497 37415 7531
rect 12992 7429 13026 7463
rect 21281 7429 21315 7463
rect 26433 7429 26467 7463
rect 4169 7361 4203 7395
rect 4436 7361 4470 7395
rect 6469 7361 6503 7395
rect 6653 7361 6687 7395
rect 7297 7361 7331 7395
rect 7564 7361 7598 7395
rect 11529 7361 11563 7395
rect 11713 7361 11747 7395
rect 12081 7361 12115 7395
rect 19257 7361 19291 7395
rect 21097 7361 21131 7395
rect 22293 7361 22327 7395
rect 22385 7361 22419 7395
rect 22477 7361 22511 7395
rect 22661 7361 22695 7395
rect 24409 7361 24443 7395
rect 25789 7361 25823 7395
rect 25973 7361 26007 7395
rect 26065 7361 26099 7395
rect 26157 7361 26191 7395
rect 27241 7361 27275 7395
rect 28825 7361 28859 7395
rect 29101 7361 29135 7395
rect 29745 7361 29779 7395
rect 29837 7361 29871 7395
rect 35826 7361 35860 7395
rect 36093 7361 36127 7395
rect 11805 7293 11839 7327
rect 11897 7293 11931 7327
rect 12725 7293 12759 7327
rect 14749 7293 14783 7327
rect 15025 7293 15059 7327
rect 18981 7293 19015 7327
rect 23121 7293 23155 7327
rect 24685 7293 24719 7327
rect 26985 7293 27019 7327
rect 29009 7293 29043 7327
rect 9229 7225 9263 7259
rect 17693 7225 17727 7259
rect 3065 7157 3099 7191
rect 6837 7157 6871 7191
rect 10241 7157 10275 7191
rect 10977 7157 11011 7191
rect 14105 7157 14139 7191
rect 16037 7157 16071 7191
rect 17049 7157 17083 7191
rect 22017 7157 22051 7191
rect 23857 7157 23891 7191
rect 28365 7157 28399 7191
rect 29101 7157 29135 7191
rect 29745 7157 29779 7191
rect 30113 7157 30147 7191
rect 7573 6953 7607 6987
rect 11621 6953 11655 6987
rect 30205 6953 30239 6987
rect 31861 6953 31895 6987
rect 5549 6817 5583 6851
rect 9137 6817 9171 6851
rect 13553 6817 13587 6851
rect 19349 6817 19383 6851
rect 19993 6817 20027 6851
rect 22109 6817 22143 6851
rect 24501 6817 24535 6851
rect 26617 6817 26651 6851
rect 30389 6817 30423 6851
rect 1777 6749 1811 6783
rect 1961 6749 1995 6783
rect 2053 6749 2087 6783
rect 2191 6749 2225 6783
rect 2881 6749 2915 6783
rect 5825 6749 5859 6783
rect 5917 6749 5951 6783
rect 6009 6749 6043 6783
rect 6193 6749 6227 6783
rect 6929 6749 6963 6783
rect 7113 6749 7147 6783
rect 7205 6749 7239 6783
rect 7297 6749 7331 6783
rect 11069 6749 11103 6783
rect 11161 6749 11195 6783
rect 11345 6749 11379 6783
rect 11437 6749 11471 6783
rect 12265 6749 12299 6783
rect 12909 6749 12943 6783
rect 14381 6749 14415 6783
rect 14657 6749 14691 6783
rect 16129 6749 16163 6783
rect 16313 6749 16347 6783
rect 16405 6749 16439 6783
rect 16497 6749 16531 6783
rect 17325 6749 17359 6783
rect 17969 6749 18003 6783
rect 19257 6749 19291 6783
rect 19441 6749 19475 6783
rect 22365 6749 22399 6783
rect 24777 6749 24811 6783
rect 26249 6749 26283 6783
rect 30205 6749 30239 6783
rect 30481 6749 30515 6783
rect 32045 6749 32079 6783
rect 32137 6749 32171 6783
rect 34897 6749 34931 6783
rect 35173 6749 35207 6783
rect 35357 6749 35391 6783
rect 68109 6749 68143 6783
rect 2421 6681 2455 6715
rect 9382 6681 9416 6715
rect 20238 6681 20272 6715
rect 26433 6681 26467 6715
rect 31861 6681 31895 6715
rect 3801 6613 3835 6647
rect 8309 6613 8343 6647
rect 10517 6613 10551 6647
rect 12725 6613 12759 6647
rect 16773 6613 16807 6647
rect 18613 6613 18647 6647
rect 21373 6613 21407 6647
rect 23489 6613 23523 6647
rect 30665 6613 30699 6647
rect 32321 6613 32355 6647
rect 34713 6613 34747 6647
rect 2145 6409 2179 6443
rect 4077 6409 4111 6443
rect 6469 6409 6503 6443
rect 9229 6409 9263 6443
rect 19349 6409 19383 6443
rect 23121 6409 23155 6443
rect 25605 6409 25639 6443
rect 27629 6409 27663 6443
rect 30573 6409 30607 6443
rect 31585 6409 31619 6443
rect 32413 6409 32447 6443
rect 34529 6409 34563 6443
rect 1777 6341 1811 6375
rect 7757 6341 7791 6375
rect 7941 6341 7975 6375
rect 8125 6341 8159 6375
rect 10885 6341 10919 6375
rect 23305 6341 23339 6375
rect 24501 6341 24535 6375
rect 28089 6341 28123 6375
rect 29438 6341 29472 6375
rect 35265 6341 35299 6375
rect 1961 6273 1995 6307
rect 2697 6273 2731 6307
rect 2964 6273 2998 6307
rect 6653 6273 6687 6307
rect 8585 6273 8619 6307
rect 8769 6273 8803 6307
rect 8861 6273 8895 6307
rect 8953 6273 8987 6307
rect 11519 6263 11553 6297
rect 11621 6273 11655 6307
rect 11732 6273 11766 6307
rect 11894 6273 11928 6307
rect 12817 6273 12851 6307
rect 14197 6273 14231 6307
rect 14289 6273 14323 6307
rect 14381 6273 14415 6307
rect 14565 6273 14599 6307
rect 15255 6273 15289 6307
rect 15393 6273 15427 6307
rect 15485 6273 15519 6307
rect 15669 6273 15703 6307
rect 16773 6273 16807 6307
rect 17029 6273 17063 6307
rect 18705 6273 18739 6307
rect 18889 6273 18923 6307
rect 18981 6273 19015 6307
rect 19073 6273 19107 6307
rect 19809 6273 19843 6307
rect 21833 6273 21867 6307
rect 22109 6273 22143 6307
rect 23489 6273 23523 6307
rect 24777 6273 24811 6307
rect 25421 6273 25455 6307
rect 28365 6273 28399 6307
rect 28454 6273 28488 6307
rect 28554 6273 28588 6307
rect 28733 6273 28767 6307
rect 29193 6273 29227 6307
rect 31217 6273 31251 6307
rect 32597 6273 32631 6307
rect 32689 6273 32723 6307
rect 33793 6273 33827 6307
rect 38393 6273 38427 6307
rect 39221 6273 39255 6307
rect 9873 6205 9907 6239
rect 12541 6205 12575 6239
rect 24593 6205 24627 6239
rect 31125 6205 31159 6239
rect 33057 6205 33091 6239
rect 33517 6205 33551 6239
rect 34989 6205 35023 6239
rect 38117 6205 38151 6239
rect 5825 6069 5859 6103
rect 7297 6069 7331 6103
rect 10425 6069 10459 6103
rect 12081 6069 12115 6103
rect 13921 6069 13955 6103
rect 15025 6069 15059 6103
rect 18153 6069 18187 6103
rect 20453 6069 20487 6103
rect 21005 6069 21039 6103
rect 24777 6069 24811 6103
rect 24961 6069 24995 6103
rect 36737 6069 36771 6103
rect 3249 5865 3283 5899
rect 9045 5865 9079 5899
rect 9689 5865 9723 5899
rect 16129 5865 16163 5899
rect 19717 5865 19751 5899
rect 28457 5865 28491 5899
rect 31953 5865 31987 5899
rect 32597 5865 32631 5899
rect 36277 5865 36311 5899
rect 37749 5865 37783 5899
rect 24685 5797 24719 5831
rect 27629 5797 27663 5831
rect 1869 5729 1903 5763
rect 6745 5729 6779 5763
rect 14841 5729 14875 5763
rect 20821 5729 20855 5763
rect 26249 5729 26283 5763
rect 31861 5729 31895 5763
rect 33057 5729 33091 5763
rect 4905 5661 4939 5695
rect 5641 5661 5675 5695
rect 5733 5661 5767 5695
rect 5825 5661 5859 5695
rect 6009 5661 6043 5695
rect 6469 5661 6503 5695
rect 8033 5661 8067 5695
rect 8125 5661 8159 5695
rect 8217 5661 8251 5695
rect 8401 5661 8435 5695
rect 10425 5661 10459 5695
rect 11161 5661 11195 5695
rect 11805 5661 11839 5695
rect 11897 5661 11931 5695
rect 12081 5661 12115 5695
rect 12173 5661 12207 5695
rect 12817 5661 12851 5695
rect 13093 5661 13127 5695
rect 14565 5661 14599 5695
rect 16313 5661 16347 5695
rect 16589 5661 16623 5695
rect 17325 5661 17359 5695
rect 17785 5661 17819 5695
rect 18429 5661 18463 5695
rect 19257 5661 19291 5695
rect 19349 5661 19383 5695
rect 19533 5661 19567 5695
rect 20177 5661 20211 5695
rect 20453 5661 20487 5695
rect 20637 5661 20671 5695
rect 24501 5661 24535 5695
rect 25421 5661 25455 5695
rect 25605 5661 25639 5695
rect 28089 5661 28123 5695
rect 28273 5661 28307 5695
rect 31677 5661 31711 5695
rect 31953 5661 31987 5695
rect 32781 5661 32815 5695
rect 32873 5661 32907 5695
rect 33149 5661 33183 5695
rect 33885 5661 33919 5695
rect 33977 5661 34011 5695
rect 36277 5661 36311 5695
rect 36461 5661 36495 5695
rect 37565 5661 37599 5695
rect 68109 5661 68143 5695
rect 2114 5593 2148 5627
rect 16497 5593 16531 5627
rect 26516 5593 26550 5627
rect 5365 5525 5399 5559
rect 7757 5525 7791 5559
rect 10241 5525 10275 5559
rect 10977 5525 11011 5559
rect 11621 5525 11655 5559
rect 12909 5525 12943 5559
rect 21281 5525 21315 5559
rect 25789 5525 25823 5559
rect 32137 5525 32171 5559
rect 34161 5525 34195 5559
rect 1869 5321 1903 5355
rect 3525 5321 3559 5355
rect 6377 5321 6411 5355
rect 7665 5321 7699 5355
rect 14197 5321 14231 5355
rect 14565 5321 14599 5355
rect 15209 5321 15243 5355
rect 15577 5321 15611 5355
rect 17509 5321 17543 5355
rect 19809 5321 19843 5355
rect 20821 5321 20855 5355
rect 22201 5321 22235 5355
rect 24041 5321 24075 5355
rect 26433 5321 26467 5355
rect 31033 5321 31067 5355
rect 34897 5321 34931 5355
rect 36185 5321 36219 5355
rect 4344 5253 4378 5287
rect 6745 5253 6779 5287
rect 7297 5253 7331 5287
rect 8401 5253 8435 5287
rect 16773 5253 16807 5287
rect 19073 5253 19107 5287
rect 24777 5253 24811 5287
rect 28549 5253 28583 5287
rect 28733 5253 28767 5287
rect 2145 5185 2179 5219
rect 2237 5185 2271 5219
rect 2329 5185 2363 5219
rect 2513 5185 2547 5219
rect 4077 5185 4111 5219
rect 6561 5185 6595 5219
rect 7481 5185 7515 5219
rect 8309 5185 8343 5219
rect 8493 5185 8527 5219
rect 8953 5185 8987 5219
rect 9137 5185 9171 5219
rect 9864 5185 9898 5219
rect 11529 5185 11563 5219
rect 11713 5185 11747 5219
rect 11989 5185 12023 5219
rect 12081 5185 12115 5219
rect 12265 5185 12299 5219
rect 13185 5185 13219 5219
rect 13277 5185 13311 5219
rect 13461 5185 13495 5219
rect 14381 5185 14415 5219
rect 14657 5185 14691 5219
rect 15117 5185 15151 5219
rect 15393 5185 15427 5219
rect 17233 5185 17267 5219
rect 20269 5185 20303 5219
rect 20545 5185 20579 5219
rect 20821 5185 20855 5219
rect 22661 5185 22695 5219
rect 22928 5185 22962 5219
rect 24593 5185 24627 5219
rect 25789 5185 25823 5219
rect 25973 5185 26007 5219
rect 26065 5185 26099 5219
rect 26157 5185 26191 5219
rect 26985 5185 27019 5219
rect 30665 5185 30699 5219
rect 33241 5185 33275 5219
rect 33517 5185 33551 5219
rect 34713 5185 34747 5219
rect 36177 5185 36211 5219
rect 36369 5185 36403 5219
rect 9597 5117 9631 5151
rect 11897 5117 11931 5151
rect 13369 5117 13403 5151
rect 17325 5117 17359 5151
rect 19533 5117 19567 5151
rect 19625 5117 19659 5151
rect 29377 5117 29411 5151
rect 30573 5117 30607 5151
rect 59461 5117 59495 5151
rect 5457 5049 5491 5083
rect 10977 5049 11011 5083
rect 13001 5049 13035 5083
rect 16773 5049 16807 5083
rect 19073 5049 19107 5083
rect 21281 5049 21315 5083
rect 60105 5049 60139 5083
rect 3065 4981 3099 5015
rect 9137 4981 9171 5015
rect 16037 4981 16071 5015
rect 18521 4981 18555 5015
rect 24961 4981 24995 5015
rect 28917 4981 28951 5015
rect 34253 4981 34287 5015
rect 58817 4981 58851 5015
rect 2145 4777 2179 4811
rect 3893 4777 3927 4811
rect 8401 4777 8435 4811
rect 10517 4777 10551 4811
rect 14105 4777 14139 4811
rect 22937 4777 22971 4811
rect 23857 4777 23891 4811
rect 31769 4777 31803 4811
rect 36369 4777 36403 4811
rect 9137 4709 9171 4743
rect 16589 4709 16623 4743
rect 18245 4709 18279 4743
rect 21189 4709 21223 4743
rect 37013 4709 37047 4743
rect 57897 4709 57931 4743
rect 59185 4709 59219 4743
rect 12081 4641 12115 4675
rect 12173 4641 12207 4675
rect 15485 4641 15519 4675
rect 20545 4641 20579 4675
rect 26801 4641 26835 4675
rect 60473 4641 60507 4675
rect 1777 4573 1811 4607
rect 1961 4573 1995 4607
rect 2973 4573 3007 4607
rect 6009 4573 6043 4607
rect 7021 4573 7055 4607
rect 7288 4573 7322 4607
rect 8953 4573 8987 4607
rect 9597 4573 9631 4607
rect 10333 4573 10367 4607
rect 11069 4573 11103 4607
rect 11805 4573 11839 4607
rect 11989 4573 12023 4607
rect 12357 4573 12391 4607
rect 17325 4573 17359 4607
rect 17693 4573 17727 4607
rect 17877 4573 17911 4607
rect 18613 4573 18647 4607
rect 19349 4573 19383 4607
rect 19533 4573 19567 4607
rect 19809 4573 19843 4607
rect 19993 4573 20027 4607
rect 22293 4573 22327 4607
rect 22456 4573 22490 4607
rect 22556 4573 22590 4607
rect 22707 4573 22741 4607
rect 24685 4573 24719 4607
rect 24777 4573 24811 4607
rect 24869 4573 24903 4607
rect 25053 4573 25087 4607
rect 25697 4573 25731 4607
rect 25881 4573 25915 4607
rect 25973 4573 26007 4607
rect 26065 4573 26099 4607
rect 27813 4573 27847 4607
rect 28641 4573 28675 4607
rect 28730 4573 28764 4607
rect 28825 4573 28859 4607
rect 29009 4573 29043 4607
rect 29561 4573 29595 4607
rect 29745 4573 29779 4607
rect 29837 4573 29871 4607
rect 29929 4573 29963 4607
rect 33149 4573 33183 4607
rect 36277 4573 36311 4607
rect 36921 4573 36955 4607
rect 57253 4573 57287 4607
rect 58541 4573 58575 4607
rect 2789 4505 2823 4539
rect 4905 4505 4939 4539
rect 10425 4505 10459 4539
rect 10609 4505 10643 4539
rect 13369 4505 13403 4539
rect 15218 4505 15252 4539
rect 26341 4505 26375 4539
rect 28365 4505 28399 4539
rect 32882 4505 32916 4539
rect 2605 4437 2639 4471
rect 5457 4437 5491 4471
rect 6561 4437 6595 4471
rect 9781 4437 9815 4471
rect 11253 4437 11287 4471
rect 12541 4437 12575 4471
rect 13461 4437 13495 4471
rect 19993 4437 20027 4471
rect 24409 4437 24443 4471
rect 30205 4437 30239 4471
rect 12081 4233 12115 4267
rect 17233 4233 17267 4267
rect 22201 4233 22235 4267
rect 24777 4233 24811 4267
rect 25789 4233 25823 4267
rect 29193 4233 29227 4267
rect 31401 4233 31435 4267
rect 33701 4233 33735 4267
rect 36001 4233 36035 4267
rect 5641 4165 5675 4199
rect 5825 4165 5859 4199
rect 8953 4165 8987 4199
rect 13194 4165 13228 4199
rect 22385 4165 22419 4199
rect 22569 4165 22603 4199
rect 23664 4165 23698 4199
rect 26157 4165 26191 4199
rect 28825 4165 28859 4199
rect 29009 4165 29043 4199
rect 2145 4097 2179 4131
rect 2237 4097 2271 4131
rect 2329 4097 2363 4131
rect 2513 4097 2547 4131
rect 2973 4097 3007 4131
rect 3229 4097 3263 4131
rect 4997 4097 5031 4131
rect 6653 4097 6687 4131
rect 6745 4097 6779 4131
rect 6837 4097 6871 4131
rect 7021 4097 7055 4131
rect 7481 4097 7515 4131
rect 8401 4097 8435 4131
rect 9689 4097 9723 4131
rect 10333 4097 10367 4131
rect 10517 4097 10551 4131
rect 10793 4097 10827 4131
rect 10977 4097 11011 4131
rect 11621 4097 11655 4131
rect 13461 4097 13495 4131
rect 13921 4097 13955 4131
rect 14933 4097 14967 4131
rect 15393 4097 15427 4131
rect 16865 4097 16899 4131
rect 16957 4097 16991 4131
rect 17233 4097 17267 4131
rect 18337 4097 18371 4131
rect 18981 4097 19015 4131
rect 19625 4097 19659 4131
rect 20269 4097 20303 4131
rect 20545 4097 20579 4131
rect 20913 4097 20947 4131
rect 21281 4097 21315 4131
rect 23397 4097 23431 4131
rect 25973 4097 26007 4131
rect 26985 4097 27019 4131
rect 27252 4097 27286 4131
rect 30288 4097 30322 4131
rect 34253 4097 34287 4131
rect 59829 4097 59863 4131
rect 1869 4029 1903 4063
rect 5457 4029 5491 4063
rect 9137 4029 9171 4063
rect 21005 4029 21039 4063
rect 30021 4029 30055 4063
rect 34529 4029 34563 4063
rect 61117 4029 61151 4063
rect 7665 3961 7699 3995
rect 9873 3961 9907 3995
rect 14749 3961 14783 3995
rect 15577 3961 15611 3995
rect 17693 3961 17727 3995
rect 58541 3961 58575 3995
rect 60473 3961 60507 3995
rect 4353 3893 4387 3927
rect 6377 3893 6411 3927
rect 8217 3893 8251 3927
rect 14105 3893 14139 3927
rect 18521 3893 18555 3927
rect 19165 3893 19199 3927
rect 19809 3893 19843 3927
rect 28365 3893 28399 3927
rect 56241 3893 56275 3927
rect 56885 3893 56919 3927
rect 57897 3893 57931 3927
rect 59185 3893 59219 3927
rect 67649 3893 67683 3927
rect 2237 3689 2271 3723
rect 2789 3689 2823 3723
rect 4721 3689 4755 3723
rect 11621 3689 11655 3723
rect 15853 3689 15887 3723
rect 7205 3621 7239 3655
rect 10977 3621 11011 3655
rect 11805 3621 11839 3655
rect 15117 3621 15151 3655
rect 19993 3621 20027 3655
rect 41797 3621 41831 3655
rect 57897 3621 57931 3655
rect 61117 3621 61151 3655
rect 12817 3553 12851 3587
rect 19441 3553 19475 3587
rect 19533 3553 19567 3587
rect 56609 3553 56643 3587
rect 58541 3553 58575 3587
rect 61761 3553 61795 3587
rect 6294 3485 6328 3519
rect 6561 3485 6595 3519
rect 7021 3485 7055 3519
rect 7849 3485 7883 3519
rect 8033 3485 8067 3519
rect 9137 3485 9171 3519
rect 9597 3485 9631 3519
rect 9864 3485 9898 3519
rect 13553 3485 13587 3519
rect 14565 3485 14599 3519
rect 15301 3485 15335 3519
rect 16313 3485 16347 3519
rect 16497 3485 16531 3519
rect 16681 3485 16715 3519
rect 16865 3485 16899 3519
rect 17141 3485 17175 3519
rect 18061 3485 18095 3519
rect 18705 3485 18739 3519
rect 20545 3485 20579 3519
rect 21649 3485 21683 3519
rect 22477 3485 22511 3519
rect 23581 3485 23615 3519
rect 24409 3485 24443 3519
rect 25237 3485 25271 3519
rect 26065 3485 26099 3519
rect 26893 3485 26927 3519
rect 27721 3485 27755 3519
rect 28825 3485 28859 3519
rect 29929 3485 29963 3519
rect 30757 3485 30791 3519
rect 31585 3485 31619 3519
rect 32413 3485 32447 3519
rect 33241 3485 33275 3519
rect 39865 3485 39899 3519
rect 40509 3485 40543 3519
rect 41153 3485 41187 3519
rect 42625 3485 42659 3519
rect 43269 3485 43303 3519
rect 45109 3485 45143 3519
rect 45753 3485 45787 3519
rect 46397 3485 46431 3519
rect 47041 3485 47075 3519
rect 47869 3485 47903 3519
rect 48973 3485 49007 3519
rect 50353 3485 50387 3519
rect 50997 3485 51031 3519
rect 51641 3485 51675 3519
rect 52837 3485 52871 3519
rect 53481 3485 53515 3519
rect 55321 3485 55355 3519
rect 55965 3485 55999 3519
rect 57253 3485 57287 3519
rect 59185 3485 59219 3519
rect 60473 3485 60507 3519
rect 11437 3417 11471 3451
rect 12633 3417 12667 3451
rect 19993 3417 20027 3451
rect 4169 3349 4203 3383
rect 5181 3349 5215 3383
rect 7665 3349 7699 3383
rect 11647 3349 11681 3383
rect 13369 3349 13403 3383
rect 14381 3349 14415 3383
rect 19257 3349 19291 3383
rect 8493 3145 8527 3179
rect 10425 3145 10459 3179
rect 14933 3145 14967 3179
rect 15577 3145 15611 3179
rect 16865 3145 16899 3179
rect 19349 3145 19383 3179
rect 21833 3145 21867 3179
rect 13820 3077 13854 3111
rect 5549 3009 5583 3043
rect 6653 3009 6687 3043
rect 7113 3009 7147 3043
rect 7380 3009 7414 3043
rect 9045 3009 9079 3043
rect 9301 3009 9335 3043
rect 11805 3009 11839 3043
rect 12265 3009 12299 3043
rect 13553 3009 13587 3043
rect 15393 3009 15427 3043
rect 16681 3009 16715 3043
rect 17693 3009 17727 3043
rect 19165 3009 19199 3043
rect 61117 3009 61151 3043
rect 3433 2941 3467 2975
rect 5089 2941 5123 2975
rect 12541 2941 12575 2975
rect 18705 2941 18739 2975
rect 21281 2941 21315 2975
rect 37933 2941 37967 2975
rect 45661 2941 45695 2975
rect 49525 2941 49559 2975
rect 53389 2941 53423 2975
rect 61761 2941 61795 2975
rect 4537 2873 4571 2907
rect 5733 2873 5767 2907
rect 6469 2873 6503 2907
rect 10977 2873 11011 2907
rect 39221 2873 39255 2907
rect 40509 2873 40543 2907
rect 43085 2873 43119 2907
rect 44373 2873 44407 2907
rect 48237 2873 48271 2907
rect 50169 2873 50203 2907
rect 51457 2873 51491 2907
rect 54033 2873 54067 2907
rect 55321 2873 55355 2907
rect 56609 2873 56643 2907
rect 58541 2873 58575 2907
rect 63049 2873 63083 2907
rect 3985 2805 4019 2839
rect 11621 2805 11655 2839
rect 17509 2805 17543 2839
rect 19993 2805 20027 2839
rect 20637 2805 20671 2839
rect 22569 2805 22603 2839
rect 23029 2805 23063 2839
rect 23857 2805 23891 2839
rect 24501 2805 24535 2839
rect 25145 2805 25179 2839
rect 25789 2805 25823 2839
rect 26433 2805 26467 2839
rect 27721 2805 27755 2839
rect 28365 2805 28399 2839
rect 29009 2805 29043 2839
rect 29653 2805 29687 2839
rect 30297 2805 30331 2839
rect 30941 2805 30975 2839
rect 31585 2805 31619 2839
rect 32873 2805 32907 2839
rect 33517 2805 33551 2839
rect 34161 2805 34195 2839
rect 34621 2805 34655 2839
rect 35449 2805 35483 2839
rect 36277 2805 36311 2839
rect 37289 2805 37323 2839
rect 38577 2805 38611 2839
rect 39865 2805 39899 2839
rect 41153 2805 41187 2839
rect 42441 2805 42475 2839
rect 43729 2805 43763 2839
rect 45017 2805 45051 2839
rect 46305 2805 46339 2839
rect 47593 2805 47627 2839
rect 48881 2805 48915 2839
rect 50813 2805 50847 2839
rect 52745 2805 52779 2839
rect 54677 2805 54711 2839
rect 55965 2805 55999 2839
rect 57897 2805 57931 2839
rect 59185 2805 59219 2839
rect 59829 2805 59863 2839
rect 60473 2805 60507 2839
rect 7849 2601 7883 2635
rect 12081 2601 12115 2635
rect 12265 2601 12299 2635
rect 16865 2601 16899 2635
rect 17601 2601 17635 2635
rect 18245 2601 18279 2635
rect 21833 2601 21867 2635
rect 55321 2601 55355 2635
rect 61117 2601 61151 2635
rect 9321 2533 9355 2567
rect 20637 2533 20671 2567
rect 22569 2533 22603 2567
rect 28365 2533 28399 2567
rect 30297 2533 30331 2567
rect 42441 2533 42475 2567
rect 46305 2533 46339 2567
rect 50169 2533 50203 2567
rect 54033 2533 54067 2567
rect 57897 2533 57931 2567
rect 58541 2533 58575 2567
rect 60473 2533 60507 2567
rect 3893 2465 3927 2499
rect 8401 2465 8435 2499
rect 25789 2465 25823 2499
rect 37933 2465 37967 2499
rect 39865 2465 39899 2499
rect 43085 2465 43119 2499
rect 45017 2465 45051 2499
rect 48237 2465 48271 2499
rect 50813 2465 50847 2499
rect 52745 2465 52779 2499
rect 56609 2465 56643 2499
rect 63693 2465 63727 2499
rect 4905 2397 4939 2431
rect 6561 2397 6595 2431
rect 7205 2397 7239 2431
rect 7389 2397 7423 2431
rect 7481 2397 7515 2431
rect 7573 2397 7607 2431
rect 9505 2397 9539 2431
rect 10241 2397 10275 2431
rect 10977 2397 11011 2431
rect 12725 2397 12759 2431
rect 13001 2397 13035 2431
rect 14381 2397 14415 2431
rect 14841 2397 14875 2431
rect 15853 2397 15887 2431
rect 16681 2397 16715 2431
rect 18429 2397 18463 2431
rect 19993 2397 20027 2431
rect 21281 2397 21315 2431
rect 23213 2397 23247 2431
rect 23857 2397 23891 2431
rect 25145 2397 25179 2431
rect 26433 2397 26467 2431
rect 27721 2397 27755 2431
rect 29009 2397 29043 2431
rect 30941 2397 30975 2431
rect 31585 2397 31619 2431
rect 32873 2397 32907 2431
rect 33517 2397 33551 2431
rect 34161 2397 34195 2431
rect 34897 2397 34931 2431
rect 35541 2397 35575 2431
rect 36001 2397 36035 2431
rect 37289 2397 37323 2431
rect 38577 2397 38611 2431
rect 40509 2397 40543 2431
rect 41153 2397 41187 2431
rect 43729 2397 43763 2431
rect 45661 2397 45695 2431
rect 47593 2397 47627 2431
rect 48881 2397 48915 2431
rect 51457 2397 51491 2431
rect 53389 2397 53423 2431
rect 55965 2397 55999 2431
rect 59185 2397 59219 2431
rect 61761 2397 61795 2431
rect 63049 2397 63083 2431
rect 67649 2397 67683 2431
rect 12127 2363 12161 2397
rect 3249 2329 3283 2363
rect 5641 2329 5675 2363
rect 6745 2329 6779 2363
rect 11897 2329 11931 2363
rect 17509 2329 17543 2363
rect 24409 2329 24443 2363
rect 4445 2261 4479 2295
rect 5089 2261 5123 2295
rect 5733 2261 5767 2295
rect 10057 2261 10091 2295
rect 10793 2261 10827 2295
rect 14197 2261 14231 2295
rect 15025 2261 15059 2295
rect 15669 2261 15703 2295
rect 19349 2261 19383 2295
<< metal1 >>
rect 1104 57690 68816 57712
rect 1104 57638 19574 57690
rect 19626 57638 19638 57690
rect 19690 57638 19702 57690
rect 19754 57638 19766 57690
rect 19818 57638 19830 57690
rect 19882 57638 50294 57690
rect 50346 57638 50358 57690
rect 50410 57638 50422 57690
rect 50474 57638 50486 57690
rect 50538 57638 50550 57690
rect 50602 57638 68816 57690
rect 1104 57616 68816 57638
rect 22094 57576 22100 57588
rect 22055 57548 22100 57576
rect 22094 57536 22100 57548
rect 22152 57536 22158 57588
rect 30558 57536 30564 57588
rect 30616 57576 30622 57588
rect 30837 57579 30895 57585
rect 30837 57576 30849 57579
rect 30616 57548 30849 57576
rect 30616 57536 30622 57548
rect 30837 57545 30849 57548
rect 30883 57545 30895 57579
rect 30837 57539 30895 57545
rect 39298 57536 39304 57588
rect 39356 57576 39362 57588
rect 40037 57579 40095 57585
rect 40037 57576 40049 57579
rect 39356 57548 40049 57576
rect 39356 57536 39362 57548
rect 40037 57545 40049 57548
rect 40083 57545 40095 57579
rect 48314 57576 48320 57588
rect 48275 57548 48320 57576
rect 40037 57539 40095 57545
rect 48314 57536 48320 57548
rect 48372 57536 48378 57588
rect 56778 57536 56784 57588
rect 56836 57576 56842 57588
rect 57057 57579 57115 57585
rect 57057 57576 57069 57579
rect 56836 57548 57069 57576
rect 56836 57536 56842 57548
rect 57057 57545 57069 57548
rect 57103 57545 57115 57579
rect 57057 57539 57115 57545
rect 65518 57536 65524 57588
rect 65576 57576 65582 57588
rect 65797 57579 65855 57585
rect 65797 57576 65809 57579
rect 65576 57548 65809 57576
rect 65576 57536 65582 57548
rect 65797 57545 65809 57548
rect 65843 57545 65855 57579
rect 65797 57539 65855 57545
rect 36814 57468 36820 57520
rect 36872 57508 36878 57520
rect 47581 57511 47639 57517
rect 47581 57508 47593 57511
rect 36872 57480 47593 57508
rect 36872 57468 36878 57480
rect 47581 57477 47593 57480
rect 47627 57508 47639 57511
rect 47627 57480 48176 57508
rect 47627 57477 47639 57480
rect 47581 57471 47639 57477
rect 4338 57400 4344 57452
rect 4396 57440 4402 57452
rect 4433 57443 4491 57449
rect 4433 57440 4445 57443
rect 4396 57412 4445 57440
rect 4396 57400 4402 57412
rect 4433 57409 4445 57412
rect 4479 57409 4491 57443
rect 4433 57403 4491 57409
rect 13078 57400 13084 57452
rect 13136 57440 13142 57452
rect 13173 57443 13231 57449
rect 13173 57440 13185 57443
rect 13136 57412 13185 57440
rect 13136 57400 13142 57412
rect 13173 57409 13185 57412
rect 13219 57409 13231 57443
rect 13173 57403 13231 57409
rect 21634 57400 21640 57452
rect 21692 57440 21698 57452
rect 21913 57443 21971 57449
rect 21913 57440 21925 57443
rect 21692 57412 21925 57440
rect 21692 57400 21698 57412
rect 21913 57409 21925 57412
rect 21959 57409 21971 57443
rect 21913 57403 21971 57409
rect 30098 57400 30104 57452
rect 30156 57440 30162 57452
rect 48148 57449 48176 57480
rect 30653 57443 30711 57449
rect 30653 57440 30665 57443
rect 30156 57412 30665 57440
rect 30156 57400 30162 57412
rect 30653 57409 30665 57412
rect 30699 57409 30711 57443
rect 39853 57443 39911 57449
rect 39853 57440 39865 57443
rect 30653 57403 30711 57409
rect 39224 57412 39865 57440
rect 39224 57248 39252 57412
rect 39853 57409 39865 57412
rect 39899 57409 39911 57443
rect 39853 57403 39911 57409
rect 48133 57443 48191 57449
rect 48133 57409 48145 57443
rect 48179 57409 48191 57443
rect 48133 57403 48191 57409
rect 56318 57400 56324 57452
rect 56376 57440 56382 57452
rect 56873 57443 56931 57449
rect 56873 57440 56885 57443
rect 56376 57412 56885 57440
rect 56376 57400 56382 57412
rect 56873 57409 56885 57412
rect 56919 57409 56931 57443
rect 65061 57443 65119 57449
rect 65061 57440 65073 57443
rect 56873 57403 56931 57409
rect 64846 57412 65073 57440
rect 39298 57332 39304 57384
rect 39356 57372 39362 57384
rect 64846 57372 64874 57412
rect 65061 57409 65073 57412
rect 65107 57440 65119 57443
rect 65613 57443 65671 57449
rect 65613 57440 65625 57443
rect 65107 57412 65625 57440
rect 65107 57409 65119 57412
rect 65061 57403 65119 57409
rect 65613 57409 65625 57412
rect 65659 57409 65671 57443
rect 67634 57440 67640 57452
rect 67595 57412 67640 57440
rect 65613 57403 65671 57409
rect 67634 57400 67640 57412
rect 67692 57400 67698 57452
rect 39356 57344 64874 57372
rect 39356 57332 39362 57344
rect 30098 57236 30104 57248
rect 30059 57208 30104 57236
rect 30098 57196 30104 57208
rect 30156 57196 30162 57248
rect 39206 57236 39212 57248
rect 39167 57208 39212 57236
rect 39206 57196 39212 57208
rect 39264 57196 39270 57248
rect 56318 57236 56324 57248
rect 56279 57208 56324 57236
rect 56318 57196 56324 57208
rect 56376 57196 56382 57248
rect 1104 57146 68816 57168
rect 1104 57094 4214 57146
rect 4266 57094 4278 57146
rect 4330 57094 4342 57146
rect 4394 57094 4406 57146
rect 4458 57094 4470 57146
rect 4522 57094 34934 57146
rect 34986 57094 34998 57146
rect 35050 57094 35062 57146
rect 35114 57094 35126 57146
rect 35178 57094 35190 57146
rect 35242 57094 65654 57146
rect 65706 57094 65718 57146
rect 65770 57094 65782 57146
rect 65834 57094 65846 57146
rect 65898 57094 65910 57146
rect 65962 57094 68816 57146
rect 1104 57072 68816 57094
rect 27154 56992 27160 57044
rect 27212 57032 27218 57044
rect 39206 57032 39212 57044
rect 27212 57004 39212 57032
rect 27212 56992 27218 57004
rect 39206 56992 39212 57004
rect 39264 56992 39270 57044
rect 21634 56652 21640 56704
rect 21692 56692 21698 56704
rect 21729 56695 21787 56701
rect 21729 56692 21741 56695
rect 21692 56664 21741 56692
rect 21692 56652 21698 56664
rect 21729 56661 21741 56664
rect 21775 56661 21787 56695
rect 21729 56655 21787 56661
rect 1104 56602 68816 56624
rect 1104 56550 19574 56602
rect 19626 56550 19638 56602
rect 19690 56550 19702 56602
rect 19754 56550 19766 56602
rect 19818 56550 19830 56602
rect 19882 56550 50294 56602
rect 50346 56550 50358 56602
rect 50410 56550 50422 56602
rect 50474 56550 50486 56602
rect 50538 56550 50550 56602
rect 50602 56550 68816 56602
rect 1104 56528 68816 56550
rect 67634 56148 67640 56160
rect 67595 56120 67640 56148
rect 67634 56108 67640 56120
rect 67692 56108 67698 56160
rect 1104 56058 68816 56080
rect 1104 56006 4214 56058
rect 4266 56006 4278 56058
rect 4330 56006 4342 56058
rect 4394 56006 4406 56058
rect 4458 56006 4470 56058
rect 4522 56006 34934 56058
rect 34986 56006 34998 56058
rect 35050 56006 35062 56058
rect 35114 56006 35126 56058
rect 35178 56006 35190 56058
rect 35242 56006 65654 56058
rect 65706 56006 65718 56058
rect 65770 56006 65782 56058
rect 65834 56006 65846 56058
rect 65898 56006 65910 56058
rect 65962 56006 68816 56058
rect 1104 55984 68816 56006
rect 1104 55514 68816 55536
rect 1104 55462 19574 55514
rect 19626 55462 19638 55514
rect 19690 55462 19702 55514
rect 19754 55462 19766 55514
rect 19818 55462 19830 55514
rect 19882 55462 50294 55514
rect 50346 55462 50358 55514
rect 50410 55462 50422 55514
rect 50474 55462 50486 55514
rect 50538 55462 50550 55514
rect 50602 55462 68816 55514
rect 1104 55440 68816 55462
rect 1104 54970 68816 54992
rect 1104 54918 4214 54970
rect 4266 54918 4278 54970
rect 4330 54918 4342 54970
rect 4394 54918 4406 54970
rect 4458 54918 4470 54970
rect 4522 54918 34934 54970
rect 34986 54918 34998 54970
rect 35050 54918 35062 54970
rect 35114 54918 35126 54970
rect 35178 54918 35190 54970
rect 35242 54918 65654 54970
rect 65706 54918 65718 54970
rect 65770 54918 65782 54970
rect 65834 54918 65846 54970
rect 65898 54918 65910 54970
rect 65962 54918 68816 54970
rect 1104 54896 68816 54918
rect 68094 54652 68100 54664
rect 68055 54624 68100 54652
rect 68094 54612 68100 54624
rect 68152 54612 68158 54664
rect 1104 54426 68816 54448
rect 1104 54374 19574 54426
rect 19626 54374 19638 54426
rect 19690 54374 19702 54426
rect 19754 54374 19766 54426
rect 19818 54374 19830 54426
rect 19882 54374 50294 54426
rect 50346 54374 50358 54426
rect 50410 54374 50422 54426
rect 50474 54374 50486 54426
rect 50538 54374 50550 54426
rect 50602 54374 68816 54426
rect 1104 54352 68816 54374
rect 1104 53882 68816 53904
rect 1104 53830 4214 53882
rect 4266 53830 4278 53882
rect 4330 53830 4342 53882
rect 4394 53830 4406 53882
rect 4458 53830 4470 53882
rect 4522 53830 34934 53882
rect 34986 53830 34998 53882
rect 35050 53830 35062 53882
rect 35114 53830 35126 53882
rect 35178 53830 35190 53882
rect 35242 53830 65654 53882
rect 65706 53830 65718 53882
rect 65770 53830 65782 53882
rect 65834 53830 65846 53882
rect 65898 53830 65910 53882
rect 65962 53830 68816 53882
rect 1104 53808 68816 53830
rect 68094 53564 68100 53576
rect 68055 53536 68100 53564
rect 68094 53524 68100 53536
rect 68152 53524 68158 53576
rect 1104 53338 68816 53360
rect 1104 53286 19574 53338
rect 19626 53286 19638 53338
rect 19690 53286 19702 53338
rect 19754 53286 19766 53338
rect 19818 53286 19830 53338
rect 19882 53286 50294 53338
rect 50346 53286 50358 53338
rect 50410 53286 50422 53338
rect 50474 53286 50486 53338
rect 50538 53286 50550 53338
rect 50602 53286 68816 53338
rect 1104 53264 68816 53286
rect 1104 52794 68816 52816
rect 1104 52742 4214 52794
rect 4266 52742 4278 52794
rect 4330 52742 4342 52794
rect 4394 52742 4406 52794
rect 4458 52742 4470 52794
rect 4522 52742 34934 52794
rect 34986 52742 34998 52794
rect 35050 52742 35062 52794
rect 35114 52742 35126 52794
rect 35178 52742 35190 52794
rect 35242 52742 65654 52794
rect 65706 52742 65718 52794
rect 65770 52742 65782 52794
rect 65834 52742 65846 52794
rect 65898 52742 65910 52794
rect 65962 52742 68816 52794
rect 1104 52720 68816 52742
rect 1104 52250 68816 52272
rect 1104 52198 19574 52250
rect 19626 52198 19638 52250
rect 19690 52198 19702 52250
rect 19754 52198 19766 52250
rect 19818 52198 19830 52250
rect 19882 52198 50294 52250
rect 50346 52198 50358 52250
rect 50410 52198 50422 52250
rect 50474 52198 50486 52250
rect 50538 52198 50550 52250
rect 50602 52198 68816 52250
rect 1104 52176 68816 52198
rect 67634 51796 67640 51808
rect 67595 51768 67640 51796
rect 67634 51756 67640 51768
rect 67692 51756 67698 51808
rect 1104 51706 68816 51728
rect 1104 51654 4214 51706
rect 4266 51654 4278 51706
rect 4330 51654 4342 51706
rect 4394 51654 4406 51706
rect 4458 51654 4470 51706
rect 4522 51654 34934 51706
rect 34986 51654 34998 51706
rect 35050 51654 35062 51706
rect 35114 51654 35126 51706
rect 35178 51654 35190 51706
rect 35242 51654 65654 51706
rect 65706 51654 65718 51706
rect 65770 51654 65782 51706
rect 65834 51654 65846 51706
rect 65898 51654 65910 51706
rect 65962 51654 68816 51706
rect 1104 51632 68816 51654
rect 1104 51162 68816 51184
rect 1104 51110 19574 51162
rect 19626 51110 19638 51162
rect 19690 51110 19702 51162
rect 19754 51110 19766 51162
rect 19818 51110 19830 51162
rect 19882 51110 50294 51162
rect 50346 51110 50358 51162
rect 50410 51110 50422 51162
rect 50474 51110 50486 51162
rect 50538 51110 50550 51162
rect 50602 51110 68816 51162
rect 1104 51088 68816 51110
rect 1104 50618 68816 50640
rect 1104 50566 4214 50618
rect 4266 50566 4278 50618
rect 4330 50566 4342 50618
rect 4394 50566 4406 50618
rect 4458 50566 4470 50618
rect 4522 50566 34934 50618
rect 34986 50566 34998 50618
rect 35050 50566 35062 50618
rect 35114 50566 35126 50618
rect 35178 50566 35190 50618
rect 35242 50566 65654 50618
rect 65706 50566 65718 50618
rect 65770 50566 65782 50618
rect 65834 50566 65846 50618
rect 65898 50566 65910 50618
rect 65962 50566 68816 50618
rect 1104 50544 68816 50566
rect 68094 50300 68100 50312
rect 68055 50272 68100 50300
rect 68094 50260 68100 50272
rect 68152 50260 68158 50312
rect 1104 50074 68816 50096
rect 1104 50022 19574 50074
rect 19626 50022 19638 50074
rect 19690 50022 19702 50074
rect 19754 50022 19766 50074
rect 19818 50022 19830 50074
rect 19882 50022 50294 50074
rect 50346 50022 50358 50074
rect 50410 50022 50422 50074
rect 50474 50022 50486 50074
rect 50538 50022 50550 50074
rect 50602 50022 68816 50074
rect 1104 50000 68816 50022
rect 1104 49530 68816 49552
rect 1104 49478 4214 49530
rect 4266 49478 4278 49530
rect 4330 49478 4342 49530
rect 4394 49478 4406 49530
rect 4458 49478 4470 49530
rect 4522 49478 34934 49530
rect 34986 49478 34998 49530
rect 35050 49478 35062 49530
rect 35114 49478 35126 49530
rect 35178 49478 35190 49530
rect 35242 49478 65654 49530
rect 65706 49478 65718 49530
rect 65770 49478 65782 49530
rect 65834 49478 65846 49530
rect 65898 49478 65910 49530
rect 65962 49478 68816 49530
rect 1104 49456 68816 49478
rect 1104 48986 68816 49008
rect 1104 48934 19574 48986
rect 19626 48934 19638 48986
rect 19690 48934 19702 48986
rect 19754 48934 19766 48986
rect 19818 48934 19830 48986
rect 19882 48934 50294 48986
rect 50346 48934 50358 48986
rect 50410 48934 50422 48986
rect 50474 48934 50486 48986
rect 50538 48934 50550 48986
rect 50602 48934 68816 48986
rect 1104 48912 68816 48934
rect 67634 48600 67640 48612
rect 67595 48572 67640 48600
rect 67634 48560 67640 48572
rect 67692 48560 67698 48612
rect 1104 48442 68816 48464
rect 1104 48390 4214 48442
rect 4266 48390 4278 48442
rect 4330 48390 4342 48442
rect 4394 48390 4406 48442
rect 4458 48390 4470 48442
rect 4522 48390 34934 48442
rect 34986 48390 34998 48442
rect 35050 48390 35062 48442
rect 35114 48390 35126 48442
rect 35178 48390 35190 48442
rect 35242 48390 65654 48442
rect 65706 48390 65718 48442
rect 65770 48390 65782 48442
rect 65834 48390 65846 48442
rect 65898 48390 65910 48442
rect 65962 48390 68816 48442
rect 1104 48368 68816 48390
rect 1104 47898 68816 47920
rect 1104 47846 19574 47898
rect 19626 47846 19638 47898
rect 19690 47846 19702 47898
rect 19754 47846 19766 47898
rect 19818 47846 19830 47898
rect 19882 47846 50294 47898
rect 50346 47846 50358 47898
rect 50410 47846 50422 47898
rect 50474 47846 50486 47898
rect 50538 47846 50550 47898
rect 50602 47846 68816 47898
rect 1104 47824 68816 47846
rect 67634 47444 67640 47456
rect 67595 47416 67640 47444
rect 67634 47404 67640 47416
rect 67692 47404 67698 47456
rect 1104 47354 68816 47376
rect 1104 47302 4214 47354
rect 4266 47302 4278 47354
rect 4330 47302 4342 47354
rect 4394 47302 4406 47354
rect 4458 47302 4470 47354
rect 4522 47302 34934 47354
rect 34986 47302 34998 47354
rect 35050 47302 35062 47354
rect 35114 47302 35126 47354
rect 35178 47302 35190 47354
rect 35242 47302 65654 47354
rect 65706 47302 65718 47354
rect 65770 47302 65782 47354
rect 65834 47302 65846 47354
rect 65898 47302 65910 47354
rect 65962 47302 68816 47354
rect 1104 47280 68816 47302
rect 1104 46810 68816 46832
rect 1104 46758 19574 46810
rect 19626 46758 19638 46810
rect 19690 46758 19702 46810
rect 19754 46758 19766 46810
rect 19818 46758 19830 46810
rect 19882 46758 50294 46810
rect 50346 46758 50358 46810
rect 50410 46758 50422 46810
rect 50474 46758 50486 46810
rect 50538 46758 50550 46810
rect 50602 46758 68816 46810
rect 1104 46736 68816 46758
rect 1104 46266 68816 46288
rect 1104 46214 4214 46266
rect 4266 46214 4278 46266
rect 4330 46214 4342 46266
rect 4394 46214 4406 46266
rect 4458 46214 4470 46266
rect 4522 46214 34934 46266
rect 34986 46214 34998 46266
rect 35050 46214 35062 46266
rect 35114 46214 35126 46266
rect 35178 46214 35190 46266
rect 35242 46214 65654 46266
rect 65706 46214 65718 46266
rect 65770 46214 65782 46266
rect 65834 46214 65846 46266
rect 65898 46214 65910 46266
rect 65962 46214 68816 46266
rect 1104 46192 68816 46214
rect 68094 45948 68100 45960
rect 68055 45920 68100 45948
rect 68094 45908 68100 45920
rect 68152 45908 68158 45960
rect 1104 45722 68816 45744
rect 1104 45670 19574 45722
rect 19626 45670 19638 45722
rect 19690 45670 19702 45722
rect 19754 45670 19766 45722
rect 19818 45670 19830 45722
rect 19882 45670 50294 45722
rect 50346 45670 50358 45722
rect 50410 45670 50422 45722
rect 50474 45670 50486 45722
rect 50538 45670 50550 45722
rect 50602 45670 68816 45722
rect 1104 45648 68816 45670
rect 1104 45178 68816 45200
rect 1104 45126 4214 45178
rect 4266 45126 4278 45178
rect 4330 45126 4342 45178
rect 4394 45126 4406 45178
rect 4458 45126 4470 45178
rect 4522 45126 34934 45178
rect 34986 45126 34998 45178
rect 35050 45126 35062 45178
rect 35114 45126 35126 45178
rect 35178 45126 35190 45178
rect 35242 45126 65654 45178
rect 65706 45126 65718 45178
rect 65770 45126 65782 45178
rect 65834 45126 65846 45178
rect 65898 45126 65910 45178
rect 65962 45126 68816 45178
rect 1104 45104 68816 45126
rect 1104 44634 68816 44656
rect 1104 44582 19574 44634
rect 19626 44582 19638 44634
rect 19690 44582 19702 44634
rect 19754 44582 19766 44634
rect 19818 44582 19830 44634
rect 19882 44582 50294 44634
rect 50346 44582 50358 44634
rect 50410 44582 50422 44634
rect 50474 44582 50486 44634
rect 50538 44582 50550 44634
rect 50602 44582 68816 44634
rect 1104 44560 68816 44582
rect 67542 44140 67548 44192
rect 67600 44180 67606 44192
rect 67637 44183 67695 44189
rect 67637 44180 67649 44183
rect 67600 44152 67649 44180
rect 67600 44140 67606 44152
rect 67637 44149 67649 44152
rect 67683 44149 67695 44183
rect 67637 44143 67695 44149
rect 1104 44090 68816 44112
rect 1104 44038 4214 44090
rect 4266 44038 4278 44090
rect 4330 44038 4342 44090
rect 4394 44038 4406 44090
rect 4458 44038 4470 44090
rect 4522 44038 34934 44090
rect 34986 44038 34998 44090
rect 35050 44038 35062 44090
rect 35114 44038 35126 44090
rect 35178 44038 35190 44090
rect 35242 44038 65654 44090
rect 65706 44038 65718 44090
rect 65770 44038 65782 44090
rect 65834 44038 65846 44090
rect 65898 44038 65910 44090
rect 65962 44038 68816 44090
rect 1104 44016 68816 44038
rect 1104 43546 68816 43568
rect 1104 43494 19574 43546
rect 19626 43494 19638 43546
rect 19690 43494 19702 43546
rect 19754 43494 19766 43546
rect 19818 43494 19830 43546
rect 19882 43494 50294 43546
rect 50346 43494 50358 43546
rect 50410 43494 50422 43546
rect 50474 43494 50486 43546
rect 50538 43494 50550 43546
rect 50602 43494 68816 43546
rect 1104 43472 68816 43494
rect 1104 43002 68816 43024
rect 1104 42950 4214 43002
rect 4266 42950 4278 43002
rect 4330 42950 4342 43002
rect 4394 42950 4406 43002
rect 4458 42950 4470 43002
rect 4522 42950 34934 43002
rect 34986 42950 34998 43002
rect 35050 42950 35062 43002
rect 35114 42950 35126 43002
rect 35178 42950 35190 43002
rect 35242 42950 65654 43002
rect 65706 42950 65718 43002
rect 65770 42950 65782 43002
rect 65834 42950 65846 43002
rect 65898 42950 65910 43002
rect 65962 42950 68816 43002
rect 1104 42928 68816 42950
rect 68094 42684 68100 42696
rect 68055 42656 68100 42684
rect 68094 42644 68100 42656
rect 68152 42644 68158 42696
rect 1104 42458 68816 42480
rect 1104 42406 19574 42458
rect 19626 42406 19638 42458
rect 19690 42406 19702 42458
rect 19754 42406 19766 42458
rect 19818 42406 19830 42458
rect 19882 42406 50294 42458
rect 50346 42406 50358 42458
rect 50410 42406 50422 42458
rect 50474 42406 50486 42458
rect 50538 42406 50550 42458
rect 50602 42406 68816 42458
rect 1104 42384 68816 42406
rect 1104 41914 68816 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 34934 41914
rect 34986 41862 34998 41914
rect 35050 41862 35062 41914
rect 35114 41862 35126 41914
rect 35178 41862 35190 41914
rect 35242 41862 65654 41914
rect 65706 41862 65718 41914
rect 65770 41862 65782 41914
rect 65834 41862 65846 41914
rect 65898 41862 65910 41914
rect 65962 41862 68816 41914
rect 1104 41840 68816 41862
rect 68094 41596 68100 41608
rect 68055 41568 68100 41596
rect 68094 41556 68100 41568
rect 68152 41556 68158 41608
rect 1104 41370 68816 41392
rect 1104 41318 19574 41370
rect 19626 41318 19638 41370
rect 19690 41318 19702 41370
rect 19754 41318 19766 41370
rect 19818 41318 19830 41370
rect 19882 41318 50294 41370
rect 50346 41318 50358 41370
rect 50410 41318 50422 41370
rect 50474 41318 50486 41370
rect 50538 41318 50550 41370
rect 50602 41318 68816 41370
rect 1104 41296 68816 41318
rect 1104 40826 68816 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 34934 40826
rect 34986 40774 34998 40826
rect 35050 40774 35062 40826
rect 35114 40774 35126 40826
rect 35178 40774 35190 40826
rect 35242 40774 65654 40826
rect 65706 40774 65718 40826
rect 65770 40774 65782 40826
rect 65834 40774 65846 40826
rect 65898 40774 65910 40826
rect 65962 40774 68816 40826
rect 1104 40752 68816 40774
rect 1104 40282 68816 40304
rect 1104 40230 19574 40282
rect 19626 40230 19638 40282
rect 19690 40230 19702 40282
rect 19754 40230 19766 40282
rect 19818 40230 19830 40282
rect 19882 40230 50294 40282
rect 50346 40230 50358 40282
rect 50410 40230 50422 40282
rect 50474 40230 50486 40282
rect 50538 40230 50550 40282
rect 50602 40230 68816 40282
rect 1104 40208 68816 40230
rect 67634 39828 67640 39840
rect 67595 39800 67640 39828
rect 67634 39788 67640 39800
rect 67692 39788 67698 39840
rect 1104 39738 68816 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 65654 39738
rect 65706 39686 65718 39738
rect 65770 39686 65782 39738
rect 65834 39686 65846 39738
rect 65898 39686 65910 39738
rect 65962 39686 68816 39738
rect 1104 39664 68816 39686
rect 1104 39194 68816 39216
rect 1104 39142 19574 39194
rect 19626 39142 19638 39194
rect 19690 39142 19702 39194
rect 19754 39142 19766 39194
rect 19818 39142 19830 39194
rect 19882 39142 50294 39194
rect 50346 39142 50358 39194
rect 50410 39142 50422 39194
rect 50474 39142 50486 39194
rect 50538 39142 50550 39194
rect 50602 39142 68816 39194
rect 1104 39120 68816 39142
rect 1104 38650 68816 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 65654 38650
rect 65706 38598 65718 38650
rect 65770 38598 65782 38650
rect 65834 38598 65846 38650
rect 65898 38598 65910 38650
rect 65962 38598 68816 38650
rect 1104 38576 68816 38598
rect 68094 38332 68100 38344
rect 68055 38304 68100 38332
rect 68094 38292 68100 38304
rect 68152 38292 68158 38344
rect 1104 38106 68816 38128
rect 1104 38054 19574 38106
rect 19626 38054 19638 38106
rect 19690 38054 19702 38106
rect 19754 38054 19766 38106
rect 19818 38054 19830 38106
rect 19882 38054 50294 38106
rect 50346 38054 50358 38106
rect 50410 38054 50422 38106
rect 50474 38054 50486 38106
rect 50538 38054 50550 38106
rect 50602 38054 68816 38106
rect 1104 38032 68816 38054
rect 1104 37562 68816 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 65654 37562
rect 65706 37510 65718 37562
rect 65770 37510 65782 37562
rect 65834 37510 65846 37562
rect 65898 37510 65910 37562
rect 65962 37510 68816 37562
rect 1104 37488 68816 37510
rect 1104 37018 68816 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 50294 37018
rect 50346 36966 50358 37018
rect 50410 36966 50422 37018
rect 50474 36966 50486 37018
rect 50538 36966 50550 37018
rect 50602 36966 68816 37018
rect 1104 36944 68816 36966
rect 67634 36632 67640 36644
rect 67595 36604 67640 36632
rect 67634 36592 67640 36604
rect 67692 36592 67698 36644
rect 1104 36474 68816 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 65654 36474
rect 65706 36422 65718 36474
rect 65770 36422 65782 36474
rect 65834 36422 65846 36474
rect 65898 36422 65910 36474
rect 65962 36422 68816 36474
rect 1104 36400 68816 36422
rect 1104 35930 68816 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 50294 35930
rect 50346 35878 50358 35930
rect 50410 35878 50422 35930
rect 50474 35878 50486 35930
rect 50538 35878 50550 35930
rect 50602 35878 68816 35930
rect 1104 35856 68816 35878
rect 67634 35476 67640 35488
rect 67595 35448 67640 35476
rect 67634 35436 67640 35448
rect 67692 35436 67698 35488
rect 1104 35386 68816 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 65654 35386
rect 65706 35334 65718 35386
rect 65770 35334 65782 35386
rect 65834 35334 65846 35386
rect 65898 35334 65910 35386
rect 65962 35334 68816 35386
rect 1104 35312 68816 35334
rect 1104 34842 68816 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 50294 34842
rect 50346 34790 50358 34842
rect 50410 34790 50422 34842
rect 50474 34790 50486 34842
rect 50538 34790 50550 34842
rect 50602 34790 68816 34842
rect 1104 34768 68816 34790
rect 1104 34298 68816 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 65654 34298
rect 65706 34246 65718 34298
rect 65770 34246 65782 34298
rect 65834 34246 65846 34298
rect 65898 34246 65910 34298
rect 65962 34246 68816 34298
rect 1104 34224 68816 34246
rect 68094 33980 68100 33992
rect 68055 33952 68100 33980
rect 68094 33940 68100 33952
rect 68152 33940 68158 33992
rect 1104 33754 68816 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 50294 33754
rect 50346 33702 50358 33754
rect 50410 33702 50422 33754
rect 50474 33702 50486 33754
rect 50538 33702 50550 33754
rect 50602 33702 68816 33754
rect 1104 33680 68816 33702
rect 1104 33210 68816 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 65654 33210
rect 65706 33158 65718 33210
rect 65770 33158 65782 33210
rect 65834 33158 65846 33210
rect 65898 33158 65910 33210
rect 65962 33158 68816 33210
rect 1104 33136 68816 33158
rect 1104 32666 68816 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 50294 32666
rect 50346 32614 50358 32666
rect 50410 32614 50422 32666
rect 50474 32614 50486 32666
rect 50538 32614 50550 32666
rect 50602 32614 68816 32666
rect 1104 32592 68816 32614
rect 67634 32212 67640 32224
rect 67595 32184 67640 32212
rect 67634 32172 67640 32184
rect 67692 32172 67698 32224
rect 1104 32122 68816 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 65654 32122
rect 65706 32070 65718 32122
rect 65770 32070 65782 32122
rect 65834 32070 65846 32122
rect 65898 32070 65910 32122
rect 65962 32070 68816 32122
rect 1104 32048 68816 32070
rect 1104 31578 68816 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 50294 31578
rect 50346 31526 50358 31578
rect 50410 31526 50422 31578
rect 50474 31526 50486 31578
rect 50538 31526 50550 31578
rect 50602 31526 68816 31578
rect 1104 31504 68816 31526
rect 1104 31034 68816 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 65654 31034
rect 65706 30982 65718 31034
rect 65770 30982 65782 31034
rect 65834 30982 65846 31034
rect 65898 30982 65910 31034
rect 65962 30982 68816 31034
rect 1104 30960 68816 30982
rect 68094 30716 68100 30728
rect 68055 30688 68100 30716
rect 68094 30676 68100 30688
rect 68152 30676 68158 30728
rect 1104 30490 68816 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 50294 30490
rect 50346 30438 50358 30490
rect 50410 30438 50422 30490
rect 50474 30438 50486 30490
rect 50538 30438 50550 30490
rect 50602 30438 68816 30490
rect 1104 30416 68816 30438
rect 7193 30243 7251 30249
rect 7193 30209 7205 30243
rect 7239 30240 7251 30243
rect 7558 30240 7564 30252
rect 7239 30212 7564 30240
rect 7239 30209 7251 30212
rect 7193 30203 7251 30209
rect 7558 30200 7564 30212
rect 7616 30200 7622 30252
rect 8021 30243 8079 30249
rect 8021 30209 8033 30243
rect 8067 30240 8079 30243
rect 30098 30240 30104 30252
rect 8067 30212 30104 30240
rect 8067 30209 8079 30212
rect 8021 30203 8079 30209
rect 30098 30200 30104 30212
rect 30156 30200 30162 30252
rect 6730 30132 6736 30184
rect 6788 30172 6794 30184
rect 6917 30175 6975 30181
rect 6917 30172 6929 30175
rect 6788 30144 6929 30172
rect 6788 30132 6794 30144
rect 6917 30141 6929 30144
rect 6963 30141 6975 30175
rect 6917 30135 6975 30141
rect 1104 29946 68816 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 65654 29946
rect 65706 29894 65718 29946
rect 65770 29894 65782 29946
rect 65834 29894 65846 29946
rect 65898 29894 65910 29946
rect 65962 29894 68816 29946
rect 1104 29872 68816 29894
rect 27154 29832 27160 29844
rect 27115 29804 27160 29832
rect 27154 29792 27160 29804
rect 27212 29792 27218 29844
rect 7291 29631 7349 29637
rect 7291 29597 7303 29631
rect 7337 29628 7349 29631
rect 7469 29631 7527 29637
rect 7337 29600 7420 29628
rect 7337 29597 7349 29600
rect 7291 29591 7349 29597
rect 7392 29560 7420 29600
rect 7469 29597 7481 29631
rect 7515 29628 7527 29631
rect 8018 29628 8024 29640
rect 7515 29600 8024 29628
rect 7515 29597 7527 29600
rect 7469 29591 7527 29597
rect 8018 29588 8024 29600
rect 8076 29588 8082 29640
rect 25774 29588 25780 29640
rect 25832 29628 25838 29640
rect 26145 29631 26203 29637
rect 26145 29628 26157 29631
rect 25832 29600 26157 29628
rect 25832 29588 25838 29600
rect 26145 29597 26157 29600
rect 26191 29597 26203 29631
rect 26418 29628 26424 29640
rect 26379 29600 26424 29628
rect 26145 29591 26203 29597
rect 26418 29588 26424 29600
rect 26476 29588 26482 29640
rect 68094 29628 68100 29640
rect 68055 29600 68100 29628
rect 68094 29588 68100 29600
rect 68152 29588 68158 29640
rect 7926 29560 7932 29572
rect 7392 29532 7932 29560
rect 7926 29520 7932 29532
rect 7984 29520 7990 29572
rect 7377 29495 7435 29501
rect 7377 29461 7389 29495
rect 7423 29492 7435 29495
rect 7558 29492 7564 29504
rect 7423 29464 7564 29492
rect 7423 29461 7435 29464
rect 7377 29455 7435 29461
rect 7558 29452 7564 29464
rect 7616 29452 7622 29504
rect 1104 29402 68816 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 50294 29402
rect 50346 29350 50358 29402
rect 50410 29350 50422 29402
rect 50474 29350 50486 29402
rect 50538 29350 50550 29402
rect 50602 29350 68816 29402
rect 1104 29328 68816 29350
rect 7926 29220 7932 29232
rect 6748 29192 7932 29220
rect 5074 29152 5080 29164
rect 5035 29124 5080 29152
rect 5074 29112 5080 29124
rect 5132 29112 5138 29164
rect 6748 29161 6776 29192
rect 7926 29180 7932 29192
rect 7984 29180 7990 29232
rect 6733 29155 6791 29161
rect 6733 29121 6745 29155
rect 6779 29121 6791 29155
rect 6733 29115 6791 29121
rect 7837 29155 7895 29161
rect 7837 29121 7849 29155
rect 7883 29121 7895 29155
rect 7837 29115 7895 29121
rect 19337 29155 19395 29161
rect 19337 29121 19349 29155
rect 19383 29152 19395 29155
rect 19886 29152 19892 29164
rect 19383 29124 19892 29152
rect 19383 29121 19395 29124
rect 19337 29115 19395 29121
rect 4801 29087 4859 29093
rect 4801 29053 4813 29087
rect 4847 29053 4859 29087
rect 4801 29047 4859 29053
rect 6549 29087 6607 29093
rect 6549 29053 6561 29087
rect 6595 29084 6607 29087
rect 7006 29084 7012 29096
rect 6595 29056 7012 29084
rect 6595 29053 6607 29056
rect 6549 29047 6607 29053
rect 4816 28960 4844 29047
rect 7006 29044 7012 29056
rect 7064 29084 7070 29096
rect 7852 29084 7880 29115
rect 19886 29112 19892 29124
rect 19944 29112 19950 29164
rect 24489 29155 24547 29161
rect 24489 29121 24501 29155
rect 24535 29152 24547 29155
rect 25038 29152 25044 29164
rect 24535 29124 25044 29152
rect 24535 29121 24547 29124
rect 24489 29115 24547 29121
rect 25038 29112 25044 29124
rect 25096 29112 25102 29164
rect 8110 29084 8116 29096
rect 7064 29056 8116 29084
rect 7064 29044 7070 29056
rect 8110 29044 8116 29056
rect 8168 29044 8174 29096
rect 19426 29084 19432 29096
rect 19387 29056 19432 29084
rect 19426 29044 19432 29056
rect 19484 29044 19490 29096
rect 5810 29016 5816 29028
rect 5771 28988 5816 29016
rect 5810 28976 5816 28988
rect 5868 28976 5874 29028
rect 7745 29019 7803 29025
rect 7745 28985 7757 29019
rect 7791 29016 7803 29019
rect 8018 29016 8024 29028
rect 7791 28988 8024 29016
rect 7791 28985 7803 28988
rect 7745 28979 7803 28985
rect 8018 28976 8024 28988
rect 8076 28976 8082 29028
rect 8297 29019 8355 29025
rect 8297 28985 8309 29019
rect 8343 28985 8355 29019
rect 18966 29016 18972 29028
rect 18927 28988 18972 29016
rect 8297 28979 8355 28985
rect 4798 28948 4804 28960
rect 4711 28920 4804 28948
rect 4798 28908 4804 28920
rect 4856 28948 4862 28960
rect 6730 28948 6736 28960
rect 4856 28920 6736 28948
rect 4856 28908 4862 28920
rect 6730 28908 6736 28920
rect 6788 28908 6794 28960
rect 6914 28948 6920 28960
rect 6875 28920 6920 28948
rect 6914 28908 6920 28920
rect 6972 28908 6978 28960
rect 7650 28908 7656 28960
rect 7708 28948 7714 28960
rect 8312 28948 8340 28979
rect 18966 28976 18972 28988
rect 19024 28976 19030 29028
rect 7708 28920 8340 28948
rect 9217 28951 9275 28957
rect 7708 28908 7714 28920
rect 9217 28917 9229 28951
rect 9263 28948 9275 28951
rect 9398 28948 9404 28960
rect 9263 28920 9404 28948
rect 9263 28917 9275 28920
rect 9217 28911 9275 28917
rect 9398 28908 9404 28920
rect 9456 28908 9462 28960
rect 24394 28948 24400 28960
rect 24355 28920 24400 28948
rect 24394 28908 24400 28920
rect 24452 28908 24458 28960
rect 1104 28858 68816 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 65654 28858
rect 65706 28806 65718 28858
rect 65770 28806 65782 28858
rect 65834 28806 65846 28858
rect 65898 28806 65910 28858
rect 65962 28806 68816 28858
rect 1104 28784 68816 28806
rect 6730 28744 6736 28756
rect 6691 28716 6736 28744
rect 6730 28704 6736 28716
rect 6788 28704 6794 28756
rect 8294 28744 8300 28756
rect 8255 28716 8300 28744
rect 8294 28704 8300 28716
rect 8352 28704 8358 28756
rect 16945 28747 17003 28753
rect 16945 28713 16957 28747
rect 16991 28744 17003 28747
rect 17773 28747 17831 28753
rect 17773 28744 17785 28747
rect 16991 28716 17785 28744
rect 16991 28713 17003 28716
rect 16945 28707 17003 28713
rect 17773 28713 17785 28716
rect 17819 28713 17831 28747
rect 17773 28707 17831 28713
rect 18233 28747 18291 28753
rect 18233 28713 18245 28747
rect 18279 28744 18291 28747
rect 18279 28716 19196 28744
rect 18279 28713 18291 28716
rect 18233 28707 18291 28713
rect 6089 28679 6147 28685
rect 6089 28676 6101 28679
rect 5460 28648 6101 28676
rect 4798 28568 4804 28620
rect 4856 28608 4862 28620
rect 4856 28580 4901 28608
rect 4856 28568 4862 28580
rect 4525 28543 4583 28549
rect 4525 28509 4537 28543
rect 4571 28509 4583 28543
rect 4525 28503 4583 28509
rect 4540 28472 4568 28503
rect 5074 28500 5080 28552
rect 5132 28540 5138 28552
rect 5460 28549 5488 28648
rect 6089 28645 6101 28648
rect 6135 28645 6147 28679
rect 6089 28639 6147 28645
rect 9674 28636 9680 28688
rect 9732 28636 9738 28688
rect 18966 28676 18972 28688
rect 16776 28648 18972 28676
rect 9309 28611 9367 28617
rect 9309 28608 9321 28611
rect 5644 28580 9321 28608
rect 5644 28549 5672 28580
rect 9309 28577 9321 28580
rect 9355 28577 9367 28611
rect 9309 28571 9367 28577
rect 5445 28543 5503 28549
rect 5445 28540 5457 28543
rect 5132 28512 5457 28540
rect 5132 28500 5138 28512
rect 5445 28509 5457 28512
rect 5491 28509 5503 28543
rect 5445 28503 5503 28509
rect 5629 28543 5687 28549
rect 5629 28509 5641 28543
rect 5675 28509 5687 28543
rect 6270 28540 6276 28552
rect 6231 28512 6276 28540
rect 5629 28503 5687 28509
rect 6270 28500 6276 28512
rect 6328 28500 6334 28552
rect 6914 28540 6920 28552
rect 6875 28512 6920 28540
rect 6914 28500 6920 28512
rect 6972 28500 6978 28552
rect 7650 28500 7656 28552
rect 7708 28540 7714 28552
rect 7929 28543 7987 28549
rect 7929 28540 7941 28543
rect 7708 28512 7941 28540
rect 7708 28500 7714 28512
rect 7929 28509 7941 28512
rect 7975 28509 7987 28543
rect 8110 28540 8116 28552
rect 8071 28512 8116 28540
rect 7929 28503 7987 28509
rect 8110 28500 8116 28512
rect 8168 28500 8174 28552
rect 9398 28500 9404 28552
rect 9456 28540 9462 28552
rect 9689 28549 9717 28636
rect 16776 28617 16804 28648
rect 18966 28636 18972 28648
rect 19024 28636 19030 28688
rect 16761 28611 16819 28617
rect 16761 28577 16773 28611
rect 16807 28577 16819 28611
rect 16761 28571 16819 28577
rect 17957 28611 18015 28617
rect 17957 28577 17969 28611
rect 18003 28608 18015 28611
rect 18598 28608 18604 28620
rect 18003 28580 18604 28608
rect 18003 28577 18015 28580
rect 17957 28571 18015 28577
rect 18598 28568 18604 28580
rect 18656 28568 18662 28620
rect 19168 28608 19196 28716
rect 19242 28704 19248 28756
rect 19300 28744 19306 28756
rect 19705 28747 19763 28753
rect 19705 28744 19717 28747
rect 19300 28716 19717 28744
rect 19300 28704 19306 28716
rect 19705 28713 19717 28716
rect 19751 28713 19763 28747
rect 23845 28747 23903 28753
rect 23845 28744 23857 28747
rect 19705 28707 19763 28713
rect 21100 28716 23857 28744
rect 19904 28648 20852 28676
rect 19904 28608 19932 28648
rect 19168 28580 19932 28608
rect 9585 28543 9643 28549
rect 9585 28540 9597 28543
rect 9456 28512 9597 28540
rect 9456 28500 9462 28512
rect 9585 28509 9597 28512
rect 9631 28509 9643 28543
rect 9585 28503 9643 28509
rect 9674 28543 9732 28549
rect 9674 28509 9686 28543
rect 9720 28509 9732 28543
rect 9674 28503 9732 28509
rect 9769 28543 9827 28549
rect 9769 28509 9781 28543
rect 9815 28540 9827 28543
rect 9965 28543 10023 28549
rect 9815 28512 9884 28540
rect 9815 28509 9827 28512
rect 9769 28503 9827 28509
rect 5537 28475 5595 28481
rect 5537 28472 5549 28475
rect 4540 28444 5549 28472
rect 5537 28441 5549 28444
rect 5583 28441 5595 28475
rect 8389 28475 8447 28481
rect 8389 28472 8401 28475
rect 5537 28435 5595 28441
rect 7944 28444 8401 28472
rect 7944 28416 7972 28444
rect 8389 28441 8401 28444
rect 8435 28441 8447 28475
rect 8389 28435 8447 28441
rect 9122 28432 9128 28484
rect 9180 28472 9186 28484
rect 9180 28444 9674 28472
rect 9180 28432 9186 28444
rect 3786 28404 3792 28416
rect 3747 28376 3792 28404
rect 3786 28364 3792 28376
rect 3844 28364 3850 28416
rect 7745 28407 7803 28413
rect 7745 28373 7757 28407
rect 7791 28404 7803 28407
rect 7834 28404 7840 28416
rect 7791 28376 7840 28404
rect 7791 28373 7803 28376
rect 7745 28367 7803 28373
rect 7834 28364 7840 28376
rect 7892 28364 7898 28416
rect 7926 28364 7932 28416
rect 7984 28364 7990 28416
rect 9646 28404 9674 28444
rect 9856 28404 9884 28512
rect 9965 28509 9977 28543
rect 10011 28540 10023 28543
rect 10226 28540 10232 28552
rect 10011 28512 10232 28540
rect 10011 28509 10023 28512
rect 9965 28503 10023 28509
rect 10226 28500 10232 28512
rect 10284 28500 10290 28552
rect 13998 28500 14004 28552
rect 14056 28540 14062 28552
rect 15565 28543 15623 28549
rect 15565 28540 15577 28543
rect 14056 28512 15577 28540
rect 14056 28500 14062 28512
rect 15565 28509 15577 28512
rect 15611 28509 15623 28543
rect 15565 28503 15623 28509
rect 16669 28543 16727 28549
rect 16669 28509 16681 28543
rect 16715 28509 16727 28543
rect 18046 28540 18052 28552
rect 18007 28512 18052 28540
rect 16669 28503 16727 28509
rect 15378 28472 15384 28484
rect 15339 28444 15384 28472
rect 15378 28432 15384 28444
rect 15436 28432 15442 28484
rect 16684 28472 16712 28503
rect 18046 28500 18052 28512
rect 18104 28500 18110 28552
rect 19334 28500 19340 28552
rect 19392 28540 19398 28552
rect 19886 28540 19892 28552
rect 19392 28512 19892 28540
rect 19392 28500 19398 28512
rect 19886 28500 19892 28512
rect 19944 28500 19950 28552
rect 19981 28543 20039 28549
rect 19981 28509 19993 28543
rect 20027 28540 20039 28543
rect 20070 28540 20076 28552
rect 20027 28512 20076 28540
rect 20027 28509 20039 28512
rect 19981 28503 20039 28509
rect 20070 28500 20076 28512
rect 20128 28500 20134 28552
rect 20824 28549 20852 28648
rect 21100 28549 21128 28716
rect 23845 28713 23857 28716
rect 23891 28744 23903 28747
rect 26050 28744 26056 28756
rect 23891 28716 26056 28744
rect 23891 28713 23903 28716
rect 23845 28707 23903 28713
rect 26050 28704 26056 28716
rect 26108 28704 26114 28756
rect 21729 28611 21787 28617
rect 21729 28608 21741 28611
rect 21652 28580 21741 28608
rect 20625 28543 20683 28549
rect 20625 28540 20637 28543
rect 20180 28512 20637 28540
rect 16758 28472 16764 28484
rect 16684 28444 16764 28472
rect 16758 28432 16764 28444
rect 16816 28432 16822 28484
rect 17770 28472 17776 28484
rect 17731 28444 17776 28472
rect 17770 28432 17776 28444
rect 17828 28432 17834 28484
rect 19705 28475 19763 28481
rect 19705 28441 19717 28475
rect 19751 28441 19763 28475
rect 19705 28435 19763 28441
rect 9646 28376 9884 28404
rect 15749 28407 15807 28413
rect 15749 28373 15761 28407
rect 15795 28404 15807 28407
rect 19426 28404 19432 28416
rect 15795 28376 19432 28404
rect 15795 28373 15807 28376
rect 15749 28367 15807 28373
rect 19426 28364 19432 28376
rect 19484 28404 19490 28416
rect 19720 28404 19748 28435
rect 20070 28404 20076 28416
rect 19484 28376 20076 28404
rect 19484 28364 19490 28376
rect 20070 28364 20076 28376
rect 20128 28364 20134 28416
rect 20180 28413 20208 28512
rect 20625 28509 20637 28512
rect 20671 28509 20683 28543
rect 20625 28503 20683 28509
rect 20809 28543 20867 28549
rect 20809 28509 20821 28543
rect 20855 28509 20867 28543
rect 20809 28503 20867 28509
rect 21085 28543 21143 28549
rect 21085 28509 21097 28543
rect 21131 28509 21143 28543
rect 21085 28503 21143 28509
rect 21652 28472 21680 28580
rect 21729 28577 21741 28580
rect 21775 28577 21787 28611
rect 21729 28571 21787 28577
rect 25682 28568 25688 28620
rect 25740 28608 25746 28620
rect 25777 28611 25835 28617
rect 25777 28608 25789 28611
rect 25740 28580 25789 28608
rect 25740 28568 25746 28580
rect 25777 28577 25789 28580
rect 25823 28577 25835 28611
rect 25777 28571 25835 28577
rect 22002 28540 22008 28552
rect 21963 28512 22008 28540
rect 22002 28500 22008 28512
rect 22060 28500 22066 28552
rect 23198 28540 23204 28552
rect 23159 28512 23204 28540
rect 23198 28500 23204 28512
rect 23256 28500 23262 28552
rect 23290 28500 23296 28552
rect 23348 28540 23354 28552
rect 23720 28543 23778 28549
rect 23348 28512 23393 28540
rect 23348 28500 23354 28512
rect 23720 28509 23732 28543
rect 23766 28540 23778 28543
rect 24394 28540 24400 28552
rect 23766 28512 24400 28540
rect 23766 28509 23778 28512
rect 23720 28503 23778 28509
rect 24394 28500 24400 28512
rect 24452 28500 24458 28552
rect 25038 28540 25044 28552
rect 24999 28512 25044 28540
rect 25038 28500 25044 28512
rect 25096 28500 25102 28552
rect 25130 28500 25136 28552
rect 25188 28540 25194 28552
rect 26050 28540 26056 28552
rect 25188 28512 25233 28540
rect 26011 28512 26056 28540
rect 25188 28500 25194 28512
rect 26050 28500 26056 28512
rect 26108 28500 26114 28552
rect 25682 28472 25688 28484
rect 21652 28444 25688 28472
rect 25682 28432 25688 28444
rect 25740 28432 25746 28484
rect 20165 28407 20223 28413
rect 20165 28373 20177 28407
rect 20211 28373 20223 28407
rect 20165 28367 20223 28373
rect 21269 28407 21327 28413
rect 21269 28373 21281 28407
rect 21315 28404 21327 28407
rect 22002 28404 22008 28416
rect 21315 28376 22008 28404
rect 21315 28373 21327 28376
rect 21269 28367 21327 28373
rect 22002 28364 22008 28376
rect 22060 28364 22066 28416
rect 22741 28407 22799 28413
rect 22741 28373 22753 28407
rect 22787 28404 22799 28407
rect 23566 28404 23572 28416
rect 22787 28376 23572 28404
rect 22787 28373 22799 28376
rect 22741 28367 22799 28373
rect 23566 28364 23572 28376
rect 23624 28364 23630 28416
rect 23661 28407 23719 28413
rect 23661 28373 23673 28407
rect 23707 28404 23719 28407
rect 25130 28404 25136 28416
rect 23707 28376 25136 28404
rect 23707 28373 23719 28376
rect 23661 28367 23719 28373
rect 25130 28364 25136 28376
rect 25188 28364 25194 28416
rect 25317 28407 25375 28413
rect 25317 28373 25329 28407
rect 25363 28404 25375 28407
rect 25590 28404 25596 28416
rect 25363 28376 25596 28404
rect 25363 28373 25375 28376
rect 25317 28367 25375 28373
rect 25590 28364 25596 28376
rect 25648 28364 25654 28416
rect 26786 28404 26792 28416
rect 26747 28376 26792 28404
rect 26786 28364 26792 28376
rect 26844 28364 26850 28416
rect 1104 28314 68816 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 50294 28314
rect 50346 28262 50358 28314
rect 50410 28262 50422 28314
rect 50474 28262 50486 28314
rect 50538 28262 50550 28314
rect 50602 28262 68816 28314
rect 1104 28240 68816 28262
rect 6270 28160 6276 28212
rect 6328 28200 6334 28212
rect 7377 28203 7435 28209
rect 7377 28200 7389 28203
rect 6328 28172 7389 28200
rect 6328 28160 6334 28172
rect 7377 28169 7389 28172
rect 7423 28169 7435 28203
rect 9122 28200 9128 28212
rect 9083 28172 9128 28200
rect 7377 28163 7435 28169
rect 9122 28160 9128 28172
rect 9180 28160 9186 28212
rect 9493 28203 9551 28209
rect 9493 28169 9505 28203
rect 9539 28200 9551 28203
rect 9674 28200 9680 28212
rect 9539 28172 9680 28200
rect 9539 28169 9551 28172
rect 9493 28163 9551 28169
rect 9674 28160 9680 28172
rect 9732 28200 9738 28212
rect 11609 28203 11667 28209
rect 11609 28200 11621 28203
rect 9732 28172 11621 28200
rect 9732 28160 9738 28172
rect 11609 28169 11621 28172
rect 11655 28169 11667 28203
rect 11609 28163 11667 28169
rect 20533 28203 20591 28209
rect 20533 28169 20545 28203
rect 20579 28200 20591 28203
rect 23198 28200 23204 28212
rect 20579 28172 23204 28200
rect 20579 28169 20591 28172
rect 20533 28163 20591 28169
rect 23198 28160 23204 28172
rect 23256 28160 23262 28212
rect 23290 28160 23296 28212
rect 23348 28200 23354 28212
rect 23937 28203 23995 28209
rect 23937 28200 23949 28203
rect 23348 28172 23949 28200
rect 23348 28160 23354 28172
rect 23937 28169 23949 28172
rect 23983 28169 23995 28203
rect 23937 28163 23995 28169
rect 25682 28160 25688 28212
rect 25740 28200 25746 28212
rect 25777 28203 25835 28209
rect 25777 28200 25789 28203
rect 25740 28172 25789 28200
rect 25740 28160 25746 28172
rect 25777 28169 25789 28172
rect 25823 28169 25835 28203
rect 25777 28163 25835 28169
rect 14001 28135 14059 28141
rect 14001 28101 14013 28135
rect 14047 28132 14059 28135
rect 15289 28135 15347 28141
rect 15289 28132 15301 28135
rect 14047 28104 15301 28132
rect 14047 28101 14059 28104
rect 14001 28095 14059 28101
rect 15289 28101 15301 28104
rect 15335 28101 15347 28135
rect 15289 28095 15347 28101
rect 7558 28064 7564 28076
rect 7519 28036 7564 28064
rect 7558 28024 7564 28036
rect 7616 28024 7622 28076
rect 7834 28064 7840 28076
rect 7795 28036 7840 28064
rect 7834 28024 7840 28036
rect 7892 28024 7898 28076
rect 8021 28067 8079 28073
rect 8021 28033 8033 28067
rect 8067 28033 8079 28067
rect 8021 28027 8079 28033
rect 8036 27996 8064 28027
rect 8570 28024 8576 28076
rect 8628 28064 8634 28076
rect 9398 28064 9404 28076
rect 8628 28036 9404 28064
rect 8628 28024 8634 28036
rect 9398 28024 9404 28036
rect 9456 28024 9462 28076
rect 11517 28067 11575 28073
rect 11517 28033 11529 28067
rect 11563 28064 11575 28067
rect 11606 28064 11612 28076
rect 11563 28036 11612 28064
rect 11563 28033 11575 28036
rect 11517 28027 11575 28033
rect 11606 28024 11612 28036
rect 11664 28024 11670 28076
rect 11701 28067 11759 28073
rect 11701 28033 11713 28067
rect 11747 28064 11759 28067
rect 12158 28064 12164 28076
rect 11747 28036 12164 28064
rect 11747 28033 11759 28036
rect 11701 28027 11759 28033
rect 12158 28024 12164 28036
rect 12216 28024 12222 28076
rect 13817 28067 13875 28073
rect 13817 28033 13829 28067
rect 13863 28033 13875 28067
rect 13817 28027 13875 28033
rect 15105 28067 15163 28073
rect 15105 28033 15117 28067
rect 15151 28033 15163 28067
rect 15105 28027 15163 28033
rect 9582 27996 9588 28008
rect 8036 27968 9588 27996
rect 9582 27956 9588 27968
rect 9640 27956 9646 28008
rect 13832 27996 13860 28027
rect 13998 27996 14004 28008
rect 13832 27968 14004 27996
rect 13998 27956 14004 27968
rect 14056 27956 14062 28008
rect 8294 27888 8300 27940
rect 8352 27928 8358 27940
rect 9125 27931 9183 27937
rect 9125 27928 9137 27931
rect 8352 27900 9137 27928
rect 8352 27888 8358 27900
rect 9125 27897 9137 27900
rect 9171 27928 9183 27931
rect 9490 27928 9496 27940
rect 9171 27900 9496 27928
rect 9171 27897 9183 27900
rect 9125 27891 9183 27897
rect 9490 27888 9496 27900
rect 9548 27888 9554 27940
rect 15120 27928 15148 28027
rect 15304 27996 15332 28095
rect 18046 28092 18052 28144
rect 18104 28132 18110 28144
rect 22370 28132 22376 28144
rect 18104 28104 22376 28132
rect 18104 28092 18110 28104
rect 22370 28092 22376 28104
rect 22428 28132 22434 28144
rect 22428 28104 23704 28132
rect 22428 28092 22434 28104
rect 18141 28067 18199 28073
rect 18141 28033 18153 28067
rect 18187 28064 18199 28067
rect 18230 28064 18236 28076
rect 18187 28036 18236 28064
rect 18187 28033 18199 28036
rect 18141 28027 18199 28033
rect 18230 28024 18236 28036
rect 18288 28024 18294 28076
rect 18325 28067 18383 28073
rect 18325 28033 18337 28067
rect 18371 28064 18383 28067
rect 19334 28064 19340 28076
rect 18371 28036 19340 28064
rect 18371 28033 18383 28036
rect 18325 28027 18383 28033
rect 18340 27996 18368 28027
rect 19334 28024 19340 28036
rect 19392 28024 19398 28076
rect 19518 28064 19524 28076
rect 19479 28036 19524 28064
rect 19518 28024 19524 28036
rect 19576 28024 19582 28076
rect 20070 28024 20076 28076
rect 20128 28064 20134 28076
rect 20165 28067 20223 28073
rect 20165 28064 20177 28067
rect 20128 28036 20177 28064
rect 20128 28024 20134 28036
rect 20165 28033 20177 28036
rect 20211 28033 20223 28067
rect 23474 28064 23480 28076
rect 23435 28036 23480 28064
rect 20165 28027 20223 28033
rect 23474 28024 23480 28036
rect 23532 28024 23538 28076
rect 23676 28073 23704 28104
rect 23661 28067 23719 28073
rect 23661 28033 23673 28067
rect 23707 28033 23719 28067
rect 23661 28027 23719 28033
rect 23753 28067 23811 28073
rect 23753 28033 23765 28067
rect 23799 28064 23811 28067
rect 24394 28064 24400 28076
rect 23799 28036 24400 28064
rect 23799 28033 23811 28036
rect 23753 28027 23811 28033
rect 24394 28024 24400 28036
rect 24452 28024 24458 28076
rect 24581 28067 24639 28073
rect 24581 28033 24593 28067
rect 24627 28064 24639 28067
rect 25130 28064 25136 28076
rect 24627 28036 25136 28064
rect 24627 28033 24639 28036
rect 24581 28027 24639 28033
rect 15304 27968 18368 27996
rect 19705 27999 19763 28005
rect 19705 27965 19717 27999
rect 19751 27996 19763 27999
rect 19978 27996 19984 28008
rect 19751 27968 19984 27996
rect 19751 27965 19763 27968
rect 19705 27959 19763 27965
rect 19978 27956 19984 27968
rect 20036 27956 20042 28008
rect 20257 27999 20315 28005
rect 20257 27965 20269 27999
rect 20303 27965 20315 27999
rect 20257 27959 20315 27965
rect 15378 27928 15384 27940
rect 15120 27900 15384 27928
rect 15378 27888 15384 27900
rect 15436 27928 15442 27940
rect 17218 27928 17224 27940
rect 15436 27900 17224 27928
rect 15436 27888 15442 27900
rect 17218 27888 17224 27900
rect 17276 27888 17282 27940
rect 18322 27888 18328 27940
rect 18380 27928 18386 27940
rect 19242 27928 19248 27940
rect 18380 27900 19248 27928
rect 18380 27888 18386 27900
rect 19242 27888 19248 27900
rect 19300 27928 19306 27940
rect 20272 27928 20300 27959
rect 24596 27928 24624 28027
rect 25130 28024 25136 28036
rect 25188 28024 25194 28076
rect 25590 28064 25596 28076
rect 25551 28036 25596 28064
rect 25590 28024 25596 28036
rect 25648 28024 25654 28076
rect 19300 27900 20300 27928
rect 23768 27900 24624 27928
rect 19300 27888 19306 27900
rect 9214 27860 9220 27872
rect 9175 27832 9220 27860
rect 9214 27820 9220 27832
rect 9272 27820 9278 27872
rect 9306 27820 9312 27872
rect 9364 27860 9370 27872
rect 10597 27863 10655 27869
rect 9364 27832 9409 27860
rect 9364 27820 9370 27832
rect 10597 27829 10609 27863
rect 10643 27860 10655 27863
rect 10870 27860 10876 27872
rect 10643 27832 10876 27860
rect 10643 27829 10655 27832
rect 10597 27823 10655 27829
rect 10870 27820 10876 27832
rect 10928 27820 10934 27872
rect 13633 27863 13691 27869
rect 13633 27829 13645 27863
rect 13679 27860 13691 27863
rect 13906 27860 13912 27872
rect 13679 27832 13912 27860
rect 13679 27829 13691 27832
rect 13633 27823 13691 27829
rect 13906 27820 13912 27832
rect 13964 27820 13970 27872
rect 14550 27820 14556 27872
rect 14608 27860 14614 27872
rect 14921 27863 14979 27869
rect 14921 27860 14933 27863
rect 14608 27832 14933 27860
rect 14608 27820 14614 27832
rect 14921 27829 14933 27832
rect 14967 27829 14979 27863
rect 17402 27860 17408 27872
rect 17363 27832 17408 27860
rect 14921 27823 14979 27829
rect 17402 27820 17408 27832
rect 17460 27820 17466 27872
rect 17954 27860 17960 27872
rect 17915 27832 17960 27860
rect 17954 27820 17960 27832
rect 18012 27820 18018 27872
rect 19518 27820 19524 27872
rect 19576 27860 19582 27872
rect 20349 27863 20407 27869
rect 20349 27860 20361 27863
rect 19576 27832 20361 27860
rect 19576 27820 19582 27832
rect 20349 27829 20361 27832
rect 20395 27860 20407 27863
rect 22462 27860 22468 27872
rect 20395 27832 22468 27860
rect 20395 27829 20407 27832
rect 20349 27823 20407 27829
rect 22462 27820 22468 27832
rect 22520 27820 22526 27872
rect 23768 27869 23796 27900
rect 23753 27863 23811 27869
rect 23753 27829 23765 27863
rect 23799 27829 23811 27863
rect 23753 27823 23811 27829
rect 24302 27820 24308 27872
rect 24360 27860 24366 27872
rect 24581 27863 24639 27869
rect 24581 27860 24593 27863
rect 24360 27832 24593 27860
rect 24360 27820 24366 27832
rect 24581 27829 24593 27832
rect 24627 27860 24639 27863
rect 26418 27860 26424 27872
rect 24627 27832 26424 27860
rect 24627 27829 24639 27832
rect 24581 27823 24639 27829
rect 26418 27820 26424 27832
rect 26476 27820 26482 27872
rect 67634 27860 67640 27872
rect 67595 27832 67640 27860
rect 67634 27820 67640 27832
rect 67692 27820 67698 27872
rect 1104 27770 68816 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 65654 27770
rect 65706 27718 65718 27770
rect 65770 27718 65782 27770
rect 65834 27718 65846 27770
rect 65898 27718 65910 27770
rect 65962 27718 68816 27770
rect 1104 27696 68816 27718
rect 3786 27616 3792 27668
rect 3844 27656 3850 27668
rect 4414 27659 4472 27665
rect 4414 27656 4426 27659
rect 3844 27628 4426 27656
rect 3844 27616 3850 27628
rect 4414 27625 4426 27628
rect 4460 27625 4472 27659
rect 4414 27619 4472 27625
rect 8389 27659 8447 27665
rect 8389 27625 8401 27659
rect 8435 27656 8447 27659
rect 9306 27656 9312 27668
rect 8435 27628 9312 27656
rect 8435 27625 8447 27628
rect 8389 27619 8447 27625
rect 9306 27616 9312 27628
rect 9364 27616 9370 27668
rect 10226 27656 10232 27668
rect 10187 27628 10232 27656
rect 10226 27616 10232 27628
rect 10284 27616 10290 27668
rect 10873 27659 10931 27665
rect 10873 27625 10885 27659
rect 10919 27625 10931 27659
rect 10873 27619 10931 27625
rect 14660 27628 17908 27656
rect 2409 27591 2467 27597
rect 2409 27557 2421 27591
rect 2455 27588 2467 27591
rect 5905 27591 5963 27597
rect 2455 27560 2774 27588
rect 2455 27557 2467 27560
rect 2409 27551 2467 27557
rect 1946 27520 1952 27532
rect 1907 27492 1952 27520
rect 1946 27480 1952 27492
rect 2004 27480 2010 27532
rect 2746 27520 2774 27560
rect 5905 27557 5917 27591
rect 5951 27588 5963 27591
rect 7006 27588 7012 27600
rect 5951 27560 7012 27588
rect 5951 27557 5963 27560
rect 5905 27551 5963 27557
rect 7006 27548 7012 27560
rect 7064 27548 7070 27600
rect 9582 27548 9588 27600
rect 9640 27588 9646 27600
rect 9861 27591 9919 27597
rect 9861 27588 9873 27591
rect 9640 27560 9873 27588
rect 9640 27548 9646 27560
rect 9861 27557 9873 27560
rect 9907 27557 9919 27591
rect 10888 27588 10916 27619
rect 9861 27551 9919 27557
rect 10060 27560 10916 27588
rect 10060 27529 10088 27560
rect 9953 27523 10011 27529
rect 9953 27520 9965 27523
rect 2746 27492 9965 27520
rect 9953 27489 9965 27492
rect 9999 27489 10011 27523
rect 9953 27483 10011 27489
rect 10045 27523 10103 27529
rect 10045 27489 10057 27523
rect 10091 27489 10103 27523
rect 10870 27520 10876 27532
rect 10831 27492 10876 27520
rect 10045 27483 10103 27489
rect 10870 27480 10876 27492
rect 10928 27480 10934 27532
rect 10965 27523 11023 27529
rect 10965 27489 10977 27523
rect 11011 27489 11023 27523
rect 10965 27483 11023 27489
rect 2041 27455 2099 27461
rect 2041 27421 2053 27455
rect 2087 27452 2099 27455
rect 2869 27455 2927 27461
rect 2869 27452 2881 27455
rect 2087 27424 2881 27452
rect 2087 27421 2099 27424
rect 2041 27415 2099 27421
rect 2869 27421 2881 27424
rect 2915 27421 2927 27455
rect 2869 27415 2927 27421
rect 2884 27316 2912 27415
rect 2958 27412 2964 27464
rect 3016 27452 3022 27464
rect 4157 27455 4215 27461
rect 4157 27452 4169 27455
rect 3016 27424 4169 27452
rect 3016 27412 3022 27424
rect 4157 27421 4169 27424
rect 4203 27421 4215 27455
rect 7742 27452 7748 27464
rect 7703 27424 7748 27452
rect 4157 27415 4215 27421
rect 7742 27412 7748 27424
rect 7800 27412 7806 27464
rect 7926 27461 7932 27464
rect 7893 27455 7932 27461
rect 7893 27421 7905 27455
rect 7893 27415 7932 27421
rect 7926 27412 7932 27415
rect 7984 27412 7990 27464
rect 8018 27412 8024 27464
rect 8076 27452 8082 27464
rect 8251 27455 8309 27461
rect 8076 27424 8121 27452
rect 8076 27412 8082 27424
rect 8251 27421 8263 27455
rect 8297 27452 8309 27455
rect 9398 27452 9404 27464
rect 8297 27424 9404 27452
rect 8297 27421 8309 27424
rect 8251 27415 8309 27421
rect 9398 27412 9404 27424
rect 9456 27412 9462 27464
rect 9766 27412 9772 27464
rect 9824 27452 9830 27464
rect 10980 27452 11008 27483
rect 13814 27480 13820 27532
rect 13872 27520 13878 27532
rect 14660 27520 14688 27628
rect 13872 27492 14688 27520
rect 13872 27480 13878 27492
rect 9824 27424 9869 27452
rect 9968 27424 11008 27452
rect 11057 27455 11115 27461
rect 9824 27412 9830 27424
rect 5166 27344 5172 27396
rect 5224 27344 5230 27396
rect 8113 27387 8171 27393
rect 8113 27384 8125 27387
rect 7208 27356 8125 27384
rect 7208 27328 7236 27356
rect 8113 27353 8125 27356
rect 8159 27353 8171 27387
rect 9968 27384 9996 27424
rect 11057 27421 11069 27455
rect 11103 27421 11115 27455
rect 11057 27415 11115 27421
rect 10686 27384 10692 27396
rect 8113 27347 8171 27353
rect 8220 27356 9996 27384
rect 10647 27356 10692 27384
rect 5718 27316 5724 27328
rect 2884 27288 5724 27316
rect 5718 27276 5724 27288
rect 5776 27276 5782 27328
rect 7190 27316 7196 27328
rect 7151 27288 7196 27316
rect 7190 27276 7196 27288
rect 7248 27276 7254 27328
rect 8018 27276 8024 27328
rect 8076 27316 8082 27328
rect 8220 27316 8248 27356
rect 8076 27288 8248 27316
rect 8076 27276 8082 27288
rect 8570 27276 8576 27328
rect 8628 27316 8634 27328
rect 9692 27325 9720 27356
rect 10686 27344 10692 27356
rect 10744 27344 10750 27396
rect 8941 27319 8999 27325
rect 8941 27316 8953 27319
rect 8628 27288 8953 27316
rect 8628 27276 8634 27288
rect 8941 27285 8953 27288
rect 8987 27285 8999 27319
rect 8941 27279 8999 27285
rect 9677 27319 9735 27325
rect 9677 27285 9689 27319
rect 9723 27285 9735 27319
rect 9677 27279 9735 27285
rect 9950 27276 9956 27328
rect 10008 27316 10014 27328
rect 11072 27316 11100 27415
rect 11514 27412 11520 27464
rect 11572 27452 11578 27464
rect 11793 27455 11851 27461
rect 11793 27452 11805 27455
rect 11572 27424 11805 27452
rect 11572 27412 11578 27424
rect 11793 27421 11805 27424
rect 11839 27421 11851 27455
rect 11793 27415 11851 27421
rect 14369 27455 14427 27461
rect 14369 27421 14381 27455
rect 14415 27421 14427 27455
rect 14550 27452 14556 27464
rect 14511 27424 14556 27452
rect 14369 27415 14427 27421
rect 12060 27387 12118 27393
rect 12060 27353 12072 27387
rect 12106 27384 12118 27387
rect 13446 27384 13452 27396
rect 12106 27356 13452 27384
rect 12106 27353 12118 27356
rect 12060 27347 12118 27353
rect 13446 27344 13452 27356
rect 13504 27344 13510 27396
rect 13078 27316 13084 27328
rect 10008 27288 13084 27316
rect 10008 27276 10014 27288
rect 13078 27276 13084 27288
rect 13136 27276 13142 27328
rect 13173 27319 13231 27325
rect 13173 27285 13185 27319
rect 13219 27316 13231 27319
rect 13998 27316 14004 27328
rect 13219 27288 14004 27316
rect 13219 27285 13231 27288
rect 13173 27279 13231 27285
rect 13998 27276 14004 27288
rect 14056 27276 14062 27328
rect 14090 27276 14096 27328
rect 14148 27316 14154 27328
rect 14384 27316 14412 27415
rect 14550 27412 14556 27424
rect 14608 27412 14614 27464
rect 14660 27461 14688 27492
rect 17880 27520 17908 27628
rect 19334 27616 19340 27668
rect 19392 27656 19398 27668
rect 21266 27656 21272 27668
rect 19392 27628 21272 27656
rect 19392 27616 19398 27628
rect 21266 27616 21272 27628
rect 21324 27616 21330 27668
rect 25038 27616 25044 27668
rect 25096 27656 25102 27668
rect 25961 27659 26019 27665
rect 25961 27656 25973 27659
rect 25096 27628 25973 27656
rect 25096 27616 25102 27628
rect 25961 27625 25973 27628
rect 26007 27625 26019 27659
rect 25961 27619 26019 27625
rect 26786 27616 26792 27668
rect 26844 27656 26850 27668
rect 27445 27659 27503 27665
rect 27445 27656 27457 27659
rect 26844 27628 27457 27656
rect 26844 27616 26850 27628
rect 27445 27625 27457 27628
rect 27491 27625 27503 27659
rect 27445 27619 27503 27625
rect 20346 27588 20352 27600
rect 19306 27560 20352 27588
rect 19306 27520 19334 27560
rect 20346 27548 20352 27560
rect 20404 27548 20410 27600
rect 17880 27492 19334 27520
rect 14645 27455 14703 27461
rect 14645 27421 14657 27455
rect 14691 27421 14703 27455
rect 14645 27415 14703 27421
rect 14734 27412 14740 27464
rect 14792 27452 14798 27464
rect 15473 27455 15531 27461
rect 14792 27424 14837 27452
rect 14792 27412 14798 27424
rect 15473 27421 15485 27455
rect 15519 27452 15531 27455
rect 16574 27452 16580 27464
rect 15519 27424 16580 27452
rect 15519 27421 15531 27424
rect 15473 27415 15531 27421
rect 16574 27412 16580 27424
rect 16632 27412 16638 27464
rect 17402 27412 17408 27464
rect 17460 27452 17466 27464
rect 17880 27461 17908 27492
rect 19794 27480 19800 27532
rect 19852 27520 19858 27532
rect 21085 27523 21143 27529
rect 21085 27520 21097 27523
rect 19852 27492 21097 27520
rect 19852 27480 19858 27492
rect 21085 27489 21097 27492
rect 21131 27489 21143 27523
rect 21085 27483 21143 27489
rect 17773 27455 17831 27461
rect 17773 27452 17785 27455
rect 17460 27424 17785 27452
rect 17460 27412 17466 27424
rect 17773 27421 17785 27424
rect 17819 27421 17831 27455
rect 17773 27415 17831 27421
rect 17865 27455 17923 27461
rect 17865 27421 17877 27455
rect 17911 27421 17923 27455
rect 17865 27415 17923 27421
rect 17954 27412 17960 27464
rect 18012 27452 18018 27464
rect 18141 27455 18199 27461
rect 18012 27424 18057 27452
rect 18012 27412 18018 27424
rect 18141 27421 18153 27455
rect 18187 27452 18199 27455
rect 19886 27452 19892 27464
rect 18187 27424 19892 27452
rect 18187 27421 18199 27424
rect 18141 27415 18199 27421
rect 15013 27387 15071 27393
rect 15013 27353 15025 27387
rect 15059 27384 15071 27387
rect 15718 27387 15776 27393
rect 15718 27384 15730 27387
rect 15059 27356 15730 27384
rect 15059 27353 15071 27356
rect 15013 27347 15071 27353
rect 15718 27353 15730 27356
rect 15764 27353 15776 27387
rect 18156 27384 18184 27415
rect 19886 27412 19892 27424
rect 19944 27412 19950 27464
rect 19978 27412 19984 27464
rect 20036 27452 20042 27464
rect 20073 27455 20131 27461
rect 20073 27452 20085 27455
rect 20036 27424 20085 27452
rect 20036 27412 20042 27424
rect 20073 27421 20085 27424
rect 20119 27421 20131 27455
rect 20073 27415 20131 27421
rect 20165 27455 20223 27461
rect 20165 27421 20177 27455
rect 20211 27421 20223 27455
rect 20165 27415 20223 27421
rect 19794 27384 19800 27396
rect 15718 27347 15776 27353
rect 15856 27356 18184 27384
rect 18248 27356 19800 27384
rect 15856 27316 15884 27356
rect 14148 27288 15884 27316
rect 16853 27319 16911 27325
rect 14148 27276 14154 27288
rect 16853 27285 16865 27319
rect 16899 27316 16911 27319
rect 17218 27316 17224 27328
rect 16899 27288 17224 27316
rect 16899 27285 16911 27288
rect 16853 27279 16911 27285
rect 17218 27276 17224 27288
rect 17276 27276 17282 27328
rect 17494 27316 17500 27328
rect 17455 27288 17500 27316
rect 17494 27276 17500 27288
rect 17552 27276 17558 27328
rect 17678 27276 17684 27328
rect 17736 27316 17742 27328
rect 18248 27316 18276 27356
rect 19794 27344 19800 27356
rect 19852 27344 19858 27396
rect 20180 27384 20208 27415
rect 20254 27412 20260 27464
rect 20312 27452 20318 27464
rect 27709 27455 27767 27461
rect 20312 27424 20357 27452
rect 20312 27412 20318 27424
rect 27709 27421 27721 27455
rect 27755 27452 27767 27455
rect 27890 27452 27896 27464
rect 27755 27424 27896 27452
rect 27755 27421 27767 27424
rect 27709 27415 27767 27421
rect 27890 27412 27896 27424
rect 27948 27412 27954 27464
rect 20346 27384 20352 27396
rect 20180 27356 20352 27384
rect 20346 27344 20352 27356
rect 20404 27344 20410 27396
rect 20533 27387 20591 27393
rect 20533 27353 20545 27387
rect 20579 27384 20591 27387
rect 21330 27387 21388 27393
rect 21330 27384 21342 27387
rect 20579 27356 21342 27384
rect 20579 27353 20591 27356
rect 20533 27347 20591 27353
rect 21330 27353 21342 27356
rect 21376 27353 21388 27387
rect 21330 27347 21388 27353
rect 26970 27344 26976 27396
rect 27028 27344 27034 27396
rect 17736 27288 18276 27316
rect 19429 27319 19487 27325
rect 17736 27276 17742 27288
rect 19429 27285 19441 27319
rect 19475 27316 19487 27319
rect 20254 27316 20260 27328
rect 19475 27288 20260 27316
rect 19475 27285 19487 27288
rect 19429 27279 19487 27285
rect 20254 27276 20260 27288
rect 20312 27276 20318 27328
rect 22462 27316 22468 27328
rect 22375 27288 22468 27316
rect 22462 27276 22468 27288
rect 22520 27316 22526 27328
rect 23198 27316 23204 27328
rect 22520 27288 23204 27316
rect 22520 27276 22526 27288
rect 23198 27276 23204 27288
rect 23256 27276 23262 27328
rect 1104 27226 68816 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 50294 27226
rect 50346 27174 50358 27226
rect 50410 27174 50422 27226
rect 50474 27174 50486 27226
rect 50538 27174 50550 27226
rect 50602 27174 68816 27226
rect 1104 27152 68816 27174
rect 1946 27072 1952 27124
rect 2004 27112 2010 27124
rect 2041 27115 2099 27121
rect 2041 27112 2053 27115
rect 2004 27084 2053 27112
rect 2004 27072 2010 27084
rect 2041 27081 2053 27084
rect 2087 27081 2099 27115
rect 4614 27112 4620 27124
rect 2041 27075 2099 27081
rect 2746 27084 4620 27112
rect 1673 26979 1731 26985
rect 1673 26945 1685 26979
rect 1719 26976 1731 26979
rect 2501 26979 2559 26985
rect 2501 26976 2513 26979
rect 1719 26948 2513 26976
rect 1719 26945 1731 26948
rect 1673 26939 1731 26945
rect 2501 26945 2513 26948
rect 2547 26976 2559 26979
rect 2746 26976 2774 27084
rect 4614 27072 4620 27084
rect 4672 27072 4678 27124
rect 5166 27072 5172 27124
rect 5224 27112 5230 27124
rect 5261 27115 5319 27121
rect 5261 27112 5273 27115
rect 5224 27084 5273 27112
rect 5224 27072 5230 27084
rect 5261 27081 5273 27084
rect 5307 27081 5319 27115
rect 8757 27115 8815 27121
rect 8757 27112 8769 27115
rect 5261 27075 5319 27081
rect 5736 27084 8769 27112
rect 4632 27044 4660 27072
rect 5736 27044 5764 27084
rect 8757 27081 8769 27084
rect 8803 27081 8815 27115
rect 8757 27075 8815 27081
rect 4632 27016 5764 27044
rect 5810 27004 5816 27056
rect 5868 27044 5874 27056
rect 6641 27047 6699 27053
rect 6641 27044 6653 27047
rect 5868 27016 6653 27044
rect 5868 27004 5874 27016
rect 6641 27013 6653 27016
rect 6687 27013 6699 27047
rect 6641 27007 6699 27013
rect 7098 27004 7104 27056
rect 7156 27004 7162 27056
rect 8772 27044 8800 27075
rect 9398 27072 9404 27124
rect 9456 27112 9462 27124
rect 9674 27112 9680 27124
rect 9456 27084 9680 27112
rect 9456 27072 9462 27084
rect 9674 27072 9680 27084
rect 9732 27112 9738 27124
rect 10686 27112 10692 27124
rect 9732 27084 10692 27112
rect 9732 27072 9738 27084
rect 10686 27072 10692 27084
rect 10744 27072 10750 27124
rect 11517 27115 11575 27121
rect 11517 27081 11529 27115
rect 11563 27112 11575 27115
rect 11606 27112 11612 27124
rect 11563 27084 11612 27112
rect 11563 27081 11575 27084
rect 11517 27075 11575 27081
rect 11606 27072 11612 27084
rect 11664 27072 11670 27124
rect 13446 27112 13452 27124
rect 13407 27084 13452 27112
rect 13446 27072 13452 27084
rect 13504 27072 13510 27124
rect 14366 27072 14372 27124
rect 14424 27112 14430 27124
rect 18230 27112 18236 27124
rect 14424 27084 18236 27112
rect 14424 27072 14430 27084
rect 18230 27072 18236 27084
rect 18288 27072 18294 27124
rect 19978 27112 19984 27124
rect 19812 27084 19984 27112
rect 14645 27047 14703 27053
rect 8772 27016 11836 27044
rect 2547 26948 2774 26976
rect 2547 26945 2559 26948
rect 2501 26939 2559 26945
rect 3142 26936 3148 26988
rect 3200 26976 3206 26988
rect 3309 26979 3367 26985
rect 3309 26976 3321 26979
rect 3200 26948 3321 26976
rect 3200 26936 3206 26948
rect 3309 26945 3321 26948
rect 3355 26945 3367 26979
rect 3309 26939 3367 26945
rect 5353 26979 5411 26985
rect 5353 26945 5365 26979
rect 5399 26976 5411 26979
rect 5718 26976 5724 26988
rect 5399 26948 5724 26976
rect 5399 26945 5411 26948
rect 5353 26939 5411 26945
rect 5718 26936 5724 26948
rect 5776 26936 5782 26988
rect 9217 26979 9275 26985
rect 9217 26945 9229 26979
rect 9263 26945 9275 26979
rect 9217 26939 9275 26945
rect 1765 26911 1823 26917
rect 1765 26877 1777 26911
rect 1811 26908 1823 26911
rect 1811 26880 2774 26908
rect 1811 26877 1823 26880
rect 1765 26871 1823 26877
rect 2746 26772 2774 26880
rect 2958 26868 2964 26920
rect 3016 26908 3022 26920
rect 3053 26911 3111 26917
rect 3053 26908 3065 26911
rect 3016 26880 3065 26908
rect 3016 26868 3022 26880
rect 3053 26877 3065 26880
rect 3099 26877 3111 26911
rect 3053 26871 3111 26877
rect 6270 26868 6276 26920
rect 6328 26908 6334 26920
rect 6365 26911 6423 26917
rect 6365 26908 6377 26911
rect 6328 26880 6377 26908
rect 6328 26868 6334 26880
rect 6365 26877 6377 26880
rect 6411 26877 6423 26911
rect 9232 26908 9260 26939
rect 6365 26871 6423 26877
rect 7668 26880 9260 26908
rect 4356 26812 6500 26840
rect 4356 26772 4384 26812
rect 2746 26744 4384 26772
rect 4433 26775 4491 26781
rect 4433 26741 4445 26775
rect 4479 26772 4491 26775
rect 4706 26772 4712 26784
rect 4479 26744 4712 26772
rect 4479 26741 4491 26744
rect 4433 26735 4491 26741
rect 4706 26732 4712 26744
rect 4764 26732 4770 26784
rect 6472 26772 6500 26812
rect 7668 26784 7696 26880
rect 7926 26800 7932 26852
rect 7984 26840 7990 26852
rect 8113 26843 8171 26849
rect 8113 26840 8125 26843
rect 7984 26812 8125 26840
rect 7984 26800 7990 26812
rect 8113 26809 8125 26812
rect 8159 26809 8171 26843
rect 8113 26803 8171 26809
rect 7650 26772 7656 26784
rect 6472 26744 7656 26772
rect 7650 26732 7656 26744
rect 7708 26732 7714 26784
rect 9324 26781 9352 27016
rect 9401 26979 9459 26985
rect 9401 26945 9413 26979
rect 9447 26976 9459 26979
rect 10042 26976 10048 26988
rect 9447 26948 10048 26976
rect 9447 26945 9459 26948
rect 9401 26939 9459 26945
rect 10042 26936 10048 26948
rect 10100 26936 10106 26988
rect 11808 26985 11836 27016
rect 14645 27013 14657 27047
rect 14691 27044 14703 27047
rect 14734 27044 14740 27056
rect 14691 27016 14740 27044
rect 14691 27013 14703 27016
rect 14645 27007 14703 27013
rect 14734 27004 14740 27016
rect 14792 27004 14798 27056
rect 17494 27004 17500 27056
rect 17552 27044 17558 27056
rect 17926 27047 17984 27053
rect 17926 27044 17938 27047
rect 17552 27016 17938 27044
rect 17552 27004 17558 27016
rect 17926 27013 17938 27016
rect 17972 27013 17984 27047
rect 17926 27007 17984 27013
rect 11793 26979 11851 26985
rect 11793 26945 11805 26979
rect 11839 26976 11851 26979
rect 13679 26979 13737 26985
rect 13679 26976 13691 26979
rect 11839 26948 12434 26976
rect 11839 26945 11851 26948
rect 11793 26939 11851 26945
rect 10060 26908 10088 26936
rect 11517 26911 11575 26917
rect 11517 26908 11529 26911
rect 10060 26880 11529 26908
rect 11517 26877 11529 26880
rect 11563 26908 11575 26911
rect 12253 26911 12311 26917
rect 12253 26908 12265 26911
rect 11563 26880 12265 26908
rect 11563 26877 11575 26880
rect 11517 26871 11575 26877
rect 12253 26877 12265 26880
rect 12299 26877 12311 26911
rect 12253 26871 12311 26877
rect 9585 26843 9643 26849
rect 9585 26809 9597 26843
rect 9631 26840 9643 26843
rect 12158 26840 12164 26852
rect 9631 26812 12164 26840
rect 9631 26809 9643 26812
rect 9585 26803 9643 26809
rect 12158 26800 12164 26812
rect 12216 26800 12222 26852
rect 12406 26840 12434 26948
rect 13004 26948 13691 26976
rect 13004 26920 13032 26948
rect 13679 26945 13691 26948
rect 13725 26945 13737 26979
rect 13814 26976 13820 26988
rect 13775 26948 13820 26976
rect 13679 26939 13737 26945
rect 13814 26936 13820 26948
rect 13872 26936 13878 26988
rect 13906 26936 13912 26988
rect 13964 26976 13970 26988
rect 13964 26948 14009 26976
rect 13964 26936 13970 26948
rect 14090 26936 14096 26988
rect 14148 26976 14154 26988
rect 17678 26976 17684 26988
rect 14148 26948 14193 26976
rect 17639 26948 17684 26976
rect 14148 26936 14154 26948
rect 17678 26936 17684 26948
rect 17736 26936 17742 26988
rect 19812 26985 19840 27084
rect 19978 27072 19984 27084
rect 20036 27072 20042 27124
rect 20901 27115 20959 27121
rect 20901 27112 20913 27115
rect 20088 27084 20913 27112
rect 20088 27044 20116 27084
rect 20901 27081 20913 27084
rect 20947 27081 20959 27115
rect 20901 27075 20959 27081
rect 25130 27072 25136 27124
rect 25188 27112 25194 27124
rect 25777 27115 25835 27121
rect 25777 27112 25789 27115
rect 25188 27084 25789 27112
rect 25188 27072 25194 27084
rect 25777 27081 25789 27084
rect 25823 27081 25835 27115
rect 25777 27075 25835 27081
rect 26970 27072 26976 27124
rect 27028 27112 27034 27124
rect 27065 27115 27123 27121
rect 27065 27112 27077 27115
rect 27028 27084 27077 27112
rect 27028 27072 27034 27084
rect 27065 27081 27077 27084
rect 27111 27081 27123 27115
rect 27065 27075 27123 27081
rect 19996 27016 20116 27044
rect 20441 27047 20499 27053
rect 19996 26985 20024 27016
rect 20441 27013 20453 27047
rect 20487 27044 20499 27047
rect 23302 27047 23360 27053
rect 23302 27044 23314 27047
rect 20487 27016 23314 27044
rect 20487 27013 20499 27016
rect 20441 27007 20499 27013
rect 23302 27013 23314 27016
rect 23348 27013 23360 27047
rect 23302 27007 23360 27013
rect 23566 27004 23572 27056
rect 23624 27044 23630 27056
rect 24305 27047 24363 27053
rect 24305 27044 24317 27047
rect 23624 27016 24317 27044
rect 23624 27004 23630 27016
rect 24305 27013 24317 27016
rect 24351 27013 24363 27047
rect 24305 27007 24363 27013
rect 25314 27004 25320 27056
rect 25372 27004 25378 27056
rect 19797 26979 19855 26985
rect 19797 26945 19809 26979
rect 19843 26945 19855 26979
rect 19797 26939 19855 26945
rect 19981 26979 20039 26985
rect 19981 26945 19993 26979
rect 20027 26945 20039 26979
rect 19981 26939 20039 26945
rect 20073 26979 20131 26985
rect 20073 26945 20085 26979
rect 20119 26945 20131 26979
rect 20073 26939 20131 26945
rect 12986 26908 12992 26920
rect 12947 26880 12992 26908
rect 12986 26868 12992 26880
rect 13044 26868 13050 26920
rect 13078 26868 13084 26920
rect 13136 26908 13142 26920
rect 14550 26908 14556 26920
rect 13136 26880 14556 26908
rect 13136 26868 13142 26880
rect 14550 26868 14556 26880
rect 14608 26908 14614 26920
rect 17126 26908 17132 26920
rect 14608 26880 17132 26908
rect 14608 26868 14614 26880
rect 17126 26868 17132 26880
rect 17184 26868 17190 26920
rect 20088 26908 20116 26939
rect 20162 26936 20168 26988
rect 20220 26976 20226 26988
rect 21085 26979 21143 26985
rect 20220 26948 20265 26976
rect 20220 26936 20226 26948
rect 21085 26945 21097 26979
rect 21131 26945 21143 26979
rect 21266 26976 21272 26988
rect 21227 26948 21272 26976
rect 21085 26939 21143 26945
rect 20346 26908 20352 26920
rect 20088 26880 20352 26908
rect 20346 26868 20352 26880
rect 20404 26868 20410 26920
rect 21100 26908 21128 26939
rect 21266 26936 21272 26948
rect 21324 26936 21330 26988
rect 25774 26936 25780 26988
rect 25832 26976 25838 26988
rect 26973 26979 27031 26985
rect 26973 26976 26985 26979
rect 25832 26948 26985 26976
rect 25832 26936 25838 26948
rect 26973 26945 26985 26948
rect 27019 26976 27031 26979
rect 27617 26979 27675 26985
rect 27617 26976 27629 26979
rect 27019 26948 27629 26976
rect 27019 26945 27031 26948
rect 26973 26939 27031 26945
rect 27617 26945 27629 26948
rect 27663 26945 27675 26979
rect 27617 26939 27675 26945
rect 23566 26908 23572 26920
rect 21100 26880 22094 26908
rect 23527 26880 23572 26908
rect 16298 26840 16304 26852
rect 12406 26812 16304 26840
rect 16298 26800 16304 26812
rect 16356 26800 16362 26852
rect 9309 26775 9367 26781
rect 9309 26741 9321 26775
rect 9355 26772 9367 26775
rect 10321 26775 10379 26781
rect 10321 26772 10333 26775
rect 9355 26744 10333 26772
rect 9355 26741 9367 26744
rect 9309 26735 9367 26741
rect 10321 26741 10333 26744
rect 10367 26741 10379 26775
rect 10870 26772 10876 26784
rect 10831 26744 10876 26772
rect 10321 26735 10379 26741
rect 10870 26732 10876 26744
rect 10928 26772 10934 26784
rect 11701 26775 11759 26781
rect 11701 26772 11713 26775
rect 10928 26744 11713 26772
rect 10928 26732 10934 26744
rect 11701 26741 11713 26744
rect 11747 26772 11759 26775
rect 14366 26772 14372 26784
rect 11747 26744 14372 26772
rect 11747 26741 11759 26744
rect 11701 26735 11759 26741
rect 14366 26732 14372 26744
rect 14424 26732 14430 26784
rect 18322 26732 18328 26784
rect 18380 26772 18386 26784
rect 18966 26772 18972 26784
rect 18380 26744 18972 26772
rect 18380 26732 18386 26744
rect 18966 26732 18972 26744
rect 19024 26772 19030 26784
rect 19061 26775 19119 26781
rect 19061 26772 19073 26775
rect 19024 26744 19073 26772
rect 19024 26732 19030 26744
rect 19061 26741 19073 26744
rect 19107 26741 19119 26775
rect 22066 26772 22094 26880
rect 23566 26868 23572 26880
rect 23624 26908 23630 26920
rect 24029 26911 24087 26917
rect 24029 26908 24041 26911
rect 23624 26880 24041 26908
rect 23624 26868 23630 26880
rect 24029 26877 24041 26880
rect 24075 26877 24087 26911
rect 24029 26871 24087 26877
rect 22189 26775 22247 26781
rect 22189 26772 22201 26775
rect 22066 26744 22201 26772
rect 19061 26735 19119 26741
rect 22189 26741 22201 26744
rect 22235 26772 22247 26775
rect 23750 26772 23756 26784
rect 22235 26744 23756 26772
rect 22235 26741 22247 26744
rect 22189 26735 22247 26741
rect 23750 26732 23756 26744
rect 23808 26732 23814 26784
rect 1104 26682 68816 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 65654 26682
rect 65706 26630 65718 26682
rect 65770 26630 65782 26682
rect 65834 26630 65846 26682
rect 65898 26630 65910 26682
rect 65962 26630 68816 26682
rect 1104 26608 68816 26630
rect 7098 26568 7104 26580
rect 7059 26540 7104 26568
rect 7098 26528 7104 26540
rect 7156 26528 7162 26580
rect 7190 26528 7196 26580
rect 7248 26568 7254 26580
rect 9493 26571 9551 26577
rect 9493 26568 9505 26571
rect 7248 26540 9505 26568
rect 7248 26528 7254 26540
rect 9493 26537 9505 26540
rect 9539 26568 9551 26571
rect 10870 26568 10876 26580
rect 9539 26540 10876 26568
rect 9539 26537 9551 26540
rect 9493 26531 9551 26537
rect 10870 26528 10876 26540
rect 10928 26528 10934 26580
rect 13357 26571 13415 26577
rect 13357 26537 13369 26571
rect 13403 26568 13415 26571
rect 14274 26568 14280 26580
rect 13403 26540 14280 26568
rect 13403 26537 13415 26540
rect 13357 26531 13415 26537
rect 14274 26528 14280 26540
rect 14332 26528 14338 26580
rect 17402 26568 17408 26580
rect 14384 26540 17408 26568
rect 4706 26460 4712 26512
rect 4764 26500 4770 26512
rect 7558 26500 7564 26512
rect 4764 26472 7564 26500
rect 4764 26460 4770 26472
rect 7558 26460 7564 26472
rect 7616 26460 7622 26512
rect 9582 26460 9588 26512
rect 9640 26500 9646 26512
rect 12897 26503 12955 26509
rect 12897 26500 12909 26503
rect 9640 26472 12909 26500
rect 9640 26460 9646 26472
rect 12897 26469 12909 26472
rect 12943 26469 12955 26503
rect 14384 26500 14412 26540
rect 17402 26528 17408 26540
rect 17460 26528 17466 26580
rect 21085 26571 21143 26577
rect 21085 26537 21097 26571
rect 21131 26568 21143 26571
rect 21266 26568 21272 26580
rect 21131 26540 21272 26568
rect 21131 26537 21143 26540
rect 21085 26531 21143 26537
rect 21266 26528 21272 26540
rect 21324 26528 21330 26580
rect 25225 26571 25283 26577
rect 25225 26537 25237 26571
rect 25271 26568 25283 26571
rect 25314 26568 25320 26580
rect 25271 26540 25320 26568
rect 25271 26537 25283 26540
rect 25225 26531 25283 26537
rect 25314 26528 25320 26540
rect 25372 26528 25378 26580
rect 36814 26568 36820 26580
rect 36775 26540 36820 26568
rect 36814 26528 36820 26540
rect 36872 26528 36878 26580
rect 17126 26500 17132 26512
rect 12897 26463 12955 26469
rect 13004 26472 14412 26500
rect 17087 26472 17132 26500
rect 11238 26432 11244 26444
rect 11072 26404 11244 26432
rect 7009 26367 7067 26373
rect 7009 26333 7021 26367
rect 7055 26333 7067 26367
rect 7009 26327 7067 26333
rect 5537 26299 5595 26305
rect 5537 26265 5549 26299
rect 5583 26296 5595 26299
rect 5718 26296 5724 26308
rect 5583 26268 5724 26296
rect 5583 26265 5595 26268
rect 5537 26259 5595 26265
rect 5718 26256 5724 26268
rect 5776 26296 5782 26308
rect 7024 26296 7052 26327
rect 7650 26324 7656 26376
rect 7708 26364 7714 26376
rect 9401 26367 9459 26373
rect 9401 26364 9413 26367
rect 7708 26336 9413 26364
rect 7708 26324 7714 26336
rect 9401 26333 9413 26336
rect 9447 26333 9459 26367
rect 10778 26364 10784 26376
rect 10739 26336 10784 26364
rect 9401 26327 9459 26333
rect 10778 26324 10784 26336
rect 10836 26324 10842 26376
rect 11072 26373 11100 26404
rect 11238 26392 11244 26404
rect 11296 26392 11302 26444
rect 11977 26435 12035 26441
rect 11977 26401 11989 26435
rect 12023 26432 12035 26435
rect 13004 26432 13032 26472
rect 17126 26460 17132 26472
rect 17184 26460 17190 26512
rect 12023 26404 13032 26432
rect 13096 26404 14044 26432
rect 12023 26401 12035 26404
rect 11977 26395 12035 26401
rect 10965 26367 11023 26373
rect 10965 26333 10977 26367
rect 11011 26333 11023 26367
rect 10965 26327 11023 26333
rect 11057 26367 11115 26373
rect 11057 26333 11069 26367
rect 11103 26333 11115 26367
rect 11057 26327 11115 26333
rect 11149 26367 11207 26373
rect 11149 26333 11161 26367
rect 11195 26364 11207 26367
rect 11992 26364 12020 26395
rect 12912 26376 12940 26404
rect 11195 26336 12020 26364
rect 11195 26333 11207 26336
rect 11149 26327 11207 26333
rect 7745 26299 7803 26305
rect 7745 26296 7757 26299
rect 5776 26268 7757 26296
rect 5776 26256 5782 26268
rect 7745 26265 7757 26268
rect 7791 26265 7803 26299
rect 7745 26259 7803 26265
rect 10042 26228 10048 26240
rect 10003 26200 10048 26228
rect 10042 26188 10048 26200
rect 10100 26188 10106 26240
rect 10980 26228 11008 26327
rect 12894 26324 12900 26376
rect 12952 26324 12958 26376
rect 13096 26373 13124 26404
rect 13081 26367 13139 26373
rect 13081 26333 13093 26367
rect 13127 26333 13139 26367
rect 13081 26327 13139 26333
rect 13173 26367 13231 26373
rect 13173 26333 13185 26367
rect 13219 26364 13231 26367
rect 13262 26364 13268 26376
rect 13219 26336 13268 26364
rect 13219 26333 13231 26336
rect 13173 26327 13231 26333
rect 13262 26324 13268 26336
rect 13320 26324 13326 26376
rect 12158 26256 12164 26308
rect 12216 26296 12222 26308
rect 13357 26299 13415 26305
rect 13357 26296 13369 26299
rect 12216 26268 13369 26296
rect 12216 26256 12222 26268
rect 13357 26265 13369 26268
rect 13403 26265 13415 26299
rect 14016 26296 14044 26404
rect 14090 26392 14096 26444
rect 14148 26432 14154 26444
rect 14645 26435 14703 26441
rect 14645 26432 14657 26435
rect 14148 26404 14657 26432
rect 14148 26392 14154 26404
rect 14645 26401 14657 26404
rect 14691 26401 14703 26435
rect 14645 26395 14703 26401
rect 33980 26404 35664 26432
rect 14182 26324 14188 26376
rect 14240 26364 14246 26376
rect 14921 26367 14979 26373
rect 14921 26364 14933 26367
rect 14240 26336 14933 26364
rect 14240 26324 14246 26336
rect 14921 26333 14933 26336
rect 14967 26364 14979 26367
rect 15562 26364 15568 26376
rect 14967 26336 15568 26364
rect 14967 26333 14979 26336
rect 14921 26327 14979 26333
rect 15562 26324 15568 26336
rect 15620 26324 15626 26376
rect 15749 26367 15807 26373
rect 15749 26333 15761 26367
rect 15795 26364 15807 26367
rect 16574 26364 16580 26376
rect 15795 26336 16580 26364
rect 15795 26333 15807 26336
rect 15749 26327 15807 26333
rect 16574 26324 16580 26336
rect 16632 26364 16638 26376
rect 17678 26364 17684 26376
rect 16632 26336 17684 26364
rect 16632 26324 16638 26336
rect 17678 26324 17684 26336
rect 17736 26324 17742 26376
rect 21269 26367 21327 26373
rect 21269 26333 21281 26367
rect 21315 26364 21327 26367
rect 21450 26364 21456 26376
rect 21315 26336 21456 26364
rect 21315 26333 21327 26336
rect 21269 26327 21327 26333
rect 21450 26324 21456 26336
rect 21508 26324 21514 26376
rect 25314 26364 25320 26376
rect 25275 26336 25320 26364
rect 25314 26324 25320 26336
rect 25372 26364 25378 26376
rect 25774 26364 25780 26376
rect 25372 26336 25780 26364
rect 25372 26324 25378 26336
rect 25774 26324 25780 26336
rect 25832 26324 25838 26376
rect 32214 26364 32220 26376
rect 32175 26336 32220 26364
rect 32214 26324 32220 26336
rect 32272 26324 32278 26376
rect 32398 26324 32404 26376
rect 32456 26364 32462 26376
rect 33980 26373 34008 26404
rect 32493 26367 32551 26373
rect 32493 26364 32505 26367
rect 32456 26336 32505 26364
rect 32456 26324 32462 26336
rect 32493 26333 32505 26336
rect 32539 26333 32551 26367
rect 32493 26327 32551 26333
rect 33965 26367 34023 26373
rect 33965 26333 33977 26367
rect 34011 26333 34023 26367
rect 33965 26327 34023 26333
rect 34977 26367 35035 26373
rect 34977 26333 34989 26367
rect 35023 26333 35035 26367
rect 35158 26364 35164 26376
rect 35119 26336 35164 26364
rect 34977 26327 35035 26333
rect 14016 26268 15792 26296
rect 13357 26259 13415 26265
rect 11054 26228 11060 26240
rect 10980 26200 11060 26228
rect 11054 26188 11060 26200
rect 11112 26188 11118 26240
rect 11422 26228 11428 26240
rect 11383 26200 11428 26228
rect 11422 26188 11428 26200
rect 11480 26188 11486 26240
rect 15764 26228 15792 26268
rect 15838 26256 15844 26308
rect 15896 26296 15902 26308
rect 15994 26299 16052 26305
rect 15994 26296 16006 26299
rect 15896 26268 16006 26296
rect 15896 26256 15902 26268
rect 15994 26265 16006 26268
rect 16040 26265 16052 26299
rect 17034 26296 17040 26308
rect 15994 26259 16052 26265
rect 16132 26268 17040 26296
rect 16132 26228 16160 26268
rect 17034 26256 17040 26268
rect 17092 26296 17098 26308
rect 19242 26296 19248 26308
rect 17092 26268 19248 26296
rect 17092 26256 17098 26268
rect 19242 26256 19248 26268
rect 19300 26256 19306 26308
rect 19705 26299 19763 26305
rect 19705 26265 19717 26299
rect 19751 26296 19763 26299
rect 20162 26296 20168 26308
rect 19751 26268 20168 26296
rect 19751 26265 19763 26268
rect 19705 26259 19763 26265
rect 20162 26256 20168 26268
rect 20220 26296 20226 26308
rect 20530 26296 20536 26308
rect 20220 26268 20536 26296
rect 20220 26256 20226 26268
rect 20530 26256 20536 26268
rect 20588 26256 20594 26308
rect 34992 26296 35020 26327
rect 35158 26324 35164 26336
rect 35216 26324 35222 26376
rect 35434 26296 35440 26308
rect 34992 26268 35440 26296
rect 35434 26256 35440 26268
rect 35492 26256 35498 26308
rect 35636 26296 35664 26404
rect 35802 26364 35808 26376
rect 35763 26336 35808 26364
rect 35802 26324 35808 26336
rect 35860 26324 35866 26376
rect 36078 26364 36084 26376
rect 36039 26336 36084 26364
rect 36078 26324 36084 26336
rect 36136 26324 36142 26376
rect 68094 26364 68100 26376
rect 68055 26336 68100 26364
rect 68094 26324 68100 26336
rect 68152 26324 68158 26376
rect 37734 26296 37740 26308
rect 35636 26268 37740 26296
rect 37734 26256 37740 26268
rect 37792 26256 37798 26308
rect 33226 26228 33232 26240
rect 15764 26200 16160 26228
rect 33187 26200 33232 26228
rect 33226 26188 33232 26200
rect 33284 26188 33290 26240
rect 34054 26228 34060 26240
rect 34015 26200 34060 26228
rect 34054 26188 34060 26200
rect 34112 26188 34118 26240
rect 35342 26228 35348 26240
rect 35303 26200 35348 26228
rect 35342 26188 35348 26200
rect 35400 26188 35406 26240
rect 1104 26138 68816 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 50294 26138
rect 50346 26086 50358 26138
rect 50410 26086 50422 26138
rect 50474 26086 50486 26138
rect 50538 26086 50550 26138
rect 50602 26086 68816 26138
rect 1104 26064 68816 26086
rect 3142 26024 3148 26036
rect 3103 25996 3148 26024
rect 3142 25984 3148 25996
rect 3200 25984 3206 26036
rect 3418 25984 3424 26036
rect 3476 25984 3482 26036
rect 7650 25984 7656 26036
rect 7708 26024 7714 26036
rect 7745 26027 7803 26033
rect 7745 26024 7757 26027
rect 7708 25996 7757 26024
rect 7708 25984 7714 25996
rect 7745 25993 7757 25996
rect 7791 25993 7803 26027
rect 7745 25987 7803 25993
rect 10686 25984 10692 26036
rect 10744 26024 10750 26036
rect 14182 26024 14188 26036
rect 10744 25996 14188 26024
rect 10744 25984 10750 25996
rect 14182 25984 14188 25996
rect 14240 25984 14246 26036
rect 19242 26024 19248 26036
rect 19203 25996 19248 26024
rect 19242 25984 19248 25996
rect 19300 25984 19306 26036
rect 34790 26024 34796 26036
rect 34703 25996 34796 26024
rect 34790 25984 34796 25996
rect 34848 26024 34854 26036
rect 35158 26024 35164 26036
rect 34848 25996 35164 26024
rect 34848 25984 34854 25996
rect 35158 25984 35164 25996
rect 35216 25984 35222 26036
rect 2685 25959 2743 25965
rect 2685 25925 2697 25959
rect 2731 25956 2743 25959
rect 3436 25956 3464 25984
rect 2731 25928 3464 25956
rect 6380 25928 8708 25956
rect 2731 25925 2743 25928
rect 2685 25919 2743 25925
rect 2314 25888 2320 25900
rect 2275 25860 2320 25888
rect 2314 25848 2320 25860
rect 2372 25848 2378 25900
rect 2498 25888 2504 25900
rect 2459 25860 2504 25888
rect 2498 25848 2504 25860
rect 2556 25848 2562 25900
rect 3397 25897 3403 25900
rect 3375 25891 3403 25897
rect 3375 25857 3387 25891
rect 3375 25851 3403 25857
rect 3397 25848 3403 25851
rect 3455 25848 3461 25900
rect 3494 25891 3552 25897
rect 3494 25857 3506 25891
rect 3540 25857 3552 25891
rect 3494 25851 3552 25857
rect 3509 25820 3537 25851
rect 3602 25848 3608 25900
rect 3660 25888 3666 25900
rect 3789 25891 3847 25897
rect 3660 25860 3705 25888
rect 3660 25848 3666 25860
rect 3789 25857 3801 25891
rect 3835 25857 3847 25891
rect 3789 25851 3847 25857
rect 3344 25792 3537 25820
rect 3344 25764 3372 25792
rect 3326 25712 3332 25764
rect 3384 25712 3390 25764
rect 3234 25644 3240 25696
rect 3292 25684 3298 25696
rect 3804 25684 3832 25851
rect 6270 25780 6276 25832
rect 6328 25820 6334 25832
rect 6380 25829 6408 25928
rect 6638 25897 6644 25900
rect 6632 25851 6644 25897
rect 6696 25888 6702 25900
rect 8680 25897 8708 25928
rect 11422 25916 11428 25968
rect 11480 25956 11486 25968
rect 11762 25959 11820 25965
rect 11762 25956 11774 25959
rect 11480 25928 11774 25956
rect 11480 25916 11486 25928
rect 11762 25925 11774 25928
rect 11808 25925 11820 25959
rect 11762 25919 11820 25925
rect 33226 25916 33232 25968
rect 33284 25956 33290 25968
rect 33321 25959 33379 25965
rect 33321 25956 33333 25959
rect 33284 25928 33333 25956
rect 33284 25916 33290 25928
rect 33321 25925 33333 25928
rect 33367 25925 33379 25959
rect 33321 25919 33379 25925
rect 34054 25916 34060 25968
rect 34112 25916 34118 25968
rect 8665 25891 8723 25897
rect 6696 25860 6732 25888
rect 6638 25848 6644 25851
rect 6696 25848 6702 25860
rect 8665 25857 8677 25891
rect 8711 25857 8723 25891
rect 8665 25851 8723 25857
rect 8754 25848 8760 25900
rect 8812 25888 8818 25900
rect 8921 25891 8979 25897
rect 8921 25888 8933 25891
rect 8812 25860 8933 25888
rect 8812 25848 8818 25860
rect 8921 25857 8933 25860
rect 8967 25857 8979 25891
rect 11514 25888 11520 25900
rect 11475 25860 11520 25888
rect 8921 25851 8979 25857
rect 11514 25848 11520 25860
rect 11572 25848 11578 25900
rect 15217 25891 15275 25897
rect 15217 25857 15229 25891
rect 15263 25888 15275 25891
rect 15378 25888 15384 25900
rect 15263 25860 15384 25888
rect 15263 25857 15275 25860
rect 15217 25851 15275 25857
rect 15378 25848 15384 25860
rect 15436 25848 15442 25900
rect 15473 25891 15531 25897
rect 15473 25857 15485 25891
rect 15519 25888 15531 25891
rect 16574 25888 16580 25900
rect 15519 25860 16580 25888
rect 15519 25857 15531 25860
rect 15473 25851 15531 25857
rect 16574 25848 16580 25860
rect 16632 25848 16638 25900
rect 16666 25848 16672 25900
rect 16724 25888 16730 25900
rect 16724 25860 16769 25888
rect 16724 25848 16730 25860
rect 17678 25848 17684 25900
rect 17736 25888 17742 25900
rect 17865 25891 17923 25897
rect 17865 25888 17877 25891
rect 17736 25860 17877 25888
rect 17736 25848 17742 25860
rect 17865 25857 17877 25860
rect 17911 25857 17923 25891
rect 17865 25851 17923 25857
rect 17954 25848 17960 25900
rect 18012 25888 18018 25900
rect 18121 25891 18179 25897
rect 18121 25888 18133 25891
rect 18012 25860 18133 25888
rect 18012 25848 18018 25860
rect 18121 25857 18133 25860
rect 18167 25857 18179 25891
rect 18121 25851 18179 25857
rect 20165 25891 20223 25897
rect 20165 25857 20177 25891
rect 20211 25888 20223 25891
rect 20346 25888 20352 25900
rect 20211 25860 20352 25888
rect 20211 25857 20223 25860
rect 20165 25851 20223 25857
rect 20346 25848 20352 25860
rect 20404 25848 20410 25900
rect 22462 25848 22468 25900
rect 22520 25888 22526 25900
rect 22934 25891 22992 25897
rect 22934 25888 22946 25891
rect 22520 25860 22946 25888
rect 22520 25848 22526 25860
rect 22934 25857 22946 25860
rect 22980 25857 22992 25891
rect 22934 25851 22992 25857
rect 23474 25848 23480 25900
rect 23532 25888 23538 25900
rect 23661 25891 23719 25897
rect 23661 25888 23673 25891
rect 23532 25860 23673 25888
rect 23532 25848 23538 25860
rect 23661 25857 23673 25860
rect 23707 25857 23719 25891
rect 23842 25888 23848 25900
rect 23803 25860 23848 25888
rect 23661 25851 23719 25857
rect 23842 25848 23848 25860
rect 23900 25848 23906 25900
rect 25130 25848 25136 25900
rect 25188 25888 25194 25900
rect 25297 25891 25355 25897
rect 25297 25888 25309 25891
rect 25188 25860 25309 25888
rect 25188 25848 25194 25860
rect 25297 25857 25309 25860
rect 25343 25857 25355 25891
rect 35342 25888 35348 25900
rect 35303 25860 35348 25888
rect 25297 25851 25355 25857
rect 35342 25848 35348 25860
rect 35400 25848 35406 25900
rect 6365 25823 6423 25829
rect 6365 25820 6377 25823
rect 6328 25792 6377 25820
rect 6328 25780 6334 25792
rect 6365 25789 6377 25792
rect 6411 25789 6423 25823
rect 6365 25783 6423 25789
rect 19889 25823 19947 25829
rect 19889 25789 19901 25823
rect 19935 25820 19947 25823
rect 19978 25820 19984 25832
rect 19935 25792 19984 25820
rect 19935 25789 19947 25792
rect 19889 25783 19947 25789
rect 19978 25780 19984 25792
rect 20036 25780 20042 25832
rect 23201 25823 23259 25829
rect 23201 25789 23213 25823
rect 23247 25820 23259 25823
rect 23566 25820 23572 25832
rect 23247 25792 23572 25820
rect 23247 25789 23259 25792
rect 23201 25783 23259 25789
rect 23566 25780 23572 25792
rect 23624 25820 23630 25832
rect 24762 25820 24768 25832
rect 23624 25792 24768 25820
rect 23624 25780 23630 25792
rect 24762 25780 24768 25792
rect 24820 25820 24826 25832
rect 25041 25823 25099 25829
rect 25041 25820 25053 25823
rect 24820 25792 25053 25820
rect 24820 25780 24826 25792
rect 25041 25789 25053 25792
rect 25087 25789 25099 25823
rect 33042 25820 33048 25832
rect 33003 25792 33048 25820
rect 25041 25783 25099 25789
rect 33042 25780 33048 25792
rect 33100 25780 33106 25832
rect 3878 25712 3884 25764
rect 3936 25752 3942 25764
rect 4341 25755 4399 25761
rect 4341 25752 4353 25755
rect 3936 25724 4353 25752
rect 3936 25712 3942 25724
rect 4341 25721 4353 25724
rect 4387 25752 4399 25755
rect 4982 25752 4988 25764
rect 4387 25724 4988 25752
rect 4387 25721 4399 25724
rect 4341 25715 4399 25721
rect 4982 25712 4988 25724
rect 5040 25712 5046 25764
rect 19242 25712 19248 25764
rect 19300 25752 19306 25764
rect 19300 25724 22094 25752
rect 19300 25712 19306 25724
rect 7650 25684 7656 25696
rect 3292 25656 7656 25684
rect 3292 25644 3298 25656
rect 7650 25644 7656 25656
rect 7708 25644 7714 25696
rect 10042 25684 10048 25696
rect 10003 25656 10048 25684
rect 10042 25644 10048 25656
rect 10100 25644 10106 25696
rect 12897 25687 12955 25693
rect 12897 25653 12909 25687
rect 12943 25684 12955 25687
rect 13262 25684 13268 25696
rect 12943 25656 13268 25684
rect 12943 25653 12955 25656
rect 12897 25647 12955 25653
rect 13262 25644 13268 25656
rect 13320 25644 13326 25696
rect 14093 25687 14151 25693
rect 14093 25653 14105 25687
rect 14139 25684 14151 25687
rect 14274 25684 14280 25696
rect 14139 25656 14280 25684
rect 14139 25653 14151 25656
rect 14093 25647 14151 25653
rect 14274 25644 14280 25656
rect 14332 25644 14338 25696
rect 15930 25644 15936 25696
rect 15988 25684 15994 25696
rect 16025 25687 16083 25693
rect 16025 25684 16037 25687
rect 15988 25656 16037 25684
rect 15988 25644 15994 25656
rect 16025 25653 16037 25656
rect 16071 25653 16083 25687
rect 16850 25684 16856 25696
rect 16811 25656 16856 25684
rect 16025 25647 16083 25653
rect 16850 25644 16856 25656
rect 16908 25644 16914 25696
rect 21821 25687 21879 25693
rect 21821 25653 21833 25687
rect 21867 25684 21879 25687
rect 21910 25684 21916 25696
rect 21867 25656 21916 25684
rect 21867 25653 21879 25656
rect 21821 25647 21879 25653
rect 21910 25644 21916 25656
rect 21968 25644 21974 25696
rect 22066 25684 22094 25724
rect 22278 25684 22284 25696
rect 22066 25656 22284 25684
rect 22278 25644 22284 25656
rect 22336 25644 22342 25696
rect 24029 25687 24087 25693
rect 24029 25653 24041 25687
rect 24075 25684 24087 25687
rect 24394 25684 24400 25696
rect 24075 25656 24400 25684
rect 24075 25653 24087 25656
rect 24029 25647 24087 25653
rect 24394 25644 24400 25656
rect 24452 25644 24458 25696
rect 24578 25684 24584 25696
rect 24539 25656 24584 25684
rect 24578 25644 24584 25656
rect 24636 25644 24642 25696
rect 26050 25644 26056 25696
rect 26108 25684 26114 25696
rect 26421 25687 26479 25693
rect 26421 25684 26433 25687
rect 26108 25656 26433 25684
rect 26108 25644 26114 25656
rect 26421 25653 26433 25656
rect 26467 25653 26479 25687
rect 26421 25647 26479 25653
rect 32214 25644 32220 25696
rect 32272 25684 32278 25696
rect 34698 25684 34704 25696
rect 32272 25656 34704 25684
rect 32272 25644 32278 25656
rect 34698 25644 34704 25656
rect 34756 25684 34762 25696
rect 35529 25687 35587 25693
rect 35529 25684 35541 25687
rect 34756 25656 35541 25684
rect 34756 25644 34762 25656
rect 35529 25653 35541 25656
rect 35575 25684 35587 25687
rect 35802 25684 35808 25696
rect 35575 25656 35808 25684
rect 35575 25653 35587 25656
rect 35529 25647 35587 25653
rect 35802 25644 35808 25656
rect 35860 25644 35866 25696
rect 1104 25594 68816 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 65654 25594
rect 65706 25542 65718 25594
rect 65770 25542 65782 25594
rect 65834 25542 65846 25594
rect 65898 25542 65910 25594
rect 65962 25542 68816 25594
rect 1104 25520 68816 25542
rect 2498 25440 2504 25492
rect 2556 25480 2562 25492
rect 2556 25452 2774 25480
rect 2556 25440 2562 25452
rect 2746 25344 2774 25452
rect 3326 25440 3332 25492
rect 3384 25480 3390 25492
rect 6549 25483 6607 25489
rect 3384 25452 6500 25480
rect 3384 25440 3390 25452
rect 2869 25347 2927 25353
rect 2869 25344 2881 25347
rect 2746 25316 2881 25344
rect 2869 25313 2881 25316
rect 2915 25344 2927 25347
rect 6472 25344 6500 25452
rect 6549 25449 6561 25483
rect 6595 25480 6607 25483
rect 6638 25480 6644 25492
rect 6595 25452 6644 25480
rect 6595 25449 6607 25452
rect 6549 25443 6607 25449
rect 6638 25440 6644 25452
rect 6696 25440 6702 25492
rect 8389 25483 8447 25489
rect 8389 25449 8401 25483
rect 8435 25480 8447 25483
rect 8754 25480 8760 25492
rect 8435 25452 8760 25480
rect 8435 25449 8447 25452
rect 8389 25443 8447 25449
rect 8754 25440 8760 25452
rect 8812 25440 8818 25492
rect 15378 25440 15384 25492
rect 15436 25480 15442 25492
rect 16209 25483 16267 25489
rect 16209 25480 16221 25483
rect 15436 25452 16221 25480
rect 15436 25440 15442 25452
rect 16209 25449 16221 25452
rect 16255 25449 16267 25483
rect 16209 25443 16267 25449
rect 17773 25483 17831 25489
rect 17773 25449 17785 25483
rect 17819 25480 17831 25483
rect 17954 25480 17960 25492
rect 17819 25452 17960 25480
rect 17819 25449 17831 25452
rect 17773 25443 17831 25449
rect 17954 25440 17960 25452
rect 18012 25440 18018 25492
rect 23842 25440 23848 25492
rect 23900 25480 23906 25492
rect 25130 25480 25136 25492
rect 23900 25452 24900 25480
rect 25091 25452 25136 25480
rect 23900 25440 23906 25452
rect 10778 25372 10784 25424
rect 10836 25412 10842 25424
rect 10836 25384 15608 25412
rect 10836 25372 10842 25384
rect 11238 25344 11244 25356
rect 2915 25316 4016 25344
rect 6472 25316 11244 25344
rect 2915 25313 2927 25316
rect 2869 25307 2927 25313
rect 2958 25236 2964 25288
rect 3016 25276 3022 25288
rect 3881 25279 3939 25285
rect 3881 25276 3893 25279
rect 3016 25248 3893 25276
rect 3016 25236 3022 25248
rect 3881 25245 3893 25248
rect 3927 25245 3939 25279
rect 3988 25276 4016 25316
rect 4706 25276 4712 25288
rect 3988 25248 4712 25276
rect 3881 25239 3939 25245
rect 4706 25236 4712 25248
rect 4764 25236 4770 25288
rect 6932 25285 6960 25316
rect 6825 25279 6883 25285
rect 6825 25245 6837 25279
rect 6871 25245 6883 25279
rect 6825 25239 6883 25245
rect 6917 25279 6975 25285
rect 6917 25245 6929 25279
rect 6963 25245 6975 25279
rect 6917 25239 6975 25245
rect 4154 25217 4160 25220
rect 4148 25171 4160 25217
rect 4212 25208 4218 25220
rect 4212 25180 4248 25208
rect 4154 25168 4160 25171
rect 4212 25168 4218 25180
rect 6840 25152 6868 25239
rect 7006 25236 7012 25288
rect 7064 25273 7070 25288
rect 7193 25279 7251 25285
rect 7064 25245 7106 25273
rect 7193 25245 7205 25279
rect 7239 25276 7251 25279
rect 7466 25276 7472 25288
rect 7239 25248 7472 25276
rect 7239 25245 7251 25248
rect 7064 25236 7070 25245
rect 7193 25239 7251 25245
rect 7466 25236 7472 25248
rect 7524 25236 7530 25288
rect 7650 25236 7656 25288
rect 7708 25276 7714 25288
rect 7745 25279 7803 25285
rect 7745 25276 7757 25279
rect 7708 25248 7757 25276
rect 7708 25236 7714 25248
rect 7745 25245 7757 25248
rect 7791 25245 7803 25279
rect 7926 25276 7932 25288
rect 7887 25248 7932 25276
rect 7745 25239 7803 25245
rect 7760 25208 7788 25239
rect 7926 25236 7932 25248
rect 7984 25236 7990 25288
rect 8036 25285 8064 25316
rect 11238 25304 11244 25316
rect 11296 25344 11302 25356
rect 12897 25347 12955 25353
rect 12897 25344 12909 25347
rect 11296 25316 12909 25344
rect 11296 25304 11302 25316
rect 12897 25313 12909 25316
rect 12943 25313 12955 25347
rect 12897 25307 12955 25313
rect 13173 25347 13231 25353
rect 13173 25313 13185 25347
rect 13219 25344 13231 25347
rect 13219 25316 14964 25344
rect 13219 25313 13231 25316
rect 13173 25307 13231 25313
rect 14936 25288 14964 25316
rect 8021 25279 8079 25285
rect 8021 25245 8033 25279
rect 8067 25245 8079 25279
rect 8021 25239 8079 25245
rect 8110 25236 8116 25288
rect 8168 25276 8174 25288
rect 9769 25279 9827 25285
rect 8168 25248 8213 25276
rect 8168 25236 8174 25248
rect 9769 25245 9781 25279
rect 9815 25276 9827 25279
rect 10134 25276 10140 25288
rect 9815 25248 10140 25276
rect 9815 25245 9827 25248
rect 9769 25239 9827 25245
rect 10134 25236 10140 25248
rect 10192 25276 10198 25288
rect 10686 25276 10692 25288
rect 10192 25248 10692 25276
rect 10192 25236 10198 25248
rect 10686 25236 10692 25248
rect 10744 25236 10750 25288
rect 10965 25279 11023 25285
rect 10965 25245 10977 25279
rect 11011 25245 11023 25279
rect 10965 25239 11023 25245
rect 14829 25279 14887 25285
rect 14829 25245 14841 25279
rect 14875 25245 14887 25279
rect 14829 25239 14887 25245
rect 10778 25208 10784 25220
rect 7760 25180 10784 25208
rect 10778 25168 10784 25180
rect 10836 25208 10842 25220
rect 10980 25208 11008 25239
rect 10836 25180 11008 25208
rect 14844 25208 14872 25239
rect 14918 25236 14924 25288
rect 14976 25276 14982 25288
rect 15580 25285 15608 25384
rect 24670 25372 24676 25424
rect 24728 25412 24734 25424
rect 24872 25412 24900 25452
rect 25130 25440 25136 25452
rect 25188 25440 25194 25492
rect 35529 25483 35587 25489
rect 35529 25449 35541 25483
rect 35575 25480 35587 25483
rect 36078 25480 36084 25492
rect 35575 25452 36084 25480
rect 35575 25449 35587 25452
rect 35529 25443 35587 25449
rect 26513 25415 26571 25421
rect 26513 25412 26525 25415
rect 24728 25384 24808 25412
rect 24872 25384 26525 25412
rect 24728 25372 24734 25384
rect 15654 25304 15660 25356
rect 15712 25344 15718 25356
rect 15712 25316 17448 25344
rect 15712 25304 15718 25316
rect 15856 25285 15884 25316
rect 15105 25279 15163 25285
rect 15105 25276 15117 25279
rect 14976 25248 15117 25276
rect 14976 25236 14982 25248
rect 15105 25245 15117 25248
rect 15151 25245 15163 25279
rect 15105 25239 15163 25245
rect 15565 25279 15623 25285
rect 15565 25245 15577 25279
rect 15611 25245 15623 25279
rect 15565 25239 15623 25245
rect 15749 25279 15807 25285
rect 15749 25245 15761 25279
rect 15795 25245 15807 25279
rect 15749 25239 15807 25245
rect 15841 25279 15899 25285
rect 15841 25245 15853 25279
rect 15887 25245 15899 25279
rect 15841 25239 15899 25245
rect 15286 25208 15292 25220
rect 14844 25180 15292 25208
rect 10836 25168 10842 25180
rect 15286 25168 15292 25180
rect 15344 25168 15350 25220
rect 5258 25100 5264 25152
rect 5316 25140 5322 25152
rect 5994 25140 6000 25152
rect 5316 25112 5361 25140
rect 5955 25112 6000 25140
rect 5316 25100 5322 25112
rect 5994 25100 6000 25112
rect 6052 25100 6058 25152
rect 6822 25100 6828 25152
rect 6880 25100 6886 25152
rect 7466 25100 7472 25152
rect 7524 25140 7530 25152
rect 8294 25140 8300 25152
rect 7524 25112 8300 25140
rect 7524 25100 7530 25112
rect 8294 25100 8300 25112
rect 8352 25140 8358 25152
rect 9539 25143 9597 25149
rect 9539 25140 9551 25143
rect 8352 25112 9551 25140
rect 8352 25100 8358 25112
rect 9539 25109 9551 25112
rect 9585 25109 9597 25143
rect 9539 25103 9597 25109
rect 13814 25100 13820 25152
rect 13872 25140 13878 25152
rect 15764 25140 15792 25239
rect 15930 25236 15936 25288
rect 15988 25276 15994 25288
rect 17126 25276 17132 25288
rect 15988 25248 16033 25276
rect 17087 25248 17132 25276
rect 15988 25236 15994 25248
rect 17126 25236 17132 25248
rect 17184 25236 17190 25288
rect 17310 25276 17316 25288
rect 17271 25248 17316 25276
rect 17310 25236 17316 25248
rect 17368 25236 17374 25288
rect 17420 25285 17448 25316
rect 19978 25304 19984 25356
rect 20036 25344 20042 25356
rect 20993 25347 21051 25353
rect 20993 25344 21005 25347
rect 20036 25316 21005 25344
rect 20036 25304 20042 25316
rect 20993 25313 21005 25316
rect 21039 25313 21051 25347
rect 20993 25307 21051 25313
rect 23845 25347 23903 25353
rect 23845 25313 23857 25347
rect 23891 25344 23903 25347
rect 23891 25316 24716 25344
rect 23891 25313 23903 25316
rect 23845 25307 23903 25313
rect 17405 25279 17463 25285
rect 17405 25245 17417 25279
rect 17451 25245 17463 25279
rect 17405 25239 17463 25245
rect 17497 25279 17555 25285
rect 17497 25245 17509 25279
rect 17543 25276 17555 25279
rect 20714 25276 20720 25288
rect 17543 25248 18368 25276
rect 20675 25248 20720 25276
rect 17543 25245 17555 25248
rect 17497 25239 17555 25245
rect 18340 25149 18368 25248
rect 20714 25236 20720 25248
rect 20772 25236 20778 25288
rect 21450 25236 21456 25288
rect 21508 25276 21514 25288
rect 21729 25279 21787 25285
rect 21729 25276 21741 25279
rect 21508 25248 21741 25276
rect 21508 25236 21514 25248
rect 21729 25245 21741 25248
rect 21775 25245 21787 25279
rect 21729 25239 21787 25245
rect 24210 25236 24216 25288
rect 24268 25276 24274 25288
rect 24688 25285 24716 25316
rect 24780 25285 24808 25384
rect 26513 25381 26525 25384
rect 26559 25381 26571 25415
rect 26513 25375 26571 25381
rect 33413 25415 33471 25421
rect 33413 25381 33425 25415
rect 33459 25412 33471 25415
rect 34790 25412 34796 25424
rect 33459 25384 34796 25412
rect 33459 25381 33471 25384
rect 33413 25375 33471 25381
rect 34790 25372 34796 25384
rect 34848 25372 34854 25424
rect 32125 25347 32183 25353
rect 32125 25313 32137 25347
rect 32171 25344 32183 25347
rect 32214 25344 32220 25356
rect 32171 25316 32220 25344
rect 32171 25313 32183 25316
rect 32125 25307 32183 25313
rect 32214 25304 32220 25316
rect 32272 25304 32278 25356
rect 33505 25347 33563 25353
rect 33505 25313 33517 25347
rect 33551 25313 33563 25347
rect 34238 25344 34244 25356
rect 34151 25316 34244 25344
rect 33505 25307 33563 25313
rect 24489 25279 24547 25285
rect 24489 25276 24501 25279
rect 24268 25248 24501 25276
rect 24268 25236 24274 25248
rect 24489 25245 24501 25248
rect 24535 25245 24547 25279
rect 24489 25239 24547 25245
rect 24673 25279 24731 25285
rect 24673 25245 24685 25279
rect 24719 25245 24731 25279
rect 24673 25239 24731 25245
rect 24765 25279 24823 25285
rect 24765 25245 24777 25279
rect 24811 25245 24823 25279
rect 24765 25239 24823 25245
rect 24857 25279 24915 25285
rect 24857 25245 24869 25279
rect 24903 25245 24915 25279
rect 27890 25276 27896 25288
rect 27803 25248 27896 25276
rect 24857 25239 24915 25245
rect 23474 25208 23480 25220
rect 22066 25180 23480 25208
rect 13872 25112 15792 25140
rect 18325 25143 18383 25149
rect 13872 25100 13878 25112
rect 18325 25109 18337 25143
rect 18371 25140 18383 25143
rect 19334 25140 19340 25152
rect 18371 25112 19340 25140
rect 18371 25109 18383 25112
rect 18325 25103 18383 25109
rect 19334 25100 19340 25112
rect 19392 25100 19398 25152
rect 21266 25100 21272 25152
rect 21324 25140 21330 25152
rect 21545 25143 21603 25149
rect 21545 25140 21557 25143
rect 21324 25112 21557 25140
rect 21324 25100 21330 25112
rect 21545 25109 21557 25112
rect 21591 25140 21603 25143
rect 22066 25140 22094 25180
rect 23474 25168 23480 25180
rect 23532 25168 23538 25220
rect 23658 25208 23664 25220
rect 23619 25180 23664 25208
rect 23658 25168 23664 25180
rect 23716 25168 23722 25220
rect 23842 25168 23848 25220
rect 23900 25208 23906 25220
rect 24578 25208 24584 25220
rect 23900 25180 24584 25208
rect 23900 25168 23906 25180
rect 24578 25168 24584 25180
rect 24636 25208 24642 25220
rect 24872 25208 24900 25239
rect 27890 25236 27896 25248
rect 27948 25276 27954 25288
rect 28350 25276 28356 25288
rect 27948 25248 28356 25276
rect 27948 25236 27954 25248
rect 28350 25236 28356 25248
rect 28408 25236 28414 25288
rect 30650 25236 30656 25288
rect 30708 25276 30714 25288
rect 31021 25279 31079 25285
rect 31021 25276 31033 25279
rect 30708 25248 31033 25276
rect 30708 25236 30714 25248
rect 31021 25245 31033 25248
rect 31067 25245 31079 25279
rect 31021 25239 31079 25245
rect 31849 25279 31907 25285
rect 31849 25245 31861 25279
rect 31895 25245 31907 25279
rect 33520 25276 33548 25307
rect 34164 25285 34192 25316
rect 34238 25304 34244 25316
rect 34296 25344 34302 25356
rect 35544 25344 35572 25443
rect 36078 25440 36084 25452
rect 36136 25440 36142 25492
rect 34296 25316 35572 25344
rect 34296 25304 34302 25316
rect 33965 25279 34023 25285
rect 33965 25276 33977 25279
rect 33520 25248 33977 25276
rect 31849 25239 31907 25245
rect 33965 25245 33977 25248
rect 34011 25245 34023 25279
rect 33965 25239 34023 25245
rect 34149 25279 34207 25285
rect 34149 25245 34161 25279
rect 34195 25245 34207 25279
rect 35342 25276 35348 25288
rect 35303 25248 35348 25276
rect 34149 25239 34207 25245
rect 24636 25180 24900 25208
rect 24636 25168 24642 25180
rect 26234 25168 26240 25220
rect 26292 25208 26298 25220
rect 27626 25211 27684 25217
rect 27626 25208 27638 25211
rect 26292 25180 27638 25208
rect 26292 25168 26298 25180
rect 27626 25177 27638 25180
rect 27672 25177 27684 25211
rect 27626 25171 27684 25177
rect 22554 25140 22560 25152
rect 21591 25112 22094 25140
rect 22515 25112 22560 25140
rect 21591 25109 21603 25112
rect 21545 25103 21603 25109
rect 22554 25100 22560 25112
rect 22612 25100 22618 25152
rect 31864 25140 31892 25239
rect 35342 25236 35348 25248
rect 35400 25236 35406 25288
rect 35894 25236 35900 25288
rect 35952 25276 35958 25288
rect 36449 25279 36507 25285
rect 36449 25276 36461 25279
rect 35952 25248 36461 25276
rect 35952 25236 35958 25248
rect 36449 25245 36461 25248
rect 36495 25245 36507 25279
rect 36449 25239 36507 25245
rect 33045 25211 33103 25217
rect 33045 25177 33057 25211
rect 33091 25208 33103 25211
rect 33502 25208 33508 25220
rect 33091 25180 33508 25208
rect 33091 25177 33103 25180
rect 33045 25171 33103 25177
rect 33502 25168 33508 25180
rect 33560 25168 33566 25220
rect 36722 25208 36728 25220
rect 36683 25180 36728 25208
rect 36722 25168 36728 25180
rect 36780 25168 36786 25220
rect 37458 25168 37464 25220
rect 37516 25168 37522 25220
rect 34057 25143 34115 25149
rect 34057 25140 34069 25143
rect 31864 25112 34069 25140
rect 34057 25109 34069 25112
rect 34103 25109 34115 25143
rect 34057 25103 34115 25109
rect 35434 25100 35440 25152
rect 35492 25140 35498 25152
rect 38197 25143 38255 25149
rect 38197 25140 38209 25143
rect 35492 25112 38209 25140
rect 35492 25100 35498 25112
rect 38197 25109 38209 25112
rect 38243 25109 38255 25143
rect 38197 25103 38255 25109
rect 1104 25050 68816 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 50294 25050
rect 50346 24998 50358 25050
rect 50410 24998 50422 25050
rect 50474 24998 50486 25050
rect 50538 24998 50550 25050
rect 50602 24998 68816 25050
rect 1104 24976 68816 24998
rect 3326 24896 3332 24948
rect 3384 24936 3390 24948
rect 7006 24936 7012 24948
rect 3384 24908 3537 24936
rect 6967 24908 7012 24936
rect 3384 24896 3390 24908
rect 2314 24828 2320 24880
rect 2372 24868 2378 24880
rect 2409 24871 2467 24877
rect 2409 24868 2421 24871
rect 2372 24840 2421 24868
rect 2372 24828 2378 24840
rect 2409 24837 2421 24840
rect 2455 24837 2467 24871
rect 2409 24831 2467 24837
rect 3509 24815 3537 24908
rect 7006 24896 7012 24908
rect 7064 24896 7070 24948
rect 7926 24896 7932 24948
rect 7984 24936 7990 24948
rect 8205 24939 8263 24945
rect 8205 24936 8217 24939
rect 7984 24908 8217 24936
rect 7984 24896 7990 24908
rect 8205 24905 8217 24908
rect 8251 24905 8263 24939
rect 8205 24899 8263 24905
rect 11900 24908 13860 24936
rect 5994 24828 6000 24880
rect 6052 24868 6058 24880
rect 8110 24868 8116 24880
rect 6052 24840 8116 24868
rect 6052 24828 6058 24840
rect 8110 24828 8116 24840
rect 8168 24828 8174 24880
rect 11900 24877 11928 24908
rect 11885 24871 11943 24877
rect 11885 24868 11897 24871
rect 8312 24840 8524 24868
rect 2593 24803 2651 24809
rect 2593 24769 2605 24803
rect 2639 24769 2651 24803
rect 3234 24800 3240 24812
rect 3195 24772 3240 24800
rect 2593 24763 2651 24769
rect 2608 24664 2636 24763
rect 3234 24760 3240 24772
rect 3292 24760 3298 24812
rect 3500 24809 3558 24815
rect 3400 24803 3458 24809
rect 3400 24800 3412 24803
rect 3344 24772 3412 24800
rect 2777 24735 2835 24741
rect 2777 24701 2789 24735
rect 2823 24732 2835 24735
rect 3344 24732 3372 24772
rect 3400 24769 3412 24772
rect 3446 24769 3458 24803
rect 3500 24775 3512 24809
rect 3546 24775 3558 24809
rect 3500 24769 3558 24775
rect 3605 24803 3663 24809
rect 3605 24769 3617 24803
rect 3651 24800 3663 24803
rect 3694 24800 3700 24812
rect 3651 24772 3700 24800
rect 3651 24769 3663 24772
rect 3400 24763 3458 24769
rect 3605 24763 3663 24769
rect 3694 24760 3700 24772
rect 3752 24760 3758 24812
rect 7190 24800 7196 24812
rect 7151 24772 7196 24800
rect 7190 24760 7196 24772
rect 7248 24760 7254 24812
rect 7377 24803 7435 24809
rect 7377 24769 7389 24803
rect 7423 24800 7435 24803
rect 8312 24800 8340 24840
rect 7423 24772 8340 24800
rect 8389 24803 8447 24809
rect 7423 24769 7435 24772
rect 7377 24763 7435 24769
rect 8389 24769 8401 24803
rect 8435 24769 8447 24803
rect 8496 24800 8524 24840
rect 9646 24840 11897 24868
rect 8573 24803 8631 24809
rect 8573 24800 8585 24803
rect 8496 24772 8585 24800
rect 8389 24763 8447 24769
rect 8573 24769 8585 24772
rect 8619 24800 8631 24803
rect 9646 24800 9674 24840
rect 11885 24837 11897 24840
rect 11931 24837 11943 24871
rect 11885 24831 11943 24837
rect 8619 24772 9674 24800
rect 11701 24803 11759 24809
rect 8619 24769 8631 24772
rect 8573 24763 8631 24769
rect 11701 24769 11713 24803
rect 11747 24769 11759 24803
rect 11701 24763 11759 24769
rect 13633 24803 13691 24809
rect 13633 24769 13645 24803
rect 13679 24800 13691 24803
rect 13832 24800 13860 24908
rect 15470 24896 15476 24948
rect 15528 24936 15534 24948
rect 15930 24936 15936 24948
rect 15528 24908 15936 24936
rect 15528 24896 15534 24908
rect 15930 24896 15936 24908
rect 15988 24896 15994 24948
rect 17310 24936 17316 24948
rect 17271 24908 17316 24936
rect 17310 24896 17316 24908
rect 17368 24896 17374 24948
rect 20438 24896 20444 24948
rect 20496 24936 20502 24948
rect 20496 24908 20576 24936
rect 20496 24896 20502 24908
rect 15286 24828 15292 24880
rect 15344 24868 15350 24880
rect 15654 24868 15660 24880
rect 15344 24840 15660 24868
rect 15344 24828 15350 24840
rect 13679 24772 13860 24800
rect 14369 24803 14427 24809
rect 13679 24769 13691 24772
rect 13633 24763 13691 24769
rect 14369 24769 14381 24803
rect 14415 24769 14427 24803
rect 14550 24800 14556 24812
rect 14511 24772 14556 24800
rect 14369 24763 14427 24769
rect 2823 24704 3372 24732
rect 3881 24735 3939 24741
rect 2823 24701 2835 24704
rect 2777 24695 2835 24701
rect 3881 24701 3893 24735
rect 3927 24732 3939 24735
rect 4154 24732 4160 24744
rect 3927 24704 4160 24732
rect 3927 24701 3939 24704
rect 3881 24695 3939 24701
rect 4154 24692 4160 24704
rect 4212 24692 4218 24744
rect 7392 24732 7420 24763
rect 5736 24704 7420 24732
rect 8404 24732 8432 24763
rect 11716 24732 11744 24763
rect 13262 24732 13268 24744
rect 8404 24704 9168 24732
rect 11716 24704 13268 24732
rect 4341 24667 4399 24673
rect 4341 24664 4353 24667
rect 2608 24636 4353 24664
rect 4341 24633 4353 24636
rect 4387 24664 4399 24667
rect 4614 24664 4620 24676
rect 4387 24636 4620 24664
rect 4387 24633 4399 24636
rect 4341 24627 4399 24633
rect 4614 24624 4620 24636
rect 4672 24664 4678 24676
rect 5258 24664 5264 24676
rect 4672 24636 5264 24664
rect 4672 24624 4678 24636
rect 5258 24624 5264 24636
rect 5316 24624 5322 24676
rect 2314 24556 2320 24608
rect 2372 24596 2378 24608
rect 5736 24596 5764 24704
rect 5813 24667 5871 24673
rect 5813 24633 5825 24667
rect 5859 24664 5871 24667
rect 7190 24664 7196 24676
rect 5859 24636 7196 24664
rect 5859 24633 5871 24636
rect 5813 24627 5871 24633
rect 7190 24624 7196 24636
rect 7248 24624 7254 24676
rect 2372 24568 5764 24596
rect 6549 24599 6607 24605
rect 2372 24556 2378 24568
rect 6549 24565 6561 24599
rect 6595 24596 6607 24599
rect 6822 24596 6828 24608
rect 6595 24568 6828 24596
rect 6595 24565 6607 24568
rect 6549 24559 6607 24565
rect 6822 24556 6828 24568
rect 6880 24596 6886 24608
rect 8662 24596 8668 24608
rect 6880 24568 8668 24596
rect 6880 24556 6886 24568
rect 8662 24556 8668 24568
rect 8720 24556 8726 24608
rect 9140 24605 9168 24704
rect 13262 24692 13268 24704
rect 13320 24692 13326 24744
rect 13909 24735 13967 24741
rect 13909 24701 13921 24735
rect 13955 24732 13967 24735
rect 13955 24704 14320 24732
rect 13955 24701 13967 24704
rect 13909 24695 13967 24701
rect 11054 24624 11060 24676
rect 11112 24664 11118 24676
rect 11517 24667 11575 24673
rect 11517 24664 11529 24667
rect 11112 24636 11529 24664
rect 11112 24624 11118 24636
rect 11517 24633 11529 24636
rect 11563 24633 11575 24667
rect 11517 24627 11575 24633
rect 9125 24599 9183 24605
rect 9125 24565 9137 24599
rect 9171 24596 9183 24599
rect 10042 24596 10048 24608
rect 9171 24568 10048 24596
rect 9171 24565 9183 24568
rect 9125 24559 9183 24565
rect 10042 24556 10048 24568
rect 10100 24596 10106 24608
rect 10962 24596 10968 24608
rect 10100 24568 10968 24596
rect 10100 24556 10106 24568
rect 10962 24556 10968 24568
rect 11020 24556 11026 24608
rect 14292 24596 14320 24704
rect 14384 24664 14412 24763
rect 14550 24760 14556 24772
rect 14608 24800 14614 24812
rect 15010 24800 15016 24812
rect 14608 24772 15016 24800
rect 14608 24760 14614 24772
rect 15010 24760 15016 24772
rect 15068 24760 15074 24812
rect 15194 24800 15200 24812
rect 15155 24772 15200 24800
rect 15194 24760 15200 24772
rect 15252 24760 15258 24812
rect 15488 24809 15516 24840
rect 15654 24828 15660 24840
rect 15712 24828 15718 24880
rect 16850 24828 16856 24880
rect 16908 24868 16914 24880
rect 16945 24871 17003 24877
rect 16945 24868 16957 24871
rect 16908 24840 16957 24868
rect 16908 24828 16914 24840
rect 16945 24837 16957 24840
rect 16991 24837 17003 24871
rect 16945 24831 17003 24837
rect 17678 24828 17684 24880
rect 17736 24868 17742 24880
rect 17736 24840 18000 24868
rect 17736 24828 17742 24840
rect 15381 24803 15439 24809
rect 15381 24769 15393 24803
rect 15427 24769 15439 24803
rect 15381 24763 15439 24769
rect 15473 24803 15531 24809
rect 15473 24769 15485 24803
rect 15519 24769 15531 24803
rect 15473 24763 15531 24769
rect 15565 24803 15623 24809
rect 15565 24769 15577 24803
rect 15611 24800 15623 24803
rect 16022 24800 16028 24812
rect 15611 24772 16028 24800
rect 15611 24769 15623 24772
rect 15565 24763 15623 24769
rect 14737 24735 14795 24741
rect 14737 24701 14749 24735
rect 14783 24732 14795 24735
rect 15396 24732 15424 24763
rect 16022 24760 16028 24772
rect 16080 24760 16086 24812
rect 17034 24760 17040 24812
rect 17092 24800 17098 24812
rect 17129 24803 17187 24809
rect 17129 24800 17141 24803
rect 17092 24772 17141 24800
rect 17092 24760 17098 24772
rect 17129 24769 17141 24772
rect 17175 24769 17187 24803
rect 17972 24800 18000 24840
rect 18322 24800 18328 24812
rect 17972 24772 18328 24800
rect 17129 24763 17187 24769
rect 18322 24760 18328 24772
rect 18380 24760 18386 24812
rect 18414 24760 18420 24812
rect 18472 24800 18478 24812
rect 18581 24803 18639 24809
rect 18581 24800 18593 24803
rect 18472 24772 18593 24800
rect 18472 24760 18478 24772
rect 18581 24769 18593 24772
rect 18627 24769 18639 24803
rect 20162 24800 20168 24812
rect 20123 24772 20168 24800
rect 18581 24763 18639 24769
rect 20162 24760 20168 24772
rect 20220 24760 20226 24812
rect 20346 24800 20352 24812
rect 20307 24772 20352 24800
rect 20346 24760 20352 24772
rect 20404 24760 20410 24812
rect 20548 24809 20576 24908
rect 24486 24896 24492 24948
rect 24544 24936 24550 24948
rect 24670 24936 24676 24948
rect 24544 24908 24676 24936
rect 24544 24896 24550 24908
rect 20714 24828 20720 24880
rect 20772 24868 20778 24880
rect 24596 24868 24624 24908
rect 24670 24896 24676 24908
rect 24728 24896 24734 24948
rect 34238 24936 34244 24948
rect 33244 24908 34244 24936
rect 33244 24868 33272 24908
rect 34238 24896 34244 24908
rect 34296 24896 34302 24948
rect 36081 24939 36139 24945
rect 36081 24905 36093 24939
rect 36127 24936 36139 24939
rect 36722 24936 36728 24948
rect 36127 24908 36728 24936
rect 36127 24905 36139 24908
rect 36081 24899 36139 24905
rect 36722 24896 36728 24908
rect 36780 24896 36786 24948
rect 34790 24868 34796 24880
rect 20772 24840 24624 24868
rect 20772 24828 20778 24840
rect 20441 24803 20499 24809
rect 20441 24769 20453 24803
rect 20487 24769 20499 24803
rect 20441 24763 20499 24769
rect 20533 24803 20591 24809
rect 20533 24769 20545 24803
rect 20579 24769 20591 24803
rect 21818 24800 21824 24812
rect 21779 24772 21824 24800
rect 20533 24763 20591 24769
rect 15838 24732 15844 24744
rect 14783 24704 15424 24732
rect 15799 24704 15844 24732
rect 14783 24701 14795 24704
rect 14737 24695 14795 24701
rect 15838 24692 15844 24704
rect 15896 24692 15902 24744
rect 15930 24692 15936 24744
rect 15988 24732 15994 24744
rect 17678 24732 17684 24744
rect 15988 24704 17684 24732
rect 15988 24692 15994 24704
rect 17052 24676 17080 24704
rect 17678 24692 17684 24704
rect 17736 24692 17742 24744
rect 20456 24732 20484 24763
rect 21818 24760 21824 24772
rect 21876 24760 21882 24812
rect 22002 24800 22008 24812
rect 21963 24772 22008 24800
rect 22002 24760 22008 24772
rect 22060 24760 22066 24812
rect 22112 24809 22140 24840
rect 22097 24803 22155 24809
rect 22097 24769 22109 24803
rect 22143 24769 22155 24803
rect 22097 24763 22155 24769
rect 22186 24760 22192 24812
rect 22244 24800 22250 24812
rect 22554 24800 22560 24812
rect 22244 24772 22560 24800
rect 22244 24760 22250 24772
rect 22554 24760 22560 24772
rect 22612 24760 22618 24812
rect 23750 24800 23756 24812
rect 23711 24772 23756 24800
rect 23750 24760 23756 24772
rect 23808 24760 23814 24812
rect 24210 24760 24216 24812
rect 24268 24800 24274 24812
rect 24305 24803 24363 24809
rect 24305 24800 24317 24803
rect 24268 24772 24317 24800
rect 24268 24760 24274 24772
rect 24305 24769 24317 24772
rect 24351 24769 24363 24803
rect 24305 24763 24363 24769
rect 24394 24760 24400 24812
rect 24452 24800 24458 24812
rect 24596 24809 24624 24840
rect 33060 24840 33272 24868
rect 33612 24840 34796 24868
rect 24489 24803 24547 24809
rect 24489 24800 24501 24803
rect 24452 24772 24501 24800
rect 24452 24760 24458 24772
rect 24489 24769 24501 24772
rect 24535 24769 24547 24803
rect 24489 24763 24547 24769
rect 24581 24803 24639 24809
rect 24581 24769 24593 24803
rect 24627 24769 24639 24803
rect 24581 24763 24639 24769
rect 24673 24803 24731 24809
rect 24673 24769 24685 24803
rect 24719 24769 24731 24803
rect 24673 24763 24731 24769
rect 20714 24732 20720 24744
rect 20456 24704 20720 24732
rect 20714 24692 20720 24704
rect 20772 24692 20778 24744
rect 20809 24735 20867 24741
rect 20809 24701 20821 24735
rect 20855 24732 20867 24735
rect 22462 24732 22468 24744
rect 20855 24704 22468 24732
rect 20855 24701 20867 24704
rect 20809 24695 20867 24701
rect 22462 24692 22468 24704
rect 22520 24692 22526 24744
rect 23661 24735 23719 24741
rect 23661 24701 23673 24735
rect 23707 24732 23719 24735
rect 23934 24732 23940 24744
rect 23707 24704 23940 24732
rect 23707 24701 23719 24704
rect 23661 24695 23719 24701
rect 23934 24692 23940 24704
rect 23992 24692 23998 24744
rect 24688 24676 24716 24763
rect 28442 24760 28448 24812
rect 28500 24800 28506 24812
rect 28609 24803 28667 24809
rect 28609 24800 28621 24803
rect 28500 24772 28621 24800
rect 28500 24760 28506 24772
rect 28609 24769 28621 24772
rect 28655 24769 28667 24803
rect 28609 24763 28667 24769
rect 32401 24803 32459 24809
rect 32401 24769 32413 24803
rect 32447 24769 32459 24803
rect 32401 24763 32459 24769
rect 32585 24803 32643 24809
rect 32585 24769 32597 24803
rect 32631 24800 32643 24803
rect 33060 24800 33088 24840
rect 32631 24772 33088 24800
rect 32631 24769 32643 24772
rect 32585 24763 32643 24769
rect 24949 24735 25007 24741
rect 24949 24701 24961 24735
rect 24995 24732 25007 24735
rect 26234 24732 26240 24744
rect 24995 24704 26240 24732
rect 24995 24701 25007 24704
rect 24949 24695 25007 24701
rect 26234 24692 26240 24704
rect 26292 24692 26298 24744
rect 28350 24732 28356 24744
rect 28311 24704 28356 24732
rect 28350 24692 28356 24704
rect 28408 24692 28414 24744
rect 32416 24732 32444 24763
rect 33134 24760 33140 24812
rect 33192 24800 33198 24812
rect 33612 24809 33640 24840
rect 34790 24828 34796 24840
rect 34848 24828 34854 24880
rect 39942 24828 39948 24880
rect 40000 24828 40006 24880
rect 33229 24803 33287 24809
rect 33229 24800 33241 24803
rect 33192 24772 33241 24800
rect 33192 24760 33198 24772
rect 33229 24769 33241 24772
rect 33275 24769 33287 24803
rect 33229 24763 33287 24769
rect 33597 24803 33655 24809
rect 33597 24769 33609 24803
rect 33643 24769 33655 24803
rect 33597 24763 33655 24769
rect 33686 24760 33692 24812
rect 33744 24800 33750 24812
rect 34149 24803 34207 24809
rect 34149 24800 34161 24803
rect 33744 24772 34161 24800
rect 33744 24760 33750 24772
rect 34149 24769 34161 24772
rect 34195 24769 34207 24803
rect 34422 24800 34428 24812
rect 34383 24772 34428 24800
rect 34149 24763 34207 24769
rect 34422 24760 34428 24772
rect 34480 24760 34486 24812
rect 34609 24803 34667 24809
rect 34609 24769 34621 24803
rect 34655 24800 34667 24803
rect 35345 24803 35403 24809
rect 35345 24800 35357 24803
rect 34655 24772 35357 24800
rect 34655 24769 34667 24772
rect 34609 24763 34667 24769
rect 35345 24769 35357 24772
rect 35391 24769 35403 24803
rect 35345 24763 35403 24769
rect 37458 24760 37464 24812
rect 37516 24800 37522 24812
rect 37645 24803 37703 24809
rect 37645 24800 37657 24803
rect 37516 24772 37657 24800
rect 37516 24760 37522 24772
rect 37645 24769 37657 24772
rect 37691 24769 37703 24803
rect 37645 24763 37703 24769
rect 37734 24760 37740 24812
rect 37792 24800 37798 24812
rect 38930 24800 38936 24812
rect 37792 24772 38936 24800
rect 37792 24760 37798 24772
rect 38930 24760 38936 24772
rect 38988 24760 38994 24812
rect 43165 24803 43223 24809
rect 43165 24769 43177 24803
rect 43211 24800 43223 24803
rect 43254 24800 43260 24812
rect 43211 24772 43260 24800
rect 43211 24769 43223 24772
rect 43165 24763 43223 24769
rect 43254 24760 43260 24772
rect 43312 24760 43318 24812
rect 32674 24732 32680 24744
rect 32416 24704 32680 24732
rect 32674 24692 32680 24704
rect 32732 24692 32738 24744
rect 34698 24692 34704 24744
rect 34756 24732 34762 24744
rect 35069 24735 35127 24741
rect 35069 24732 35081 24735
rect 34756 24704 35081 24732
rect 34756 24692 34762 24704
rect 35069 24701 35081 24704
rect 35115 24701 35127 24735
rect 35069 24695 35127 24701
rect 36262 24692 36268 24744
rect 36320 24732 36326 24744
rect 37752 24732 37780 24760
rect 36320 24704 37780 24732
rect 36320 24692 36326 24704
rect 38654 24692 38660 24744
rect 38712 24732 38718 24744
rect 39025 24735 39083 24741
rect 39025 24732 39037 24735
rect 38712 24704 39037 24732
rect 38712 24692 38718 24704
rect 39025 24701 39037 24704
rect 39071 24701 39083 24735
rect 39025 24695 39083 24701
rect 39301 24735 39359 24741
rect 39301 24701 39313 24735
rect 39347 24732 39359 24735
rect 41782 24732 41788 24744
rect 39347 24704 41788 24732
rect 39347 24701 39359 24704
rect 39301 24695 39359 24701
rect 41782 24692 41788 24704
rect 41840 24692 41846 24744
rect 42886 24732 42892 24744
rect 42847 24704 42892 24732
rect 42886 24692 42892 24704
rect 42944 24692 42950 24744
rect 16206 24664 16212 24676
rect 14384 24636 16212 24664
rect 16206 24624 16212 24636
rect 16264 24624 16270 24676
rect 17034 24624 17040 24676
rect 17092 24624 17098 24676
rect 19334 24624 19340 24676
rect 19392 24664 19398 24676
rect 24670 24664 24676 24676
rect 19392 24636 24676 24664
rect 19392 24624 19398 24636
rect 24670 24624 24676 24636
rect 24728 24624 24734 24676
rect 32398 24664 32404 24676
rect 32359 24636 32404 24664
rect 32398 24624 32404 24636
rect 32456 24624 32462 24676
rect 67634 24664 67640 24676
rect 67595 24636 67640 24664
rect 67634 24624 67640 24636
rect 67692 24624 67698 24676
rect 16666 24596 16672 24608
rect 14292 24568 16672 24596
rect 16666 24556 16672 24568
rect 16724 24556 16730 24608
rect 19426 24556 19432 24608
rect 19484 24596 19490 24608
rect 19705 24599 19763 24605
rect 19705 24596 19717 24599
rect 19484 24568 19717 24596
rect 19484 24556 19490 24568
rect 19705 24565 19717 24568
rect 19751 24565 19763 24599
rect 19705 24559 19763 24565
rect 20162 24556 20168 24608
rect 20220 24596 20226 24608
rect 21818 24596 21824 24608
rect 20220 24568 21824 24596
rect 20220 24556 20226 24568
rect 21818 24556 21824 24568
rect 21876 24556 21882 24608
rect 22462 24596 22468 24608
rect 22423 24568 22468 24596
rect 22462 24556 22468 24568
rect 22520 24556 22526 24608
rect 22738 24556 22744 24608
rect 22796 24596 22802 24608
rect 23382 24596 23388 24608
rect 22796 24568 23388 24596
rect 22796 24556 22802 24568
rect 23382 24556 23388 24568
rect 23440 24556 23446 24608
rect 23658 24556 23664 24608
rect 23716 24596 23722 24608
rect 23753 24599 23811 24605
rect 23753 24596 23765 24599
rect 23716 24568 23765 24596
rect 23716 24556 23722 24568
rect 23753 24565 23765 24568
rect 23799 24596 23811 24599
rect 26050 24596 26056 24608
rect 23799 24568 26056 24596
rect 23799 24565 23811 24568
rect 23753 24559 23811 24565
rect 26050 24556 26056 24568
rect 26108 24556 26114 24608
rect 29730 24596 29736 24608
rect 29691 24568 29736 24596
rect 29730 24556 29736 24568
rect 29788 24556 29794 24608
rect 32766 24556 32772 24608
rect 32824 24596 32830 24608
rect 33045 24599 33103 24605
rect 33045 24596 33057 24599
rect 32824 24568 33057 24596
rect 32824 24556 32830 24568
rect 33045 24565 33057 24568
rect 33091 24565 33103 24599
rect 33502 24596 33508 24608
rect 33415 24568 33508 24596
rect 33045 24559 33103 24565
rect 33502 24556 33508 24568
rect 33560 24596 33566 24608
rect 35434 24596 35440 24608
rect 33560 24568 35440 24596
rect 33560 24556 33566 24568
rect 35434 24556 35440 24568
rect 35492 24556 35498 24608
rect 40773 24599 40831 24605
rect 40773 24565 40785 24599
rect 40819 24596 40831 24599
rect 41138 24596 41144 24608
rect 40819 24568 41144 24596
rect 40819 24565 40831 24568
rect 40773 24559 40831 24565
rect 41138 24556 41144 24568
rect 41196 24556 41202 24608
rect 43901 24599 43959 24605
rect 43901 24565 43913 24599
rect 43947 24596 43959 24599
rect 56318 24596 56324 24608
rect 43947 24568 56324 24596
rect 43947 24565 43959 24568
rect 43901 24559 43959 24565
rect 56318 24556 56324 24568
rect 56376 24556 56382 24608
rect 1104 24506 68816 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 65654 24506
rect 65706 24454 65718 24506
rect 65770 24454 65782 24506
rect 65834 24454 65846 24506
rect 65898 24454 65910 24506
rect 65962 24454 68816 24506
rect 1104 24432 68816 24454
rect 5626 24352 5632 24404
rect 5684 24392 5690 24404
rect 6641 24395 6699 24401
rect 6641 24392 6653 24395
rect 5684 24364 6653 24392
rect 5684 24352 5690 24364
rect 6641 24361 6653 24364
rect 6687 24361 6699 24395
rect 8018 24392 8024 24404
rect 7979 24364 8024 24392
rect 6641 24355 6699 24361
rect 8018 24352 8024 24364
rect 8076 24352 8082 24404
rect 13078 24392 13084 24404
rect 13039 24364 13084 24392
rect 13078 24352 13084 24364
rect 13136 24352 13142 24404
rect 15286 24352 15292 24404
rect 15344 24392 15350 24404
rect 15473 24395 15531 24401
rect 15473 24392 15485 24395
rect 15344 24364 15485 24392
rect 15344 24352 15350 24364
rect 15473 24361 15485 24364
rect 15519 24392 15531 24395
rect 15930 24392 15936 24404
rect 15519 24364 15936 24392
rect 15519 24361 15531 24364
rect 15473 24355 15531 24361
rect 15930 24352 15936 24364
rect 15988 24352 15994 24404
rect 16022 24352 16028 24404
rect 16080 24392 16086 24404
rect 17402 24392 17408 24404
rect 16080 24364 17408 24392
rect 16080 24352 16086 24364
rect 17402 24352 17408 24364
rect 17460 24392 17466 24404
rect 17957 24395 18015 24401
rect 17460 24364 17816 24392
rect 17460 24352 17466 24364
rect 9766 24324 9772 24336
rect 7221 24296 9772 24324
rect 2958 24216 2964 24268
rect 3016 24256 3022 24268
rect 5261 24259 5319 24265
rect 5261 24256 5273 24259
rect 3016 24228 5273 24256
rect 3016 24216 3022 24228
rect 5261 24225 5273 24228
rect 5307 24225 5319 24259
rect 5261 24219 5319 24225
rect 5276 24188 5304 24219
rect 6270 24188 6276 24200
rect 5276 24160 6276 24188
rect 6270 24148 6276 24160
rect 6328 24148 6334 24200
rect 5534 24129 5540 24132
rect 5528 24083 5540 24129
rect 5592 24120 5598 24132
rect 5592 24092 5628 24120
rect 5534 24080 5540 24083
rect 5592 24080 5598 24092
rect 3145 24055 3203 24061
rect 3145 24021 3157 24055
rect 3191 24052 3203 24055
rect 3694 24052 3700 24064
rect 3191 24024 3700 24052
rect 3191 24021 3203 24024
rect 3145 24015 3203 24021
rect 3694 24012 3700 24024
rect 3752 24052 3758 24064
rect 4709 24055 4767 24061
rect 4709 24052 4721 24055
rect 3752 24024 4721 24052
rect 3752 24012 3758 24024
rect 4709 24021 4721 24024
rect 4755 24052 4767 24055
rect 5258 24052 5264 24064
rect 4755 24024 5264 24052
rect 4755 24021 4767 24024
rect 4709 24015 4767 24021
rect 5258 24012 5264 24024
rect 5316 24052 5322 24064
rect 7221 24052 7249 24296
rect 9766 24284 9772 24296
rect 9824 24284 9830 24336
rect 15654 24284 15660 24336
rect 15712 24324 15718 24336
rect 16482 24324 16488 24336
rect 15712 24296 16488 24324
rect 15712 24284 15718 24296
rect 16482 24284 16488 24296
rect 16540 24324 16546 24336
rect 16540 24296 17632 24324
rect 16540 24284 16546 24296
rect 7300 24228 9168 24256
rect 7300 24197 7328 24228
rect 9140 24200 9168 24228
rect 11514 24216 11520 24268
rect 11572 24256 11578 24268
rect 11701 24259 11759 24265
rect 11701 24256 11713 24259
rect 11572 24228 11713 24256
rect 11572 24216 11578 24228
rect 11701 24225 11713 24228
rect 11747 24225 11759 24259
rect 11701 24219 11759 24225
rect 16853 24259 16911 24265
rect 16853 24225 16865 24259
rect 16899 24256 16911 24259
rect 16899 24228 17540 24256
rect 16899 24225 16911 24228
rect 16853 24219 16911 24225
rect 7285 24191 7343 24197
rect 7285 24157 7297 24191
rect 7331 24157 7343 24191
rect 7285 24151 7343 24157
rect 7469 24191 7527 24197
rect 7469 24157 7481 24191
rect 7515 24188 7527 24191
rect 7926 24188 7932 24200
rect 7515 24160 7932 24188
rect 7515 24157 7527 24160
rect 7469 24151 7527 24157
rect 7926 24148 7932 24160
rect 7984 24148 7990 24200
rect 8110 24188 8116 24200
rect 8071 24160 8116 24188
rect 8110 24148 8116 24160
rect 8168 24148 8174 24200
rect 8941 24191 8999 24197
rect 8941 24157 8953 24191
rect 8987 24188 8999 24191
rect 8987 24160 9076 24188
rect 8987 24157 8999 24160
rect 8941 24151 8999 24157
rect 7466 24052 7472 24064
rect 5316 24024 7249 24052
rect 7427 24024 7472 24052
rect 5316 24012 5322 24024
rect 7466 24012 7472 24024
rect 7524 24012 7530 24064
rect 8846 24012 8852 24064
rect 8904 24052 8910 24064
rect 8941 24055 8999 24061
rect 8941 24052 8953 24055
rect 8904 24024 8953 24052
rect 8904 24012 8910 24024
rect 8941 24021 8953 24024
rect 8987 24021 8999 24055
rect 9048 24052 9076 24160
rect 9122 24148 9128 24200
rect 9180 24188 9186 24200
rect 9180 24160 9225 24188
rect 9180 24148 9186 24160
rect 9582 24148 9588 24200
rect 9640 24188 9646 24200
rect 9769 24191 9827 24197
rect 9769 24188 9781 24191
rect 9640 24160 9781 24188
rect 9640 24148 9646 24160
rect 9769 24157 9781 24160
rect 9815 24157 9827 24191
rect 11716 24188 11744 24219
rect 14093 24191 14151 24197
rect 14093 24188 14105 24191
rect 11716 24160 14105 24188
rect 9769 24151 9827 24157
rect 14093 24157 14105 24160
rect 14139 24188 14151 24191
rect 14642 24188 14648 24200
rect 14139 24160 14648 24188
rect 14139 24157 14151 24160
rect 14093 24151 14151 24157
rect 14642 24148 14648 24160
rect 14700 24148 14706 24200
rect 16206 24148 16212 24200
rect 16264 24188 16270 24200
rect 16485 24191 16543 24197
rect 16485 24188 16497 24191
rect 16264 24160 16497 24188
rect 16264 24148 16270 24160
rect 16485 24157 16497 24160
rect 16531 24188 16543 24191
rect 16758 24188 16764 24200
rect 16531 24160 16764 24188
rect 16531 24157 16543 24160
rect 16485 24151 16543 24157
rect 16758 24148 16764 24160
rect 16816 24148 16822 24200
rect 17218 24148 17224 24200
rect 17276 24188 17282 24200
rect 17512 24197 17540 24228
rect 17604 24197 17632 24296
rect 17678 24284 17684 24336
rect 17736 24284 17742 24336
rect 17788 24324 17816 24364
rect 17957 24361 17969 24395
rect 18003 24392 18015 24395
rect 18414 24392 18420 24404
rect 18003 24364 18420 24392
rect 18003 24361 18015 24364
rect 17957 24355 18015 24361
rect 18414 24352 18420 24364
rect 18472 24352 18478 24404
rect 19889 24395 19947 24401
rect 19889 24361 19901 24395
rect 19935 24392 19947 24395
rect 20346 24392 20352 24404
rect 19935 24364 20352 24392
rect 19935 24361 19947 24364
rect 19889 24355 19947 24361
rect 20346 24352 20352 24364
rect 20404 24352 20410 24404
rect 20438 24352 20444 24404
rect 20496 24392 20502 24404
rect 21637 24395 21695 24401
rect 20496 24364 20541 24392
rect 20496 24352 20502 24364
rect 21637 24361 21649 24395
rect 21683 24392 21695 24395
rect 22002 24392 22008 24404
rect 21683 24364 22008 24392
rect 21683 24361 21695 24364
rect 21637 24355 21695 24361
rect 22002 24352 22008 24364
rect 22060 24352 22066 24404
rect 24489 24395 24547 24401
rect 24489 24361 24501 24395
rect 24535 24392 24547 24395
rect 24670 24392 24676 24404
rect 24535 24364 24676 24392
rect 24535 24361 24547 24364
rect 24489 24355 24547 24361
rect 24670 24352 24676 24364
rect 24728 24352 24734 24404
rect 32674 24352 32680 24404
rect 32732 24392 32738 24404
rect 32769 24395 32827 24401
rect 32769 24392 32781 24395
rect 32732 24364 32781 24392
rect 32732 24352 32738 24364
rect 32769 24361 32781 24364
rect 32815 24392 32827 24395
rect 34422 24392 34428 24404
rect 32815 24364 34428 24392
rect 32815 24361 32827 24364
rect 32769 24355 32827 24361
rect 34422 24352 34428 24364
rect 34480 24352 34486 24404
rect 35342 24392 35348 24404
rect 35303 24364 35348 24392
rect 35342 24352 35348 24364
rect 35400 24352 35406 24404
rect 39942 24392 39948 24404
rect 39903 24364 39948 24392
rect 39942 24352 39948 24364
rect 40000 24352 40006 24404
rect 41782 24392 41788 24404
rect 41743 24364 41788 24392
rect 41782 24352 41788 24364
rect 41840 24352 41846 24404
rect 43254 24392 43260 24404
rect 43215 24364 43260 24392
rect 43254 24352 43260 24364
rect 43312 24352 43318 24404
rect 20456 24324 20484 24352
rect 22186 24324 22192 24336
rect 17788 24296 20484 24324
rect 20548 24296 22192 24324
rect 17696 24256 17724 24284
rect 20070 24256 20076 24268
rect 17696 24228 20076 24256
rect 20070 24216 20076 24228
rect 20128 24216 20134 24268
rect 17313 24191 17371 24197
rect 17313 24188 17325 24191
rect 17276 24160 17325 24188
rect 17276 24148 17282 24160
rect 17313 24157 17325 24160
rect 17359 24157 17371 24191
rect 17313 24151 17371 24157
rect 17497 24191 17555 24197
rect 17497 24157 17509 24191
rect 17543 24157 17555 24191
rect 17497 24151 17555 24157
rect 17589 24191 17647 24197
rect 17589 24157 17601 24191
rect 17635 24157 17647 24191
rect 17589 24151 17647 24157
rect 17678 24148 17684 24200
rect 17736 24188 17742 24200
rect 17736 24160 17781 24188
rect 17736 24148 17742 24160
rect 17862 24148 17868 24200
rect 17920 24188 17926 24200
rect 19797 24191 19855 24197
rect 19797 24188 19809 24191
rect 17920 24160 19809 24188
rect 17920 24148 17926 24160
rect 19797 24157 19809 24160
rect 19843 24157 19855 24191
rect 19797 24151 19855 24157
rect 19978 24148 19984 24200
rect 20036 24188 20042 24200
rect 20162 24188 20168 24200
rect 20036 24160 20168 24188
rect 20036 24148 20042 24160
rect 20162 24148 20168 24160
rect 20220 24148 20226 24200
rect 9398 24080 9404 24132
rect 9456 24120 9462 24132
rect 10014 24123 10072 24129
rect 10014 24120 10026 24123
rect 9456 24092 10026 24120
rect 9456 24080 9462 24092
rect 10014 24089 10026 24092
rect 10060 24089 10072 24123
rect 10014 24083 10072 24089
rect 11790 24080 11796 24132
rect 11848 24120 11854 24132
rect 11946 24123 12004 24129
rect 11946 24120 11958 24123
rect 11848 24092 11958 24120
rect 11848 24080 11854 24092
rect 11946 24089 11958 24092
rect 11992 24089 12004 24123
rect 11946 24083 12004 24089
rect 13538 24080 13544 24132
rect 13596 24120 13602 24132
rect 14338 24123 14396 24129
rect 14338 24120 14350 24123
rect 13596 24092 14350 24120
rect 13596 24080 13602 24092
rect 14338 24089 14350 24092
rect 14384 24089 14396 24123
rect 14338 24083 14396 24089
rect 16669 24123 16727 24129
rect 16669 24089 16681 24123
rect 16715 24120 16727 24123
rect 19426 24120 19432 24132
rect 16715 24092 19432 24120
rect 16715 24089 16727 24092
rect 16669 24083 16727 24089
rect 19426 24080 19432 24092
rect 19484 24080 19490 24132
rect 9674 24052 9680 24064
rect 9048 24024 9680 24052
rect 8941 24015 8999 24021
rect 9674 24012 9680 24024
rect 9732 24012 9738 24064
rect 11146 24052 11152 24064
rect 11107 24024 11152 24052
rect 11146 24012 11152 24024
rect 11204 24012 11210 24064
rect 16574 24012 16580 24064
rect 16632 24052 16638 24064
rect 17218 24052 17224 24064
rect 16632 24024 17224 24052
rect 16632 24012 16638 24024
rect 17218 24012 17224 24024
rect 17276 24012 17282 24064
rect 17678 24012 17684 24064
rect 17736 24052 17742 24064
rect 18417 24055 18475 24061
rect 18417 24052 18429 24055
rect 17736 24024 18429 24052
rect 17736 24012 17742 24024
rect 18417 24021 18429 24024
rect 18463 24052 18475 24055
rect 20548 24052 20576 24296
rect 22186 24284 22192 24296
rect 22244 24284 22250 24336
rect 35253 24327 35311 24333
rect 35253 24293 35265 24327
rect 35299 24324 35311 24327
rect 35434 24324 35440 24336
rect 35299 24296 35440 24324
rect 35299 24293 35311 24296
rect 35253 24287 35311 24293
rect 35434 24284 35440 24296
rect 35492 24284 35498 24336
rect 20622 24216 20628 24268
rect 20680 24256 20686 24268
rect 20680 24228 22094 24256
rect 20680 24216 20686 24228
rect 21266 24188 21272 24200
rect 21227 24160 21272 24188
rect 21266 24148 21272 24160
rect 21324 24148 21330 24200
rect 21453 24123 21511 24129
rect 21453 24089 21465 24123
rect 21499 24120 21511 24123
rect 22066 24120 22094 24228
rect 34790 24216 34796 24268
rect 34848 24256 34854 24268
rect 34885 24259 34943 24265
rect 34885 24256 34897 24259
rect 34848 24228 34897 24256
rect 34848 24216 34854 24228
rect 34885 24225 34897 24228
rect 34931 24225 34943 24259
rect 34885 24219 34943 24225
rect 22462 24148 22468 24200
rect 22520 24188 22526 24200
rect 23210 24191 23268 24197
rect 23210 24188 23222 24191
rect 22520 24160 23222 24188
rect 22520 24148 22526 24160
rect 23210 24157 23222 24160
rect 23256 24157 23268 24191
rect 23210 24151 23268 24157
rect 23477 24191 23535 24197
rect 23477 24157 23489 24191
rect 23523 24188 23535 24191
rect 24762 24188 24768 24200
rect 23523 24160 24768 24188
rect 23523 24157 23535 24160
rect 23477 24151 23535 24157
rect 24762 24148 24768 24160
rect 24820 24188 24826 24200
rect 24949 24191 25007 24197
rect 24949 24188 24961 24191
rect 24820 24160 24961 24188
rect 24820 24148 24826 24160
rect 24949 24157 24961 24160
rect 24995 24188 25007 24191
rect 26789 24191 26847 24197
rect 26789 24188 26801 24191
rect 24995 24160 26801 24188
rect 24995 24157 25007 24160
rect 24949 24151 25007 24157
rect 26789 24157 26801 24160
rect 26835 24188 26847 24191
rect 28350 24188 28356 24200
rect 26835 24160 28356 24188
rect 26835 24157 26847 24160
rect 26789 24151 26847 24157
rect 28350 24148 28356 24160
rect 28408 24188 28414 24200
rect 29362 24188 29368 24200
rect 28408 24160 29368 24188
rect 28408 24148 28414 24160
rect 29362 24148 29368 24160
rect 29420 24188 29426 24200
rect 29825 24191 29883 24197
rect 29825 24188 29837 24191
rect 29420 24160 29837 24188
rect 29420 24148 29426 24160
rect 29825 24157 29837 24160
rect 29871 24157 29883 24191
rect 29825 24151 29883 24157
rect 31018 24148 31024 24200
rect 31076 24188 31082 24200
rect 32677 24191 32735 24197
rect 32677 24188 32689 24191
rect 31076 24160 32689 24188
rect 31076 24148 31082 24160
rect 32677 24157 32689 24160
rect 32723 24157 32735 24191
rect 32677 24151 32735 24157
rect 32766 24148 32772 24200
rect 32824 24188 32830 24200
rect 38654 24188 38660 24200
rect 32824 24160 32869 24188
rect 38615 24160 38660 24188
rect 32824 24148 32830 24160
rect 38654 24148 38660 24160
rect 38712 24148 38718 24200
rect 38930 24148 38936 24200
rect 38988 24188 38994 24200
rect 39853 24191 39911 24197
rect 39853 24188 39865 24191
rect 38988 24160 39865 24188
rect 38988 24148 38994 24160
rect 39853 24157 39865 24160
rect 39899 24188 39911 24191
rect 40034 24188 40040 24200
rect 39899 24160 40040 24188
rect 39899 24157 39911 24160
rect 39853 24151 39911 24157
rect 40034 24148 40040 24160
rect 40092 24148 40098 24200
rect 41138 24188 41144 24200
rect 41099 24160 41144 24188
rect 41138 24148 41144 24160
rect 41196 24148 41202 24200
rect 42518 24188 42524 24200
rect 42479 24160 42524 24188
rect 42518 24148 42524 24160
rect 42576 24148 42582 24200
rect 42797 24191 42855 24197
rect 42797 24157 42809 24191
rect 42843 24188 42855 24191
rect 42886 24188 42892 24200
rect 42843 24160 42892 24188
rect 42843 24157 42855 24160
rect 42797 24151 42855 24157
rect 42886 24148 42892 24160
rect 42944 24148 42950 24200
rect 43254 24188 43260 24200
rect 43215 24160 43260 24188
rect 43254 24148 43260 24160
rect 43312 24148 43318 24200
rect 24118 24120 24124 24132
rect 21499 24092 21772 24120
rect 22066 24092 24124 24120
rect 21499 24089 21511 24092
rect 21453 24083 21511 24089
rect 21744 24064 21772 24092
rect 24118 24080 24124 24092
rect 24176 24120 24182 24132
rect 24670 24120 24676 24132
rect 24176 24092 24676 24120
rect 24176 24080 24182 24092
rect 24670 24080 24676 24092
rect 24728 24080 24734 24132
rect 24854 24080 24860 24132
rect 24912 24120 24918 24132
rect 27062 24129 27068 24132
rect 25194 24123 25252 24129
rect 25194 24120 25206 24123
rect 24912 24092 25206 24120
rect 24912 24080 24918 24092
rect 25194 24089 25206 24092
rect 25240 24089 25252 24123
rect 25194 24083 25252 24089
rect 27056 24083 27068 24129
rect 27120 24120 27126 24132
rect 30092 24123 30150 24129
rect 27120 24092 27156 24120
rect 27062 24080 27068 24083
rect 27120 24080 27126 24092
rect 30092 24089 30104 24123
rect 30138 24120 30150 24123
rect 30282 24120 30288 24132
rect 30138 24092 30288 24120
rect 30138 24089 30150 24092
rect 30092 24083 30150 24089
rect 30282 24080 30288 24092
rect 30340 24080 30346 24132
rect 32214 24080 32220 24132
rect 32272 24120 32278 24132
rect 32493 24123 32551 24129
rect 32493 24120 32505 24123
rect 32272 24092 32505 24120
rect 32272 24080 32278 24092
rect 32493 24089 32505 24092
rect 32539 24120 32551 24123
rect 33229 24123 33287 24129
rect 33229 24120 33241 24123
rect 32539 24092 33241 24120
rect 32539 24089 32551 24092
rect 32493 24083 32551 24089
rect 33229 24089 33241 24092
rect 33275 24089 33287 24123
rect 33229 24083 33287 24089
rect 37918 24080 37924 24132
rect 37976 24120 37982 24132
rect 38390 24123 38448 24129
rect 38390 24120 38402 24123
rect 37976 24092 38402 24120
rect 37976 24080 37982 24092
rect 38390 24089 38402 24092
rect 38436 24089 38448 24123
rect 38390 24083 38448 24089
rect 18463 24024 20576 24052
rect 18463 24021 18475 24024
rect 18417 24015 18475 24021
rect 21726 24012 21732 24064
rect 21784 24052 21790 24064
rect 22097 24055 22155 24061
rect 22097 24052 22109 24055
rect 21784 24024 22109 24052
rect 21784 24012 21790 24024
rect 22097 24021 22109 24024
rect 22143 24021 22155 24055
rect 22097 24015 22155 24021
rect 25958 24012 25964 24064
rect 26016 24052 26022 24064
rect 26329 24055 26387 24061
rect 26329 24052 26341 24055
rect 26016 24024 26341 24052
rect 26016 24012 26022 24024
rect 26329 24021 26341 24024
rect 26375 24021 26387 24055
rect 26329 24015 26387 24021
rect 27798 24012 27804 24064
rect 27856 24052 27862 24064
rect 28169 24055 28227 24061
rect 28169 24052 28181 24055
rect 27856 24024 28181 24052
rect 27856 24012 27862 24024
rect 28169 24021 28181 24024
rect 28215 24021 28227 24055
rect 28169 24015 28227 24021
rect 29914 24012 29920 24064
rect 29972 24052 29978 24064
rect 31205 24055 31263 24061
rect 31205 24052 31217 24055
rect 29972 24024 31217 24052
rect 29972 24012 29978 24024
rect 31205 24021 31217 24024
rect 31251 24021 31263 24055
rect 31205 24015 31263 24021
rect 36446 24012 36452 24064
rect 36504 24052 36510 24064
rect 37277 24055 37335 24061
rect 37277 24052 37289 24055
rect 36504 24024 37289 24052
rect 36504 24012 36510 24024
rect 37277 24021 37289 24024
rect 37323 24021 37335 24055
rect 37277 24015 37335 24021
rect 41233 24055 41291 24061
rect 41233 24021 41245 24055
rect 41279 24052 41291 24055
rect 42426 24052 42432 24064
rect 41279 24024 42432 24052
rect 41279 24021 41291 24024
rect 41233 24015 41291 24021
rect 42426 24012 42432 24024
rect 42484 24012 42490 24064
rect 1104 23962 68816 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 50294 23962
rect 50346 23910 50358 23962
rect 50410 23910 50422 23962
rect 50474 23910 50486 23962
rect 50538 23910 50550 23962
rect 50602 23910 68816 23962
rect 1104 23888 68816 23910
rect 3418 23808 3424 23860
rect 3476 23848 3482 23860
rect 4338 23848 4344 23860
rect 3476 23820 4344 23848
rect 3476 23808 3482 23820
rect 4338 23808 4344 23820
rect 4396 23808 4402 23860
rect 5534 23848 5540 23860
rect 5495 23820 5540 23848
rect 5534 23808 5540 23820
rect 5592 23808 5598 23860
rect 9398 23848 9404 23860
rect 8772 23820 9168 23848
rect 9359 23820 9404 23848
rect 1857 23783 1915 23789
rect 1857 23749 1869 23783
rect 1903 23780 1915 23783
rect 3206 23783 3264 23789
rect 3206 23780 3218 23783
rect 1903 23752 3218 23780
rect 1903 23749 1915 23752
rect 1857 23743 1915 23749
rect 3206 23749 3218 23752
rect 3252 23749 3264 23783
rect 3206 23743 3264 23749
rect 7466 23740 7472 23792
rect 7524 23780 7530 23792
rect 7524 23752 8156 23780
rect 7524 23740 7530 23752
rect 2130 23712 2136 23724
rect 2091 23684 2136 23712
rect 2130 23672 2136 23684
rect 2188 23672 2194 23724
rect 2225 23715 2283 23721
rect 2225 23681 2237 23715
rect 2271 23681 2283 23715
rect 2225 23675 2283 23681
rect 2240 23644 2268 23675
rect 2314 23672 2320 23724
rect 2372 23712 2378 23724
rect 2372 23684 2417 23712
rect 2372 23672 2378 23684
rect 2498 23672 2504 23724
rect 2556 23712 2562 23724
rect 4890 23712 4896 23724
rect 2556 23684 2601 23712
rect 4851 23684 4896 23712
rect 2556 23672 2562 23684
rect 4890 23672 4896 23684
rect 4948 23672 4954 23724
rect 5074 23712 5080 23724
rect 5035 23684 5080 23712
rect 5074 23672 5080 23684
rect 5132 23672 5138 23724
rect 5172 23715 5230 23721
rect 5172 23681 5184 23715
rect 5218 23681 5230 23715
rect 5172 23675 5230 23681
rect 2682 23644 2688 23656
rect 2240 23616 2688 23644
rect 2682 23604 2688 23616
rect 2740 23604 2746 23656
rect 2958 23644 2964 23656
rect 2919 23616 2964 23644
rect 2958 23604 2964 23616
rect 3016 23604 3022 23656
rect 5184 23576 5212 23675
rect 5258 23672 5264 23724
rect 5316 23712 5322 23724
rect 5316 23684 5361 23712
rect 5316 23672 5322 23684
rect 7834 23672 7840 23724
rect 7892 23721 7898 23724
rect 8128 23721 8156 23752
rect 7892 23715 7941 23721
rect 7892 23681 7895 23715
rect 7929 23681 7941 23715
rect 7892 23675 7941 23681
rect 8021 23715 8079 23721
rect 8021 23681 8033 23715
rect 8067 23681 8079 23715
rect 8021 23675 8079 23681
rect 8113 23715 8171 23721
rect 8113 23681 8125 23715
rect 8159 23681 8171 23715
rect 8294 23712 8300 23724
rect 8255 23684 8300 23712
rect 8113 23675 8171 23681
rect 7892 23672 7898 23675
rect 8036 23644 8064 23675
rect 8294 23672 8300 23684
rect 8352 23672 8358 23724
rect 8478 23672 8484 23724
rect 8536 23712 8542 23724
rect 8772 23721 8800 23820
rect 9140 23780 9168 23820
rect 9398 23808 9404 23820
rect 9456 23808 9462 23860
rect 9674 23808 9680 23860
rect 9732 23848 9738 23860
rect 10689 23851 10747 23857
rect 10689 23848 10701 23851
rect 9732 23820 10701 23848
rect 9732 23808 9738 23820
rect 10689 23817 10701 23820
rect 10735 23817 10747 23851
rect 10689 23811 10747 23817
rect 13449 23851 13507 23857
rect 13449 23817 13461 23851
rect 13495 23848 13507 23851
rect 13814 23848 13820 23860
rect 13495 23820 13820 23848
rect 13495 23817 13507 23820
rect 13449 23811 13507 23817
rect 13814 23808 13820 23820
rect 13872 23808 13878 23860
rect 17865 23851 17923 23857
rect 17865 23848 17877 23851
rect 17052 23820 17877 23848
rect 9858 23780 9864 23792
rect 9140 23752 9864 23780
rect 9858 23740 9864 23752
rect 9916 23740 9922 23792
rect 16482 23740 16488 23792
rect 16540 23780 16546 23792
rect 16540 23752 16988 23780
rect 16540 23740 16546 23752
rect 8757 23715 8815 23721
rect 8757 23712 8769 23715
rect 8536 23684 8769 23712
rect 8536 23672 8542 23684
rect 8757 23681 8769 23684
rect 8803 23681 8815 23715
rect 8757 23675 8815 23681
rect 8846 23672 8852 23724
rect 8904 23712 8910 23724
rect 8941 23715 8999 23721
rect 8941 23712 8953 23715
rect 8904 23684 8953 23712
rect 8904 23672 8910 23684
rect 8941 23681 8953 23684
rect 8987 23681 8999 23715
rect 8941 23675 8999 23681
rect 9033 23672 9039 23724
rect 9091 23721 9097 23724
rect 9091 23715 9110 23721
rect 9098 23681 9110 23715
rect 9091 23675 9110 23681
rect 9171 23715 9229 23721
rect 9171 23681 9183 23715
rect 9217 23712 9229 23715
rect 10781 23715 10839 23721
rect 9217 23684 9720 23712
rect 9217 23681 9229 23684
rect 9171 23675 9229 23681
rect 9091 23672 9097 23675
rect 8036 23616 8294 23644
rect 5258 23576 5264 23588
rect 5184 23548 5264 23576
rect 5258 23536 5264 23548
rect 5316 23536 5322 23588
rect 7650 23508 7656 23520
rect 7611 23480 7656 23508
rect 7650 23468 7656 23480
rect 7708 23468 7714 23520
rect 8266 23508 8294 23616
rect 8662 23604 8668 23656
rect 8720 23644 8726 23656
rect 9186 23644 9214 23675
rect 8720 23616 9214 23644
rect 8720 23604 8726 23616
rect 9692 23576 9720 23684
rect 10781 23681 10793 23715
rect 10827 23712 10839 23715
rect 11146 23712 11152 23724
rect 10827 23684 11152 23712
rect 10827 23681 10839 23684
rect 10781 23675 10839 23681
rect 11146 23672 11152 23684
rect 11204 23672 11210 23724
rect 13633 23715 13691 23721
rect 13633 23681 13645 23715
rect 13679 23681 13691 23715
rect 13633 23675 13691 23681
rect 13817 23715 13875 23721
rect 13817 23681 13829 23715
rect 13863 23712 13875 23715
rect 16206 23712 16212 23724
rect 13863 23684 16212 23712
rect 13863 23681 13875 23684
rect 13817 23675 13875 23681
rect 9766 23604 9772 23656
rect 9824 23644 9830 23656
rect 12713 23647 12771 23653
rect 12713 23644 12725 23647
rect 9824 23616 12725 23644
rect 9824 23604 9830 23616
rect 12713 23613 12725 23616
rect 12759 23644 12771 23647
rect 12986 23644 12992 23656
rect 12759 23616 12992 23644
rect 12759 23613 12771 23616
rect 12713 23607 12771 23613
rect 12986 23604 12992 23616
rect 13044 23644 13050 23656
rect 13354 23644 13360 23656
rect 13044 23616 13360 23644
rect 13044 23604 13050 23616
rect 13354 23604 13360 23616
rect 13412 23604 13418 23656
rect 13648 23644 13676 23675
rect 16206 23672 16212 23684
rect 16264 23672 16270 23724
rect 16574 23672 16580 23724
rect 16632 23712 16638 23724
rect 16669 23715 16727 23721
rect 16669 23712 16681 23715
rect 16632 23684 16681 23712
rect 16632 23672 16638 23684
rect 16669 23681 16681 23684
rect 16715 23681 16727 23715
rect 16850 23712 16856 23724
rect 16811 23684 16856 23712
rect 16669 23675 16727 23681
rect 16850 23672 16856 23684
rect 16908 23672 16914 23724
rect 16960 23721 16988 23752
rect 17052 23721 17080 23820
rect 17865 23817 17877 23820
rect 17911 23848 17923 23851
rect 20622 23848 20628 23860
rect 17911 23820 20628 23848
rect 17911 23817 17923 23820
rect 17865 23811 17923 23817
rect 20622 23808 20628 23820
rect 20680 23808 20686 23860
rect 22370 23848 22376 23860
rect 22331 23820 22376 23848
rect 22370 23808 22376 23820
rect 22428 23808 22434 23860
rect 24854 23848 24860 23860
rect 24815 23820 24860 23848
rect 24854 23808 24860 23820
rect 24912 23808 24918 23860
rect 30098 23848 30104 23860
rect 29932 23820 30104 23848
rect 21634 23780 21640 23792
rect 18800 23752 21640 23780
rect 18800 23724 18828 23752
rect 21634 23740 21640 23752
rect 21692 23780 21698 23792
rect 21910 23780 21916 23792
rect 21692 23752 21916 23780
rect 21692 23740 21698 23752
rect 21910 23740 21916 23752
rect 21968 23740 21974 23792
rect 23385 23783 23443 23789
rect 23385 23749 23397 23783
rect 23431 23780 23443 23783
rect 23474 23780 23480 23792
rect 23431 23752 23480 23780
rect 23431 23749 23443 23752
rect 23385 23743 23443 23749
rect 23474 23740 23480 23752
rect 23532 23740 23538 23792
rect 23753 23783 23811 23789
rect 23753 23749 23765 23783
rect 23799 23780 23811 23783
rect 23799 23752 24440 23780
rect 23799 23749 23811 23752
rect 23753 23743 23811 23749
rect 16945 23715 17003 23721
rect 16945 23681 16957 23715
rect 16991 23681 17003 23715
rect 16945 23675 17003 23681
rect 17037 23715 17095 23721
rect 17037 23681 17049 23715
rect 17083 23681 17095 23715
rect 18782 23712 18788 23724
rect 18695 23684 18788 23712
rect 17037 23675 17095 23681
rect 14274 23644 14280 23656
rect 13648 23616 14280 23644
rect 14274 23604 14280 23616
rect 14332 23604 14338 23656
rect 15194 23604 15200 23656
rect 15252 23644 15258 23656
rect 15381 23647 15439 23653
rect 15381 23644 15393 23647
rect 15252 23616 15393 23644
rect 15252 23604 15258 23616
rect 15381 23613 15393 23616
rect 15427 23613 15439 23647
rect 15381 23607 15439 23613
rect 15396 23576 15424 23607
rect 15562 23604 15568 23656
rect 15620 23644 15626 23656
rect 15657 23647 15715 23653
rect 15657 23644 15669 23647
rect 15620 23616 15669 23644
rect 15620 23604 15626 23616
rect 15657 23613 15669 23616
rect 15703 23644 15715 23647
rect 15703 23616 16712 23644
rect 15703 23613 15715 23616
rect 15657 23607 15715 23613
rect 16684 23588 16712 23616
rect 16574 23576 16580 23588
rect 9692 23548 9996 23576
rect 15396 23548 16580 23576
rect 8754 23508 8760 23520
rect 8266 23480 8760 23508
rect 8754 23468 8760 23480
rect 8812 23468 8818 23520
rect 9968 23517 9996 23548
rect 16574 23536 16580 23548
rect 16632 23536 16638 23588
rect 16666 23536 16672 23588
rect 16724 23536 16730 23588
rect 16942 23536 16948 23588
rect 17000 23576 17006 23588
rect 17052 23576 17080 23675
rect 18782 23672 18788 23684
rect 18840 23672 18846 23724
rect 19334 23672 19340 23724
rect 19392 23712 19398 23724
rect 19429 23715 19487 23721
rect 19429 23712 19441 23715
rect 19392 23684 19441 23712
rect 19392 23672 19398 23684
rect 19429 23681 19441 23684
rect 19475 23681 19487 23715
rect 19429 23675 19487 23681
rect 19613 23715 19671 23721
rect 19613 23681 19625 23715
rect 19659 23681 19671 23715
rect 19613 23675 19671 23681
rect 19705 23715 19763 23721
rect 19705 23681 19717 23715
rect 19751 23681 19763 23715
rect 19705 23675 19763 23681
rect 19797 23715 19855 23721
rect 19797 23681 19809 23715
rect 19843 23712 19855 23715
rect 20622 23712 20628 23724
rect 19843 23684 20628 23712
rect 19843 23681 19855 23684
rect 19797 23675 19855 23681
rect 17678 23576 17684 23588
rect 17000 23548 17080 23576
rect 17236 23548 17684 23576
rect 17000 23536 17006 23548
rect 9953 23511 10011 23517
rect 9953 23477 9965 23511
rect 9999 23508 10011 23511
rect 12066 23508 12072 23520
rect 9999 23480 12072 23508
rect 9999 23477 10011 23480
rect 9953 23471 10011 23477
rect 12066 23468 12072 23480
rect 12124 23468 12130 23520
rect 14366 23508 14372 23520
rect 14327 23480 14372 23508
rect 14366 23468 14372 23480
rect 14424 23468 14430 23520
rect 15930 23468 15936 23520
rect 15988 23508 15994 23520
rect 17236 23508 17264 23548
rect 17678 23536 17684 23548
rect 17736 23536 17742 23588
rect 19628 23576 19656 23675
rect 19720 23644 19748 23675
rect 20622 23672 20628 23684
rect 20680 23672 20686 23724
rect 22186 23712 22192 23724
rect 22099 23684 22192 23712
rect 22186 23672 22192 23684
rect 22244 23712 22250 23724
rect 23290 23712 23296 23724
rect 22244 23684 23296 23712
rect 22244 23672 22250 23684
rect 23290 23672 23296 23684
rect 23348 23672 23354 23724
rect 23569 23715 23627 23721
rect 23569 23681 23581 23715
rect 23615 23681 23627 23715
rect 24210 23712 24216 23724
rect 24171 23684 24216 23712
rect 23569 23675 23627 23681
rect 20162 23644 20168 23656
rect 19720 23616 20168 23644
rect 20162 23604 20168 23616
rect 20220 23604 20226 23656
rect 22097 23647 22155 23653
rect 22097 23613 22109 23647
rect 22143 23644 22155 23647
rect 23584 23644 23612 23675
rect 24210 23672 24216 23684
rect 24268 23672 24274 23724
rect 24412 23721 24440 23752
rect 24397 23715 24455 23721
rect 24397 23681 24409 23715
rect 24443 23681 24455 23715
rect 24397 23675 24455 23681
rect 24486 23672 24492 23724
rect 24544 23712 24550 23724
rect 24670 23721 24676 23724
rect 24627 23715 24676 23721
rect 24544 23684 24589 23712
rect 24544 23672 24550 23684
rect 24627 23681 24639 23715
rect 24673 23681 24676 23715
rect 24627 23675 24676 23681
rect 24670 23672 24676 23675
rect 24728 23712 24734 23724
rect 25317 23715 25375 23721
rect 25317 23712 25329 23715
rect 24728 23684 25329 23712
rect 24728 23672 24734 23684
rect 25317 23681 25329 23684
rect 25363 23681 25375 23715
rect 29638 23712 29644 23724
rect 29599 23684 29644 23712
rect 25317 23675 25375 23681
rect 29638 23672 29644 23684
rect 29696 23672 29702 23724
rect 29822 23712 29828 23724
rect 29783 23684 29828 23712
rect 29822 23672 29828 23684
rect 29880 23672 29886 23724
rect 29932 23721 29960 23820
rect 30098 23808 30104 23820
rect 30156 23808 30162 23860
rect 30282 23848 30288 23860
rect 30243 23820 30288 23848
rect 30282 23808 30288 23820
rect 30340 23808 30346 23860
rect 37918 23848 37924 23860
rect 37879 23820 37924 23848
rect 37918 23808 37924 23820
rect 37976 23808 37982 23860
rect 42613 23851 42671 23857
rect 42613 23817 42625 23851
rect 42659 23848 42671 23851
rect 42794 23848 42800 23860
rect 42659 23820 42800 23848
rect 42659 23817 42671 23820
rect 42613 23811 42671 23817
rect 42794 23808 42800 23820
rect 42852 23848 42858 23860
rect 43254 23848 43260 23860
rect 42852 23820 43260 23848
rect 42852 23808 42858 23820
rect 43254 23808 43260 23820
rect 43312 23808 43318 23860
rect 30024 23752 37688 23780
rect 30024 23721 30052 23752
rect 37660 23724 37688 23752
rect 29917 23715 29975 23721
rect 29917 23681 29929 23715
rect 29963 23681 29975 23715
rect 29917 23675 29975 23681
rect 30009 23715 30067 23721
rect 30009 23681 30021 23715
rect 30055 23681 30067 23715
rect 34054 23712 34060 23724
rect 34015 23684 34060 23712
rect 30009 23675 30067 23681
rect 25958 23644 25964 23656
rect 22143 23616 25964 23644
rect 22143 23613 22155 23616
rect 22097 23607 22155 23613
rect 25958 23604 25964 23616
rect 26016 23604 26022 23656
rect 30024 23644 30052 23675
rect 34054 23672 34060 23684
rect 34112 23672 34118 23724
rect 34241 23715 34299 23721
rect 34241 23681 34253 23715
rect 34287 23712 34299 23715
rect 36265 23715 36323 23721
rect 36265 23712 36277 23715
rect 34287 23684 36277 23712
rect 34287 23681 34299 23684
rect 34241 23675 34299 23681
rect 36265 23681 36277 23684
rect 36311 23681 36323 23715
rect 36446 23712 36452 23724
rect 36407 23684 36452 23712
rect 36265 23675 36323 23681
rect 29472 23616 30052 23644
rect 23106 23576 23112 23588
rect 19628 23548 23112 23576
rect 23106 23536 23112 23548
rect 23164 23536 23170 23588
rect 29472 23520 29500 23616
rect 33870 23604 33876 23656
rect 33928 23644 33934 23656
rect 34256 23644 34284 23675
rect 36446 23672 36452 23684
rect 36504 23672 36510 23724
rect 37274 23712 37280 23724
rect 37235 23684 37280 23712
rect 37274 23672 37280 23684
rect 37332 23672 37338 23724
rect 37440 23715 37498 23721
rect 37440 23712 37452 23715
rect 37384 23684 37452 23712
rect 33928 23616 34284 23644
rect 36633 23647 36691 23653
rect 33928 23604 33934 23616
rect 36633 23613 36645 23647
rect 36679 23644 36691 23647
rect 37384 23644 37412 23684
rect 37440 23681 37452 23684
rect 37486 23681 37498 23715
rect 37440 23675 37498 23681
rect 37556 23715 37614 23721
rect 37556 23681 37568 23715
rect 37602 23681 37614 23715
rect 37556 23675 37614 23681
rect 37571 23644 37599 23675
rect 37642 23672 37648 23724
rect 37700 23712 37706 23724
rect 41693 23715 41751 23721
rect 37700 23684 37793 23712
rect 37700 23672 37706 23684
rect 41693 23681 41705 23715
rect 41739 23681 41751 23715
rect 42426 23712 42432 23724
rect 42387 23684 42432 23712
rect 41693 23675 41751 23681
rect 36679 23616 37412 23644
rect 37476 23616 37599 23644
rect 36679 23613 36691 23616
rect 36633 23607 36691 23613
rect 37476 23588 37504 23616
rect 41598 23604 41604 23656
rect 41656 23644 41662 23656
rect 41708 23644 41736 23675
rect 42426 23672 42432 23684
rect 42484 23672 42490 23724
rect 42613 23715 42671 23721
rect 42613 23681 42625 23715
rect 42659 23681 42671 23715
rect 42613 23675 42671 23681
rect 42628 23644 42656 23675
rect 41656 23616 42656 23644
rect 41656 23604 41662 23616
rect 37458 23536 37464 23588
rect 37516 23536 37522 23588
rect 15988 23480 17264 23508
rect 17313 23511 17371 23517
rect 15988 23468 15994 23480
rect 17313 23477 17325 23511
rect 17359 23508 17371 23511
rect 17586 23508 17592 23520
rect 17359 23480 17592 23508
rect 17359 23477 17371 23480
rect 17313 23471 17371 23477
rect 17586 23468 17592 23480
rect 17644 23468 17650 23520
rect 17862 23468 17868 23520
rect 17920 23508 17926 23520
rect 18877 23511 18935 23517
rect 18877 23508 18889 23511
rect 17920 23480 18889 23508
rect 17920 23468 17926 23480
rect 18877 23477 18889 23480
rect 18923 23477 18935 23511
rect 20070 23508 20076 23520
rect 20031 23480 20076 23508
rect 18877 23471 18935 23477
rect 20070 23468 20076 23480
rect 20128 23468 20134 23520
rect 21726 23468 21732 23520
rect 21784 23508 21790 23520
rect 21913 23511 21971 23517
rect 21913 23508 21925 23511
rect 21784 23480 21925 23508
rect 21784 23468 21790 23480
rect 21913 23477 21925 23480
rect 21959 23477 21971 23511
rect 21913 23471 21971 23477
rect 27985 23511 28043 23517
rect 27985 23477 27997 23511
rect 28031 23508 28043 23511
rect 28258 23508 28264 23520
rect 28031 23480 28264 23508
rect 28031 23477 28043 23480
rect 27985 23471 28043 23477
rect 28258 23468 28264 23480
rect 28316 23468 28322 23520
rect 29181 23511 29239 23517
rect 29181 23477 29193 23511
rect 29227 23508 29239 23511
rect 29454 23508 29460 23520
rect 29227 23480 29460 23508
rect 29227 23477 29239 23480
rect 29181 23471 29239 23477
rect 29454 23468 29460 23480
rect 29512 23468 29518 23520
rect 33413 23511 33471 23517
rect 33413 23477 33425 23511
rect 33459 23508 33471 23511
rect 33778 23508 33784 23520
rect 33459 23480 33784 23508
rect 33459 23477 33471 23480
rect 33413 23471 33471 23477
rect 33778 23468 33784 23480
rect 33836 23468 33842 23520
rect 33873 23511 33931 23517
rect 33873 23477 33885 23511
rect 33919 23508 33931 23511
rect 33962 23508 33968 23520
rect 33919 23480 33968 23508
rect 33919 23477 33931 23480
rect 33873 23471 33931 23477
rect 33962 23468 33968 23480
rect 34020 23468 34026 23520
rect 41690 23468 41696 23520
rect 41748 23508 41754 23520
rect 41785 23511 41843 23517
rect 41785 23508 41797 23511
rect 41748 23480 41797 23508
rect 41748 23468 41754 23480
rect 41785 23477 41797 23480
rect 41831 23477 41843 23511
rect 41785 23471 41843 23477
rect 67542 23468 67548 23520
rect 67600 23508 67606 23520
rect 67637 23511 67695 23517
rect 67637 23508 67649 23511
rect 67600 23480 67649 23508
rect 67600 23468 67606 23480
rect 67637 23477 67649 23480
rect 67683 23477 67695 23511
rect 67637 23471 67695 23477
rect 1104 23418 68816 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 65654 23418
rect 65706 23366 65718 23418
rect 65770 23366 65782 23418
rect 65834 23366 65846 23418
rect 65898 23366 65910 23418
rect 65962 23366 68816 23418
rect 1104 23344 68816 23366
rect 2133 23307 2191 23313
rect 2133 23273 2145 23307
rect 2179 23304 2191 23307
rect 2314 23304 2320 23316
rect 2179 23276 2320 23304
rect 2179 23273 2191 23276
rect 2133 23267 2191 23273
rect 2314 23264 2320 23276
rect 2372 23264 2378 23316
rect 5074 23264 5080 23316
rect 5132 23304 5138 23316
rect 5169 23307 5227 23313
rect 5169 23304 5181 23307
rect 5132 23276 5181 23304
rect 5132 23264 5138 23276
rect 5169 23273 5181 23276
rect 5215 23273 5227 23307
rect 5626 23304 5632 23316
rect 5587 23276 5632 23304
rect 5169 23267 5227 23273
rect 5626 23264 5632 23276
rect 5684 23264 5690 23316
rect 9030 23304 9036 23316
rect 6288 23276 9036 23304
rect 5258 23196 5264 23248
rect 5316 23236 5322 23248
rect 6288 23236 6316 23276
rect 9030 23264 9036 23276
rect 9088 23304 9094 23316
rect 11790 23304 11796 23316
rect 9088 23276 9260 23304
rect 11751 23276 11796 23304
rect 9088 23264 9094 23276
rect 5316 23208 6316 23236
rect 5316 23196 5322 23208
rect 6270 23168 6276 23180
rect 6231 23140 6276 23168
rect 6270 23128 6276 23140
rect 6328 23128 6334 23180
rect 8938 23168 8944 23180
rect 8899 23140 8944 23168
rect 8938 23128 8944 23140
rect 8996 23168 9002 23180
rect 9122 23168 9128 23180
rect 8996 23140 9128 23168
rect 8996 23128 9002 23140
rect 9122 23128 9128 23140
rect 9180 23128 9186 23180
rect 9232 23177 9260 23276
rect 11790 23264 11796 23276
rect 11848 23264 11854 23316
rect 13538 23304 13544 23316
rect 13499 23276 13544 23304
rect 13538 23264 13544 23276
rect 13596 23264 13602 23316
rect 16577 23307 16635 23313
rect 16577 23273 16589 23307
rect 16623 23304 16635 23307
rect 16850 23304 16856 23316
rect 16623 23276 16856 23304
rect 16623 23273 16635 23276
rect 16577 23267 16635 23273
rect 16850 23264 16856 23276
rect 16908 23264 16914 23316
rect 19334 23304 19340 23316
rect 16960 23276 19340 23304
rect 9217 23171 9275 23177
rect 9217 23137 9229 23171
rect 9263 23137 9275 23171
rect 12342 23168 12348 23180
rect 9217 23131 9275 23137
rect 12176 23140 12348 23168
rect 2317 23103 2375 23109
rect 2317 23069 2329 23103
rect 2363 23100 2375 23103
rect 3418 23100 3424 23112
rect 2363 23072 3424 23100
rect 2363 23069 2375 23072
rect 2317 23063 2375 23069
rect 3418 23060 3424 23072
rect 3476 23060 3482 23112
rect 4801 23103 4859 23109
rect 4801 23069 4813 23103
rect 4847 23100 4859 23103
rect 6362 23100 6368 23112
rect 4847 23072 6368 23100
rect 4847 23069 4859 23072
rect 4801 23063 4859 23069
rect 2222 22992 2228 23044
rect 2280 23032 2286 23044
rect 2501 23035 2559 23041
rect 2501 23032 2513 23035
rect 2280 23004 2513 23032
rect 2280 22992 2286 23004
rect 2501 23001 2513 23004
rect 2547 23032 2559 23035
rect 4816 23032 4844 23063
rect 6362 23060 6368 23072
rect 6420 23060 6426 23112
rect 6540 23103 6598 23109
rect 6540 23069 6552 23103
rect 6586 23100 6598 23103
rect 7650 23100 7656 23112
rect 6586 23072 7656 23100
rect 6586 23069 6598 23072
rect 6540 23063 6598 23069
rect 7650 23060 7656 23072
rect 7708 23060 7714 23112
rect 8202 23060 8208 23112
rect 8260 23100 8266 23112
rect 11330 23100 11336 23112
rect 8260 23072 11336 23100
rect 8260 23060 8266 23072
rect 11330 23060 11336 23072
rect 11388 23060 11394 23112
rect 12176 23109 12204 23140
rect 12342 23128 12348 23140
rect 12400 23168 12406 23180
rect 12618 23168 12624 23180
rect 12400 23140 12624 23168
rect 12400 23128 12406 23140
rect 12618 23128 12624 23140
rect 12676 23128 12682 23180
rect 12802 23128 12808 23180
rect 12860 23168 12866 23180
rect 16960 23168 16988 23276
rect 19334 23264 19340 23276
rect 19392 23264 19398 23316
rect 21361 23307 21419 23313
rect 21361 23273 21373 23307
rect 21407 23304 21419 23307
rect 21910 23304 21916 23316
rect 21407 23276 21916 23304
rect 21407 23273 21419 23276
rect 21361 23267 21419 23273
rect 21910 23264 21916 23276
rect 21968 23304 21974 23316
rect 22186 23304 22192 23316
rect 21968 23276 22192 23304
rect 21968 23264 21974 23276
rect 22186 23264 22192 23276
rect 22244 23264 22250 23316
rect 23106 23304 23112 23316
rect 23067 23276 23112 23304
rect 23106 23264 23112 23276
rect 23164 23264 23170 23316
rect 26973 23307 27031 23313
rect 26973 23273 26985 23307
rect 27019 23304 27031 23307
rect 27062 23304 27068 23316
rect 27019 23276 27068 23304
rect 27019 23273 27031 23276
rect 26973 23267 27031 23273
rect 27062 23264 27068 23276
rect 27120 23264 27126 23316
rect 29822 23264 29828 23316
rect 29880 23304 29886 23316
rect 29917 23307 29975 23313
rect 29917 23304 29929 23307
rect 29880 23276 29929 23304
rect 29880 23264 29886 23276
rect 29917 23273 29929 23276
rect 29963 23273 29975 23307
rect 34054 23304 34060 23316
rect 29917 23267 29975 23273
rect 31726 23276 34060 23304
rect 26326 23196 26332 23248
rect 26384 23236 26390 23248
rect 31481 23239 31539 23245
rect 31481 23236 31493 23239
rect 26384 23208 31493 23236
rect 26384 23196 26390 23208
rect 31481 23205 31493 23208
rect 31527 23236 31539 23239
rect 31726 23236 31754 23276
rect 34054 23264 34060 23276
rect 34112 23264 34118 23316
rect 36078 23304 36084 23316
rect 34164 23276 36084 23304
rect 31527 23208 31754 23236
rect 31527 23205 31539 23208
rect 31481 23199 31539 23205
rect 33502 23196 33508 23248
rect 33560 23236 33566 23248
rect 34164 23236 34192 23276
rect 36078 23264 36084 23276
rect 36136 23304 36142 23316
rect 36265 23307 36323 23313
rect 36265 23304 36277 23307
rect 36136 23276 36277 23304
rect 36136 23264 36142 23276
rect 36265 23273 36277 23276
rect 36311 23273 36323 23307
rect 37642 23304 37648 23316
rect 37603 23276 37648 23304
rect 36265 23267 36323 23273
rect 37642 23264 37648 23276
rect 37700 23264 37706 23316
rect 41598 23304 41604 23316
rect 41559 23276 41604 23304
rect 41598 23264 41604 23276
rect 41656 23264 41662 23316
rect 33560 23208 34192 23236
rect 42613 23239 42671 23245
rect 33560 23196 33566 23208
rect 42613 23205 42625 23239
rect 42659 23205 42671 23239
rect 42613 23199 42671 23205
rect 12860 23140 13216 23168
rect 12860 23128 12866 23140
rect 12069 23103 12127 23109
rect 12069 23069 12081 23103
rect 12115 23069 12127 23103
rect 12069 23063 12127 23069
rect 12158 23103 12216 23109
rect 12158 23069 12170 23103
rect 12204 23069 12216 23103
rect 12158 23063 12216 23069
rect 2547 23004 4844 23032
rect 4985 23035 5043 23041
rect 2547 23001 2559 23004
rect 2501 22995 2559 23001
rect 4985 23001 4997 23035
rect 5031 23032 5043 23035
rect 5626 23032 5632 23044
rect 5031 23004 5632 23032
rect 5031 23001 5043 23004
rect 4985 22995 5043 23001
rect 5626 22992 5632 23004
rect 5684 23032 5690 23044
rect 5810 23032 5816 23044
rect 5684 23004 5816 23032
rect 5684 22992 5690 23004
rect 5810 22992 5816 23004
rect 5868 22992 5874 23044
rect 7834 22992 7840 23044
rect 7892 23032 7898 23044
rect 11348 23032 11376 23060
rect 12084 23032 12112 23063
rect 12250 23060 12256 23112
rect 12308 23109 12314 23112
rect 12308 23100 12316 23109
rect 12308 23072 12353 23100
rect 12308 23063 12316 23072
rect 12308 23060 12314 23063
rect 12434 23060 12440 23112
rect 12492 23100 12498 23112
rect 12897 23103 12955 23109
rect 12897 23100 12909 23103
rect 12492 23072 12909 23100
rect 12492 23060 12498 23072
rect 12897 23069 12909 23072
rect 12943 23069 12955 23103
rect 13078 23100 13084 23112
rect 13039 23072 13084 23100
rect 12897 23063 12955 23069
rect 7892 23004 8432 23032
rect 11348 23004 12112 23032
rect 12912 23032 12940 23063
rect 13078 23060 13084 23072
rect 13136 23060 13142 23112
rect 13188 23106 13216 23140
rect 13464 23140 16988 23168
rect 13354 23109 13360 23112
rect 13176 23100 13234 23106
rect 13176 23066 13188 23100
rect 13222 23066 13234 23100
rect 13176 23060 13234 23066
rect 13311 23103 13360 23109
rect 13311 23069 13323 23103
rect 13357 23069 13360 23103
rect 13311 23063 13360 23069
rect 13354 23060 13360 23063
rect 13412 23060 13418 23112
rect 13464 23032 13492 23140
rect 18322 23128 18328 23180
rect 18380 23168 18386 23180
rect 19981 23171 20039 23177
rect 19981 23168 19993 23171
rect 18380 23140 19993 23168
rect 18380 23128 18386 23140
rect 19981 23137 19993 23140
rect 20027 23137 20039 23171
rect 19981 23131 20039 23137
rect 21818 23128 21824 23180
rect 21876 23168 21882 23180
rect 22373 23171 22431 23177
rect 22373 23168 22385 23171
rect 21876 23140 22385 23168
rect 21876 23128 21882 23140
rect 22373 23137 22385 23140
rect 22419 23168 22431 23171
rect 24210 23168 24216 23180
rect 22419 23140 24216 23168
rect 22419 23137 22431 23140
rect 22373 23131 22431 23137
rect 24210 23128 24216 23140
rect 24268 23128 24274 23180
rect 32861 23171 32919 23177
rect 32861 23137 32873 23171
rect 32907 23168 32919 23171
rect 33042 23168 33048 23180
rect 32907 23140 33048 23168
rect 32907 23137 32919 23140
rect 32861 23131 32919 23137
rect 33042 23128 33048 23140
rect 33100 23168 33106 23180
rect 34885 23171 34943 23177
rect 34885 23168 34897 23171
rect 33100 23140 34897 23168
rect 33100 23128 33106 23140
rect 34885 23137 34897 23140
rect 34931 23137 34943 23171
rect 34885 23131 34943 23137
rect 40129 23171 40187 23177
rect 40129 23137 40141 23171
rect 40175 23168 40187 23171
rect 42628 23168 42656 23199
rect 40175 23140 42656 23168
rect 40175 23137 40187 23140
rect 40129 23131 40187 23137
rect 14366 23060 14372 23112
rect 14424 23100 14430 23112
rect 14461 23103 14519 23109
rect 14461 23100 14473 23103
rect 14424 23072 14473 23100
rect 14424 23060 14430 23072
rect 14461 23069 14473 23072
rect 14507 23069 14519 23103
rect 14461 23063 14519 23069
rect 14642 23060 14648 23112
rect 14700 23100 14706 23112
rect 15102 23100 15108 23112
rect 14700 23072 15108 23100
rect 14700 23060 14706 23072
rect 15102 23060 15108 23072
rect 15160 23100 15166 23112
rect 15289 23103 15347 23109
rect 15289 23100 15301 23103
rect 15160 23072 15301 23100
rect 15160 23060 15166 23072
rect 15289 23069 15301 23072
rect 15335 23100 15347 23103
rect 17313 23103 17371 23109
rect 17313 23100 17325 23103
rect 15335 23072 17325 23100
rect 15335 23069 15347 23072
rect 15289 23063 15347 23069
rect 17313 23069 17325 23072
rect 17359 23100 17371 23103
rect 18340 23100 18368 23128
rect 17359 23072 18368 23100
rect 17359 23069 17371 23072
rect 17313 23063 17371 23069
rect 20070 23060 20076 23112
rect 20128 23100 20134 23112
rect 20237 23103 20295 23109
rect 20237 23100 20249 23103
rect 20128 23072 20249 23100
rect 20128 23060 20134 23072
rect 20237 23069 20249 23072
rect 20283 23069 20295 23103
rect 20237 23063 20295 23069
rect 22649 23103 22707 23109
rect 22649 23069 22661 23103
rect 22695 23100 22707 23103
rect 24857 23103 24915 23109
rect 24857 23100 24869 23103
rect 22695 23072 24869 23100
rect 22695 23069 22707 23072
rect 22649 23063 22707 23069
rect 24857 23069 24869 23072
rect 24903 23069 24915 23103
rect 24857 23063 24915 23069
rect 26513 23103 26571 23109
rect 26513 23069 26525 23103
rect 26559 23100 26571 23103
rect 27246 23100 27252 23112
rect 26559 23072 27252 23100
rect 26559 23069 26571 23072
rect 26513 23063 26571 23069
rect 16206 23032 16212 23044
rect 12912 23004 13492 23032
rect 16167 23004 16212 23032
rect 7892 22992 7898 23004
rect 2130 22924 2136 22976
rect 2188 22964 2194 22976
rect 3053 22967 3111 22973
rect 3053 22964 3065 22967
rect 2188 22936 3065 22964
rect 2188 22924 2194 22936
rect 3053 22933 3065 22936
rect 3099 22964 3111 22967
rect 3326 22964 3332 22976
rect 3099 22936 3332 22964
rect 3099 22933 3111 22936
rect 3053 22927 3111 22933
rect 3326 22924 3332 22936
rect 3384 22964 3390 22976
rect 5994 22964 6000 22976
rect 3384 22936 6000 22964
rect 3384 22924 3390 22936
rect 5994 22924 6000 22936
rect 6052 22924 6058 22976
rect 7374 22924 7380 22976
rect 7432 22964 7438 22976
rect 7653 22967 7711 22973
rect 7653 22964 7665 22967
rect 7432 22936 7665 22964
rect 7432 22924 7438 22936
rect 7653 22933 7665 22936
rect 7699 22964 7711 22967
rect 8110 22964 8116 22976
rect 7699 22936 8116 22964
rect 7699 22933 7711 22936
rect 7653 22927 7711 22933
rect 8110 22924 8116 22936
rect 8168 22924 8174 22976
rect 8404 22973 8432 23004
rect 16206 22992 16212 23004
rect 16264 22992 16270 23044
rect 17586 23041 17592 23044
rect 16393 23035 16451 23041
rect 16393 23001 16405 23035
rect 16439 23001 16451 23035
rect 17580 23032 17592 23041
rect 17547 23004 17592 23032
rect 16393 22995 16451 23001
rect 17580 22995 17592 23004
rect 8389 22967 8447 22973
rect 8389 22933 8401 22967
rect 8435 22964 8447 22967
rect 8662 22964 8668 22976
rect 8435 22936 8668 22964
rect 8435 22933 8447 22936
rect 8389 22927 8447 22933
rect 8662 22924 8668 22936
rect 8720 22924 8726 22976
rect 16408 22964 16436 22995
rect 17586 22992 17592 22995
rect 17644 22992 17650 23044
rect 19978 22992 19984 23044
rect 20036 23032 20042 23044
rect 20438 23032 20444 23044
rect 20036 23004 20444 23032
rect 20036 22992 20042 23004
rect 20438 22992 20444 23004
rect 20496 23032 20502 23044
rect 22664 23032 22692 23063
rect 27246 23060 27252 23072
rect 27304 23060 27310 23112
rect 27338 23100 27396 23106
rect 27338 23066 27350 23100
rect 27384 23066 27396 23100
rect 27338 23060 27396 23066
rect 27430 23060 27436 23112
rect 27488 23100 27494 23112
rect 27488 23072 27530 23100
rect 27488 23060 27494 23072
rect 27614 23060 27620 23112
rect 27672 23100 27678 23112
rect 28626 23100 28632 23112
rect 27672 23072 28632 23100
rect 27672 23060 27678 23072
rect 28626 23060 28632 23072
rect 28684 23060 28690 23112
rect 29086 23060 29092 23112
rect 29144 23100 29150 23112
rect 29733 23103 29791 23109
rect 29733 23100 29745 23103
rect 29144 23072 29745 23100
rect 29144 23060 29150 23072
rect 29733 23069 29745 23072
rect 29779 23100 29791 23103
rect 29914 23100 29920 23112
rect 29779 23072 29920 23100
rect 29779 23069 29791 23072
rect 29733 23063 29791 23069
rect 29914 23060 29920 23072
rect 29972 23060 29978 23112
rect 33778 23100 33784 23112
rect 33739 23072 33784 23100
rect 33778 23060 33784 23072
rect 33836 23060 33842 23112
rect 33873 23103 33931 23109
rect 33873 23069 33885 23103
rect 33919 23069 33931 23103
rect 33873 23063 33931 23069
rect 23290 23032 23296 23044
rect 20496 23004 22692 23032
rect 23251 23004 23296 23032
rect 20496 22992 20502 23004
rect 23290 22992 23296 23004
rect 23348 22992 23354 23044
rect 23474 23032 23480 23044
rect 23435 23004 23480 23032
rect 23474 22992 23480 23004
rect 23532 22992 23538 23044
rect 25038 23032 25044 23044
rect 24999 23004 25044 23032
rect 25038 22992 25044 23004
rect 25096 22992 25102 23044
rect 27356 23032 27384 23060
rect 27264 23004 27384 23032
rect 28077 23035 28135 23041
rect 17954 22964 17960 22976
rect 16408 22936 17960 22964
rect 17954 22924 17960 22936
rect 18012 22964 18018 22976
rect 18693 22967 18751 22973
rect 18693 22964 18705 22967
rect 18012 22936 18705 22964
rect 18012 22924 18018 22936
rect 18693 22933 18705 22936
rect 18739 22933 18751 22967
rect 18693 22927 18751 22933
rect 23382 22924 23388 22976
rect 23440 22964 23446 22976
rect 27154 22964 27160 22976
rect 23440 22936 27160 22964
rect 23440 22924 23446 22936
rect 27154 22924 27160 22936
rect 27212 22924 27218 22976
rect 27264 22964 27292 23004
rect 28077 23001 28089 23035
rect 28123 23032 28135 23035
rect 28258 23032 28264 23044
rect 28123 23004 28264 23032
rect 28123 23001 28135 23004
rect 28077 22995 28135 23001
rect 28258 22992 28264 23004
rect 28316 22992 28322 23044
rect 28905 23035 28963 23041
rect 28905 23001 28917 23035
rect 28951 23032 28963 23035
rect 29362 23032 29368 23044
rect 28951 23004 29368 23032
rect 28951 23001 28963 23004
rect 28905 22995 28963 23001
rect 29362 22992 29368 23004
rect 29420 22992 29426 23044
rect 29549 23035 29607 23041
rect 29549 23001 29561 23035
rect 29595 23032 29607 23035
rect 30377 23035 30435 23041
rect 30377 23032 30389 23035
rect 29595 23004 30389 23032
rect 29595 23001 29607 23004
rect 29549 22995 29607 23001
rect 29932 22976 29960 23004
rect 30377 23001 30389 23004
rect 30423 23001 30435 23035
rect 30377 22995 30435 23001
rect 30466 22992 30472 23044
rect 30524 23032 30530 23044
rect 30561 23035 30619 23041
rect 30561 23032 30573 23035
rect 30524 23004 30573 23032
rect 30524 22992 30530 23004
rect 30561 23001 30573 23004
rect 30607 23001 30619 23035
rect 30561 22995 30619 23001
rect 32616 23035 32674 23041
rect 32616 23001 32628 23035
rect 32662 23032 32674 23035
rect 33505 23035 33563 23041
rect 33505 23032 33517 23035
rect 32662 23004 33517 23032
rect 32662 23001 32674 23004
rect 32616 22995 32674 23001
rect 33505 23001 33517 23004
rect 33551 23001 33563 23035
rect 33888 23032 33916 23063
rect 33962 23060 33968 23112
rect 34020 23100 34026 23112
rect 34020 23072 34065 23100
rect 34020 23060 34026 23072
rect 34146 23060 34152 23112
rect 34204 23100 34210 23112
rect 34900 23100 34928 23131
rect 35894 23100 35900 23112
rect 34204 23072 34249 23100
rect 34900 23072 35900 23100
rect 34204 23060 34210 23072
rect 35894 23060 35900 23072
rect 35952 23100 35958 23112
rect 38654 23100 38660 23112
rect 35952 23072 38660 23100
rect 35952 23060 35958 23072
rect 38654 23060 38660 23072
rect 38712 23100 38718 23112
rect 39850 23100 39856 23112
rect 38712 23072 39856 23100
rect 38712 23060 38718 23072
rect 39850 23060 39856 23072
rect 39908 23060 39914 23112
rect 43346 23100 43352 23112
rect 43307 23072 43352 23100
rect 43346 23060 43352 23072
rect 43404 23060 43410 23112
rect 43622 23100 43628 23112
rect 43583 23072 43628 23100
rect 43622 23060 43628 23072
rect 43680 23060 43686 23112
rect 34422 23032 34428 23044
rect 33888 23004 34428 23032
rect 33505 22995 33563 23001
rect 34422 22992 34428 23004
rect 34480 22992 34486 23044
rect 34790 22992 34796 23044
rect 34848 23032 34854 23044
rect 35130 23035 35188 23041
rect 35130 23032 35142 23035
rect 34848 23004 35142 23032
rect 34848 22992 34854 23004
rect 35130 23001 35142 23004
rect 35176 23001 35188 23035
rect 35130 22995 35188 23001
rect 35618 22992 35624 23044
rect 35676 23032 35682 23044
rect 36725 23035 36783 23041
rect 36725 23032 36737 23035
rect 35676 23004 36737 23032
rect 35676 22992 35682 23004
rect 36725 23001 36737 23004
rect 36771 23001 36783 23035
rect 36906 23032 36912 23044
rect 36867 23004 36912 23032
rect 36725 22995 36783 23001
rect 36906 22992 36912 23004
rect 36964 22992 36970 23044
rect 40126 22992 40132 23044
rect 40184 23032 40190 23044
rect 40184 23004 40618 23032
rect 40184 22992 40190 23004
rect 27982 22964 27988 22976
rect 27264 22936 27988 22964
rect 27982 22924 27988 22936
rect 28040 22924 28046 22976
rect 29914 22924 29920 22976
rect 29972 22924 29978 22976
rect 30006 22924 30012 22976
rect 30064 22964 30070 22976
rect 30745 22967 30803 22973
rect 30745 22964 30757 22967
rect 30064 22936 30757 22964
rect 30064 22924 30070 22936
rect 30745 22933 30757 22936
rect 30791 22933 30803 22967
rect 30745 22927 30803 22933
rect 33594 22924 33600 22976
rect 33652 22964 33658 22976
rect 34146 22964 34152 22976
rect 33652 22936 34152 22964
rect 33652 22924 33658 22936
rect 34146 22924 34152 22936
rect 34204 22924 34210 22976
rect 37093 22967 37151 22973
rect 37093 22933 37105 22967
rect 37139 22964 37151 22967
rect 37366 22964 37372 22976
rect 37139 22936 37372 22964
rect 37139 22933 37151 22936
rect 37093 22927 37151 22933
rect 37366 22924 37372 22936
rect 37424 22924 37430 22976
rect 1104 22874 68816 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 50294 22874
rect 50346 22822 50358 22874
rect 50410 22822 50422 22874
rect 50474 22822 50486 22874
rect 50538 22822 50550 22874
rect 50602 22822 68816 22874
rect 1104 22800 68816 22822
rect 3145 22763 3203 22769
rect 3145 22729 3157 22763
rect 3191 22760 3203 22763
rect 3418 22760 3424 22772
rect 3191 22732 3424 22760
rect 3191 22729 3203 22732
rect 3145 22723 3203 22729
rect 3418 22720 3424 22732
rect 3476 22720 3482 22772
rect 12161 22763 12219 22769
rect 12161 22729 12173 22763
rect 12207 22760 12219 22763
rect 12250 22760 12256 22772
rect 12207 22732 12256 22760
rect 12207 22729 12219 22732
rect 12161 22723 12219 22729
rect 12250 22720 12256 22732
rect 12308 22720 12314 22772
rect 12710 22760 12716 22772
rect 12360 22732 12716 22760
rect 2222 22692 2228 22704
rect 2183 22664 2228 22692
rect 2222 22652 2228 22664
rect 2280 22652 2286 22704
rect 2682 22652 2688 22704
rect 2740 22692 2746 22704
rect 5258 22692 5264 22704
rect 2740 22664 5264 22692
rect 2740 22652 2746 22664
rect 5258 22652 5264 22664
rect 5316 22692 5322 22704
rect 5316 22664 5580 22692
rect 5316 22652 5322 22664
rect 2409 22627 2467 22633
rect 2409 22593 2421 22627
rect 2455 22624 2467 22627
rect 2455 22596 3740 22624
rect 2455 22593 2467 22596
rect 2409 22587 2467 22593
rect 2590 22420 2596 22432
rect 2551 22392 2596 22420
rect 2590 22380 2596 22392
rect 2648 22380 2654 22432
rect 3712 22429 3740 22596
rect 5074 22584 5080 22636
rect 5132 22624 5138 22636
rect 5552 22633 5580 22664
rect 6270 22652 6276 22704
rect 6328 22692 6334 22704
rect 8849 22695 8907 22701
rect 8849 22692 8861 22695
rect 6328 22664 8861 22692
rect 6328 22652 6334 22664
rect 8849 22661 8861 22664
rect 8895 22692 8907 22695
rect 9582 22692 9588 22704
rect 8895 22664 9588 22692
rect 8895 22661 8907 22664
rect 8849 22655 8907 22661
rect 9582 22652 9588 22664
rect 9640 22692 9646 22704
rect 12360 22701 12388 22732
rect 12710 22720 12716 22732
rect 12768 22760 12774 22772
rect 12986 22760 12992 22772
rect 12768 22732 12992 22760
rect 12768 22720 12774 22732
rect 12986 22720 12992 22732
rect 13044 22720 13050 22772
rect 13078 22720 13084 22772
rect 13136 22760 13142 22772
rect 14093 22763 14151 22769
rect 14093 22760 14105 22763
rect 13136 22732 14105 22760
rect 13136 22720 13142 22732
rect 14093 22729 14105 22732
rect 14139 22729 14151 22763
rect 14093 22723 14151 22729
rect 14274 22720 14280 22772
rect 14332 22760 14338 22772
rect 17770 22760 17776 22772
rect 14332 22732 17540 22760
rect 17731 22732 17776 22760
rect 14332 22720 14338 22732
rect 12345 22695 12403 22701
rect 9640 22664 11008 22692
rect 9640 22652 9646 22664
rect 5445 22627 5503 22633
rect 5445 22624 5457 22627
rect 5132 22596 5457 22624
rect 5132 22584 5138 22596
rect 5445 22593 5457 22596
rect 5491 22593 5503 22627
rect 5445 22587 5503 22593
rect 5537 22627 5595 22633
rect 5537 22593 5549 22627
rect 5583 22593 5595 22627
rect 5537 22587 5595 22593
rect 5460 22556 5488 22587
rect 5626 22584 5632 22636
rect 5684 22624 5690 22636
rect 5813 22627 5871 22633
rect 5684 22596 5729 22624
rect 5684 22584 5690 22596
rect 5813 22593 5825 22627
rect 5859 22624 5871 22627
rect 5902 22624 5908 22636
rect 5859 22596 5908 22624
rect 5859 22593 5871 22596
rect 5813 22587 5871 22593
rect 5902 22584 5908 22596
rect 5960 22624 5966 22636
rect 7466 22624 7472 22636
rect 5960 22596 7472 22624
rect 5960 22584 5966 22596
rect 7466 22584 7472 22596
rect 7524 22584 7530 22636
rect 7653 22627 7711 22633
rect 7653 22593 7665 22627
rect 7699 22624 7711 22627
rect 8113 22627 8171 22633
rect 8113 22624 8125 22627
rect 7699 22596 8125 22624
rect 7699 22593 7711 22596
rect 7653 22587 7711 22593
rect 8113 22593 8125 22596
rect 8159 22624 8171 22627
rect 9398 22624 9404 22636
rect 8159 22596 9404 22624
rect 8159 22593 8171 22596
rect 8113 22587 8171 22593
rect 9398 22584 9404 22596
rect 9456 22584 9462 22636
rect 10709 22627 10767 22633
rect 10709 22593 10721 22627
rect 10755 22624 10767 22627
rect 10870 22624 10876 22636
rect 10755 22596 10876 22624
rect 10755 22593 10767 22596
rect 10709 22587 10767 22593
rect 10870 22584 10876 22596
rect 10928 22584 10934 22636
rect 10980 22633 11008 22664
rect 12345 22661 12357 22695
rect 12391 22661 12403 22695
rect 14461 22695 14519 22701
rect 14461 22692 14473 22695
rect 12345 22655 12403 22661
rect 12544 22664 14473 22692
rect 12544 22636 12572 22664
rect 14461 22661 14473 22664
rect 14507 22692 14519 22695
rect 15289 22695 15347 22701
rect 15289 22692 15301 22695
rect 14507 22664 15301 22692
rect 14507 22661 14519 22664
rect 14461 22655 14519 22661
rect 15289 22661 15301 22664
rect 15335 22661 15347 22695
rect 15289 22655 15347 22661
rect 16117 22695 16175 22701
rect 16117 22661 16129 22695
rect 16163 22692 16175 22695
rect 17405 22695 17463 22701
rect 17405 22692 17417 22695
rect 16163 22664 17417 22692
rect 16163 22661 16175 22664
rect 16117 22655 16175 22661
rect 17405 22661 17417 22664
rect 17451 22661 17463 22695
rect 17512 22692 17540 22732
rect 17770 22720 17776 22732
rect 17828 22720 17834 22772
rect 17880 22732 22094 22760
rect 17880 22692 17908 22732
rect 17512 22664 17908 22692
rect 17405 22655 17463 22661
rect 10965 22627 11023 22633
rect 10965 22593 10977 22627
rect 11011 22593 11023 22627
rect 12526 22624 12532 22636
rect 12487 22596 12532 22624
rect 10965 22587 11023 22593
rect 12526 22584 12532 22596
rect 12584 22584 12590 22636
rect 14277 22627 14335 22633
rect 14277 22593 14289 22627
rect 14323 22593 14335 22627
rect 14277 22587 14335 22593
rect 15105 22627 15163 22633
rect 15105 22593 15117 22627
rect 15151 22624 15163 22627
rect 15194 22624 15200 22636
rect 15151 22596 15200 22624
rect 15151 22593 15163 22596
rect 15105 22587 15163 22593
rect 6365 22559 6423 22565
rect 6365 22556 6377 22559
rect 5460 22528 6377 22556
rect 6365 22525 6377 22528
rect 6411 22556 6423 22559
rect 14292 22556 14320 22587
rect 15194 22584 15200 22596
rect 15252 22584 15258 22636
rect 15562 22584 15568 22636
rect 15620 22624 15626 22636
rect 15749 22627 15807 22633
rect 15749 22624 15761 22627
rect 15620 22596 15761 22624
rect 15620 22584 15626 22596
rect 15749 22593 15761 22596
rect 15795 22593 15807 22627
rect 15749 22587 15807 22593
rect 15838 22584 15844 22636
rect 15896 22624 15902 22636
rect 15933 22627 15991 22633
rect 15933 22624 15945 22627
rect 15896 22596 15945 22624
rect 15896 22584 15902 22596
rect 15933 22593 15945 22596
rect 15979 22593 15991 22627
rect 17126 22624 17132 22636
rect 17087 22596 17132 22624
rect 15933 22587 15991 22593
rect 17126 22584 17132 22596
rect 17184 22584 17190 22636
rect 17218 22584 17224 22636
rect 17276 22624 17282 22636
rect 17276 22596 17321 22624
rect 17276 22584 17282 22596
rect 17494 22584 17500 22636
rect 17552 22624 17558 22636
rect 17635 22627 17693 22633
rect 17552 22596 17597 22624
rect 17552 22584 17558 22596
rect 17635 22593 17647 22627
rect 17681 22624 17693 22627
rect 17862 22624 17868 22636
rect 17681 22596 17868 22624
rect 17681 22593 17693 22596
rect 17635 22587 17693 22593
rect 17862 22584 17868 22596
rect 17920 22584 17926 22636
rect 19334 22584 19340 22636
rect 19392 22624 19398 22636
rect 19705 22627 19763 22633
rect 19705 22624 19717 22627
rect 19392 22596 19717 22624
rect 19392 22584 19398 22596
rect 19705 22593 19717 22596
rect 19751 22593 19763 22627
rect 19978 22624 19984 22636
rect 19939 22596 19984 22624
rect 19705 22587 19763 22593
rect 19978 22584 19984 22596
rect 20036 22584 20042 22636
rect 15286 22556 15292 22568
rect 6411 22528 9674 22556
rect 14292 22528 15292 22556
rect 6411 22525 6423 22528
rect 6365 22519 6423 22525
rect 9646 22488 9674 22528
rect 15286 22516 15292 22528
rect 15344 22516 15350 22568
rect 22066 22556 22094 22732
rect 22830 22720 22836 22772
rect 22888 22760 22894 22772
rect 22888 22732 23980 22760
rect 22888 22720 22894 22732
rect 23952 22704 23980 22732
rect 24026 22720 24032 22772
rect 24084 22760 24090 22772
rect 27341 22763 27399 22769
rect 24084 22732 25084 22760
rect 24084 22720 24090 22732
rect 22278 22652 22284 22704
rect 22336 22692 22342 22704
rect 22741 22695 22799 22701
rect 22741 22692 22753 22695
rect 22336 22664 22753 22692
rect 22336 22652 22342 22664
rect 22741 22661 22753 22664
rect 22787 22661 22799 22695
rect 23845 22695 23903 22701
rect 23845 22692 23857 22695
rect 22741 22655 22799 22661
rect 22940 22664 23857 22692
rect 22646 22633 22652 22636
rect 22644 22624 22652 22633
rect 22607 22596 22652 22624
rect 22644 22587 22652 22596
rect 22646 22584 22652 22587
rect 22704 22584 22710 22636
rect 22830 22624 22836 22636
rect 22791 22596 22836 22624
rect 22830 22584 22836 22596
rect 22888 22584 22894 22636
rect 22940 22556 22968 22664
rect 23845 22661 23857 22664
rect 23891 22661 23903 22695
rect 23845 22655 23903 22661
rect 23934 22652 23940 22704
rect 23992 22692 23998 22704
rect 24854 22692 24860 22704
rect 23992 22664 24085 22692
rect 24135 22664 24860 22692
rect 23992 22652 23998 22664
rect 23016 22627 23074 22633
rect 23016 22593 23028 22627
rect 23062 22593 23074 22627
rect 23016 22587 23074 22593
rect 23109 22627 23167 22633
rect 23109 22593 23121 22627
rect 23155 22593 23167 22627
rect 23109 22587 23167 22593
rect 22066 22528 22968 22556
rect 9646 22460 9720 22488
rect 3697 22423 3755 22429
rect 3697 22389 3709 22423
rect 3743 22420 3755 22423
rect 4614 22420 4620 22432
rect 3743 22392 4620 22420
rect 3743 22389 3755 22392
rect 3697 22383 3755 22389
rect 4614 22380 4620 22392
rect 4672 22380 4678 22432
rect 5166 22420 5172 22432
rect 5127 22392 5172 22420
rect 5166 22380 5172 22392
rect 5224 22380 5230 22432
rect 9306 22380 9312 22432
rect 9364 22420 9370 22432
rect 9585 22423 9643 22429
rect 9585 22420 9597 22423
rect 9364 22392 9597 22420
rect 9364 22380 9370 22392
rect 9585 22389 9597 22392
rect 9631 22389 9643 22423
rect 9692 22420 9720 22460
rect 11330 22448 11336 22500
rect 11388 22488 11394 22500
rect 20254 22488 20260 22500
rect 11388 22460 20260 22488
rect 11388 22448 11394 22460
rect 20254 22448 20260 22460
rect 20312 22448 20318 22500
rect 11054 22420 11060 22432
rect 9692 22392 11060 22420
rect 9585 22383 9643 22389
rect 11054 22380 11060 22392
rect 11112 22380 11118 22432
rect 12802 22380 12808 22432
rect 12860 22420 12866 22432
rect 14921 22423 14979 22429
rect 14921 22420 14933 22423
rect 12860 22392 14933 22420
rect 12860 22380 12866 22392
rect 14921 22389 14933 22392
rect 14967 22389 14979 22423
rect 14921 22383 14979 22389
rect 22465 22423 22523 22429
rect 22465 22389 22477 22423
rect 22511 22420 22523 22423
rect 22830 22420 22836 22432
rect 22511 22392 22836 22420
rect 22511 22389 22523 22392
rect 22465 22383 22523 22389
rect 22830 22380 22836 22392
rect 22888 22380 22894 22432
rect 23032 22420 23060 22587
rect 23124 22556 23152 22587
rect 23474 22584 23480 22636
rect 23532 22624 23538 22636
rect 24135 22633 24163 22664
rect 24854 22652 24860 22664
rect 24912 22652 24918 22704
rect 23707 22627 23765 22633
rect 23707 22624 23719 22627
rect 23532 22596 23719 22624
rect 23532 22584 23538 22596
rect 23707 22593 23719 22596
rect 23753 22593 23765 22627
rect 23707 22587 23765 22593
rect 24120 22627 24178 22633
rect 24120 22593 24132 22627
rect 24166 22593 24178 22627
rect 24120 22587 24178 22593
rect 24213 22627 24271 22633
rect 24213 22593 24225 22627
rect 24259 22593 24271 22627
rect 24213 22587 24271 22593
rect 24228 22556 24256 22587
rect 24762 22584 24768 22636
rect 24820 22624 24826 22636
rect 25056 22633 25084 22732
rect 27341 22729 27353 22763
rect 27387 22760 27399 22763
rect 27430 22760 27436 22772
rect 27387 22732 27436 22760
rect 27387 22729 27399 22732
rect 27341 22723 27399 22729
rect 27430 22720 27436 22732
rect 27488 22720 27494 22772
rect 28353 22763 28411 22769
rect 28353 22729 28365 22763
rect 28399 22760 28411 22763
rect 28442 22760 28448 22772
rect 28399 22732 28448 22760
rect 28399 22729 28411 22732
rect 28353 22723 28411 22729
rect 28442 22720 28448 22732
rect 28500 22720 28506 22772
rect 28902 22720 28908 22772
rect 28960 22760 28966 22772
rect 29546 22760 29552 22772
rect 28960 22732 29552 22760
rect 28960 22720 28966 22732
rect 29546 22720 29552 22732
rect 29604 22720 29610 22772
rect 34790 22760 34796 22772
rect 34751 22732 34796 22760
rect 34790 22720 34796 22732
rect 34848 22720 34854 22772
rect 35802 22720 35808 22772
rect 35860 22760 35866 22772
rect 36906 22760 36912 22772
rect 35860 22732 36912 22760
rect 35860 22720 35866 22732
rect 36906 22720 36912 22732
rect 36964 22760 36970 22772
rect 37645 22763 37703 22769
rect 37645 22760 37657 22763
rect 36964 22732 37657 22760
rect 36964 22720 36970 22732
rect 37645 22729 37657 22732
rect 37691 22729 37703 22763
rect 40126 22760 40132 22772
rect 40087 22732 40132 22760
rect 37645 22723 37703 22729
rect 40126 22720 40132 22732
rect 40184 22720 40190 22772
rect 41785 22763 41843 22769
rect 41785 22729 41797 22763
rect 41831 22760 41843 22763
rect 42886 22760 42892 22772
rect 41831 22732 42892 22760
rect 41831 22729 41843 22732
rect 41785 22723 41843 22729
rect 42886 22720 42892 22732
rect 42944 22760 42950 22772
rect 43622 22760 43628 22772
rect 42944 22732 43628 22760
rect 42944 22720 42950 22732
rect 43622 22720 43628 22732
rect 43680 22720 43686 22772
rect 26050 22692 26056 22704
rect 26011 22664 26056 22692
rect 26050 22652 26056 22664
rect 26108 22652 26114 22704
rect 27154 22692 27160 22704
rect 27115 22664 27160 22692
rect 27154 22652 27160 22664
rect 27212 22692 27218 22704
rect 27798 22692 27804 22704
rect 27212 22664 27804 22692
rect 27212 22652 27218 22664
rect 27798 22652 27804 22664
rect 27856 22652 27862 22704
rect 27982 22652 27988 22704
rect 28040 22692 28046 22704
rect 29178 22692 29184 22704
rect 28040 22664 29184 22692
rect 28040 22652 28046 22664
rect 24949 22627 25007 22633
rect 24949 22624 24961 22627
rect 24820 22596 24961 22624
rect 24820 22584 24826 22596
rect 24949 22593 24961 22596
rect 24995 22593 25007 22627
rect 24949 22587 25007 22593
rect 25041 22627 25099 22633
rect 25041 22593 25053 22627
rect 25087 22593 25099 22627
rect 25041 22587 25099 22593
rect 25130 22584 25136 22636
rect 25188 22624 25194 22636
rect 25317 22627 25375 22633
rect 25188 22596 25233 22624
rect 25188 22584 25194 22596
rect 25317 22593 25329 22627
rect 25363 22624 25375 22627
rect 25774 22624 25780 22636
rect 25363 22596 25780 22624
rect 25363 22593 25375 22596
rect 25317 22587 25375 22593
rect 25774 22584 25780 22596
rect 25832 22584 25838 22636
rect 25866 22584 25872 22636
rect 25924 22624 25930 22636
rect 25961 22627 26019 22633
rect 25961 22624 25973 22627
rect 25924 22596 25973 22624
rect 25924 22584 25930 22596
rect 25961 22593 25973 22596
rect 26007 22593 26019 22627
rect 26142 22624 26148 22636
rect 26103 22596 26148 22624
rect 25961 22587 26019 22593
rect 26142 22584 26148 22596
rect 26200 22584 26206 22636
rect 26326 22584 26332 22636
rect 26384 22624 26390 22636
rect 26970 22624 26976 22636
rect 26384 22596 26429 22624
rect 26931 22596 26976 22624
rect 26384 22584 26390 22596
rect 26970 22584 26976 22596
rect 27028 22584 27034 22636
rect 28736 22633 28764 22664
rect 29178 22652 29184 22664
rect 29236 22692 29242 22704
rect 29236 22664 30144 22692
rect 29236 22652 29242 22664
rect 30116 22636 30144 22664
rect 35894 22652 35900 22704
rect 35952 22692 35958 22704
rect 36173 22695 36231 22701
rect 36173 22692 36185 22695
rect 35952 22664 36185 22692
rect 35952 22652 35958 22664
rect 36173 22661 36185 22664
rect 36219 22661 36231 22695
rect 36173 22655 36231 22661
rect 38654 22652 38660 22704
rect 38712 22692 38718 22704
rect 38712 22664 39068 22692
rect 38712 22652 38718 22664
rect 28609 22627 28667 22633
rect 28609 22593 28621 22627
rect 28655 22593 28667 22627
rect 28609 22587 28667 22593
rect 28721 22627 28779 22633
rect 28721 22593 28733 22627
rect 28767 22593 28779 22627
rect 28721 22587 28779 22593
rect 28813 22627 28871 22633
rect 28813 22593 28825 22627
rect 28859 22593 28871 22627
rect 28994 22624 29000 22636
rect 28955 22596 29000 22624
rect 28813 22587 28871 22593
rect 23124 22528 24072 22556
rect 24228 22528 24900 22556
rect 24044 22488 24072 22528
rect 24765 22491 24823 22497
rect 24765 22488 24777 22491
rect 24044 22460 24777 22488
rect 24765 22457 24777 22460
rect 24811 22457 24823 22491
rect 24872 22488 24900 22528
rect 25777 22491 25835 22497
rect 25777 22488 25789 22491
rect 24872 22460 25789 22488
rect 24765 22451 24823 22457
rect 25777 22457 25789 22460
rect 25823 22457 25835 22491
rect 25777 22451 25835 22457
rect 23382 22420 23388 22432
rect 23032 22392 23388 22420
rect 23382 22380 23388 22392
rect 23440 22380 23446 22432
rect 23566 22420 23572 22432
rect 23527 22392 23572 22420
rect 23566 22380 23572 22392
rect 23624 22380 23630 22432
rect 27893 22423 27951 22429
rect 27893 22389 27905 22423
rect 27939 22420 27951 22423
rect 28624 22420 28652 22587
rect 28828 22556 28856 22587
rect 28994 22584 29000 22596
rect 29052 22584 29058 22636
rect 29825 22627 29883 22633
rect 29825 22593 29837 22627
rect 29871 22593 29883 22627
rect 30006 22624 30012 22636
rect 29967 22596 30012 22624
rect 29825 22587 29883 22593
rect 29546 22556 29552 22568
rect 28828 22528 29552 22556
rect 29546 22516 29552 22528
rect 29604 22516 29610 22568
rect 29638 22516 29644 22568
rect 29696 22556 29702 22568
rect 29840 22556 29868 22587
rect 30006 22584 30012 22596
rect 30064 22584 30070 22636
rect 30098 22584 30104 22636
rect 30156 22624 30162 22636
rect 30282 22633 30288 22636
rect 30239 22627 30288 22633
rect 30156 22596 30201 22624
rect 30156 22584 30162 22596
rect 30239 22593 30251 22627
rect 30285 22593 30288 22627
rect 30239 22587 30288 22593
rect 30282 22584 30288 22587
rect 30340 22584 30346 22636
rect 33502 22624 33508 22636
rect 33463 22596 33508 22624
rect 33502 22584 33508 22596
rect 33560 22584 33566 22636
rect 33689 22627 33747 22633
rect 33689 22593 33701 22627
rect 33735 22624 33747 22627
rect 33870 22624 33876 22636
rect 33735 22596 33876 22624
rect 33735 22593 33747 22596
rect 33689 22587 33747 22593
rect 33870 22584 33876 22596
rect 33928 22584 33934 22636
rect 34146 22624 34152 22636
rect 34107 22596 34152 22624
rect 34146 22584 34152 22596
rect 34204 22584 34210 22636
rect 34312 22627 34370 22633
rect 34312 22624 34324 22627
rect 34256 22596 34324 22624
rect 29696 22528 29868 22556
rect 33321 22559 33379 22565
rect 29696 22516 29702 22528
rect 33321 22525 33333 22559
rect 33367 22556 33379 22559
rect 34256 22556 34284 22596
rect 34312 22593 34324 22596
rect 34358 22593 34370 22627
rect 34312 22587 34370 22593
rect 34422 22584 34428 22636
rect 34480 22624 34486 22636
rect 34563 22627 34621 22633
rect 34480 22596 34525 22624
rect 34480 22584 34486 22596
rect 34563 22593 34575 22627
rect 34609 22624 34621 22627
rect 34790 22624 34796 22636
rect 34609 22596 34796 22624
rect 34609 22593 34621 22596
rect 34563 22587 34621 22593
rect 34790 22584 34796 22596
rect 34848 22584 34854 22636
rect 35342 22584 35348 22636
rect 35400 22624 35406 22636
rect 35437 22627 35495 22633
rect 35437 22624 35449 22627
rect 35400 22596 35449 22624
rect 35400 22584 35406 22596
rect 35437 22593 35449 22596
rect 35483 22593 35495 22627
rect 38746 22624 38752 22636
rect 38804 22633 38810 22636
rect 39040 22633 39068 22664
rect 38716 22596 38752 22624
rect 35437 22587 35495 22593
rect 38746 22584 38752 22596
rect 38804 22587 38816 22633
rect 39025 22627 39083 22633
rect 39025 22593 39037 22627
rect 39071 22593 39083 22627
rect 40034 22624 40040 22636
rect 39995 22596 40040 22624
rect 39025 22587 39083 22593
rect 38804 22584 38810 22587
rect 40034 22584 40040 22596
rect 40092 22584 40098 22636
rect 41690 22624 41696 22636
rect 41651 22596 41696 22624
rect 41690 22584 41696 22596
rect 41748 22584 41754 22636
rect 41874 22584 41880 22636
rect 41932 22624 41938 22636
rect 42426 22624 42432 22636
rect 41932 22596 42432 22624
rect 41932 22584 41938 22596
rect 42426 22584 42432 22596
rect 42484 22584 42490 22636
rect 42610 22624 42616 22636
rect 42571 22596 42616 22624
rect 42610 22584 42616 22596
rect 42668 22584 42674 22636
rect 42794 22624 42800 22636
rect 42755 22596 42800 22624
rect 42794 22584 42800 22596
rect 42852 22584 42858 22636
rect 33367 22528 34284 22556
rect 33367 22525 33379 22528
rect 33321 22519 33379 22525
rect 30103 22460 33824 22488
rect 30103 22420 30131 22460
rect 33796 22432 33824 22460
rect 33870 22448 33876 22500
rect 33928 22488 33934 22500
rect 35618 22488 35624 22500
rect 33928 22460 35624 22488
rect 33928 22448 33934 22460
rect 35618 22448 35624 22460
rect 35676 22448 35682 22500
rect 27939 22392 30131 22420
rect 30469 22423 30527 22429
rect 27939 22389 27951 22392
rect 27893 22383 27951 22389
rect 30469 22389 30481 22423
rect 30515 22420 30527 22423
rect 32122 22420 32128 22432
rect 30515 22392 32128 22420
rect 30515 22389 30527 22392
rect 30469 22383 30527 22389
rect 32122 22380 32128 22392
rect 32180 22380 32186 22432
rect 33778 22380 33784 22432
rect 33836 22420 33842 22432
rect 36630 22420 36636 22432
rect 33836 22392 36636 22420
rect 33836 22380 33842 22392
rect 36630 22380 36636 22392
rect 36688 22380 36694 22432
rect 42058 22380 42064 22432
rect 42116 22420 42122 22432
rect 42429 22423 42487 22429
rect 42429 22420 42441 22423
rect 42116 22392 42441 22420
rect 42116 22380 42122 22392
rect 42429 22389 42441 22392
rect 42475 22389 42487 22423
rect 42429 22383 42487 22389
rect 1104 22330 68816 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 65654 22330
rect 65706 22278 65718 22330
rect 65770 22278 65782 22330
rect 65834 22278 65846 22330
rect 65898 22278 65910 22330
rect 65962 22278 68816 22330
rect 1104 22256 68816 22278
rect 5626 22176 5632 22228
rect 5684 22216 5690 22228
rect 5997 22219 6055 22225
rect 5997 22216 6009 22219
rect 5684 22188 6009 22216
rect 5684 22176 5690 22188
rect 5997 22185 6009 22188
rect 6043 22185 6055 22219
rect 5997 22179 6055 22185
rect 8294 22176 8300 22228
rect 8352 22216 8358 22228
rect 9030 22216 9036 22228
rect 8352 22188 9036 22216
rect 8352 22176 8358 22188
rect 9030 22176 9036 22188
rect 9088 22216 9094 22228
rect 10870 22216 10876 22228
rect 9088 22188 9674 22216
rect 10831 22188 10876 22216
rect 9088 22176 9094 22188
rect 2590 22108 2596 22160
rect 2648 22108 2654 22160
rect 2682 22108 2688 22160
rect 2740 22108 2746 22160
rect 2406 22012 2412 22024
rect 2367 21984 2412 22012
rect 2406 21972 2412 21984
rect 2464 21972 2470 22024
rect 2608 22021 2636 22108
rect 2700 22021 2728 22108
rect 2958 22040 2964 22092
rect 3016 22080 3022 22092
rect 4157 22083 4215 22089
rect 4157 22080 4169 22083
rect 3016 22052 4169 22080
rect 3016 22040 3022 22052
rect 4157 22049 4169 22052
rect 4203 22049 4215 22083
rect 7926 22080 7932 22092
rect 4157 22043 4215 22049
rect 6196 22052 7932 22080
rect 2572 22015 2636 22021
rect 2572 21981 2584 22015
rect 2618 21984 2636 22015
rect 2672 22015 2730 22021
rect 2618 21981 2630 21984
rect 2572 21975 2630 21981
rect 2672 21981 2684 22015
rect 2718 21981 2730 22015
rect 2672 21975 2730 21981
rect 2823 22015 2881 22021
rect 2823 21981 2835 22015
rect 2869 22012 2881 22015
rect 3234 22012 3240 22024
rect 2869 21984 3240 22012
rect 2869 21981 2881 21984
rect 2823 21975 2881 21981
rect 3234 21972 3240 21984
rect 3292 21972 3298 22024
rect 4424 22015 4482 22021
rect 4424 21981 4436 22015
rect 4470 22012 4482 22015
rect 5166 22012 5172 22024
rect 4470 21984 5172 22012
rect 4470 21981 4482 21984
rect 4424 21975 4482 21981
rect 5166 21972 5172 21984
rect 5224 21972 5230 22024
rect 6196 22021 6224 22052
rect 7926 22040 7932 22052
rect 7984 22040 7990 22092
rect 8938 22040 8944 22092
rect 8996 22080 9002 22092
rect 9646 22080 9674 22188
rect 10870 22176 10876 22188
rect 10928 22176 10934 22228
rect 11054 22176 11060 22228
rect 11112 22216 11118 22228
rect 13446 22216 13452 22228
rect 11112 22188 13452 22216
rect 11112 22176 11118 22188
rect 13446 22176 13452 22188
rect 13504 22176 13510 22228
rect 14734 22216 14740 22228
rect 13556 22188 14740 22216
rect 12802 22148 12808 22160
rect 12728 22120 12808 22148
rect 12728 22080 12756 22120
rect 12802 22108 12808 22120
rect 12860 22108 12866 22160
rect 13170 22080 13176 22092
rect 8996 22052 9041 22080
rect 9646 22052 10272 22080
rect 8996 22040 9002 22052
rect 6181 22015 6239 22021
rect 6181 21981 6193 22015
rect 6227 21981 6239 22015
rect 6181 21975 6239 21981
rect 7377 22015 7435 22021
rect 7377 21981 7389 22015
rect 7423 22012 7435 22015
rect 8294 22012 8300 22024
rect 7423 21984 8300 22012
rect 7423 21981 7435 21984
rect 7377 21975 7435 21981
rect 3053 21879 3111 21885
rect 3053 21845 3065 21879
rect 3099 21876 3111 21879
rect 3142 21876 3148 21888
rect 3099 21848 3148 21876
rect 3099 21845 3111 21848
rect 3053 21839 3111 21845
rect 3142 21836 3148 21848
rect 3200 21836 3206 21888
rect 5537 21879 5595 21885
rect 5537 21845 5549 21879
rect 5583 21876 5595 21879
rect 6196 21876 6224 21975
rect 8294 21972 8300 21984
rect 8352 21972 8358 22024
rect 8754 21972 8760 22024
rect 8812 22012 8818 22024
rect 10244 22021 10272 22052
rect 12636 22052 12756 22080
rect 12820 22052 13176 22080
rect 9217 22015 9275 22021
rect 9217 22012 9229 22015
rect 8812 21984 9229 22012
rect 8812 21972 8818 21984
rect 9217 21981 9229 21984
rect 9263 21981 9275 22015
rect 9217 21975 9275 21981
rect 10229 22015 10287 22021
rect 10229 21981 10241 22015
rect 10275 21981 10287 22015
rect 10229 21975 10287 21981
rect 10413 22015 10471 22021
rect 10413 21981 10425 22015
rect 10459 21981 10471 22015
rect 10413 21975 10471 21981
rect 10505 22015 10563 22021
rect 10505 21981 10517 22015
rect 10551 21981 10563 22015
rect 10505 21975 10563 21981
rect 6362 21944 6368 21956
rect 6323 21916 6368 21944
rect 6362 21904 6368 21916
rect 6420 21904 6426 21956
rect 7561 21947 7619 21953
rect 7561 21913 7573 21947
rect 7607 21944 7619 21947
rect 8021 21947 8079 21953
rect 8021 21944 8033 21947
rect 7607 21916 8033 21944
rect 7607 21913 7619 21916
rect 7561 21907 7619 21913
rect 8021 21913 8033 21916
rect 8067 21944 8079 21947
rect 8110 21944 8116 21956
rect 8067 21916 8116 21944
rect 8067 21913 8079 21916
rect 8021 21907 8079 21913
rect 8110 21904 8116 21916
rect 8168 21904 8174 21956
rect 8205 21947 8263 21953
rect 8205 21913 8217 21947
rect 8251 21913 8263 21947
rect 8205 21907 8263 21913
rect 8389 21947 8447 21953
rect 8389 21913 8401 21947
rect 8435 21944 8447 21947
rect 10428 21944 10456 21975
rect 8435 21916 10456 21944
rect 8435 21913 8447 21916
rect 8389 21907 8447 21913
rect 7190 21876 7196 21888
rect 5583 21848 6224 21876
rect 7151 21848 7196 21876
rect 5583 21845 5595 21848
rect 5537 21839 5595 21845
rect 7190 21836 7196 21848
rect 7248 21836 7254 21888
rect 8220 21876 8248 21907
rect 8478 21876 8484 21888
rect 8220 21848 8484 21876
rect 8478 21836 8484 21848
rect 8536 21836 8542 21888
rect 8938 21836 8944 21888
rect 8996 21876 9002 21888
rect 10520 21876 10548 21975
rect 10594 21972 10600 22024
rect 10652 22012 10658 22024
rect 10652 21984 10697 22012
rect 10652 21972 10658 21984
rect 12434 21972 12440 22024
rect 12492 22012 12498 22024
rect 12529 22015 12587 22021
rect 12529 22012 12541 22015
rect 12492 21984 12541 22012
rect 12492 21972 12498 21984
rect 12529 21981 12541 21984
rect 12575 21981 12587 22015
rect 12636 22012 12664 22052
rect 12820 22021 12848 22052
rect 13170 22040 13176 22052
rect 13228 22040 13234 22092
rect 12692 22015 12750 22021
rect 12692 22012 12704 22015
rect 12636 21984 12704 22012
rect 12529 21975 12587 21981
rect 12692 21981 12704 21984
rect 12738 21981 12750 22015
rect 12692 21975 12750 21981
rect 12805 22015 12863 22021
rect 12805 21981 12817 22015
rect 12851 21981 12863 22015
rect 12805 21975 12863 21981
rect 12897 22015 12955 22021
rect 12897 21981 12909 22015
rect 12943 22012 12955 22015
rect 13556 22012 13584 22188
rect 14734 22176 14740 22188
rect 14792 22176 14798 22228
rect 15010 22176 15016 22228
rect 15068 22176 15074 22228
rect 18049 22219 18107 22225
rect 18049 22185 18061 22219
rect 18095 22216 18107 22219
rect 19426 22216 19432 22228
rect 18095 22188 19432 22216
rect 18095 22185 18107 22188
rect 18049 22179 18107 22185
rect 19426 22176 19432 22188
rect 19484 22216 19490 22228
rect 20070 22216 20076 22228
rect 19484 22188 20076 22216
rect 19484 22176 19490 22188
rect 20070 22176 20076 22188
rect 20128 22176 20134 22228
rect 22646 22176 22652 22228
rect 22704 22216 22710 22228
rect 23474 22216 23480 22228
rect 22704 22188 23480 22216
rect 22704 22176 22710 22188
rect 23474 22176 23480 22188
rect 23532 22176 23538 22228
rect 35802 22216 35808 22228
rect 35763 22188 35808 22216
rect 35802 22176 35808 22188
rect 35860 22176 35866 22228
rect 35912 22188 36124 22216
rect 15028 22148 15056 22176
rect 25685 22151 25743 22157
rect 25685 22148 25697 22151
rect 15028 22120 15148 22148
rect 15120 22080 15148 22120
rect 19904 22120 25697 22148
rect 17865 22083 17923 22089
rect 15120 22052 17724 22080
rect 12943 21984 13584 22012
rect 14093 22015 14151 22021
rect 12943 21981 12955 21984
rect 12897 21975 12955 21981
rect 14093 21981 14105 22015
rect 14139 22012 14151 22015
rect 15102 22012 15108 22024
rect 14139 21984 15108 22012
rect 14139 21981 14151 21984
rect 14093 21975 14151 21981
rect 12066 21944 12072 21956
rect 11979 21916 12072 21944
rect 12066 21904 12072 21916
rect 12124 21944 12130 21956
rect 12342 21944 12348 21956
rect 12124 21916 12348 21944
rect 12124 21904 12130 21916
rect 12342 21904 12348 21916
rect 12400 21944 12406 21956
rect 12912 21944 12940 21975
rect 15102 21972 15108 21984
rect 15160 21972 15166 22024
rect 16206 22012 16212 22024
rect 16167 21984 16212 22012
rect 16206 21972 16212 21984
rect 16264 21972 16270 22024
rect 16301 22015 16359 22021
rect 16301 21981 16313 22015
rect 16347 21981 16359 22015
rect 16301 21975 16359 21981
rect 12400 21916 12940 21944
rect 13173 21947 13231 21953
rect 12400 21904 12406 21916
rect 13173 21913 13185 21947
rect 13219 21944 13231 21947
rect 14338 21947 14396 21953
rect 14338 21944 14350 21947
rect 13219 21916 14350 21944
rect 13219 21913 13231 21916
rect 13173 21907 13231 21913
rect 14338 21913 14350 21916
rect 14384 21913 14396 21947
rect 14338 21907 14396 21913
rect 14918 21904 14924 21956
rect 14976 21944 14982 21956
rect 16316 21944 16344 21975
rect 16390 21972 16396 22024
rect 16448 22012 16454 22024
rect 16574 22012 16580 22024
rect 16448 21984 16493 22012
rect 16535 21984 16580 22012
rect 16448 21972 16454 21984
rect 16574 21972 16580 21984
rect 16632 21972 16638 22024
rect 17586 21972 17592 22024
rect 17644 21972 17650 22024
rect 17604 21944 17632 21972
rect 14976 21916 17632 21944
rect 14976 21904 14982 21916
rect 8996 21848 10548 21876
rect 8996 21836 9002 21848
rect 15194 21836 15200 21888
rect 15252 21876 15258 21888
rect 15473 21879 15531 21885
rect 15473 21876 15485 21879
rect 15252 21848 15485 21876
rect 15252 21836 15258 21848
rect 15473 21845 15485 21848
rect 15519 21876 15531 21879
rect 15746 21876 15752 21888
rect 15519 21848 15752 21876
rect 15519 21845 15531 21848
rect 15473 21839 15531 21845
rect 15746 21836 15752 21848
rect 15804 21836 15810 21888
rect 15930 21876 15936 21888
rect 15891 21848 15936 21876
rect 15930 21836 15936 21848
rect 15988 21836 15994 21888
rect 17586 21876 17592 21888
rect 17547 21848 17592 21876
rect 17586 21836 17592 21848
rect 17644 21836 17650 21888
rect 17696 21876 17724 22052
rect 17865 22049 17877 22083
rect 17911 22080 17923 22083
rect 17954 22080 17960 22092
rect 17911 22052 17960 22080
rect 17911 22049 17923 22052
rect 17865 22043 17923 22049
rect 17954 22040 17960 22052
rect 18012 22080 18018 22092
rect 18012 22052 19564 22080
rect 18012 22040 18018 22052
rect 17773 22015 17831 22021
rect 17773 21981 17785 22015
rect 17819 22012 17831 22015
rect 18874 22012 18880 22024
rect 17819 21984 18880 22012
rect 17819 21981 17831 21984
rect 17773 21975 17831 21981
rect 18874 21972 18880 21984
rect 18932 21972 18938 22024
rect 19426 22021 19432 22024
rect 19424 22012 19432 22021
rect 19387 21984 19432 22012
rect 19424 21975 19432 21984
rect 19426 21972 19432 21975
rect 19484 21972 19490 22024
rect 19536 22021 19564 22052
rect 19904 22021 19932 22120
rect 25685 22117 25697 22120
rect 25731 22117 25743 22151
rect 25685 22111 25743 22117
rect 26970 22108 26976 22160
rect 27028 22148 27034 22160
rect 29914 22148 29920 22160
rect 27028 22120 29920 22148
rect 27028 22108 27034 22120
rect 29914 22108 29920 22120
rect 29972 22108 29978 22160
rect 27709 22083 27767 22089
rect 27709 22049 27721 22083
rect 27755 22080 27767 22083
rect 28166 22080 28172 22092
rect 27755 22052 28172 22080
rect 27755 22049 27767 22052
rect 27709 22043 27767 22049
rect 28166 22040 28172 22052
rect 28224 22040 28230 22092
rect 29546 22080 29552 22092
rect 29507 22052 29552 22080
rect 29546 22040 29552 22052
rect 29604 22040 29610 22092
rect 34057 22083 34115 22089
rect 34057 22049 34069 22083
rect 34103 22080 34115 22083
rect 34790 22080 34796 22092
rect 34103 22052 34796 22080
rect 34103 22049 34115 22052
rect 34057 22043 34115 22049
rect 34790 22040 34796 22052
rect 34848 22080 34854 22092
rect 35434 22080 35440 22092
rect 34848 22052 35440 22080
rect 34848 22040 34854 22052
rect 35434 22040 35440 22052
rect 35492 22040 35498 22092
rect 35912 22089 35940 22188
rect 35986 22108 35992 22160
rect 36044 22108 36050 22160
rect 35897 22083 35955 22089
rect 35897 22080 35909 22083
rect 35807 22052 35909 22080
rect 35897 22049 35909 22052
rect 35943 22049 35955 22083
rect 35897 22043 35955 22049
rect 19521 22015 19579 22021
rect 19521 21981 19533 22015
rect 19567 21981 19579 22015
rect 19521 21975 19579 21981
rect 19796 22015 19854 22021
rect 19796 21981 19808 22015
rect 19842 21981 19854 22015
rect 19796 21975 19854 21981
rect 19889 22015 19947 22021
rect 19889 21981 19901 22015
rect 19935 21981 19947 22015
rect 19889 21975 19947 21981
rect 18049 21947 18107 21953
rect 18049 21913 18061 21947
rect 18095 21944 18107 21947
rect 19334 21944 19340 21956
rect 18095 21916 19340 21944
rect 18095 21913 18107 21916
rect 18049 21907 18107 21913
rect 18064 21876 18092 21907
rect 19334 21904 19340 21916
rect 19392 21904 19398 21956
rect 19613 21947 19671 21953
rect 19613 21913 19625 21947
rect 19659 21913 19671 21947
rect 19812 21944 19840 21975
rect 19978 21972 19984 22024
rect 20036 22012 20042 22024
rect 20530 22012 20536 22024
rect 20036 21984 20536 22012
rect 20036 21972 20042 21984
rect 20530 21972 20536 21984
rect 20588 21972 20594 22024
rect 21818 22012 21824 22024
rect 21779 21984 21824 22012
rect 21818 21972 21824 21984
rect 21876 21972 21882 22024
rect 21910 21972 21916 22024
rect 21968 22012 21974 22024
rect 22186 22012 22192 22024
rect 21968 21984 22013 22012
rect 22147 21984 22192 22012
rect 21968 21972 21974 21984
rect 22186 21972 22192 21984
rect 22244 21972 22250 22024
rect 22833 22015 22891 22021
rect 22833 21981 22845 22015
rect 22879 22012 22891 22015
rect 22922 22012 22928 22024
rect 22879 21984 22928 22012
rect 22879 21981 22891 21984
rect 22833 21975 22891 21981
rect 22922 21972 22928 21984
rect 22980 21972 22986 22024
rect 23014 21972 23020 22024
rect 23072 22012 23078 22024
rect 23201 22015 23259 22021
rect 23072 21984 23117 22012
rect 23072 21972 23078 21984
rect 23201 21981 23213 22015
rect 23247 21981 23259 22015
rect 23201 21975 23259 21981
rect 20990 21944 20996 21956
rect 19812 21916 20996 21944
rect 19613 21907 19671 21913
rect 17696 21848 18092 21876
rect 18506 21836 18512 21888
rect 18564 21876 18570 21888
rect 19245 21879 19303 21885
rect 19245 21876 19257 21879
rect 18564 21848 19257 21876
rect 18564 21836 18570 21848
rect 19245 21845 19257 21848
rect 19291 21845 19303 21879
rect 19628 21876 19656 21907
rect 20990 21904 20996 21916
rect 21048 21904 21054 21956
rect 22005 21947 22063 21953
rect 22005 21913 22017 21947
rect 22051 21944 22063 21947
rect 22462 21944 22468 21956
rect 22051 21916 22468 21944
rect 22051 21913 22063 21916
rect 22005 21907 22063 21913
rect 22462 21904 22468 21916
rect 22520 21904 22526 21956
rect 23109 21947 23167 21953
rect 23109 21913 23121 21947
rect 23155 21913 23167 21947
rect 23216 21944 23244 21975
rect 24762 21972 24768 22024
rect 24820 22012 24826 22024
rect 25866 22012 25872 22024
rect 24820 21984 25872 22012
rect 24820 21972 24826 21984
rect 25866 21972 25872 21984
rect 25924 21972 25930 22024
rect 25958 21972 25964 22024
rect 26016 22012 26022 22024
rect 26237 22015 26295 22021
rect 26016 21984 26061 22012
rect 26016 21972 26022 21984
rect 26237 21981 26249 22015
rect 26283 21981 26295 22015
rect 27982 22012 27988 22024
rect 27943 21984 27988 22012
rect 26237 21975 26295 21981
rect 24780 21944 24808 21972
rect 23216 21916 24808 21944
rect 23109 21907 23167 21913
rect 20254 21876 20260 21888
rect 19628 21848 20260 21876
rect 19245 21839 19303 21845
rect 20254 21836 20260 21848
rect 20312 21836 20318 21888
rect 21542 21836 21548 21888
rect 21600 21876 21606 21888
rect 21637 21879 21695 21885
rect 21637 21876 21649 21879
rect 21600 21848 21649 21876
rect 21600 21836 21606 21848
rect 21637 21845 21649 21848
rect 21683 21845 21695 21879
rect 23124 21876 23152 21907
rect 25130 21904 25136 21956
rect 25188 21944 25194 21956
rect 26053 21947 26111 21953
rect 26053 21944 26065 21947
rect 25188 21916 26065 21944
rect 25188 21904 25194 21916
rect 26053 21913 26065 21916
rect 26099 21944 26111 21947
rect 26142 21944 26148 21956
rect 26099 21916 26148 21944
rect 26099 21913 26111 21916
rect 26053 21907 26111 21913
rect 26142 21904 26148 21916
rect 26200 21904 26206 21956
rect 23198 21876 23204 21888
rect 23124 21848 23204 21876
rect 21637 21839 21695 21845
rect 23198 21836 23204 21848
rect 23256 21836 23262 21888
rect 23385 21879 23443 21885
rect 23385 21845 23397 21879
rect 23431 21876 23443 21879
rect 23658 21876 23664 21888
rect 23431 21848 23664 21876
rect 23431 21845 23443 21848
rect 23385 21839 23443 21845
rect 23658 21836 23664 21848
rect 23716 21836 23722 21888
rect 24486 21876 24492 21888
rect 24447 21848 24492 21876
rect 24486 21836 24492 21848
rect 24544 21836 24550 21888
rect 26252 21876 26280 21975
rect 27982 21972 27988 21984
rect 28040 21972 28046 22024
rect 29914 22012 29920 22024
rect 29875 21984 29920 22012
rect 29914 21972 29920 21984
rect 29972 21972 29978 22024
rect 30282 21972 30288 22024
rect 30340 22012 30346 22024
rect 30469 22015 30527 22021
rect 30469 22012 30481 22015
rect 30340 21984 30481 22012
rect 30340 21972 30346 21984
rect 30469 21981 30481 21984
rect 30515 22012 30527 22015
rect 31662 22012 31668 22024
rect 30515 21984 31668 22012
rect 30515 21981 30527 21984
rect 30469 21975 30527 21981
rect 31662 21972 31668 21984
rect 31720 21972 31726 22024
rect 32122 22012 32128 22024
rect 32180 22021 32186 22024
rect 32092 21984 32128 22012
rect 32122 21972 32128 21984
rect 32180 21975 32192 22021
rect 32398 22012 32404 22024
rect 32359 21984 32404 22012
rect 32180 21972 32186 21975
rect 32398 21972 32404 21984
rect 32456 21972 32462 22024
rect 35912 22012 35940 22043
rect 36004 22021 36032 22108
rect 36096 22080 36124 22188
rect 68094 22148 68100 22160
rect 68055 22120 68100 22148
rect 68094 22108 68100 22120
rect 68152 22108 68158 22160
rect 36446 22080 36452 22092
rect 36096 22052 36452 22080
rect 36446 22040 36452 22052
rect 36504 22040 36510 22092
rect 37829 22083 37887 22089
rect 37829 22049 37841 22083
rect 37875 22080 37887 22083
rect 38746 22080 38752 22092
rect 37875 22052 38752 22080
rect 37875 22049 37887 22052
rect 37829 22043 37887 22049
rect 38746 22040 38752 22052
rect 38804 22040 38810 22092
rect 39850 22080 39856 22092
rect 39811 22052 39856 22080
rect 39850 22040 39856 22052
rect 39908 22040 39914 22092
rect 35452 21984 35940 22012
rect 35989 22015 36047 22021
rect 27614 21904 27620 21956
rect 27672 21944 27678 21956
rect 29730 21944 29736 21956
rect 27672 21916 29736 21944
rect 27672 21904 27678 21916
rect 29730 21904 29736 21916
rect 29788 21904 29794 21956
rect 35452 21944 35480 21984
rect 35989 21981 36001 22015
rect 36035 21981 36047 22015
rect 35989 21975 36047 21981
rect 37185 22015 37243 22021
rect 37185 21981 37197 22015
rect 37231 21981 37243 22015
rect 37366 22012 37372 22024
rect 37327 21984 37372 22012
rect 37185 21975 37243 21981
rect 29840 21916 35480 21944
rect 29840 21876 29868 21916
rect 35526 21904 35532 21956
rect 35584 21944 35590 21956
rect 35713 21947 35771 21953
rect 35713 21944 35725 21947
rect 35584 21916 35725 21944
rect 35584 21904 35590 21916
rect 35713 21913 35725 21916
rect 35759 21944 35771 21947
rect 36633 21947 36691 21953
rect 36633 21944 36645 21947
rect 35759 21916 36645 21944
rect 35759 21913 35771 21916
rect 35713 21907 35771 21913
rect 36633 21913 36645 21916
rect 36679 21913 36691 21947
rect 37200 21944 37228 21975
rect 37366 21972 37372 21984
rect 37424 21972 37430 22024
rect 37458 21972 37464 22024
rect 37516 22012 37522 22024
rect 37599 22015 37657 22021
rect 37516 21984 37561 22012
rect 37516 21972 37522 21984
rect 37599 21981 37611 22015
rect 37645 22012 37657 22015
rect 38289 22015 38347 22021
rect 38289 22012 38301 22015
rect 37645 21984 38301 22012
rect 37645 21981 37657 21984
rect 37599 21975 37657 21981
rect 38289 21981 38301 21984
rect 38335 22012 38347 22015
rect 38378 22012 38384 22024
rect 38335 21984 38384 22012
rect 38335 21981 38347 21984
rect 38289 21975 38347 21981
rect 38378 21972 38384 21984
rect 38436 21972 38442 22024
rect 42058 22012 42064 22024
rect 42019 21984 42064 22012
rect 42058 21972 42064 21984
rect 42116 21972 42122 22024
rect 37274 21944 37280 21956
rect 37200 21916 37280 21944
rect 36633 21907 36691 21913
rect 37274 21904 37280 21916
rect 37332 21904 37338 21956
rect 38194 21904 38200 21956
rect 38252 21944 38258 21956
rect 40098 21947 40156 21953
rect 40098 21944 40110 21947
rect 38252 21916 40110 21944
rect 38252 21904 38258 21916
rect 40098 21913 40110 21916
rect 40144 21913 40156 21947
rect 40098 21907 40156 21913
rect 26252 21848 29868 21876
rect 30466 21836 30472 21888
rect 30524 21876 30530 21888
rect 31021 21879 31079 21885
rect 31021 21876 31033 21879
rect 30524 21848 31033 21876
rect 30524 21836 30530 21848
rect 31021 21845 31033 21848
rect 31067 21845 31079 21879
rect 31021 21839 31079 21845
rect 35253 21879 35311 21885
rect 35253 21845 35265 21879
rect 35299 21876 35311 21879
rect 35342 21876 35348 21888
rect 35299 21848 35348 21876
rect 35299 21845 35311 21848
rect 35253 21839 35311 21845
rect 35342 21836 35348 21848
rect 35400 21836 35406 21888
rect 36173 21879 36231 21885
rect 36173 21845 36185 21879
rect 36219 21876 36231 21879
rect 36538 21876 36544 21888
rect 36219 21848 36544 21876
rect 36219 21845 36231 21848
rect 36173 21839 36231 21845
rect 36538 21836 36544 21848
rect 36596 21836 36602 21888
rect 41233 21879 41291 21885
rect 41233 21845 41245 21879
rect 41279 21876 41291 21879
rect 41782 21876 41788 21888
rect 41279 21848 41788 21876
rect 41279 21845 41291 21848
rect 41233 21839 41291 21845
rect 41782 21836 41788 21848
rect 41840 21836 41846 21888
rect 42245 21879 42303 21885
rect 42245 21845 42257 21879
rect 42291 21876 42303 21879
rect 42518 21876 42524 21888
rect 42291 21848 42524 21876
rect 42291 21845 42303 21848
rect 42245 21839 42303 21845
rect 42518 21836 42524 21848
rect 42576 21836 42582 21888
rect 1104 21786 68816 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 50294 21786
rect 50346 21734 50358 21786
rect 50410 21734 50422 21786
rect 50474 21734 50486 21786
rect 50538 21734 50550 21786
rect 50602 21734 68816 21786
rect 1104 21712 68816 21734
rect 5810 21632 5816 21684
rect 5868 21672 5874 21684
rect 10502 21672 10508 21684
rect 5868 21644 10508 21672
rect 5868 21632 5874 21644
rect 10502 21632 10508 21644
rect 10560 21632 10566 21684
rect 10594 21632 10600 21684
rect 10652 21672 10658 21684
rect 12618 21672 12624 21684
rect 10652 21644 12624 21672
rect 10652 21632 10658 21644
rect 12618 21632 12624 21644
rect 12676 21672 12682 21684
rect 16206 21672 16212 21684
rect 12676 21644 16212 21672
rect 12676 21632 12682 21644
rect 16206 21632 16212 21644
rect 16264 21632 16270 21684
rect 16390 21632 16396 21684
rect 16448 21672 16454 21684
rect 17037 21675 17095 21681
rect 17037 21672 17049 21675
rect 16448 21644 17049 21672
rect 16448 21632 16454 21644
rect 17037 21641 17049 21644
rect 17083 21641 17095 21675
rect 17037 21635 17095 21641
rect 17678 21632 17684 21684
rect 17736 21672 17742 21684
rect 17865 21675 17923 21681
rect 17865 21672 17877 21675
rect 17736 21644 17877 21672
rect 17736 21632 17742 21644
rect 17865 21641 17877 21644
rect 17911 21641 17923 21675
rect 17865 21635 17923 21641
rect 20162 21632 20168 21684
rect 20220 21672 20226 21684
rect 20901 21675 20959 21681
rect 20901 21672 20913 21675
rect 20220 21644 20913 21672
rect 20220 21632 20226 21644
rect 20901 21641 20913 21644
rect 20947 21641 20959 21675
rect 20901 21635 20959 21641
rect 20990 21632 20996 21684
rect 21048 21672 21054 21684
rect 29086 21672 29092 21684
rect 21048 21644 29092 21672
rect 21048 21632 21054 21644
rect 8573 21607 8631 21613
rect 8573 21573 8585 21607
rect 8619 21604 8631 21607
rect 12250 21604 12256 21616
rect 8619 21576 9168 21604
rect 8619 21573 8631 21576
rect 8573 21567 8631 21573
rect 2869 21539 2927 21545
rect 2869 21505 2881 21539
rect 2915 21536 2927 21539
rect 2958 21536 2964 21548
rect 2915 21508 2964 21536
rect 2915 21505 2927 21508
rect 2869 21499 2927 21505
rect 2958 21496 2964 21508
rect 3016 21496 3022 21548
rect 3142 21545 3148 21548
rect 3136 21536 3148 21545
rect 3103 21508 3148 21536
rect 3136 21499 3148 21508
rect 3142 21496 3148 21499
rect 3200 21496 3206 21548
rect 6638 21545 6644 21548
rect 6632 21499 6644 21545
rect 6696 21536 6702 21548
rect 8202 21536 8208 21548
rect 6696 21508 6732 21536
rect 8163 21508 8208 21536
rect 6638 21496 6644 21499
rect 6696 21496 6702 21508
rect 8202 21496 8208 21508
rect 8260 21496 8266 21548
rect 8294 21496 8300 21548
rect 8352 21536 8358 21548
rect 8389 21539 8447 21545
rect 8389 21536 8401 21539
rect 8352 21508 8401 21536
rect 8352 21496 8358 21508
rect 8389 21505 8401 21508
rect 8435 21505 8447 21539
rect 9030 21536 9036 21548
rect 8991 21508 9036 21536
rect 8389 21499 8447 21505
rect 9030 21496 9036 21508
rect 9088 21496 9094 21548
rect 9140 21536 9168 21576
rect 11913 21576 12256 21604
rect 11913 21548 11941 21576
rect 12250 21564 12256 21576
rect 12308 21604 12314 21616
rect 12713 21607 12771 21613
rect 12308 21576 12572 21604
rect 12308 21564 12314 21576
rect 9217 21539 9275 21545
rect 9217 21536 9229 21539
rect 9140 21508 9229 21536
rect 9217 21505 9229 21508
rect 9263 21505 9275 21539
rect 9217 21499 9275 21505
rect 9309 21539 9367 21545
rect 9309 21505 9321 21539
rect 9355 21505 9367 21539
rect 9309 21499 9367 21505
rect 9401 21539 9459 21545
rect 9401 21505 9413 21539
rect 9447 21536 9459 21539
rect 10226 21536 10232 21548
rect 9447 21508 10232 21536
rect 9447 21505 9459 21508
rect 9401 21499 9459 21505
rect 5534 21428 5540 21480
rect 5592 21468 5598 21480
rect 6365 21471 6423 21477
rect 6365 21468 6377 21471
rect 5592 21440 6377 21468
rect 5592 21428 5598 21440
rect 6365 21437 6377 21440
rect 6411 21437 6423 21471
rect 6365 21431 6423 21437
rect 7834 21428 7840 21480
rect 7892 21468 7898 21480
rect 8754 21468 8760 21480
rect 7892 21440 8760 21468
rect 7892 21428 7898 21440
rect 8754 21428 8760 21440
rect 8812 21468 8818 21480
rect 9324 21468 9352 21499
rect 10226 21496 10232 21508
rect 10284 21496 10290 21548
rect 11698 21496 11704 21548
rect 11756 21545 11762 21548
rect 11756 21539 11805 21545
rect 11756 21505 11759 21539
rect 11793 21505 11805 21539
rect 11756 21499 11805 21505
rect 11898 21542 11956 21548
rect 11898 21508 11910 21542
rect 11944 21508 11956 21542
rect 11898 21502 11956 21508
rect 11998 21539 12056 21545
rect 11998 21505 12010 21539
rect 12044 21536 12056 21539
rect 12161 21539 12219 21545
rect 12044 21508 12112 21536
rect 12044 21505 12056 21508
rect 11998 21499 12056 21505
rect 11756 21496 11762 21499
rect 9674 21468 9680 21480
rect 8812 21440 9352 21468
rect 9416 21440 9680 21468
rect 8812 21428 8818 21440
rect 9416 21400 9444 21440
rect 9674 21428 9680 21440
rect 9732 21428 9738 21480
rect 12084 21468 12112 21508
rect 12161 21505 12173 21539
rect 12207 21536 12219 21539
rect 12434 21536 12440 21548
rect 12207 21508 12440 21536
rect 12207 21505 12219 21508
rect 12161 21499 12219 21505
rect 12434 21496 12440 21508
rect 12492 21496 12498 21548
rect 12544 21536 12572 21576
rect 12713 21573 12725 21607
rect 12759 21604 12771 21607
rect 12894 21604 12900 21616
rect 12759 21576 12900 21604
rect 12759 21573 12771 21576
rect 12713 21567 12771 21573
rect 12894 21564 12900 21576
rect 12952 21564 12958 21616
rect 15657 21607 15715 21613
rect 15657 21573 15669 21607
rect 15703 21604 15715 21607
rect 17218 21604 17224 21616
rect 15703 21576 17224 21604
rect 15703 21573 15715 21576
rect 15657 21567 15715 21573
rect 17218 21564 17224 21576
rect 17276 21564 17282 21616
rect 18509 21607 18567 21613
rect 18509 21604 18521 21607
rect 17880 21576 18521 21604
rect 17880 21548 17908 21576
rect 18509 21573 18521 21576
rect 18555 21604 18567 21607
rect 19794 21604 19800 21616
rect 18555 21576 19800 21604
rect 18555 21573 18567 21576
rect 18509 21567 18567 21573
rect 19794 21564 19800 21576
rect 19852 21564 19858 21616
rect 20070 21604 20076 21616
rect 20031 21576 20076 21604
rect 20070 21564 20076 21576
rect 20128 21564 20134 21616
rect 23382 21604 23388 21616
rect 20363 21576 23388 21604
rect 13170 21536 13176 21548
rect 12544 21508 13176 21536
rect 13170 21496 13176 21508
rect 13228 21496 13234 21548
rect 15562 21536 15568 21548
rect 15475 21508 15568 21536
rect 15562 21496 15568 21508
rect 15620 21496 15626 21548
rect 15746 21496 15752 21548
rect 15804 21536 15810 21548
rect 16022 21536 16028 21548
rect 15804 21508 16028 21536
rect 15804 21496 15810 21508
rect 16022 21496 16028 21508
rect 16080 21496 16086 21548
rect 16669 21539 16727 21545
rect 16669 21505 16681 21539
rect 16715 21536 16727 21539
rect 16758 21536 16764 21548
rect 16715 21508 16764 21536
rect 16715 21505 16727 21508
rect 16669 21499 16727 21505
rect 16758 21496 16764 21508
rect 16816 21496 16822 21548
rect 16861 21539 16919 21545
rect 16861 21505 16873 21539
rect 16907 21536 16919 21539
rect 17862 21536 17868 21548
rect 16907 21508 17264 21536
rect 17823 21508 17868 21536
rect 16907 21505 16919 21508
rect 16861 21499 16919 21505
rect 12250 21468 12256 21480
rect 12084 21440 12256 21468
rect 12250 21428 12256 21440
rect 12308 21428 12314 21480
rect 15580 21468 15608 21496
rect 17236 21480 17264 21508
rect 17862 21496 17868 21508
rect 17920 21496 17926 21548
rect 18049 21539 18107 21545
rect 18049 21505 18061 21539
rect 18095 21536 18107 21539
rect 19058 21536 19064 21548
rect 18095 21508 19064 21536
rect 18095 21505 18107 21508
rect 18049 21499 18107 21505
rect 19058 21496 19064 21508
rect 19116 21496 19122 21548
rect 19426 21496 19432 21548
rect 19484 21536 19490 21548
rect 19935 21539 19993 21545
rect 19935 21536 19947 21539
rect 19484 21508 19947 21536
rect 19484 21496 19490 21508
rect 19935 21505 19947 21508
rect 19981 21505 19993 21539
rect 19935 21499 19993 21505
rect 20165 21539 20223 21545
rect 20165 21505 20177 21539
rect 20211 21536 20223 21539
rect 20254 21536 20260 21548
rect 20211 21508 20260 21536
rect 20211 21505 20223 21508
rect 20165 21499 20223 21505
rect 20254 21496 20260 21508
rect 20312 21496 20318 21548
rect 20363 21545 20391 21576
rect 23382 21564 23388 21576
rect 23440 21564 23446 21616
rect 23474 21564 23480 21616
rect 23532 21604 23538 21616
rect 23934 21604 23940 21616
rect 23532 21576 23940 21604
rect 23532 21564 23538 21576
rect 23934 21564 23940 21576
rect 23992 21604 23998 21616
rect 24397 21607 24455 21613
rect 24397 21604 24409 21607
rect 23992 21576 24409 21604
rect 23992 21564 23998 21576
rect 24397 21573 24409 21576
rect 24443 21573 24455 21607
rect 25590 21604 25596 21616
rect 24397 21567 24455 21573
rect 24596 21576 25596 21604
rect 20348 21539 20406 21545
rect 20348 21505 20360 21539
rect 20394 21505 20406 21539
rect 20348 21499 20406 21505
rect 20438 21496 20444 21548
rect 20496 21536 20502 21548
rect 20898 21536 20904 21548
rect 20496 21508 20541 21536
rect 20859 21508 20904 21536
rect 20496 21496 20502 21508
rect 20898 21496 20904 21508
rect 20956 21496 20962 21548
rect 21085 21539 21143 21545
rect 21085 21505 21097 21539
rect 21131 21536 21143 21539
rect 22370 21536 22376 21548
rect 21131 21508 22376 21536
rect 21131 21505 21143 21508
rect 21085 21499 21143 21505
rect 16574 21468 16580 21480
rect 15580 21440 16580 21468
rect 16574 21428 16580 21440
rect 16632 21428 16638 21480
rect 17218 21428 17224 21480
rect 17276 21428 17282 21480
rect 19150 21428 19156 21480
rect 19208 21468 19214 21480
rect 21100 21468 21128 21499
rect 22370 21496 22376 21508
rect 22428 21496 22434 21548
rect 22833 21539 22891 21545
rect 22833 21505 22845 21539
rect 22879 21536 22891 21539
rect 23014 21536 23020 21548
rect 22879 21508 23020 21536
rect 22879 21505 22891 21508
rect 22833 21499 22891 21505
rect 23014 21496 23020 21508
rect 23072 21496 23078 21548
rect 23566 21496 23572 21548
rect 23624 21536 23630 21548
rect 24167 21539 24225 21545
rect 24167 21536 24179 21539
rect 23624 21508 24179 21536
rect 23624 21496 23630 21508
rect 24167 21505 24179 21508
rect 24213 21505 24225 21539
rect 24302 21536 24308 21548
rect 24263 21508 24308 21536
rect 24167 21499 24225 21505
rect 24302 21496 24308 21508
rect 24360 21496 24366 21548
rect 24596 21545 24624 21576
rect 25590 21564 25596 21576
rect 25648 21564 25654 21616
rect 27249 21607 27307 21613
rect 27249 21573 27261 21607
rect 27295 21604 27307 21607
rect 27890 21604 27896 21616
rect 27295 21576 27896 21604
rect 27295 21573 27307 21576
rect 27249 21567 27307 21573
rect 27890 21564 27896 21576
rect 27948 21564 27954 21616
rect 24580 21539 24638 21545
rect 24580 21505 24592 21539
rect 24626 21505 24638 21539
rect 24580 21499 24638 21505
rect 24670 21496 24676 21548
rect 24728 21536 24734 21548
rect 24728 21508 24773 21536
rect 24728 21496 24734 21508
rect 24854 21496 24860 21548
rect 24912 21536 24918 21548
rect 25608 21536 25636 21564
rect 27706 21536 27712 21548
rect 24912 21508 25544 21536
rect 25608 21508 27712 21536
rect 24912 21496 24918 21508
rect 19208 21440 21128 21468
rect 19208 21428 19214 21440
rect 22462 21428 22468 21480
rect 22520 21468 22526 21480
rect 22557 21471 22615 21477
rect 22557 21468 22569 21471
rect 22520 21440 22569 21468
rect 22520 21428 22526 21440
rect 22557 21437 22569 21440
rect 22603 21437 22615 21471
rect 24320 21468 24348 21496
rect 25133 21471 25191 21477
rect 25133 21468 25145 21471
rect 24320 21440 25145 21468
rect 22557 21431 22615 21437
rect 25133 21437 25145 21440
rect 25179 21437 25191 21471
rect 25516 21468 25544 21508
rect 27706 21496 27712 21508
rect 27764 21496 27770 21548
rect 28000 21545 28028 21644
rect 29086 21632 29092 21644
rect 29144 21632 29150 21684
rect 32490 21632 32496 21684
rect 32548 21672 32554 21684
rect 34701 21675 34759 21681
rect 34701 21672 34713 21675
rect 32548 21644 34713 21672
rect 32548 21632 32554 21644
rect 34701 21641 34713 21644
rect 34747 21672 34759 21675
rect 35986 21672 35992 21684
rect 34747 21644 35992 21672
rect 34747 21641 34759 21644
rect 34701 21635 34759 21641
rect 35986 21632 35992 21644
rect 36044 21632 36050 21684
rect 38194 21672 38200 21684
rect 38155 21644 38200 21672
rect 38194 21632 38200 21644
rect 38252 21632 38258 21684
rect 41693 21675 41751 21681
rect 41693 21641 41705 21675
rect 41739 21672 41751 21675
rect 42610 21672 42616 21684
rect 41739 21644 42616 21672
rect 41739 21641 41751 21644
rect 41693 21635 41751 21641
rect 42610 21632 42616 21644
rect 42668 21632 42674 21684
rect 43073 21675 43131 21681
rect 43073 21641 43085 21675
rect 43119 21672 43131 21675
rect 43346 21672 43352 21684
rect 43119 21644 43352 21672
rect 43119 21641 43131 21644
rect 43073 21635 43131 21641
rect 43346 21632 43352 21644
rect 43404 21632 43410 21684
rect 29273 21607 29331 21613
rect 29273 21573 29285 21607
rect 29319 21604 29331 21607
rect 30438 21607 30496 21613
rect 30438 21604 30450 21607
rect 29319 21576 30450 21604
rect 29319 21573 29331 21576
rect 29273 21567 29331 21573
rect 30438 21573 30450 21576
rect 30484 21573 30496 21607
rect 30438 21567 30496 21573
rect 32950 21564 32956 21616
rect 33008 21604 33014 21616
rect 33566 21607 33624 21613
rect 33566 21604 33578 21607
rect 33008 21576 33578 21604
rect 33008 21564 33014 21576
rect 33566 21573 33578 21576
rect 33612 21573 33624 21607
rect 33566 21567 33624 21573
rect 37476 21576 37872 21604
rect 37476 21548 37504 21576
rect 27985 21539 28043 21545
rect 27985 21505 27997 21539
rect 28031 21505 28043 21539
rect 28626 21536 28632 21548
rect 28587 21508 28632 21536
rect 27985 21499 28043 21505
rect 28626 21496 28632 21508
rect 28684 21496 28690 21548
rect 28718 21496 28724 21548
rect 28776 21539 28782 21548
rect 28813 21542 28871 21548
rect 28813 21539 28825 21542
rect 28776 21511 28825 21539
rect 28776 21496 28782 21511
rect 28813 21508 28825 21511
rect 28859 21508 28871 21542
rect 28813 21502 28871 21508
rect 28905 21539 28963 21545
rect 28905 21505 28917 21539
rect 28951 21505 28963 21539
rect 28905 21499 28963 21505
rect 27614 21468 27620 21480
rect 25516 21440 27620 21468
rect 25133 21431 25191 21437
rect 27614 21428 27620 21440
rect 27672 21468 27678 21480
rect 27801 21471 27859 21477
rect 27801 21468 27813 21471
rect 27672 21440 27813 21468
rect 27672 21428 27678 21440
rect 27801 21437 27813 21440
rect 27847 21437 27859 21471
rect 28920 21468 28948 21499
rect 28994 21496 29000 21548
rect 29052 21545 29058 21548
rect 29052 21539 29101 21545
rect 29052 21505 29055 21539
rect 29089 21505 29101 21539
rect 29052 21499 29101 21505
rect 29052 21496 29058 21499
rect 29362 21496 29368 21548
rect 29420 21536 29426 21548
rect 30193 21539 30251 21545
rect 30193 21536 30205 21539
rect 29420 21508 30205 21536
rect 29420 21496 29426 21508
rect 30193 21505 30205 21508
rect 30239 21505 30251 21539
rect 30193 21499 30251 21505
rect 30282 21496 30288 21548
rect 30340 21536 30346 21548
rect 32306 21536 32312 21548
rect 30340 21508 32312 21536
rect 30340 21496 30346 21508
rect 32306 21496 32312 21508
rect 32364 21496 32370 21548
rect 32398 21496 32404 21548
rect 32456 21536 32462 21548
rect 33042 21536 33048 21548
rect 32456 21508 33048 21536
rect 32456 21496 32462 21508
rect 33042 21496 33048 21508
rect 33100 21536 33106 21548
rect 33321 21539 33379 21545
rect 33321 21536 33333 21539
rect 33100 21508 33333 21536
rect 33100 21496 33106 21508
rect 33321 21505 33333 21508
rect 33367 21505 33379 21539
rect 33321 21499 33379 21505
rect 34422 21496 34428 21548
rect 34480 21536 34486 21548
rect 35437 21539 35495 21545
rect 35437 21536 35449 21539
rect 34480 21508 35449 21536
rect 34480 21496 34486 21508
rect 35437 21505 35449 21508
rect 35483 21536 35495 21539
rect 37458 21536 37464 21548
rect 35483 21508 37464 21536
rect 35483 21505 35495 21508
rect 35437 21499 35495 21505
rect 37458 21496 37464 21508
rect 37516 21496 37522 21548
rect 37553 21539 37611 21545
rect 37553 21505 37565 21539
rect 37599 21505 37611 21539
rect 37734 21536 37740 21548
rect 37695 21508 37740 21536
rect 37553 21499 37611 21505
rect 29178 21468 29184 21480
rect 28920 21440 29184 21468
rect 27801 21431 27859 21437
rect 29178 21428 29184 21440
rect 29236 21428 29242 21480
rect 34698 21428 34704 21480
rect 34756 21468 34762 21480
rect 35161 21471 35219 21477
rect 35161 21468 35173 21471
rect 34756 21440 35173 21468
rect 34756 21428 34762 21440
rect 35161 21437 35173 21440
rect 35207 21437 35219 21471
rect 37274 21468 37280 21480
rect 35161 21431 35219 21437
rect 36280 21440 37280 21468
rect 7300 21372 9444 21400
rect 7300 21344 7328 21372
rect 9582 21360 9588 21412
rect 9640 21400 9646 21412
rect 17586 21400 17592 21412
rect 9640 21372 11836 21400
rect 9640 21360 9646 21372
rect 4249 21335 4307 21341
rect 4249 21301 4261 21335
rect 4295 21332 4307 21335
rect 4614 21332 4620 21344
rect 4295 21304 4620 21332
rect 4295 21301 4307 21304
rect 4249 21295 4307 21301
rect 4614 21292 4620 21304
rect 4672 21292 4678 21344
rect 7282 21292 7288 21344
rect 7340 21292 7346 21344
rect 7745 21335 7803 21341
rect 7745 21301 7757 21335
rect 7791 21332 7803 21335
rect 8386 21332 8392 21344
rect 7791 21304 8392 21332
rect 7791 21301 7803 21304
rect 7745 21295 7803 21301
rect 8386 21292 8392 21304
rect 8444 21292 8450 21344
rect 9674 21332 9680 21344
rect 9635 21304 9680 21332
rect 9674 21292 9680 21304
rect 9732 21292 9738 21344
rect 10226 21332 10232 21344
rect 10187 21304 10232 21332
rect 10226 21292 10232 21304
rect 10284 21292 10290 21344
rect 11517 21335 11575 21341
rect 11517 21301 11529 21335
rect 11563 21332 11575 21335
rect 11698 21332 11704 21344
rect 11563 21304 11704 21332
rect 11563 21301 11575 21304
rect 11517 21295 11575 21301
rect 11698 21292 11704 21304
rect 11756 21292 11762 21344
rect 11808 21332 11836 21372
rect 12075 21372 17592 21400
rect 12075 21332 12103 21372
rect 17586 21360 17592 21372
rect 17644 21360 17650 21412
rect 19334 21360 19340 21412
rect 19392 21400 19398 21412
rect 20254 21400 20260 21412
rect 19392 21372 20260 21400
rect 19392 21360 19398 21372
rect 20254 21360 20260 21372
rect 20312 21360 20318 21412
rect 22186 21360 22192 21412
rect 22244 21400 22250 21412
rect 30098 21400 30104 21412
rect 22244 21372 30104 21400
rect 22244 21360 22250 21372
rect 30098 21360 30104 21372
rect 30156 21360 30162 21412
rect 11808 21304 12103 21332
rect 14826 21292 14832 21344
rect 14884 21332 14890 21344
rect 15838 21332 15844 21344
rect 14884 21304 15844 21332
rect 14884 21292 14890 21304
rect 15838 21292 15844 21304
rect 15896 21292 15902 21344
rect 16574 21292 16580 21344
rect 16632 21332 16638 21344
rect 17310 21332 17316 21344
rect 16632 21304 17316 21332
rect 16632 21292 16638 21304
rect 17310 21292 17316 21304
rect 17368 21292 17374 21344
rect 19797 21335 19855 21341
rect 19797 21301 19809 21335
rect 19843 21332 19855 21335
rect 20070 21332 20076 21344
rect 19843 21304 20076 21332
rect 19843 21301 19855 21304
rect 19797 21295 19855 21301
rect 20070 21292 20076 21304
rect 20128 21292 20134 21344
rect 21910 21292 21916 21344
rect 21968 21332 21974 21344
rect 22097 21335 22155 21341
rect 22097 21332 22109 21335
rect 21968 21304 22109 21332
rect 21968 21292 21974 21304
rect 22097 21301 22109 21304
rect 22143 21301 22155 21335
rect 24026 21332 24032 21344
rect 23987 21304 24032 21332
rect 22097 21295 22155 21301
rect 24026 21292 24032 21304
rect 24084 21292 24090 21344
rect 27798 21332 27804 21344
rect 27759 21304 27804 21332
rect 27798 21292 27804 21304
rect 27856 21292 27862 21344
rect 28169 21335 28227 21341
rect 28169 21301 28181 21335
rect 28215 21332 28227 21335
rect 30834 21332 30840 21344
rect 28215 21304 30840 21332
rect 28215 21301 28227 21304
rect 28169 21295 28227 21301
rect 30834 21292 30840 21304
rect 30892 21292 30898 21344
rect 30926 21292 30932 21344
rect 30984 21332 30990 21344
rect 31573 21335 31631 21341
rect 31573 21332 31585 21335
rect 30984 21304 31585 21332
rect 30984 21292 30990 21304
rect 31573 21301 31585 21304
rect 31619 21301 31631 21335
rect 31573 21295 31631 21301
rect 32493 21335 32551 21341
rect 32493 21301 32505 21335
rect 32539 21332 32551 21335
rect 32766 21332 32772 21344
rect 32539 21304 32772 21332
rect 32539 21301 32551 21304
rect 32493 21295 32551 21301
rect 32766 21292 32772 21304
rect 32824 21292 32830 21344
rect 33594 21292 33600 21344
rect 33652 21332 33658 21344
rect 36280 21332 36308 21440
rect 37274 21428 37280 21440
rect 37332 21468 37338 21480
rect 37568 21468 37596 21499
rect 37734 21496 37740 21508
rect 37792 21496 37798 21548
rect 37844 21545 37872 21576
rect 42518 21564 42524 21616
rect 42576 21604 42582 21616
rect 42576 21576 42932 21604
rect 42576 21564 42582 21576
rect 37829 21539 37887 21545
rect 37829 21505 37841 21539
rect 37875 21505 37887 21539
rect 37829 21499 37887 21505
rect 37921 21539 37979 21545
rect 37921 21505 37933 21539
rect 37967 21505 37979 21539
rect 41230 21536 41236 21548
rect 41191 21508 41236 21536
rect 37921 21499 37979 21505
rect 37936 21468 37964 21499
rect 41230 21496 41236 21508
rect 41288 21496 41294 21548
rect 41509 21539 41567 21545
rect 41509 21505 41521 21539
rect 41555 21536 41567 21539
rect 41598 21536 41604 21548
rect 41555 21508 41604 21536
rect 41555 21505 41567 21508
rect 41509 21499 41567 21505
rect 41598 21496 41604 21508
rect 41656 21496 41662 21548
rect 42426 21536 42432 21548
rect 42387 21508 42432 21536
rect 42426 21496 42432 21508
rect 42484 21496 42490 21548
rect 42613 21539 42671 21545
rect 42613 21505 42625 21539
rect 42659 21536 42671 21539
rect 42794 21536 42800 21548
rect 42659 21508 42800 21536
rect 42659 21505 42671 21508
rect 42613 21499 42671 21505
rect 42794 21496 42800 21508
rect 42852 21496 42858 21548
rect 42904 21545 42932 21576
rect 42889 21539 42947 21545
rect 42889 21505 42901 21539
rect 42935 21505 42947 21539
rect 42889 21499 42947 21505
rect 41414 21468 41420 21480
rect 37332 21440 37596 21468
rect 37844 21440 37964 21468
rect 41375 21440 41420 21468
rect 37332 21428 37338 21440
rect 37844 21400 37872 21440
rect 41414 21428 41420 21440
rect 41472 21428 41478 21480
rect 36648 21372 37872 21400
rect 33652 21304 36308 21332
rect 33652 21292 33658 21304
rect 36354 21292 36360 21344
rect 36412 21332 36418 21344
rect 36648 21341 36676 21372
rect 36633 21335 36691 21341
rect 36633 21332 36645 21335
rect 36412 21304 36645 21332
rect 36412 21292 36418 21304
rect 36633 21301 36645 21304
rect 36679 21301 36691 21335
rect 36633 21295 36691 21301
rect 37826 21292 37832 21344
rect 37884 21332 37890 21344
rect 38657 21335 38715 21341
rect 38657 21332 38669 21335
rect 37884 21304 38669 21332
rect 37884 21292 37890 21304
rect 38657 21301 38669 21304
rect 38703 21301 38715 21335
rect 38657 21295 38715 21301
rect 41509 21335 41567 21341
rect 41509 21301 41521 21335
rect 41555 21332 41567 21335
rect 41598 21332 41604 21344
rect 41555 21304 41604 21332
rect 41555 21301 41567 21304
rect 41509 21295 41567 21301
rect 41598 21292 41604 21304
rect 41656 21332 41662 21344
rect 41874 21332 41880 21344
rect 41656 21304 41880 21332
rect 41656 21292 41662 21304
rect 41874 21292 41880 21304
rect 41932 21292 41938 21344
rect 1104 21242 68816 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 65654 21242
rect 65706 21190 65718 21242
rect 65770 21190 65782 21242
rect 65834 21190 65846 21242
rect 65898 21190 65910 21242
rect 65962 21190 68816 21242
rect 1104 21168 68816 21190
rect 2603 21131 2661 21137
rect 2603 21097 2615 21131
rect 2649 21128 2661 21131
rect 6546 21128 6552 21140
rect 2649 21100 6552 21128
rect 2649 21097 2661 21100
rect 2603 21091 2661 21097
rect 6546 21088 6552 21100
rect 6604 21088 6610 21140
rect 6638 21088 6644 21140
rect 6696 21128 6702 21140
rect 6825 21131 6883 21137
rect 6825 21128 6837 21131
rect 6696 21100 6837 21128
rect 6696 21088 6702 21100
rect 6825 21097 6837 21100
rect 6871 21097 6883 21131
rect 6825 21091 6883 21097
rect 7742 21088 7748 21140
rect 7800 21128 7806 21140
rect 7929 21131 7987 21137
rect 7929 21128 7941 21131
rect 7800 21100 7941 21128
rect 7800 21088 7806 21100
rect 7929 21097 7941 21100
rect 7975 21097 7987 21131
rect 7929 21091 7987 21097
rect 8389 21131 8447 21137
rect 8389 21097 8401 21131
rect 8435 21097 8447 21131
rect 8389 21091 8447 21097
rect 3234 21060 3240 21072
rect 3147 21032 3240 21060
rect 3234 21020 3240 21032
rect 3292 21060 3298 21072
rect 3418 21060 3424 21072
rect 3292 21032 3424 21060
rect 3292 21020 3298 21032
rect 3418 21020 3424 21032
rect 3476 21060 3482 21072
rect 7282 21060 7288 21072
rect 3476 21032 7288 21060
rect 3476 21020 3482 21032
rect 7282 21020 7288 21032
rect 7340 21020 7346 21072
rect 8404 21060 8432 21091
rect 8754 21088 8760 21140
rect 8812 21128 8818 21140
rect 16669 21131 16727 21137
rect 8812 21100 16620 21128
rect 8812 21088 8818 21100
rect 8478 21060 8484 21072
rect 8391 21032 8484 21060
rect 8478 21020 8484 21032
rect 8536 21060 8542 21072
rect 9306 21060 9312 21072
rect 8536 21032 9312 21060
rect 8536 21020 8542 21032
rect 9306 21020 9312 21032
rect 9364 21020 9370 21072
rect 16592 21060 16620 21100
rect 16669 21097 16681 21131
rect 16715 21128 16727 21131
rect 16850 21128 16856 21140
rect 16715 21100 16856 21128
rect 16715 21097 16727 21100
rect 16669 21091 16727 21097
rect 16850 21088 16856 21100
rect 16908 21088 16914 21140
rect 17126 21088 17132 21140
rect 17184 21128 17190 21140
rect 17681 21131 17739 21137
rect 17681 21128 17693 21131
rect 17184 21100 17693 21128
rect 17184 21088 17190 21100
rect 17681 21097 17693 21100
rect 17727 21097 17739 21131
rect 17681 21091 17739 21097
rect 20438 21088 20444 21140
rect 20496 21128 20502 21140
rect 21453 21131 21511 21137
rect 21453 21128 21465 21131
rect 20496 21100 21465 21128
rect 20496 21088 20502 21100
rect 21453 21097 21465 21100
rect 21499 21097 21511 21131
rect 27706 21128 27712 21140
rect 21453 21091 21511 21097
rect 22066 21100 27292 21128
rect 27667 21100 27712 21128
rect 21358 21060 21364 21072
rect 16592 21032 21364 21060
rect 21358 21020 21364 21032
rect 21416 21020 21422 21072
rect 21910 21020 21916 21072
rect 21968 21060 21974 21072
rect 22066 21060 22094 21100
rect 21968 21032 22094 21060
rect 24397 21063 24455 21069
rect 21968 21020 21974 21032
rect 24397 21029 24409 21063
rect 24443 21060 24455 21063
rect 24670 21060 24676 21072
rect 24443 21032 24676 21060
rect 24443 21029 24455 21032
rect 24397 21023 24455 21029
rect 24670 21020 24676 21032
rect 24728 21020 24734 21072
rect 27264 21060 27292 21100
rect 27706 21088 27712 21100
rect 27764 21088 27770 21140
rect 28261 21131 28319 21137
rect 28261 21097 28273 21131
rect 28307 21128 28319 21131
rect 28718 21128 28724 21140
rect 28307 21100 28724 21128
rect 28307 21097 28319 21100
rect 28261 21091 28319 21097
rect 28718 21088 28724 21100
rect 28776 21088 28782 21140
rect 28902 21088 28908 21140
rect 28960 21128 28966 21140
rect 29914 21128 29920 21140
rect 28960 21100 29920 21128
rect 28960 21088 28966 21100
rect 29914 21088 29920 21100
rect 29972 21088 29978 21140
rect 30101 21131 30159 21137
rect 30101 21097 30113 21131
rect 30147 21128 30159 21131
rect 30561 21131 30619 21137
rect 30561 21128 30573 21131
rect 30147 21100 30573 21128
rect 30147 21097 30159 21100
rect 30101 21091 30159 21097
rect 30561 21097 30573 21100
rect 30607 21097 30619 21131
rect 30561 21091 30619 21097
rect 31021 21131 31079 21137
rect 31021 21097 31033 21131
rect 31067 21128 31079 21131
rect 33686 21128 33692 21140
rect 31067 21100 33692 21128
rect 31067 21097 31079 21100
rect 31021 21091 31079 21097
rect 33686 21088 33692 21100
rect 33744 21088 33750 21140
rect 34054 21088 34060 21140
rect 34112 21128 34118 21140
rect 35713 21131 35771 21137
rect 35713 21128 35725 21131
rect 34112 21100 35725 21128
rect 34112 21088 34118 21100
rect 35713 21097 35725 21100
rect 35759 21097 35771 21131
rect 35713 21091 35771 21097
rect 37553 21131 37611 21137
rect 37553 21097 37565 21131
rect 37599 21128 37611 21131
rect 37734 21128 37740 21140
rect 37599 21100 37740 21128
rect 37599 21097 37611 21100
rect 37553 21091 37611 21097
rect 37734 21088 37740 21100
rect 37792 21088 37798 21140
rect 38010 21088 38016 21140
rect 38068 21128 38074 21140
rect 38289 21131 38347 21137
rect 38289 21128 38301 21131
rect 38068 21100 38301 21128
rect 38068 21088 38074 21100
rect 38289 21097 38301 21100
rect 38335 21097 38347 21131
rect 38289 21091 38347 21097
rect 38657 21131 38715 21137
rect 38657 21097 38669 21131
rect 38703 21128 38715 21131
rect 42426 21128 42432 21140
rect 38703 21100 42432 21128
rect 38703 21097 38715 21100
rect 38657 21091 38715 21097
rect 42426 21088 42432 21100
rect 42484 21088 42490 21140
rect 35526 21060 35532 21072
rect 27264 21032 35532 21060
rect 35526 21020 35532 21032
rect 35584 21060 35590 21072
rect 36173 21063 36231 21069
rect 35584 21032 36124 21060
rect 35584 21020 35590 21032
rect 4614 20952 4620 21004
rect 4672 20992 4678 21004
rect 6914 20992 6920 21004
rect 4672 20964 6920 20992
rect 4672 20952 4678 20964
rect 6914 20952 6920 20964
rect 6972 20952 6978 21004
rect 9030 20992 9036 21004
rect 7484 20964 9036 20992
rect 1486 20884 1492 20936
rect 1544 20924 1550 20936
rect 1581 20927 1639 20933
rect 1581 20924 1593 20927
rect 1544 20896 1593 20924
rect 1544 20884 1550 20896
rect 1581 20893 1593 20896
rect 1627 20893 1639 20927
rect 1854 20924 1860 20936
rect 1815 20896 1860 20924
rect 1581 20887 1639 20893
rect 1854 20884 1860 20896
rect 1912 20884 1918 20936
rect 7081 20927 7139 20933
rect 7081 20924 7093 20927
rect 7024 20896 7093 20924
rect 5534 20748 5540 20800
rect 5592 20788 5598 20800
rect 5629 20791 5687 20797
rect 5629 20788 5641 20791
rect 5592 20760 5641 20788
rect 5592 20748 5598 20760
rect 5629 20757 5641 20760
rect 5675 20788 5687 20791
rect 5718 20788 5724 20800
rect 5675 20760 5724 20788
rect 5675 20757 5687 20760
rect 5629 20751 5687 20757
rect 5718 20748 5724 20760
rect 5776 20748 5782 20800
rect 6365 20791 6423 20797
rect 6365 20757 6377 20791
rect 6411 20788 6423 20791
rect 7024 20788 7052 20896
rect 7081 20893 7093 20896
rect 7127 20893 7139 20927
rect 7081 20887 7139 20893
rect 7193 20927 7251 20933
rect 7193 20893 7205 20927
rect 7239 20893 7251 20927
rect 7193 20887 7251 20893
rect 7221 20856 7249 20887
rect 7282 20884 7288 20936
rect 7340 20933 7346 20936
rect 7484 20933 7512 20964
rect 9030 20952 9036 20964
rect 9088 20952 9094 21004
rect 18782 20992 18788 21004
rect 17880 20964 18788 20992
rect 7340 20924 7348 20933
rect 7469 20927 7527 20933
rect 7340 20896 7385 20924
rect 7340 20887 7348 20896
rect 7469 20893 7481 20927
rect 7515 20893 7527 20927
rect 8110 20924 8116 20936
rect 8071 20896 8116 20924
rect 7469 20887 7527 20893
rect 7340 20884 7346 20887
rect 8110 20884 8116 20896
rect 8168 20884 8174 20936
rect 8205 20927 8263 20933
rect 8205 20893 8217 20927
rect 8251 20924 8263 20927
rect 8294 20924 8300 20936
rect 8251 20896 8300 20924
rect 8251 20893 8263 20896
rect 8205 20887 8263 20893
rect 7834 20856 7840 20868
rect 7221 20828 7840 20856
rect 7834 20816 7840 20828
rect 7892 20816 7898 20868
rect 7742 20788 7748 20800
rect 6411 20760 7748 20788
rect 6411 20757 6423 20760
rect 6365 20751 6423 20757
rect 7742 20748 7748 20760
rect 7800 20748 7806 20800
rect 8220 20788 8248 20887
rect 8294 20884 8300 20896
rect 8352 20884 8358 20936
rect 8662 20884 8668 20936
rect 8720 20924 8726 20936
rect 9585 20927 9643 20933
rect 9585 20924 9597 20927
rect 8720 20896 9597 20924
rect 8720 20884 8726 20896
rect 9585 20893 9597 20896
rect 9631 20893 9643 20927
rect 9585 20887 9643 20893
rect 9674 20884 9680 20936
rect 9732 20924 9738 20936
rect 9841 20927 9899 20933
rect 9841 20924 9853 20927
rect 9732 20896 9853 20924
rect 9732 20884 9738 20896
rect 9841 20893 9853 20896
rect 9887 20893 9899 20927
rect 11606 20924 11612 20936
rect 11567 20896 11612 20924
rect 9841 20887 9899 20893
rect 11606 20884 11612 20896
rect 11664 20884 11670 20936
rect 11698 20884 11704 20936
rect 11756 20924 11762 20936
rect 11865 20927 11923 20933
rect 11865 20924 11877 20927
rect 11756 20896 11877 20924
rect 11756 20884 11762 20896
rect 11865 20893 11877 20896
rect 11911 20893 11923 20927
rect 11865 20887 11923 20893
rect 13998 20884 14004 20936
rect 14056 20924 14062 20936
rect 14093 20927 14151 20933
rect 14093 20924 14105 20927
rect 14056 20896 14105 20924
rect 14056 20884 14062 20896
rect 14093 20893 14105 20896
rect 14139 20893 14151 20927
rect 14369 20927 14427 20933
rect 14369 20924 14381 20927
rect 14093 20887 14151 20893
rect 14200 20896 14381 20924
rect 8386 20856 8392 20868
rect 8299 20828 8392 20856
rect 8386 20816 8392 20828
rect 8444 20856 8450 20868
rect 8846 20856 8852 20868
rect 8444 20828 8852 20856
rect 8444 20816 8450 20828
rect 8846 20816 8852 20828
rect 8904 20816 8910 20868
rect 8956 20828 10456 20856
rect 8956 20788 8984 20828
rect 10428 20800 10456 20828
rect 10502 20816 10508 20868
rect 10560 20856 10566 20868
rect 13449 20859 13507 20865
rect 13449 20856 13461 20859
rect 10560 20828 13461 20856
rect 10560 20816 10566 20828
rect 13449 20825 13461 20828
rect 13495 20856 13507 20859
rect 14200 20856 14228 20896
rect 14369 20893 14381 20896
rect 14415 20893 14427 20927
rect 14369 20887 14427 20893
rect 14461 20927 14519 20933
rect 14461 20893 14473 20927
rect 14507 20924 14519 20927
rect 14642 20924 14648 20936
rect 14507 20896 14648 20924
rect 14507 20893 14519 20896
rect 14461 20887 14519 20893
rect 14642 20884 14648 20896
rect 14700 20884 14706 20936
rect 15286 20924 15292 20936
rect 15247 20896 15292 20924
rect 15286 20884 15292 20896
rect 15344 20884 15350 20936
rect 15556 20927 15614 20933
rect 15556 20893 15568 20927
rect 15602 20924 15614 20927
rect 15930 20924 15936 20936
rect 15602 20896 15936 20924
rect 15602 20893 15614 20896
rect 15556 20887 15614 20893
rect 15930 20884 15936 20896
rect 15988 20884 15994 20936
rect 17880 20933 17908 20964
rect 18782 20952 18788 20964
rect 18840 20952 18846 21004
rect 18874 20952 18880 21004
rect 18932 20992 18938 21004
rect 18932 20964 19564 20992
rect 18932 20952 18938 20964
rect 17865 20927 17923 20933
rect 17865 20893 17877 20927
rect 17911 20893 17923 20927
rect 17865 20887 17923 20893
rect 17954 20884 17960 20936
rect 18012 20924 18018 20936
rect 18138 20924 18144 20936
rect 18012 20896 18057 20924
rect 18099 20896 18144 20924
rect 18012 20884 18018 20896
rect 18138 20884 18144 20896
rect 18196 20884 18202 20936
rect 18230 20884 18236 20936
rect 18288 20924 18294 20936
rect 19426 20933 19432 20936
rect 19424 20924 19432 20933
rect 18288 20896 18333 20924
rect 19387 20896 19432 20924
rect 18288 20884 18294 20896
rect 19424 20887 19432 20896
rect 19426 20884 19432 20887
rect 19484 20884 19490 20936
rect 19536 20933 19564 20964
rect 20162 20952 20168 21004
rect 20220 20992 20226 21004
rect 20622 20992 20628 21004
rect 20220 20964 20628 20992
rect 20220 20952 20226 20964
rect 20622 20952 20628 20964
rect 20680 20952 20686 21004
rect 21818 20992 21824 21004
rect 21652 20964 21824 20992
rect 19521 20927 19579 20933
rect 19521 20893 19533 20927
rect 19567 20893 19579 20927
rect 19521 20887 19579 20893
rect 19796 20927 19854 20933
rect 19796 20893 19808 20927
rect 19842 20893 19854 20927
rect 19796 20887 19854 20893
rect 19889 20927 19947 20933
rect 19889 20893 19901 20927
rect 19935 20924 19947 20927
rect 21542 20924 21548 20936
rect 19935 20896 21548 20924
rect 19935 20893 19947 20896
rect 19889 20887 19947 20893
rect 13495 20828 14228 20856
rect 14277 20859 14335 20865
rect 13495 20825 13507 20828
rect 13449 20819 13507 20825
rect 14277 20825 14289 20859
rect 14323 20856 14335 20859
rect 19150 20856 19156 20868
rect 14323 20828 19156 20856
rect 14323 20825 14335 20828
rect 14277 20819 14335 20825
rect 19150 20816 19156 20828
rect 19208 20816 19214 20868
rect 19334 20816 19340 20868
rect 19392 20856 19398 20868
rect 19613 20859 19671 20865
rect 19613 20856 19625 20859
rect 19392 20828 19625 20856
rect 19392 20816 19398 20828
rect 19613 20825 19625 20828
rect 19659 20825 19671 20859
rect 19812 20856 19840 20887
rect 21542 20884 21548 20896
rect 21600 20884 21606 20936
rect 21652 20933 21680 20964
rect 21818 20952 21824 20964
rect 21876 20992 21882 21004
rect 22649 20995 22707 21001
rect 22649 20992 22661 20995
rect 21876 20964 22661 20992
rect 21876 20952 21882 20964
rect 22649 20961 22661 20964
rect 22695 20961 22707 20995
rect 22649 20955 22707 20961
rect 22925 20995 22983 21001
rect 22925 20961 22937 20995
rect 22971 20992 22983 20995
rect 24762 20992 24768 21004
rect 22971 20964 24768 20992
rect 22971 20961 22983 20964
rect 22925 20955 22983 20961
rect 21637 20927 21695 20933
rect 21637 20893 21649 20927
rect 21683 20893 21695 20927
rect 21637 20887 21695 20893
rect 20622 20856 20628 20868
rect 19812 20828 20628 20856
rect 19613 20819 19671 20825
rect 20622 20816 20628 20828
rect 20680 20816 20686 20868
rect 8220 20760 8984 20788
rect 9033 20791 9091 20797
rect 9033 20757 9045 20791
rect 9079 20788 9091 20791
rect 9398 20788 9404 20800
rect 9079 20760 9404 20788
rect 9079 20757 9091 20760
rect 9033 20751 9091 20757
rect 9398 20748 9404 20760
rect 9456 20748 9462 20800
rect 10410 20748 10416 20800
rect 10468 20788 10474 20800
rect 10965 20791 11023 20797
rect 10965 20788 10977 20791
rect 10468 20760 10977 20788
rect 10468 20748 10474 20760
rect 10965 20757 10977 20760
rect 11011 20757 11023 20791
rect 12986 20788 12992 20800
rect 12947 20760 12992 20788
rect 10965 20751 11023 20757
rect 12986 20748 12992 20760
rect 13044 20748 13050 20800
rect 14645 20791 14703 20797
rect 14645 20757 14657 20791
rect 14691 20788 14703 20791
rect 15010 20788 15016 20800
rect 14691 20760 15016 20788
rect 14691 20757 14703 20760
rect 14645 20751 14703 20757
rect 15010 20748 15016 20760
rect 15068 20748 15074 20800
rect 17126 20788 17132 20800
rect 17087 20760 17132 20788
rect 17126 20748 17132 20760
rect 17184 20748 17190 20800
rect 18414 20748 18420 20800
rect 18472 20788 18478 20800
rect 19245 20791 19303 20797
rect 19245 20788 19257 20791
rect 18472 20760 19257 20788
rect 18472 20748 18478 20760
rect 19245 20757 19257 20760
rect 19291 20757 19303 20791
rect 19245 20751 19303 20757
rect 19794 20748 19800 20800
rect 19852 20788 19858 20800
rect 20717 20791 20775 20797
rect 20717 20788 20729 20791
rect 19852 20760 20729 20788
rect 19852 20748 19858 20760
rect 20717 20757 20729 20760
rect 20763 20788 20775 20791
rect 20898 20788 20904 20800
rect 20763 20760 20904 20788
rect 20763 20757 20775 20760
rect 20717 20751 20775 20757
rect 20898 20748 20904 20760
rect 20956 20748 20962 20800
rect 21652 20788 21680 20887
rect 21726 20884 21732 20936
rect 21784 20924 21790 20936
rect 22002 20924 22008 20936
rect 21784 20896 21829 20924
rect 21963 20896 22008 20924
rect 21784 20884 21790 20896
rect 22002 20884 22008 20896
rect 22060 20884 22066 20936
rect 24540 20933 24568 20964
rect 24762 20952 24768 20964
rect 24820 20952 24826 21004
rect 27338 20952 27344 21004
rect 27396 20992 27402 21004
rect 30466 20992 30472 21004
rect 27396 20964 29684 20992
rect 27396 20952 27402 20964
rect 24535 20927 24593 20933
rect 24535 20893 24547 20927
rect 24581 20893 24593 20927
rect 24535 20887 24593 20893
rect 24949 20927 25007 20933
rect 24949 20893 24961 20927
rect 24995 20924 25007 20927
rect 26234 20924 26240 20936
rect 24995 20896 26240 20924
rect 24995 20893 25007 20896
rect 24949 20887 25007 20893
rect 26234 20884 26240 20896
rect 26292 20884 26298 20936
rect 26329 20927 26387 20933
rect 26329 20893 26341 20927
rect 26375 20924 26387 20927
rect 28166 20924 28172 20936
rect 26375 20896 26924 20924
rect 28127 20896 28172 20924
rect 26375 20893 26387 20896
rect 26329 20887 26387 20893
rect 21821 20859 21879 20865
rect 21821 20825 21833 20859
rect 21867 20856 21879 20859
rect 22462 20856 22468 20868
rect 21867 20828 22468 20856
rect 21867 20825 21879 20828
rect 21821 20819 21879 20825
rect 22462 20816 22468 20828
rect 22520 20816 22526 20868
rect 23750 20816 23756 20868
rect 23808 20856 23814 20868
rect 24673 20859 24731 20865
rect 24673 20856 24685 20859
rect 23808 20828 24685 20856
rect 23808 20816 23814 20828
rect 24673 20825 24685 20828
rect 24719 20825 24731 20859
rect 24673 20819 24731 20825
rect 24765 20859 24823 20865
rect 24765 20825 24777 20859
rect 24811 20856 24823 20859
rect 25130 20856 25136 20868
rect 24811 20828 25136 20856
rect 24811 20825 24823 20828
rect 24765 20819 24823 20825
rect 21726 20788 21732 20800
rect 21652 20760 21732 20788
rect 21726 20748 21732 20760
rect 21784 20748 21790 20800
rect 23014 20748 23020 20800
rect 23072 20788 23078 20800
rect 24780 20788 24808 20819
rect 25130 20816 25136 20828
rect 25188 20816 25194 20868
rect 25406 20856 25412 20868
rect 25367 20828 25412 20856
rect 25406 20816 25412 20828
rect 25464 20816 25470 20868
rect 25590 20856 25596 20868
rect 25551 20828 25596 20856
rect 25590 20816 25596 20828
rect 25648 20816 25654 20868
rect 26142 20816 26148 20868
rect 26200 20856 26206 20868
rect 26574 20859 26632 20865
rect 26574 20856 26586 20859
rect 26200 20828 26586 20856
rect 26200 20816 26206 20828
rect 26574 20825 26586 20828
rect 26620 20825 26632 20859
rect 26896 20856 26924 20896
rect 28166 20884 28172 20896
rect 28224 20884 28230 20936
rect 28353 20927 28411 20933
rect 28353 20893 28365 20927
rect 28399 20924 28411 20927
rect 28902 20924 28908 20936
rect 28399 20896 28908 20924
rect 28399 20893 28411 20896
rect 28353 20887 28411 20893
rect 28902 20884 28908 20896
rect 28960 20884 28966 20936
rect 28997 20927 29055 20933
rect 28997 20893 29009 20927
rect 29043 20924 29055 20927
rect 29086 20924 29092 20936
rect 29043 20896 29092 20924
rect 29043 20893 29055 20896
rect 28997 20887 29055 20893
rect 29086 20884 29092 20896
rect 29144 20884 29150 20936
rect 29546 20924 29552 20936
rect 29507 20896 29552 20924
rect 29546 20884 29552 20896
rect 29604 20884 29610 20936
rect 29656 20933 29684 20964
rect 29840 20964 30472 20992
rect 29840 20933 29868 20964
rect 30466 20952 30472 20964
rect 30524 20952 30530 21004
rect 30742 20992 30748 21004
rect 30703 20964 30748 20992
rect 30742 20952 30748 20964
rect 30800 20952 30806 21004
rect 32232 20964 33732 20992
rect 29641 20927 29699 20933
rect 29641 20893 29653 20927
rect 29687 20924 29699 20927
rect 29825 20927 29883 20933
rect 29687 20896 29776 20924
rect 29687 20893 29699 20896
rect 29641 20887 29699 20893
rect 28442 20856 28448 20868
rect 26896 20828 28448 20856
rect 26574 20819 26632 20825
rect 28442 20816 28448 20828
rect 28500 20816 28506 20868
rect 29748 20856 29776 20896
rect 29825 20893 29837 20927
rect 29871 20893 29883 20927
rect 29825 20887 29883 20893
rect 29914 20884 29920 20936
rect 29972 20924 29978 20936
rect 29972 20896 30017 20924
rect 29972 20884 29978 20896
rect 30098 20884 30104 20936
rect 30156 20924 30162 20936
rect 30834 20924 30840 20936
rect 30156 20896 30696 20924
rect 30795 20896 30840 20924
rect 30156 20884 30162 20896
rect 30374 20856 30380 20868
rect 29748 20828 30380 20856
rect 30374 20816 30380 20828
rect 30432 20816 30438 20868
rect 30558 20856 30564 20868
rect 30519 20828 30564 20856
rect 30558 20816 30564 20828
rect 30616 20816 30622 20868
rect 30668 20856 30696 20896
rect 30834 20884 30840 20896
rect 30892 20884 30898 20936
rect 32122 20884 32128 20936
rect 32180 20924 32186 20936
rect 32232 20933 32260 20964
rect 33704 20936 33732 20964
rect 34330 20952 34336 21004
rect 34388 20992 34394 21004
rect 35710 20992 35716 21004
rect 34388 20964 35716 20992
rect 34388 20952 34394 20964
rect 35710 20952 35716 20964
rect 35768 20992 35774 21004
rect 35805 20995 35863 21001
rect 35805 20992 35817 20995
rect 35768 20964 35817 20992
rect 35768 20952 35774 20964
rect 35805 20961 35817 20964
rect 35851 20961 35863 20995
rect 36096 20992 36124 21032
rect 36173 21029 36185 21063
rect 36219 21060 36231 21063
rect 41414 21060 41420 21072
rect 36219 21032 41420 21060
rect 36219 21029 36231 21032
rect 36173 21023 36231 21029
rect 41414 21020 41420 21032
rect 41472 21020 41478 21072
rect 36096 20964 36492 20992
rect 35805 20955 35863 20961
rect 32217 20927 32275 20933
rect 32217 20924 32229 20927
rect 32180 20896 32229 20924
rect 32180 20884 32186 20896
rect 32217 20893 32229 20896
rect 32263 20893 32275 20927
rect 32217 20887 32275 20893
rect 32401 20927 32459 20933
rect 32401 20893 32413 20927
rect 32447 20924 32459 20927
rect 32490 20924 32496 20936
rect 32447 20896 32496 20924
rect 32447 20893 32459 20896
rect 32401 20887 32459 20893
rect 32416 20856 32444 20887
rect 32490 20884 32496 20896
rect 32548 20884 32554 20936
rect 33318 20924 33324 20936
rect 33279 20896 33324 20924
rect 33318 20884 33324 20896
rect 33376 20884 33382 20936
rect 33594 20924 33600 20936
rect 33555 20896 33600 20924
rect 33594 20884 33600 20896
rect 33652 20884 33658 20936
rect 33686 20884 33692 20936
rect 33744 20924 33750 20936
rect 34701 20927 34759 20933
rect 34701 20924 34713 20927
rect 33744 20896 34713 20924
rect 33744 20884 33750 20896
rect 34701 20893 34713 20896
rect 34747 20893 34759 20927
rect 34701 20887 34759 20893
rect 35989 20927 36047 20933
rect 35989 20893 36001 20927
rect 36035 20924 36047 20927
rect 36078 20924 36084 20936
rect 36035 20896 36084 20924
rect 36035 20893 36047 20896
rect 35989 20887 36047 20893
rect 36078 20884 36084 20896
rect 36136 20884 36142 20936
rect 36464 20924 36492 20964
rect 36538 20952 36544 21004
rect 36596 20992 36602 21004
rect 38381 20995 38439 21001
rect 38381 20992 38393 20995
rect 36596 20964 38393 20992
rect 36596 20952 36602 20964
rect 38381 20961 38393 20964
rect 38427 20992 38439 20995
rect 40126 20992 40132 21004
rect 38427 20964 40132 20992
rect 38427 20961 38439 20964
rect 38381 20955 38439 20961
rect 40126 20952 40132 20964
rect 40184 20952 40190 21004
rect 41690 20952 41696 21004
rect 41748 20992 41754 21004
rect 41785 20995 41843 21001
rect 41785 20992 41797 20995
rect 41748 20964 41797 20992
rect 41748 20952 41754 20964
rect 41785 20961 41797 20964
rect 41831 20961 41843 20995
rect 41785 20955 41843 20961
rect 37369 20927 37427 20933
rect 37369 20924 37381 20927
rect 36464 20896 37381 20924
rect 37369 20893 37381 20896
rect 37415 20893 37427 20927
rect 38286 20924 38292 20936
rect 38247 20896 38292 20924
rect 37369 20887 37427 20893
rect 30668 20828 32444 20856
rect 35713 20859 35771 20865
rect 35713 20825 35725 20859
rect 35759 20856 35771 20859
rect 35802 20856 35808 20868
rect 35759 20828 35808 20856
rect 35759 20825 35771 20828
rect 35713 20819 35771 20825
rect 35802 20816 35808 20828
rect 35860 20816 35866 20868
rect 37185 20859 37243 20865
rect 37185 20856 37197 20859
rect 35912 20828 37197 20856
rect 23072 20760 24808 20788
rect 23072 20748 23078 20760
rect 25682 20748 25688 20800
rect 25740 20788 25746 20800
rect 25777 20791 25835 20797
rect 25777 20788 25789 20791
rect 25740 20760 25789 20788
rect 25740 20748 25746 20760
rect 25777 20757 25789 20760
rect 25823 20757 25835 20791
rect 25777 20751 25835 20757
rect 31665 20791 31723 20797
rect 31665 20757 31677 20791
rect 31711 20788 31723 20791
rect 31754 20788 31760 20800
rect 31711 20760 31760 20788
rect 31711 20757 31723 20760
rect 31665 20751 31723 20757
rect 31754 20748 31760 20760
rect 31812 20748 31818 20800
rect 32490 20748 32496 20800
rect 32548 20788 32554 20800
rect 32585 20791 32643 20797
rect 32585 20788 32597 20791
rect 32548 20760 32597 20788
rect 32548 20748 32554 20760
rect 32585 20757 32597 20760
rect 32631 20757 32643 20791
rect 32585 20751 32643 20757
rect 34885 20791 34943 20797
rect 34885 20757 34897 20791
rect 34931 20788 34943 20791
rect 35618 20788 35624 20800
rect 34931 20760 35624 20788
rect 34931 20757 34943 20760
rect 34885 20751 34943 20757
rect 35618 20748 35624 20760
rect 35676 20788 35682 20800
rect 35912 20788 35940 20828
rect 37185 20825 37197 20828
rect 37231 20825 37243 20859
rect 37384 20856 37412 20887
rect 38286 20884 38292 20896
rect 38344 20884 38350 20936
rect 41506 20924 41512 20936
rect 41467 20896 41512 20924
rect 41506 20884 41512 20896
rect 41564 20884 41570 20936
rect 41598 20884 41604 20936
rect 41656 20924 41662 20936
rect 41877 20927 41935 20933
rect 41656 20896 41701 20924
rect 41656 20884 41662 20896
rect 41877 20893 41889 20927
rect 41923 20893 41935 20927
rect 41877 20887 41935 20893
rect 39117 20859 39175 20865
rect 39117 20856 39129 20859
rect 37384 20828 39129 20856
rect 37185 20819 37243 20825
rect 39117 20825 39129 20828
rect 39163 20856 39175 20859
rect 40773 20859 40831 20865
rect 40773 20856 40785 20859
rect 39163 20828 40785 20856
rect 39163 20825 39175 20828
rect 39117 20819 39175 20825
rect 40773 20825 40785 20828
rect 40819 20856 40831 20859
rect 41782 20856 41788 20868
rect 40819 20828 41788 20856
rect 40819 20825 40831 20828
rect 40773 20819 40831 20825
rect 41782 20816 41788 20828
rect 41840 20856 41846 20868
rect 41892 20856 41920 20887
rect 41840 20828 41920 20856
rect 41840 20816 41846 20828
rect 35676 20760 35940 20788
rect 35676 20748 35682 20760
rect 35986 20748 35992 20800
rect 36044 20788 36050 20800
rect 36633 20791 36691 20797
rect 36633 20788 36645 20791
rect 36044 20760 36645 20788
rect 36044 20748 36050 20760
rect 36633 20757 36645 20760
rect 36679 20757 36691 20791
rect 41322 20788 41328 20800
rect 41283 20760 41328 20788
rect 36633 20751 36691 20757
rect 41322 20748 41328 20760
rect 41380 20748 41386 20800
rect 1104 20698 68816 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 50294 20698
rect 50346 20646 50358 20698
rect 50410 20646 50422 20698
rect 50474 20646 50486 20698
rect 50538 20646 50550 20698
rect 50602 20646 68816 20698
rect 1104 20624 68816 20646
rect 7469 20587 7527 20593
rect 7469 20553 7481 20587
rect 7515 20584 7527 20587
rect 7558 20584 7564 20596
rect 7515 20556 7564 20584
rect 7515 20553 7527 20556
rect 7469 20547 7527 20553
rect 7558 20544 7564 20556
rect 7616 20584 7622 20596
rect 8110 20584 8116 20596
rect 7616 20556 8116 20584
rect 7616 20544 7622 20556
rect 8110 20544 8116 20556
rect 8168 20544 8174 20596
rect 12161 20587 12219 20593
rect 12161 20553 12173 20587
rect 12207 20584 12219 20587
rect 12250 20584 12256 20596
rect 12207 20556 12256 20584
rect 12207 20553 12219 20556
rect 12161 20547 12219 20553
rect 12250 20544 12256 20556
rect 12308 20544 12314 20596
rect 12986 20584 12992 20596
rect 12360 20556 12992 20584
rect 5445 20519 5503 20525
rect 5445 20516 5457 20519
rect 4186 20488 5457 20516
rect 5445 20485 5457 20488
rect 5491 20485 5503 20519
rect 5445 20479 5503 20485
rect 7929 20519 7987 20525
rect 7929 20485 7941 20519
rect 7975 20516 7987 20519
rect 9398 20516 9404 20528
rect 7975 20488 9404 20516
rect 7975 20485 7987 20488
rect 7929 20479 7987 20485
rect 9398 20476 9404 20488
rect 9456 20476 9462 20528
rect 12360 20525 12388 20556
rect 12986 20544 12992 20556
rect 13044 20544 13050 20596
rect 15289 20587 15347 20593
rect 15289 20553 15301 20587
rect 15335 20584 15347 20587
rect 17773 20587 17831 20593
rect 15335 20556 16896 20584
rect 15335 20553 15347 20556
rect 15289 20547 15347 20553
rect 12345 20519 12403 20525
rect 12345 20485 12357 20519
rect 12391 20485 12403 20519
rect 12526 20516 12532 20528
rect 12439 20488 12532 20516
rect 12345 20479 12403 20485
rect 12526 20476 12532 20488
rect 12584 20516 12590 20528
rect 14093 20519 14151 20525
rect 14093 20516 14105 20519
rect 12584 20488 14105 20516
rect 12584 20476 12590 20488
rect 14093 20485 14105 20488
rect 14139 20516 14151 20519
rect 15194 20516 15200 20528
rect 14139 20488 15200 20516
rect 14139 20485 14151 20488
rect 14093 20479 14151 20485
rect 15194 20476 15200 20488
rect 15252 20476 15258 20528
rect 15378 20516 15384 20528
rect 15304 20488 15384 20516
rect 1394 20408 1400 20460
rect 1452 20448 1458 20460
rect 1949 20451 2007 20457
rect 1949 20448 1961 20451
rect 1452 20420 1961 20448
rect 1452 20408 1458 20420
rect 1949 20417 1961 20420
rect 1995 20417 2007 20451
rect 5534 20448 5540 20460
rect 5495 20420 5540 20448
rect 1949 20411 2007 20417
rect 5534 20408 5540 20420
rect 5592 20408 5598 20460
rect 6549 20451 6607 20457
rect 6549 20417 6561 20451
rect 6595 20448 6607 20451
rect 8202 20448 8208 20460
rect 6595 20420 8208 20448
rect 6595 20417 6607 20420
rect 6549 20411 6607 20417
rect 8202 20408 8208 20420
rect 8260 20408 8266 20460
rect 10134 20448 10140 20460
rect 10095 20420 10140 20448
rect 10134 20408 10140 20420
rect 10192 20408 10198 20460
rect 14277 20451 14335 20457
rect 14277 20417 14289 20451
rect 14323 20448 14335 20451
rect 15304 20448 15332 20488
rect 15378 20476 15384 20488
rect 15436 20476 15442 20528
rect 16666 20516 16672 20528
rect 16627 20488 16672 20516
rect 16666 20476 16672 20488
rect 16724 20476 16730 20528
rect 16868 20516 16896 20556
rect 17773 20553 17785 20587
rect 17819 20584 17831 20587
rect 17954 20584 17960 20596
rect 17819 20556 17960 20584
rect 17819 20553 17831 20556
rect 17773 20547 17831 20553
rect 17954 20544 17960 20556
rect 18012 20544 18018 20596
rect 19058 20544 19064 20596
rect 19116 20584 19122 20596
rect 21818 20584 21824 20596
rect 19116 20556 21824 20584
rect 19116 20544 19122 20556
rect 21818 20544 21824 20556
rect 21876 20544 21882 20596
rect 22005 20587 22063 20593
rect 22005 20553 22017 20587
rect 22051 20584 22063 20587
rect 22278 20584 22284 20596
rect 22051 20556 22284 20584
rect 22051 20553 22063 20556
rect 22005 20547 22063 20553
rect 22278 20544 22284 20556
rect 22336 20544 22342 20596
rect 23566 20584 23572 20596
rect 23170 20556 23572 20584
rect 18598 20516 18604 20528
rect 16868 20488 18604 20516
rect 18598 20476 18604 20488
rect 18656 20476 18662 20528
rect 19334 20476 19340 20528
rect 19392 20516 19398 20528
rect 20346 20516 20352 20528
rect 19392 20488 20352 20516
rect 19392 20476 19398 20488
rect 20346 20476 20352 20488
rect 20404 20476 20410 20528
rect 21634 20476 21640 20528
rect 21692 20516 21698 20528
rect 22189 20519 22247 20525
rect 22189 20516 22201 20519
rect 21692 20488 22201 20516
rect 21692 20476 21698 20488
rect 22189 20485 22201 20488
rect 22235 20485 22247 20519
rect 22189 20479 22247 20485
rect 15470 20448 15476 20460
rect 14323 20420 15332 20448
rect 15431 20420 15476 20448
rect 14323 20417 14335 20420
rect 14277 20411 14335 20417
rect 15470 20408 15476 20420
rect 15528 20408 15534 20460
rect 15746 20448 15752 20460
rect 15707 20420 15752 20448
rect 15746 20408 15752 20420
rect 15804 20408 15810 20460
rect 16853 20451 16911 20457
rect 16853 20417 16865 20451
rect 16899 20448 16911 20451
rect 17126 20448 17132 20460
rect 16899 20420 17132 20448
rect 16899 20417 16911 20420
rect 16853 20411 16911 20417
rect 17126 20408 17132 20420
rect 17184 20408 17190 20460
rect 17218 20408 17224 20460
rect 17276 20448 17282 20460
rect 17494 20448 17500 20460
rect 17276 20420 17500 20448
rect 17276 20408 17282 20420
rect 17494 20408 17500 20420
rect 17552 20448 17558 20460
rect 17681 20451 17739 20457
rect 17681 20448 17693 20451
rect 17552 20420 17693 20448
rect 17552 20408 17558 20420
rect 17681 20417 17693 20420
rect 17727 20417 17739 20451
rect 17681 20411 17739 20417
rect 19426 20408 19432 20460
rect 19484 20448 19490 20460
rect 20165 20451 20223 20457
rect 20165 20448 20177 20451
rect 19484 20420 20177 20448
rect 19484 20408 19490 20420
rect 20165 20417 20177 20420
rect 20211 20417 20223 20451
rect 20165 20411 20223 20417
rect 20254 20408 20260 20460
rect 20312 20448 20318 20460
rect 20530 20448 20536 20460
rect 20312 20420 20357 20448
rect 20491 20420 20536 20448
rect 20312 20408 20318 20420
rect 20530 20408 20536 20420
rect 20588 20408 20594 20460
rect 21821 20451 21879 20457
rect 21821 20417 21833 20451
rect 21867 20417 21879 20451
rect 21821 20411 21879 20417
rect 1486 20340 1492 20392
rect 1544 20380 1550 20392
rect 1673 20383 1731 20389
rect 1673 20380 1685 20383
rect 1544 20352 1685 20380
rect 1544 20340 1550 20352
rect 1673 20349 1685 20352
rect 1719 20349 1731 20383
rect 4617 20383 4675 20389
rect 4617 20380 4629 20383
rect 1673 20343 1731 20349
rect 2700 20352 4629 20380
rect 2700 20321 2728 20352
rect 4617 20349 4629 20352
rect 4663 20349 4675 20383
rect 4890 20380 4896 20392
rect 4851 20352 4896 20380
rect 4617 20343 4675 20349
rect 4890 20340 4896 20352
rect 4948 20380 4954 20392
rect 5442 20380 5448 20392
rect 4948 20352 5448 20380
rect 4948 20340 4954 20352
rect 5442 20340 5448 20352
rect 5500 20340 5506 20392
rect 6914 20340 6920 20392
rect 6972 20380 6978 20392
rect 7926 20380 7932 20392
rect 6972 20352 7932 20380
rect 6972 20340 6978 20352
rect 7926 20340 7932 20352
rect 7984 20340 7990 20392
rect 8662 20380 8668 20392
rect 8623 20352 8668 20380
rect 8662 20340 8668 20352
rect 8720 20340 8726 20392
rect 9861 20383 9919 20389
rect 9861 20380 9873 20383
rect 9646 20352 9873 20380
rect 2685 20315 2743 20321
rect 2685 20281 2697 20315
rect 2731 20281 2743 20315
rect 2685 20275 2743 20281
rect 8478 20272 8484 20324
rect 8536 20312 8542 20324
rect 9646 20312 9674 20352
rect 9861 20349 9873 20352
rect 9907 20349 9919 20383
rect 9861 20343 9919 20349
rect 12986 20340 12992 20392
rect 13044 20380 13050 20392
rect 15654 20380 15660 20392
rect 13044 20352 15660 20380
rect 13044 20340 13050 20352
rect 15654 20340 15660 20352
rect 15712 20340 15718 20392
rect 16298 20340 16304 20392
rect 16356 20380 16362 20392
rect 18325 20383 18383 20389
rect 18325 20380 18337 20383
rect 16356 20352 18337 20380
rect 16356 20340 16362 20352
rect 18325 20349 18337 20352
rect 18371 20349 18383 20383
rect 21836 20380 21864 20411
rect 21910 20408 21916 20460
rect 21968 20448 21974 20460
rect 21968 20420 22013 20448
rect 21968 20408 21974 20420
rect 22094 20408 22100 20460
rect 22152 20448 22158 20460
rect 22281 20451 22339 20457
rect 22152 20420 22197 20448
rect 22152 20408 22158 20420
rect 22281 20417 22293 20451
rect 22327 20448 22339 20451
rect 22370 20448 22376 20460
rect 22327 20420 22376 20448
rect 22327 20417 22339 20420
rect 22281 20411 22339 20417
rect 22370 20408 22376 20420
rect 22428 20408 22434 20460
rect 22922 20408 22928 20460
rect 22980 20448 22986 20460
rect 23170 20457 23198 20556
rect 23566 20544 23572 20556
rect 23624 20544 23630 20596
rect 24581 20587 24639 20593
rect 24581 20553 24593 20587
rect 24627 20584 24639 20587
rect 25406 20584 25412 20596
rect 24627 20556 25412 20584
rect 24627 20553 24639 20556
rect 24581 20547 24639 20553
rect 25406 20544 25412 20556
rect 25464 20544 25470 20596
rect 26234 20544 26240 20596
rect 26292 20584 26298 20596
rect 32950 20584 32956 20596
rect 26292 20556 32812 20584
rect 32911 20556 32956 20584
rect 26292 20544 26298 20556
rect 26970 20476 26976 20528
rect 27028 20516 27034 20528
rect 27249 20519 27307 20525
rect 27249 20516 27261 20519
rect 27028 20488 27261 20516
rect 27028 20476 27034 20488
rect 27249 20485 27261 20488
rect 27295 20485 27307 20519
rect 29546 20516 29552 20528
rect 27249 20479 27307 20485
rect 27448 20488 29552 20516
rect 27448 20460 27476 20488
rect 29546 20476 29552 20488
rect 29604 20476 29610 20528
rect 32398 20476 32404 20528
rect 32456 20516 32462 20528
rect 32784 20516 32812 20556
rect 32950 20544 32956 20556
rect 33008 20544 33014 20596
rect 35710 20544 35716 20596
rect 35768 20584 35774 20596
rect 36449 20587 36507 20593
rect 36449 20584 36461 20587
rect 35768 20556 36461 20584
rect 35768 20544 35774 20556
rect 36449 20553 36461 20556
rect 36495 20553 36507 20587
rect 36449 20547 36507 20553
rect 38013 20587 38071 20593
rect 38013 20553 38025 20587
rect 38059 20584 38071 20587
rect 38286 20584 38292 20596
rect 38059 20556 38292 20584
rect 38059 20553 38071 20556
rect 38013 20547 38071 20553
rect 38286 20544 38292 20556
rect 38344 20544 38350 20596
rect 41233 20587 41291 20593
rect 41233 20553 41245 20587
rect 41279 20584 41291 20587
rect 41322 20584 41328 20596
rect 41279 20556 41328 20584
rect 41279 20553 41291 20556
rect 41233 20547 41291 20553
rect 41322 20544 41328 20556
rect 41380 20544 41386 20596
rect 42794 20544 42800 20596
rect 42852 20584 42858 20596
rect 42889 20587 42947 20593
rect 42889 20584 42901 20587
rect 42852 20556 42901 20584
rect 42852 20544 42858 20556
rect 42889 20553 42901 20556
rect 42935 20553 42947 20587
rect 42889 20547 42947 20553
rect 34330 20516 34336 20528
rect 32456 20488 32615 20516
rect 32784 20488 34336 20516
rect 32456 20476 32462 20488
rect 23157 20451 23215 20457
rect 23157 20448 23169 20451
rect 22980 20420 23169 20448
rect 22980 20408 22986 20420
rect 23157 20417 23169 20420
rect 23203 20417 23215 20451
rect 23157 20411 23215 20417
rect 23293 20451 23351 20457
rect 23293 20417 23305 20451
rect 23339 20417 23351 20451
rect 23293 20411 23351 20417
rect 23308 20380 23336 20411
rect 23382 20408 23388 20460
rect 23440 20448 23446 20460
rect 23568 20451 23626 20457
rect 23440 20420 23485 20448
rect 23440 20408 23446 20420
rect 23568 20417 23580 20451
rect 23614 20417 23626 20451
rect 23568 20411 23626 20417
rect 18325 20343 18383 20349
rect 19996 20352 21864 20380
rect 21928 20352 23336 20380
rect 23584 20380 23612 20411
rect 23658 20408 23664 20460
rect 23716 20448 23722 20460
rect 24394 20448 24400 20460
rect 23716 20420 23761 20448
rect 24307 20420 24400 20448
rect 23716 20408 23722 20420
rect 24394 20408 24400 20420
rect 24452 20448 24458 20460
rect 26602 20448 26608 20460
rect 24452 20420 26608 20448
rect 24452 20408 24458 20420
rect 26602 20408 26608 20420
rect 26660 20408 26666 20460
rect 27430 20448 27436 20460
rect 27391 20420 27436 20448
rect 27430 20408 27436 20420
rect 27488 20408 27494 20460
rect 28258 20448 28264 20460
rect 28219 20420 28264 20448
rect 28258 20408 28264 20420
rect 28316 20408 28322 20460
rect 31481 20451 31539 20457
rect 31481 20448 31493 20451
rect 28368 20420 31493 20448
rect 25130 20380 25136 20392
rect 23584 20352 25136 20380
rect 19996 20321 20024 20352
rect 8536 20284 9674 20312
rect 19981 20315 20039 20321
rect 8536 20272 8542 20284
rect 19981 20281 19993 20315
rect 20027 20281 20039 20315
rect 21928 20312 21956 20352
rect 25130 20340 25136 20352
rect 25188 20340 25194 20392
rect 25314 20380 25320 20392
rect 25275 20352 25320 20380
rect 25314 20340 25320 20352
rect 25372 20340 25378 20392
rect 28074 20340 28080 20392
rect 28132 20380 28138 20392
rect 28368 20380 28396 20420
rect 31481 20417 31493 20420
rect 31527 20417 31539 20451
rect 31481 20411 31539 20417
rect 28132 20352 28396 20380
rect 28132 20340 28138 20352
rect 28442 20340 28448 20392
rect 28500 20380 28506 20392
rect 28997 20383 29055 20389
rect 28997 20380 29009 20383
rect 28500 20352 29009 20380
rect 28500 20340 28506 20352
rect 28997 20349 29009 20352
rect 29043 20349 29055 20383
rect 31496 20380 31524 20411
rect 32030 20408 32036 20460
rect 32088 20448 32094 20460
rect 32490 20457 32496 20460
rect 32309 20451 32367 20457
rect 32309 20448 32321 20451
rect 32088 20420 32321 20448
rect 32088 20408 32094 20420
rect 32309 20417 32321 20420
rect 32355 20417 32367 20451
rect 32488 20448 32496 20457
rect 32451 20420 32496 20448
rect 32309 20411 32367 20417
rect 32488 20411 32496 20420
rect 32490 20408 32496 20411
rect 32548 20408 32554 20460
rect 32587 20457 32615 20488
rect 34330 20476 34336 20488
rect 34388 20476 34394 20528
rect 35894 20516 35900 20528
rect 35084 20488 35900 20516
rect 32585 20451 32643 20457
rect 32585 20417 32597 20451
rect 32631 20417 32643 20451
rect 32585 20411 32643 20417
rect 32697 20451 32755 20457
rect 32697 20417 32709 20451
rect 32743 20448 32755 20451
rect 33505 20451 33563 20457
rect 32743 20420 32812 20448
rect 32743 20417 32755 20420
rect 32697 20411 32755 20417
rect 31496 20352 32536 20380
rect 28997 20343 29055 20349
rect 19981 20275 20039 20281
rect 21192 20284 21956 20312
rect 3142 20244 3148 20256
rect 3103 20216 3148 20244
rect 3142 20204 3148 20216
rect 3200 20204 3206 20256
rect 6362 20244 6368 20256
rect 6323 20216 6368 20244
rect 6362 20204 6368 20216
rect 6420 20204 6426 20256
rect 14461 20247 14519 20253
rect 14461 20213 14473 20247
rect 14507 20244 14519 20247
rect 14550 20244 14556 20256
rect 14507 20216 14556 20244
rect 14507 20213 14519 20216
rect 14461 20207 14519 20213
rect 14550 20204 14556 20216
rect 14608 20204 14614 20256
rect 15378 20204 15384 20256
rect 15436 20244 15442 20256
rect 15473 20247 15531 20253
rect 15473 20244 15485 20247
rect 15436 20216 15485 20244
rect 15436 20204 15442 20216
rect 15473 20213 15485 20216
rect 15519 20213 15531 20247
rect 15473 20207 15531 20213
rect 18046 20204 18052 20256
rect 18104 20244 18110 20256
rect 21192 20253 21220 20284
rect 22094 20272 22100 20324
rect 22152 20312 22158 20324
rect 29730 20312 29736 20324
rect 22152 20284 29736 20312
rect 22152 20272 22158 20284
rect 29730 20272 29736 20284
rect 29788 20272 29794 20324
rect 32508 20312 32536 20352
rect 32784 20312 32812 20420
rect 33505 20417 33517 20451
rect 33551 20448 33563 20451
rect 33686 20448 33692 20460
rect 33551 20420 33692 20448
rect 33551 20417 33563 20420
rect 33505 20411 33563 20417
rect 33686 20408 33692 20420
rect 33744 20408 33750 20460
rect 35084 20457 35112 20488
rect 35894 20476 35900 20488
rect 35952 20476 35958 20528
rect 37553 20519 37611 20525
rect 37553 20485 37565 20519
rect 37599 20516 37611 20519
rect 38102 20516 38108 20528
rect 37599 20488 38108 20516
rect 37599 20485 37611 20488
rect 37553 20479 37611 20485
rect 38102 20476 38108 20488
rect 38160 20476 38166 20528
rect 41414 20476 41420 20528
rect 41472 20516 41478 20528
rect 41472 20488 42748 20516
rect 41472 20476 41478 20488
rect 34517 20451 34575 20457
rect 34517 20448 34529 20451
rect 34164 20420 34529 20448
rect 33778 20380 33784 20392
rect 33691 20352 33784 20380
rect 33704 20321 33732 20352
rect 33778 20340 33784 20352
rect 33836 20380 33842 20392
rect 34164 20380 34192 20420
rect 34517 20417 34529 20420
rect 34563 20417 34575 20451
rect 34517 20411 34575 20417
rect 35069 20451 35127 20457
rect 35069 20417 35081 20451
rect 35115 20417 35127 20451
rect 35325 20451 35383 20457
rect 35325 20448 35337 20451
rect 35069 20411 35127 20417
rect 35176 20420 35337 20448
rect 33836 20352 34192 20380
rect 33836 20340 33842 20352
rect 34238 20340 34244 20392
rect 34296 20380 34302 20392
rect 35176 20380 35204 20420
rect 35325 20417 35337 20420
rect 35371 20417 35383 20451
rect 37829 20451 37887 20457
rect 37829 20448 37841 20451
rect 35325 20411 35383 20417
rect 37752 20420 37841 20448
rect 37642 20380 37648 20392
rect 34296 20352 35204 20380
rect 37603 20352 37648 20380
rect 34296 20340 34302 20352
rect 37642 20340 37648 20352
rect 37700 20340 37706 20392
rect 30944 20284 31616 20312
rect 32508 20284 32812 20312
rect 33689 20315 33747 20321
rect 21177 20247 21235 20253
rect 21177 20244 21189 20247
rect 18104 20216 21189 20244
rect 18104 20204 18110 20216
rect 21177 20213 21189 20216
rect 21223 20213 21235 20247
rect 21177 20207 21235 20213
rect 21818 20204 21824 20256
rect 21876 20244 21882 20256
rect 22922 20244 22928 20256
rect 21876 20216 22928 20244
rect 21876 20204 21882 20216
rect 22922 20204 22928 20216
rect 22980 20204 22986 20256
rect 23017 20247 23075 20253
rect 23017 20213 23029 20247
rect 23063 20244 23075 20247
rect 23290 20244 23296 20256
rect 23063 20216 23296 20244
rect 23063 20213 23075 20216
rect 23017 20207 23075 20213
rect 23290 20204 23296 20216
rect 23348 20204 23354 20256
rect 25222 20204 25228 20256
rect 25280 20244 25286 20256
rect 25547 20247 25605 20253
rect 25547 20244 25559 20247
rect 25280 20216 25559 20244
rect 25280 20204 25286 20216
rect 25547 20213 25559 20216
rect 25593 20244 25605 20247
rect 25866 20244 25872 20256
rect 25593 20216 25872 20244
rect 25593 20213 25605 20216
rect 25547 20207 25605 20213
rect 25866 20204 25872 20216
rect 25924 20204 25930 20256
rect 27617 20247 27675 20253
rect 27617 20213 27629 20247
rect 27663 20244 27675 20247
rect 27890 20244 27896 20256
rect 27663 20216 27896 20244
rect 27663 20213 27675 20216
rect 27617 20207 27675 20213
rect 27890 20204 27896 20216
rect 27948 20204 27954 20256
rect 30190 20204 30196 20256
rect 30248 20244 30254 20256
rect 30944 20253 30972 20284
rect 30929 20247 30987 20253
rect 30929 20244 30941 20247
rect 30248 20216 30941 20244
rect 30248 20204 30254 20216
rect 30929 20213 30941 20216
rect 30975 20213 30987 20247
rect 31588 20244 31616 20284
rect 33689 20281 33701 20315
rect 33735 20281 33747 20315
rect 33689 20275 33747 20281
rect 37366 20272 37372 20324
rect 37424 20312 37430 20324
rect 37752 20312 37780 20420
rect 37829 20417 37841 20420
rect 37875 20417 37887 20451
rect 37829 20411 37887 20417
rect 37918 20408 37924 20460
rect 37976 20448 37982 20460
rect 39097 20451 39155 20457
rect 39097 20448 39109 20451
rect 37976 20420 39109 20448
rect 37976 20408 37982 20420
rect 39097 20417 39109 20420
rect 39143 20417 39155 20451
rect 39097 20411 39155 20417
rect 41601 20451 41659 20457
rect 41601 20417 41613 20451
rect 41647 20448 41659 20451
rect 41782 20448 41788 20460
rect 41647 20420 41788 20448
rect 41647 20417 41659 20420
rect 41601 20411 41659 20417
rect 41782 20408 41788 20420
rect 41840 20408 41846 20460
rect 42426 20448 42432 20460
rect 42387 20420 42432 20448
rect 42426 20408 42432 20420
rect 42484 20408 42490 20460
rect 42720 20457 42748 20488
rect 42705 20451 42763 20457
rect 42705 20417 42717 20451
rect 42751 20417 42763 20451
rect 42705 20411 42763 20417
rect 38838 20380 38844 20392
rect 38799 20352 38844 20380
rect 38838 20340 38844 20352
rect 38896 20340 38902 20392
rect 40218 20340 40224 20392
rect 40276 20380 40282 20392
rect 40681 20383 40739 20389
rect 40681 20380 40693 20383
rect 40276 20352 40693 20380
rect 40276 20340 40282 20352
rect 40681 20349 40693 20352
rect 40727 20349 40739 20383
rect 40681 20343 40739 20349
rect 41690 20340 41696 20392
rect 41748 20380 41754 20392
rect 41877 20383 41935 20389
rect 41748 20352 41793 20380
rect 41748 20340 41754 20352
rect 41877 20349 41889 20383
rect 41923 20380 41935 20383
rect 42521 20383 42579 20389
rect 42521 20380 42533 20383
rect 41923 20352 42533 20380
rect 41923 20349 41935 20352
rect 41877 20343 41935 20349
rect 42521 20349 42533 20352
rect 42567 20349 42579 20383
rect 42521 20343 42579 20349
rect 37424 20284 37780 20312
rect 37424 20272 37430 20284
rect 32214 20244 32220 20256
rect 31588 20216 32220 20244
rect 30929 20207 30987 20213
rect 32214 20204 32220 20216
rect 32272 20204 32278 20256
rect 34146 20244 34152 20256
rect 34107 20216 34152 20244
rect 34146 20204 34152 20216
rect 34204 20204 34210 20256
rect 37734 20244 37740 20256
rect 37695 20216 37740 20244
rect 37734 20204 37740 20216
rect 37792 20204 37798 20256
rect 39482 20204 39488 20256
rect 39540 20244 39546 20256
rect 40221 20247 40279 20253
rect 40221 20244 40233 20247
rect 39540 20216 40233 20244
rect 39540 20204 39546 20216
rect 40221 20213 40233 20216
rect 40267 20213 40279 20247
rect 40221 20207 40279 20213
rect 41782 20204 41788 20256
rect 41840 20244 41846 20256
rect 42429 20247 42487 20253
rect 42429 20244 42441 20247
rect 41840 20216 42441 20244
rect 41840 20204 41846 20216
rect 42429 20213 42441 20216
rect 42475 20213 42487 20247
rect 67634 20244 67640 20256
rect 67595 20216 67640 20244
rect 42429 20207 42487 20213
rect 67634 20204 67640 20216
rect 67692 20204 67698 20256
rect 1104 20154 68816 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 65654 20154
rect 65706 20102 65718 20154
rect 65770 20102 65782 20154
rect 65834 20102 65846 20154
rect 65898 20102 65910 20154
rect 65962 20102 68816 20154
rect 1104 20080 68816 20102
rect 7282 20000 7288 20052
rect 7340 20040 7346 20052
rect 8110 20040 8116 20052
rect 7340 20012 7420 20040
rect 8071 20012 8116 20040
rect 7340 20000 7346 20012
rect 7392 19904 7420 20012
rect 8110 20000 8116 20012
rect 8168 20000 8174 20052
rect 8389 20043 8447 20049
rect 8389 20009 8401 20043
rect 8435 20040 8447 20043
rect 9214 20040 9220 20052
rect 8435 20012 9220 20040
rect 8435 20009 8447 20012
rect 8389 20003 8447 20009
rect 9214 20000 9220 20012
rect 9272 20000 9278 20052
rect 11054 20000 11060 20052
rect 11112 20040 11118 20052
rect 18046 20040 18052 20052
rect 11112 20012 18052 20040
rect 11112 20000 11118 20012
rect 18046 20000 18052 20012
rect 18104 20000 18110 20052
rect 22186 20040 22192 20052
rect 18156 20012 22192 20040
rect 7834 19932 7840 19984
rect 7892 19972 7898 19984
rect 7892 19944 9260 19972
rect 7892 19932 7898 19944
rect 8018 19904 8024 19916
rect 7300 19876 7420 19904
rect 7979 19876 8024 19904
rect 2222 19796 2228 19848
rect 2280 19836 2286 19848
rect 2317 19839 2375 19845
rect 2317 19836 2329 19839
rect 2280 19808 2329 19836
rect 2280 19796 2286 19808
rect 2317 19805 2329 19808
rect 2363 19805 2375 19839
rect 2317 19799 2375 19805
rect 4614 19796 4620 19848
rect 4672 19836 4678 19848
rect 4890 19836 4896 19848
rect 4672 19808 4896 19836
rect 4672 19796 4678 19808
rect 4890 19796 4896 19808
rect 4948 19836 4954 19848
rect 4985 19839 5043 19845
rect 4985 19836 4997 19839
rect 4948 19808 4997 19836
rect 4948 19796 4954 19808
rect 4985 19805 4997 19808
rect 5031 19805 5043 19839
rect 7098 19836 7104 19848
rect 7059 19808 7104 19836
rect 4985 19799 5043 19805
rect 7098 19796 7104 19808
rect 7156 19796 7162 19848
rect 7300 19845 7328 19876
rect 8018 19864 8024 19876
rect 8076 19864 8082 19916
rect 8478 19904 8484 19916
rect 8128 19876 8484 19904
rect 7193 19839 7251 19845
rect 7193 19805 7205 19839
rect 7239 19805 7251 19839
rect 7193 19799 7251 19805
rect 7285 19839 7343 19845
rect 7285 19805 7297 19839
rect 7331 19805 7343 19839
rect 7466 19836 7472 19848
rect 7427 19808 7472 19836
rect 7285 19799 7343 19805
rect 5252 19771 5310 19777
rect 5252 19737 5264 19771
rect 5298 19768 5310 19771
rect 6825 19771 6883 19777
rect 6825 19768 6837 19771
rect 5298 19740 6837 19768
rect 5298 19737 5310 19740
rect 5252 19731 5310 19737
rect 6825 19737 6837 19740
rect 6871 19737 6883 19771
rect 6825 19731 6883 19737
rect 1486 19660 1492 19712
rect 1544 19700 1550 19712
rect 2133 19703 2191 19709
rect 2133 19700 2145 19703
rect 1544 19672 2145 19700
rect 1544 19660 1550 19672
rect 2133 19669 2145 19672
rect 2179 19669 2191 19703
rect 2133 19663 2191 19669
rect 6365 19703 6423 19709
rect 6365 19669 6377 19703
rect 6411 19700 6423 19703
rect 6914 19700 6920 19712
rect 6411 19672 6920 19700
rect 6411 19669 6423 19672
rect 6365 19663 6423 19669
rect 6914 19660 6920 19672
rect 6972 19660 6978 19712
rect 7208 19700 7236 19799
rect 7466 19796 7472 19808
rect 7524 19836 7530 19848
rect 8128 19836 8156 19876
rect 8478 19864 8484 19876
rect 8536 19904 8542 19916
rect 8536 19876 8984 19904
rect 8536 19864 8542 19876
rect 8956 19845 8984 19876
rect 9232 19845 9260 19944
rect 9766 19904 9772 19916
rect 9324 19876 9772 19904
rect 9324 19845 9352 19876
rect 9766 19864 9772 19876
rect 9824 19864 9830 19916
rect 13262 19864 13268 19916
rect 13320 19904 13326 19916
rect 16666 19904 16672 19916
rect 13320 19876 16160 19904
rect 13320 19864 13326 19876
rect 7524 19808 8156 19836
rect 8205 19839 8263 19845
rect 7524 19796 7530 19808
rect 8205 19805 8217 19839
rect 8251 19805 8263 19839
rect 8205 19799 8263 19805
rect 8941 19839 8999 19845
rect 8941 19805 8953 19839
rect 8987 19805 8999 19839
rect 9101 19833 9107 19845
rect 9062 19805 9107 19833
rect 8941 19799 8999 19805
rect 7926 19768 7932 19780
rect 7887 19740 7932 19768
rect 7926 19728 7932 19740
rect 7984 19728 7990 19780
rect 7834 19700 7840 19712
rect 7208 19672 7840 19700
rect 7834 19660 7840 19672
rect 7892 19660 7898 19712
rect 8220 19700 8248 19799
rect 9101 19793 9107 19805
rect 9159 19793 9165 19845
rect 9217 19839 9275 19845
rect 9217 19805 9229 19839
rect 9263 19805 9275 19839
rect 9217 19799 9275 19805
rect 9309 19839 9367 19845
rect 9309 19805 9321 19839
rect 9355 19805 9367 19839
rect 9309 19799 9367 19805
rect 9398 19796 9404 19848
rect 9456 19836 9462 19848
rect 11425 19839 11483 19845
rect 9456 19808 11284 19836
rect 9456 19796 9462 19808
rect 9585 19771 9643 19777
rect 9585 19737 9597 19771
rect 9631 19768 9643 19771
rect 11158 19771 11216 19777
rect 11158 19768 11170 19771
rect 9631 19740 11170 19768
rect 9631 19737 9643 19740
rect 9585 19731 9643 19737
rect 11158 19737 11170 19740
rect 11204 19737 11216 19771
rect 11256 19768 11284 19808
rect 11425 19805 11437 19839
rect 11471 19836 11483 19839
rect 11606 19836 11612 19848
rect 11471 19808 11612 19836
rect 11471 19805 11483 19808
rect 11425 19799 11483 19805
rect 11606 19796 11612 19808
rect 11664 19836 11670 19848
rect 12158 19836 12164 19848
rect 11664 19808 12164 19836
rect 11664 19796 11670 19808
rect 12158 19796 12164 19808
rect 12216 19796 12222 19848
rect 15654 19796 15660 19848
rect 15712 19836 15718 19848
rect 16132 19845 16160 19876
rect 16224 19876 16672 19904
rect 16224 19845 16252 19876
rect 16666 19864 16672 19876
rect 16724 19904 16730 19916
rect 16724 19876 17540 19904
rect 16724 19864 16730 19876
rect 15841 19839 15899 19845
rect 15841 19836 15853 19839
rect 15712 19808 15853 19836
rect 15712 19796 15718 19808
rect 15841 19805 15853 19808
rect 15887 19805 15899 19839
rect 15841 19799 15899 19805
rect 16117 19839 16175 19845
rect 16117 19805 16129 19839
rect 16163 19805 16175 19839
rect 16117 19799 16175 19805
rect 16209 19839 16267 19845
rect 16209 19805 16221 19839
rect 16255 19805 16267 19839
rect 16209 19799 16267 19805
rect 17034 19796 17040 19848
rect 17092 19836 17098 19848
rect 17512 19845 17540 19876
rect 18156 19845 18184 20012
rect 22186 20000 22192 20012
rect 22244 20000 22250 20052
rect 22557 20043 22615 20049
rect 22557 20009 22569 20043
rect 22603 20040 22615 20043
rect 24394 20040 24400 20052
rect 22603 20012 24400 20040
rect 22603 20009 22615 20012
rect 22557 20003 22615 20009
rect 24394 20000 24400 20012
rect 24452 20000 24458 20052
rect 24670 20040 24676 20052
rect 24631 20012 24676 20040
rect 24670 20000 24676 20012
rect 24728 20000 24734 20052
rect 26142 20040 26148 20052
rect 26103 20012 26148 20040
rect 26142 20000 26148 20012
rect 26200 20000 26206 20052
rect 26789 20043 26847 20049
rect 26789 20009 26801 20043
rect 26835 20040 26847 20043
rect 26970 20040 26976 20052
rect 26835 20012 26976 20040
rect 26835 20009 26847 20012
rect 26789 20003 26847 20009
rect 26970 20000 26976 20012
rect 27028 20000 27034 20052
rect 30193 20043 30251 20049
rect 30193 20009 30205 20043
rect 30239 20040 30251 20043
rect 30558 20040 30564 20052
rect 30239 20012 30564 20040
rect 30239 20009 30251 20012
rect 30193 20003 30251 20009
rect 30558 20000 30564 20012
rect 30616 20000 30622 20052
rect 32122 20040 32128 20052
rect 32083 20012 32128 20040
rect 32122 20000 32128 20012
rect 32180 20000 32186 20052
rect 34149 20043 34207 20049
rect 34149 20009 34161 20043
rect 34195 20040 34207 20043
rect 34238 20040 34244 20052
rect 34195 20012 34244 20040
rect 34195 20009 34207 20012
rect 34149 20003 34207 20009
rect 34238 20000 34244 20012
rect 34296 20000 34302 20052
rect 37918 20040 37924 20052
rect 37879 20012 37924 20040
rect 37918 20000 37924 20012
rect 37976 20000 37982 20052
rect 40129 20043 40187 20049
rect 40129 20009 40141 20043
rect 40175 20040 40187 20043
rect 40218 20040 40224 20052
rect 40175 20012 40224 20040
rect 40175 20009 40187 20012
rect 40129 20003 40187 20009
rect 19334 19972 19340 19984
rect 18248 19944 19340 19972
rect 17129 19839 17187 19845
rect 17129 19836 17141 19839
rect 17092 19808 17141 19836
rect 17092 19796 17098 19808
rect 17129 19805 17141 19808
rect 17175 19805 17187 19839
rect 17405 19839 17463 19845
rect 17405 19836 17417 19839
rect 17129 19799 17187 19805
rect 17236 19808 17417 19836
rect 13541 19771 13599 19777
rect 13541 19768 13553 19771
rect 11256 19740 13553 19768
rect 11158 19731 11216 19737
rect 13541 19737 13553 19740
rect 13587 19768 13599 19771
rect 14458 19768 14464 19780
rect 13587 19740 14464 19768
rect 13587 19737 13599 19740
rect 13541 19731 13599 19737
rect 14458 19728 14464 19740
rect 14516 19768 14522 19780
rect 15102 19768 15108 19780
rect 14516 19740 15108 19768
rect 14516 19728 14522 19740
rect 15102 19728 15108 19740
rect 15160 19728 15166 19780
rect 15286 19728 15292 19780
rect 15344 19768 15350 19780
rect 15562 19768 15568 19780
rect 15344 19740 15568 19768
rect 15344 19728 15350 19740
rect 15562 19728 15568 19740
rect 15620 19728 15626 19780
rect 15746 19728 15752 19780
rect 15804 19768 15810 19780
rect 16025 19771 16083 19777
rect 16025 19768 16037 19771
rect 15804 19740 16037 19768
rect 15804 19728 15810 19740
rect 16025 19737 16037 19740
rect 16071 19737 16083 19771
rect 16025 19731 16083 19737
rect 16298 19728 16304 19780
rect 16356 19768 16362 19780
rect 17236 19768 17264 19808
rect 17405 19805 17417 19808
rect 17451 19805 17463 19839
rect 17405 19799 17463 19805
rect 17497 19839 17555 19845
rect 17497 19805 17509 19839
rect 17543 19836 17555 19839
rect 18141 19839 18199 19845
rect 17543 19808 17816 19836
rect 17543 19805 17555 19808
rect 17497 19799 17555 19805
rect 16356 19740 17264 19768
rect 17313 19771 17371 19777
rect 16356 19728 16362 19740
rect 17313 19737 17325 19771
rect 17359 19737 17371 19771
rect 17313 19731 17371 19737
rect 10045 19703 10103 19709
rect 10045 19700 10057 19703
rect 8220 19672 10057 19700
rect 10045 19669 10057 19672
rect 10091 19700 10103 19703
rect 10134 19700 10140 19712
rect 10091 19672 10140 19700
rect 10091 19669 10103 19672
rect 10045 19663 10103 19669
rect 10134 19660 10140 19672
rect 10192 19660 10198 19712
rect 14366 19660 14372 19712
rect 14424 19700 14430 19712
rect 15304 19700 15332 19728
rect 14424 19672 15332 19700
rect 16393 19703 16451 19709
rect 14424 19660 14430 19672
rect 16393 19669 16405 19703
rect 16439 19700 16451 19703
rect 16482 19700 16488 19712
rect 16439 19672 16488 19700
rect 16439 19669 16451 19672
rect 16393 19663 16451 19669
rect 16482 19660 16488 19672
rect 16540 19660 16546 19712
rect 17328 19700 17356 19731
rect 17494 19700 17500 19712
rect 17328 19672 17500 19700
rect 17494 19660 17500 19672
rect 17552 19660 17558 19712
rect 17678 19700 17684 19712
rect 17639 19672 17684 19700
rect 17678 19660 17684 19672
rect 17736 19660 17742 19712
rect 17788 19700 17816 19808
rect 18141 19805 18153 19839
rect 18187 19805 18199 19839
rect 18248 19836 18276 19944
rect 19334 19932 19340 19944
rect 19392 19932 19398 19984
rect 20622 19932 20628 19984
rect 20680 19972 20686 19984
rect 27430 19972 27436 19984
rect 20680 19944 27436 19972
rect 20680 19932 20686 19944
rect 27430 19932 27436 19944
rect 27488 19932 27494 19984
rect 27706 19932 27712 19984
rect 27764 19972 27770 19984
rect 28350 19972 28356 19984
rect 27764 19944 28356 19972
rect 27764 19932 27770 19944
rect 28350 19932 28356 19944
rect 28408 19972 28414 19984
rect 29638 19972 29644 19984
rect 28408 19944 29644 19972
rect 28408 19932 28414 19944
rect 29638 19932 29644 19944
rect 29696 19932 29702 19984
rect 29730 19932 29736 19984
rect 29788 19972 29794 19984
rect 29788 19944 31984 19972
rect 29788 19932 29794 19944
rect 18322 19864 18328 19916
rect 18380 19904 18386 19916
rect 19426 19904 19432 19916
rect 18380 19876 18460 19904
rect 18380 19864 18386 19876
rect 18432 19845 18460 19876
rect 18524 19876 19432 19904
rect 18524 19845 18552 19876
rect 19426 19864 19432 19876
rect 19484 19904 19490 19916
rect 19521 19907 19579 19913
rect 19521 19904 19533 19907
rect 19484 19876 19533 19904
rect 19484 19864 19490 19876
rect 19521 19873 19533 19876
rect 19567 19873 19579 19907
rect 19521 19867 19579 19873
rect 20533 19907 20591 19913
rect 20533 19873 20545 19907
rect 20579 19904 20591 19907
rect 23017 19907 23075 19913
rect 23017 19904 23029 19907
rect 20579 19876 23029 19904
rect 20579 19873 20591 19876
rect 20533 19867 20591 19873
rect 18417 19839 18475 19845
rect 18248 19808 18368 19836
rect 18141 19799 18199 19805
rect 18340 19777 18368 19808
rect 18417 19805 18429 19839
rect 18463 19805 18475 19839
rect 18417 19799 18475 19805
rect 18509 19839 18567 19845
rect 18509 19805 18521 19839
rect 18555 19805 18567 19839
rect 18509 19799 18567 19805
rect 18874 19796 18880 19848
rect 18932 19836 18938 19848
rect 19245 19839 19303 19845
rect 19245 19836 19257 19839
rect 18932 19808 19257 19836
rect 18932 19796 18938 19808
rect 19245 19805 19257 19808
rect 19291 19805 19303 19839
rect 19245 19799 19303 19805
rect 20346 19796 20352 19848
rect 20404 19836 20410 19848
rect 22388 19845 22416 19876
rect 23017 19873 23029 19876
rect 23063 19904 23075 19907
rect 23382 19904 23388 19916
rect 23063 19876 23388 19904
rect 23063 19873 23075 19876
rect 23017 19867 23075 19873
rect 23382 19864 23388 19876
rect 23440 19864 23446 19916
rect 25314 19864 25320 19916
rect 25372 19904 25378 19916
rect 28166 19904 28172 19916
rect 25372 19876 28172 19904
rect 25372 19864 25378 19876
rect 20809 19839 20867 19845
rect 20809 19836 20821 19839
rect 20404 19808 20821 19836
rect 20404 19796 20410 19808
rect 20809 19805 20821 19808
rect 20855 19805 20867 19839
rect 22189 19839 22247 19845
rect 22189 19836 22201 19839
rect 20809 19799 20867 19805
rect 22066 19808 22201 19836
rect 18325 19771 18383 19777
rect 18325 19737 18337 19771
rect 18371 19737 18383 19771
rect 18892 19768 18920 19796
rect 18325 19731 18383 19737
rect 18432 19740 18920 19768
rect 18432 19700 18460 19740
rect 21818 19728 21824 19780
rect 21876 19768 21882 19780
rect 22066 19768 22094 19808
rect 22189 19805 22201 19808
rect 22235 19805 22247 19839
rect 22189 19799 22247 19805
rect 22373 19839 22431 19845
rect 22373 19805 22385 19839
rect 22419 19805 22431 19839
rect 22373 19799 22431 19805
rect 23293 19839 23351 19845
rect 23293 19805 23305 19839
rect 23339 19836 23351 19839
rect 23474 19836 23480 19848
rect 23339 19808 23480 19836
rect 23339 19805 23351 19808
rect 23293 19799 23351 19805
rect 23474 19796 23480 19808
rect 23532 19836 23538 19848
rect 24578 19836 24584 19848
rect 23532 19808 24584 19836
rect 23532 19796 23538 19808
rect 24578 19796 24584 19808
rect 24636 19796 24642 19848
rect 25038 19796 25044 19848
rect 25096 19836 25102 19848
rect 25501 19839 25559 19845
rect 25501 19836 25513 19839
rect 25096 19808 25513 19836
rect 25096 19796 25102 19808
rect 25501 19805 25513 19808
rect 25547 19805 25559 19839
rect 25682 19836 25688 19848
rect 25643 19808 25688 19836
rect 25501 19799 25559 19805
rect 25682 19796 25688 19808
rect 25740 19796 25746 19848
rect 25777 19839 25835 19845
rect 25777 19805 25789 19839
rect 25823 19805 25835 19839
rect 25777 19799 25835 19805
rect 25869 19839 25927 19845
rect 25869 19805 25881 19839
rect 25915 19836 25927 19839
rect 25958 19836 25964 19848
rect 25915 19808 25964 19836
rect 25915 19805 25927 19808
rect 25869 19799 25927 19805
rect 24946 19768 24952 19780
rect 21876 19740 22094 19768
rect 24907 19740 24952 19768
rect 21876 19728 21882 19740
rect 24946 19728 24952 19740
rect 25004 19728 25010 19780
rect 25792 19768 25820 19799
rect 25958 19796 25964 19808
rect 26016 19796 26022 19848
rect 26602 19836 26608 19848
rect 26563 19808 26608 19836
rect 26602 19796 26608 19808
rect 26660 19796 26666 19848
rect 27706 19836 27712 19848
rect 27667 19808 27712 19836
rect 27706 19796 27712 19808
rect 27764 19796 27770 19848
rect 27890 19836 27896 19848
rect 27851 19808 27896 19836
rect 27890 19796 27896 19808
rect 27948 19796 27954 19848
rect 28000 19845 28028 19876
rect 28166 19864 28172 19876
rect 28224 19864 28230 19916
rect 30282 19864 30288 19916
rect 30340 19904 30346 19916
rect 30561 19907 30619 19913
rect 30561 19904 30573 19907
rect 30340 19876 30573 19904
rect 30340 19864 30346 19876
rect 30561 19873 30573 19876
rect 30607 19873 30619 19907
rect 31018 19904 31024 19916
rect 30561 19867 30619 19873
rect 30668 19876 31024 19904
rect 30668 19848 30696 19876
rect 31018 19864 31024 19876
rect 31076 19864 31082 19916
rect 31754 19864 31760 19916
rect 31812 19904 31818 19916
rect 31812 19876 31857 19904
rect 31812 19864 31818 19876
rect 27985 19839 28043 19845
rect 27985 19805 27997 19839
rect 28031 19805 28043 19839
rect 27985 19799 28043 19805
rect 28074 19796 28080 19848
rect 28132 19836 28138 19848
rect 28132 19808 28177 19836
rect 28132 19796 28138 19808
rect 29730 19796 29736 19848
rect 29788 19836 29794 19848
rect 30190 19836 30196 19848
rect 29788 19808 30196 19836
rect 29788 19796 29794 19808
rect 30190 19796 30196 19808
rect 30248 19836 30254 19848
rect 30469 19839 30527 19845
rect 30469 19836 30481 19839
rect 30248 19808 30481 19836
rect 30248 19796 30254 19808
rect 30469 19805 30481 19808
rect 30515 19805 30527 19839
rect 30650 19836 30656 19848
rect 30611 19808 30656 19836
rect 30469 19799 30527 19805
rect 30650 19796 30656 19808
rect 30708 19796 30714 19848
rect 30926 19836 30932 19848
rect 30887 19808 30932 19836
rect 30926 19796 30932 19808
rect 30984 19796 30990 19848
rect 31956 19845 31984 19944
rect 37734 19932 37740 19984
rect 37792 19972 37798 19984
rect 40144 19972 40172 20003
rect 40218 20000 40224 20012
rect 40276 20000 40282 20052
rect 40589 20043 40647 20049
rect 40589 20009 40601 20043
rect 40635 20040 40647 20043
rect 41230 20040 41236 20052
rect 40635 20012 41236 20040
rect 40635 20009 40647 20012
rect 40589 20003 40647 20009
rect 41230 20000 41236 20012
rect 41288 20000 41294 20052
rect 41874 20000 41880 20052
rect 41932 20040 41938 20052
rect 42153 20043 42211 20049
rect 42153 20040 42165 20043
rect 41932 20012 42165 20040
rect 41932 20000 41938 20012
rect 42153 20009 42165 20012
rect 42199 20009 42211 20043
rect 42153 20003 42211 20009
rect 37792 19944 40172 19972
rect 37792 19932 37798 19944
rect 34146 19904 34152 19916
rect 33704 19876 34152 19904
rect 31941 19839 31999 19845
rect 31941 19805 31953 19839
rect 31987 19836 31999 19839
rect 32585 19839 32643 19845
rect 32585 19836 32597 19839
rect 31987 19808 32597 19836
rect 31987 19805 31999 19808
rect 31941 19799 31999 19805
rect 32585 19805 32597 19808
rect 32631 19805 32643 19839
rect 32766 19836 32772 19848
rect 32727 19808 32772 19836
rect 32585 19799 32643 19805
rect 32766 19796 32772 19808
rect 32824 19796 32830 19848
rect 33502 19836 33508 19848
rect 33463 19808 33508 19836
rect 33502 19796 33508 19808
rect 33560 19796 33566 19848
rect 33704 19845 33732 19876
rect 34146 19864 34152 19876
rect 34204 19864 34210 19916
rect 36078 19864 36084 19916
rect 36136 19904 36142 19916
rect 36265 19907 36323 19913
rect 36265 19904 36277 19907
rect 36136 19876 36277 19904
rect 36136 19864 36142 19876
rect 36265 19873 36277 19876
rect 36311 19904 36323 19907
rect 38838 19904 38844 19916
rect 36311 19876 38844 19904
rect 36311 19873 36323 19876
rect 36265 19867 36323 19873
rect 38838 19864 38844 19876
rect 38896 19864 38902 19916
rect 40221 19907 40279 19913
rect 40221 19904 40233 19907
rect 38948 19876 40233 19904
rect 33689 19839 33747 19845
rect 33689 19805 33701 19839
rect 33735 19805 33747 19839
rect 33689 19799 33747 19805
rect 33781 19839 33839 19845
rect 33781 19805 33793 19839
rect 33827 19805 33839 19839
rect 33781 19799 33839 19805
rect 25792 19740 25912 19768
rect 25884 19712 25912 19740
rect 27614 19728 27620 19780
rect 27672 19768 27678 19780
rect 28258 19768 28264 19780
rect 27672 19740 28264 19768
rect 27672 19728 27678 19740
rect 28258 19728 28264 19740
rect 28316 19768 28322 19780
rect 28810 19768 28816 19780
rect 28316 19740 28816 19768
rect 28316 19728 28322 19740
rect 28810 19728 28816 19740
rect 28868 19728 28874 19780
rect 33796 19768 33824 19799
rect 33870 19796 33876 19848
rect 33928 19836 33934 19848
rect 33928 19808 33973 19836
rect 33928 19796 33934 19808
rect 36722 19796 36728 19848
rect 36780 19836 36786 19848
rect 37277 19839 37335 19845
rect 37277 19836 37289 19839
rect 36780 19808 37289 19836
rect 36780 19796 36786 19808
rect 37277 19805 37289 19808
rect 37323 19805 37335 19839
rect 37440 19839 37498 19845
rect 37440 19836 37452 19839
rect 37277 19799 37335 19805
rect 37384 19808 37452 19836
rect 34790 19768 34796 19780
rect 33796 19740 34796 19768
rect 34790 19728 34796 19740
rect 34848 19728 34854 19780
rect 35342 19768 35348 19780
rect 34900 19740 35348 19768
rect 34900 19712 34928 19740
rect 35342 19728 35348 19740
rect 35400 19768 35406 19780
rect 35437 19771 35495 19777
rect 35437 19768 35449 19771
rect 35400 19740 35449 19768
rect 35400 19728 35406 19740
rect 35437 19737 35449 19740
rect 35483 19737 35495 19771
rect 35437 19731 35495 19737
rect 37090 19728 37096 19780
rect 37148 19768 37154 19780
rect 37384 19768 37412 19808
rect 37440 19805 37452 19808
rect 37486 19805 37498 19839
rect 37440 19799 37498 19805
rect 37550 19796 37556 19848
rect 37608 19836 37614 19848
rect 37691 19839 37749 19845
rect 37608 19808 37653 19836
rect 37608 19796 37614 19808
rect 37691 19805 37703 19839
rect 37737 19836 37749 19839
rect 38194 19836 38200 19848
rect 37737 19808 38200 19836
rect 37737 19805 37749 19808
rect 37691 19799 37749 19805
rect 38194 19796 38200 19808
rect 38252 19836 38258 19848
rect 38381 19839 38439 19845
rect 38381 19836 38393 19839
rect 38252 19808 38393 19836
rect 38252 19796 38258 19808
rect 38381 19805 38393 19808
rect 38427 19805 38439 19839
rect 38381 19799 38439 19805
rect 37148 19740 37412 19768
rect 37148 19728 37154 19740
rect 38286 19728 38292 19780
rect 38344 19768 38350 19780
rect 38948 19777 38976 19876
rect 40221 19873 40233 19876
rect 40267 19904 40279 19907
rect 41049 19907 41107 19913
rect 41049 19904 41061 19907
rect 40267 19876 41061 19904
rect 40267 19873 40279 19876
rect 40221 19867 40279 19873
rect 41049 19873 41061 19876
rect 41095 19873 41107 19907
rect 41049 19867 41107 19873
rect 40126 19836 40132 19848
rect 40087 19808 40132 19836
rect 40126 19796 40132 19808
rect 40184 19796 40190 19848
rect 40405 19839 40463 19845
rect 40405 19805 40417 19839
rect 40451 19805 40463 19839
rect 40405 19799 40463 19805
rect 38933 19771 38991 19777
rect 38933 19768 38945 19771
rect 38344 19740 38945 19768
rect 38344 19728 38350 19740
rect 38933 19737 38945 19740
rect 38979 19737 38991 19771
rect 38933 19731 38991 19737
rect 39482 19728 39488 19780
rect 39540 19768 39546 19780
rect 40420 19768 40448 19799
rect 41601 19771 41659 19777
rect 41601 19768 41613 19771
rect 39540 19740 41613 19768
rect 39540 19728 39546 19740
rect 41601 19737 41613 19740
rect 41647 19737 41659 19771
rect 41601 19731 41659 19737
rect 17788 19672 18460 19700
rect 18693 19703 18751 19709
rect 18693 19669 18705 19703
rect 18739 19700 18751 19703
rect 20346 19700 20352 19712
rect 18739 19672 20352 19700
rect 18739 19669 18751 19672
rect 18693 19663 18751 19669
rect 20346 19660 20352 19672
rect 20404 19660 20410 19712
rect 25866 19660 25872 19712
rect 25924 19660 25930 19712
rect 28353 19703 28411 19709
rect 28353 19669 28365 19703
rect 28399 19700 28411 19703
rect 28626 19700 28632 19712
rect 28399 19672 28632 19700
rect 28399 19669 28411 19672
rect 28353 19663 28411 19669
rect 28626 19660 28632 19672
rect 28684 19660 28690 19712
rect 30837 19703 30895 19709
rect 30837 19669 30849 19703
rect 30883 19700 30895 19703
rect 31110 19700 31116 19712
rect 30883 19672 31116 19700
rect 30883 19669 30895 19672
rect 30837 19663 30895 19669
rect 31110 19660 31116 19672
rect 31168 19660 31174 19712
rect 32398 19660 32404 19712
rect 32456 19700 32462 19712
rect 32769 19703 32827 19709
rect 32769 19700 32781 19703
rect 32456 19672 32781 19700
rect 32456 19660 32462 19672
rect 32769 19669 32781 19672
rect 32815 19700 32827 19703
rect 34698 19700 34704 19712
rect 32815 19672 34704 19700
rect 32815 19669 32827 19672
rect 32769 19663 32827 19669
rect 34698 19660 34704 19672
rect 34756 19660 34762 19712
rect 34882 19700 34888 19712
rect 34843 19672 34888 19700
rect 34882 19660 34888 19672
rect 34940 19660 34946 19712
rect 1104 19610 68816 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 50294 19610
rect 50346 19558 50358 19610
rect 50410 19558 50422 19610
rect 50474 19558 50486 19610
rect 50538 19558 50550 19610
rect 50602 19558 68816 19610
rect 1104 19536 68816 19558
rect 2222 19496 2228 19508
rect 2183 19468 2228 19496
rect 2222 19456 2228 19468
rect 2280 19456 2286 19508
rect 8018 19456 8024 19508
rect 8076 19496 8082 19508
rect 8757 19499 8815 19505
rect 8076 19468 8524 19496
rect 8076 19456 8082 19468
rect 6362 19428 6368 19440
rect 6323 19400 6368 19428
rect 6362 19388 6368 19400
rect 6420 19388 6426 19440
rect 7834 19388 7840 19440
rect 7892 19428 7898 19440
rect 8202 19428 8208 19440
rect 7892 19400 8208 19428
rect 7892 19388 7898 19400
rect 8202 19388 8208 19400
rect 8260 19428 8266 19440
rect 8389 19431 8447 19437
rect 8389 19428 8401 19431
rect 8260 19400 8401 19428
rect 8260 19388 8266 19400
rect 8389 19397 8401 19400
rect 8435 19397 8447 19431
rect 8496 19428 8524 19468
rect 8757 19465 8769 19499
rect 8803 19496 8815 19499
rect 9122 19496 9128 19508
rect 8803 19468 9128 19496
rect 8803 19465 8815 19468
rect 8757 19459 8815 19465
rect 9122 19456 9128 19468
rect 9180 19456 9186 19508
rect 13541 19499 13599 19505
rect 13541 19465 13553 19499
rect 13587 19496 13599 19499
rect 13587 19468 14780 19496
rect 13587 19465 13599 19468
rect 13541 19459 13599 19465
rect 10042 19428 10048 19440
rect 8496 19400 10048 19428
rect 8389 19391 8447 19397
rect 10042 19388 10048 19400
rect 10100 19388 10106 19440
rect 14366 19428 14372 19440
rect 12176 19400 14372 19428
rect 12176 19372 12204 19400
rect 14366 19388 14372 19400
rect 14424 19388 14430 19440
rect 14752 19428 14780 19468
rect 15194 19456 15200 19508
rect 15252 19496 15258 19508
rect 15473 19499 15531 19505
rect 15473 19496 15485 19499
rect 15252 19468 15485 19496
rect 15252 19456 15258 19468
rect 15473 19465 15485 19468
rect 15519 19465 15531 19499
rect 15473 19459 15531 19465
rect 16669 19499 16727 19505
rect 16669 19465 16681 19499
rect 16715 19496 16727 19499
rect 16758 19496 16764 19508
rect 16715 19468 16764 19496
rect 16715 19465 16727 19468
rect 16669 19459 16727 19465
rect 16758 19456 16764 19468
rect 16816 19456 16822 19508
rect 18233 19499 18291 19505
rect 16865 19468 16988 19496
rect 15286 19428 15292 19440
rect 14752 19400 15292 19428
rect 15286 19388 15292 19400
rect 15344 19388 15350 19440
rect 16865 19428 16893 19468
rect 16960 19440 16988 19468
rect 18233 19465 18245 19499
rect 18279 19496 18291 19499
rect 18322 19496 18328 19508
rect 18279 19468 18328 19496
rect 18279 19465 18291 19468
rect 18233 19459 18291 19465
rect 18322 19456 18328 19468
rect 18380 19456 18386 19508
rect 24765 19499 24823 19505
rect 24765 19465 24777 19499
rect 24811 19496 24823 19499
rect 25314 19496 25320 19508
rect 24811 19468 25320 19496
rect 24811 19465 24823 19468
rect 24765 19459 24823 19465
rect 25314 19456 25320 19468
rect 25372 19456 25378 19508
rect 29546 19456 29552 19508
rect 29604 19496 29610 19508
rect 29733 19499 29791 19505
rect 29733 19496 29745 19499
rect 29604 19468 29745 19496
rect 29604 19456 29610 19468
rect 29733 19465 29745 19468
rect 29779 19465 29791 19499
rect 29733 19459 29791 19465
rect 36004 19468 36952 19496
rect 36004 19440 36032 19468
rect 15488 19400 16893 19428
rect 2409 19363 2467 19369
rect 2409 19329 2421 19363
rect 2455 19360 2467 19363
rect 2866 19360 2872 19372
rect 2455 19332 2872 19360
rect 2455 19329 2467 19332
rect 2409 19323 2467 19329
rect 2866 19320 2872 19332
rect 2924 19320 2930 19372
rect 6549 19363 6607 19369
rect 6549 19329 6561 19363
rect 6595 19360 6607 19363
rect 6914 19360 6920 19372
rect 6595 19332 6920 19360
rect 6595 19329 6607 19332
rect 6549 19323 6607 19329
rect 6914 19320 6920 19332
rect 6972 19360 6978 19372
rect 8110 19360 8116 19372
rect 6972 19332 8116 19360
rect 6972 19320 6978 19332
rect 8110 19320 8116 19332
rect 8168 19320 8174 19372
rect 8573 19363 8631 19369
rect 8573 19329 8585 19363
rect 8619 19360 8631 19363
rect 10134 19360 10140 19372
rect 8619 19332 10140 19360
rect 8619 19329 8631 19332
rect 8573 19323 8631 19329
rect 10134 19320 10140 19332
rect 10192 19320 10198 19372
rect 12158 19360 12164 19372
rect 12119 19332 12164 19360
rect 12158 19320 12164 19332
rect 12216 19320 12222 19372
rect 12428 19363 12486 19369
rect 12428 19329 12440 19363
rect 12474 19360 12486 19363
rect 14090 19360 14096 19372
rect 12474 19332 14096 19360
rect 12474 19329 12486 19332
rect 12428 19323 12486 19329
rect 14090 19320 14096 19332
rect 14148 19320 14154 19372
rect 15488 19360 15516 19400
rect 16942 19388 16948 19440
rect 17000 19388 17006 19440
rect 25590 19428 25596 19440
rect 23492 19400 25596 19428
rect 15654 19360 15660 19372
rect 15028 19332 15516 19360
rect 15615 19332 15660 19360
rect 2593 19295 2651 19301
rect 2593 19261 2605 19295
rect 2639 19292 2651 19295
rect 2774 19292 2780 19304
rect 2639 19264 2780 19292
rect 2639 19261 2651 19264
rect 2593 19255 2651 19261
rect 2774 19252 2780 19264
rect 2832 19292 2838 19304
rect 3142 19292 3148 19304
rect 2832 19264 3148 19292
rect 2832 19252 2838 19264
rect 3142 19252 3148 19264
rect 3200 19252 3206 19304
rect 6733 19295 6791 19301
rect 6733 19261 6745 19295
rect 6779 19292 6791 19295
rect 7282 19292 7288 19304
rect 6779 19264 7288 19292
rect 6779 19261 6791 19264
rect 6733 19255 6791 19261
rect 7282 19252 7288 19264
rect 7340 19252 7346 19304
rect 9766 19292 9772 19304
rect 9727 19264 9772 19292
rect 9766 19252 9772 19264
rect 9824 19292 9830 19304
rect 11974 19292 11980 19304
rect 9824 19264 11980 19292
rect 9824 19252 9830 19264
rect 11974 19252 11980 19264
rect 12032 19252 12038 19304
rect 13170 19252 13176 19304
rect 13228 19292 13234 19304
rect 14458 19292 14464 19304
rect 13228 19264 14464 19292
rect 13228 19252 13234 19264
rect 14458 19252 14464 19264
rect 14516 19292 14522 19304
rect 15028 19301 15056 19332
rect 15654 19320 15660 19332
rect 15712 19320 15718 19372
rect 16666 19320 16672 19372
rect 16724 19360 16730 19372
rect 16853 19363 16911 19369
rect 16853 19360 16865 19363
rect 16724 19332 16865 19360
rect 16724 19320 16730 19332
rect 16853 19329 16865 19332
rect 16899 19329 16911 19363
rect 16960 19360 16988 19388
rect 23492 19372 23520 19400
rect 17497 19363 17555 19369
rect 17497 19360 17509 19363
rect 16960 19332 17509 19360
rect 16853 19323 16911 19329
rect 17497 19329 17509 19332
rect 17543 19329 17555 19363
rect 17497 19323 17555 19329
rect 17681 19363 17739 19369
rect 17681 19329 17693 19363
rect 17727 19360 17739 19363
rect 17954 19360 17960 19372
rect 17727 19332 17960 19360
rect 17727 19329 17739 19332
rect 17681 19323 17739 19329
rect 17954 19320 17960 19332
rect 18012 19320 18018 19372
rect 18782 19320 18788 19372
rect 18840 19360 18846 19372
rect 20441 19363 20499 19369
rect 20441 19360 20453 19363
rect 18840 19332 20453 19360
rect 18840 19320 18846 19332
rect 20441 19329 20453 19332
rect 20487 19329 20499 19363
rect 20441 19323 20499 19329
rect 22097 19363 22155 19369
rect 22097 19329 22109 19363
rect 22143 19360 22155 19363
rect 22370 19360 22376 19372
rect 22143 19332 22376 19360
rect 22143 19329 22155 19332
rect 22097 19323 22155 19329
rect 22370 19320 22376 19332
rect 22428 19320 22434 19372
rect 23474 19360 23480 19372
rect 23435 19332 23480 19360
rect 23474 19320 23480 19332
rect 23532 19320 23538 19372
rect 24578 19360 24584 19372
rect 24539 19332 24584 19360
rect 24578 19320 24584 19332
rect 24636 19320 24642 19372
rect 25516 19369 25544 19400
rect 25590 19388 25596 19400
rect 25648 19388 25654 19440
rect 28626 19437 28632 19440
rect 28620 19428 28632 19437
rect 28587 19400 28632 19428
rect 28620 19391 28632 19400
rect 28626 19388 28632 19391
rect 28684 19388 28690 19440
rect 31846 19428 31852 19440
rect 31036 19400 31852 19428
rect 24765 19363 24823 19369
rect 24765 19329 24777 19363
rect 24811 19329 24823 19363
rect 24765 19323 24823 19329
rect 25501 19363 25559 19369
rect 25501 19329 25513 19363
rect 25547 19329 25559 19363
rect 25682 19360 25688 19372
rect 25643 19332 25688 19360
rect 25501 19323 25559 19329
rect 14737 19295 14795 19301
rect 14737 19292 14749 19295
rect 14516 19264 14749 19292
rect 14516 19252 14522 19264
rect 14737 19261 14749 19264
rect 14783 19261 14795 19295
rect 14737 19255 14795 19261
rect 15013 19295 15071 19301
rect 15013 19261 15025 19295
rect 15059 19261 15071 19295
rect 15013 19255 15071 19261
rect 16758 19252 16764 19304
rect 16816 19292 16822 19304
rect 17037 19295 17095 19301
rect 17037 19292 17049 19295
rect 16816 19264 17049 19292
rect 16816 19252 16822 19264
rect 17037 19261 17049 19264
rect 17083 19261 17095 19295
rect 17037 19255 17095 19261
rect 17126 19252 17132 19304
rect 17184 19292 17190 19304
rect 18874 19292 18880 19304
rect 17184 19264 17724 19292
rect 18835 19264 18880 19292
rect 17184 19252 17190 19264
rect 7282 19156 7288 19168
rect 7243 19128 7288 19156
rect 7282 19116 7288 19128
rect 7340 19116 7346 19168
rect 7837 19159 7895 19165
rect 7837 19125 7849 19159
rect 7883 19156 7895 19159
rect 7926 19156 7932 19168
rect 7883 19128 7932 19156
rect 7883 19125 7895 19128
rect 7837 19119 7895 19125
rect 7926 19116 7932 19128
rect 7984 19116 7990 19168
rect 13906 19116 13912 19168
rect 13964 19156 13970 19168
rect 15838 19156 15844 19168
rect 13964 19128 15844 19156
rect 13964 19116 13970 19128
rect 15838 19116 15844 19128
rect 15896 19156 15902 19168
rect 16666 19156 16672 19168
rect 15896 19128 16672 19156
rect 15896 19116 15902 19128
rect 16666 19116 16672 19128
rect 16724 19116 16730 19168
rect 17126 19116 17132 19168
rect 17184 19156 17190 19168
rect 17589 19159 17647 19165
rect 17589 19156 17601 19159
rect 17184 19128 17601 19156
rect 17184 19116 17190 19128
rect 17589 19125 17601 19128
rect 17635 19125 17647 19159
rect 17696 19156 17724 19264
rect 18874 19252 18880 19264
rect 18932 19252 18938 19304
rect 19058 19252 19064 19304
rect 19116 19292 19122 19304
rect 19153 19295 19211 19301
rect 19153 19292 19165 19295
rect 19116 19264 19165 19292
rect 19116 19252 19122 19264
rect 19153 19261 19165 19264
rect 19199 19261 19211 19295
rect 19153 19255 19211 19261
rect 20165 19295 20223 19301
rect 20165 19261 20177 19295
rect 20211 19261 20223 19295
rect 20165 19255 20223 19261
rect 20180 19224 20208 19255
rect 20990 19252 20996 19304
rect 21048 19292 21054 19304
rect 21726 19292 21732 19304
rect 21048 19264 21732 19292
rect 21048 19252 21054 19264
rect 21726 19252 21732 19264
rect 21784 19292 21790 19304
rect 21821 19295 21879 19301
rect 21821 19292 21833 19295
rect 21784 19264 21833 19292
rect 21784 19252 21790 19264
rect 21821 19261 21833 19264
rect 21867 19261 21879 19295
rect 21821 19255 21879 19261
rect 23201 19295 23259 19301
rect 23201 19261 23213 19295
rect 23247 19261 23259 19295
rect 23201 19255 23259 19261
rect 20438 19224 20444 19236
rect 20180 19196 20444 19224
rect 20438 19184 20444 19196
rect 20496 19224 20502 19236
rect 23216 19224 23244 19255
rect 23566 19252 23572 19304
rect 23624 19292 23630 19304
rect 24780 19292 24808 19323
rect 25682 19320 25688 19332
rect 25740 19320 25746 19372
rect 25777 19363 25835 19369
rect 25777 19329 25789 19363
rect 25823 19360 25835 19363
rect 25915 19363 25973 19369
rect 25823 19332 25857 19360
rect 25823 19329 25835 19332
rect 25777 19323 25835 19329
rect 25915 19329 25927 19363
rect 25961 19360 25973 19363
rect 28353 19363 28411 19369
rect 25961 19332 27108 19360
rect 25961 19329 25973 19332
rect 25915 19323 25973 19329
rect 23624 19264 24808 19292
rect 23624 19252 23630 19264
rect 25222 19252 25228 19304
rect 25280 19292 25286 19304
rect 25792 19292 25820 19323
rect 25280 19264 25820 19292
rect 25280 19252 25286 19264
rect 27080 19233 27108 19332
rect 28353 19329 28365 19363
rect 28399 19360 28411 19363
rect 28442 19360 28448 19372
rect 28399 19332 28448 19360
rect 28399 19329 28411 19332
rect 28353 19323 28411 19329
rect 28442 19320 28448 19332
rect 28500 19320 28506 19372
rect 30466 19320 30472 19372
rect 30524 19360 30530 19372
rect 31036 19369 31064 19400
rect 31846 19388 31852 19400
rect 31904 19388 31910 19440
rect 33778 19388 33784 19440
rect 33836 19428 33842 19440
rect 35986 19428 35992 19440
rect 33836 19400 35992 19428
rect 33836 19388 33842 19400
rect 35986 19388 35992 19400
rect 36044 19388 36050 19440
rect 36173 19431 36231 19437
rect 36173 19397 36185 19431
rect 36219 19428 36231 19431
rect 36814 19428 36820 19440
rect 36219 19400 36820 19428
rect 36219 19397 36231 19400
rect 36173 19391 36231 19397
rect 36814 19388 36820 19400
rect 36872 19388 36878 19440
rect 36924 19428 36952 19468
rect 37090 19456 37096 19508
rect 37148 19496 37154 19508
rect 37277 19499 37335 19505
rect 37277 19496 37289 19499
rect 37148 19468 37289 19496
rect 37148 19456 37154 19468
rect 37277 19465 37289 19468
rect 37323 19465 37335 19499
rect 37277 19459 37335 19465
rect 37645 19431 37703 19437
rect 37645 19428 37657 19431
rect 36924 19400 37657 19428
rect 37645 19397 37657 19400
rect 37691 19428 37703 19431
rect 38105 19431 38163 19437
rect 38105 19428 38117 19431
rect 37691 19400 38117 19428
rect 37691 19397 37703 19400
rect 37645 19391 37703 19397
rect 38105 19397 38117 19400
rect 38151 19397 38163 19431
rect 38933 19431 38991 19437
rect 38933 19428 38945 19431
rect 38105 19391 38163 19397
rect 38212 19400 38945 19428
rect 31021 19363 31079 19369
rect 31021 19360 31033 19363
rect 30524 19332 31033 19360
rect 30524 19320 30530 19332
rect 31021 19329 31033 19332
rect 31067 19329 31079 19363
rect 31021 19323 31079 19329
rect 31110 19320 31116 19372
rect 31168 19360 31174 19372
rect 32582 19360 32588 19372
rect 31168 19332 31213 19360
rect 32543 19332 32588 19360
rect 31168 19320 31174 19332
rect 32582 19320 32588 19332
rect 32640 19320 32646 19372
rect 33502 19320 33508 19372
rect 33560 19360 33566 19372
rect 33689 19363 33747 19369
rect 33689 19360 33701 19363
rect 33560 19332 33701 19360
rect 33560 19320 33566 19332
rect 33689 19329 33701 19332
rect 33735 19360 33747 19363
rect 34606 19360 34612 19372
rect 33735 19332 34612 19360
rect 33735 19329 33747 19332
rect 33689 19323 33747 19329
rect 34606 19320 34612 19332
rect 34664 19320 34670 19372
rect 34790 19320 34796 19372
rect 34848 19360 34854 19372
rect 34977 19363 35035 19369
rect 34977 19360 34989 19363
rect 34848 19332 34989 19360
rect 34848 19320 34854 19332
rect 34977 19329 34989 19332
rect 35023 19329 35035 19363
rect 36262 19360 36268 19372
rect 36223 19332 36268 19360
rect 34977 19323 35035 19329
rect 36262 19320 36268 19332
rect 36320 19320 36326 19372
rect 37366 19320 37372 19372
rect 37424 19360 37430 19372
rect 37461 19363 37519 19369
rect 37461 19360 37473 19363
rect 37424 19332 37473 19360
rect 37424 19320 37430 19332
rect 37461 19329 37473 19332
rect 37507 19360 37519 19363
rect 38212 19360 38240 19400
rect 38933 19397 38945 19400
rect 38979 19428 38991 19431
rect 39482 19428 39488 19440
rect 38979 19400 39488 19428
rect 38979 19397 38991 19400
rect 38933 19391 38991 19397
rect 39482 19388 39488 19400
rect 39540 19388 39546 19440
rect 40218 19388 40224 19440
rect 40276 19428 40282 19440
rect 40276 19400 40816 19428
rect 40276 19388 40282 19400
rect 37507 19332 38240 19360
rect 37507 19329 37519 19332
rect 37461 19323 37519 19329
rect 38286 19320 38292 19372
rect 38344 19360 38350 19372
rect 40788 19369 40816 19400
rect 40037 19363 40095 19369
rect 40037 19360 40049 19363
rect 38344 19332 40049 19360
rect 38344 19320 38350 19332
rect 40037 19329 40049 19332
rect 40083 19360 40095 19363
rect 40773 19363 40831 19369
rect 40083 19332 40724 19360
rect 40083 19329 40095 19332
rect 40037 19323 40095 19329
rect 31294 19252 31300 19304
rect 31352 19292 31358 19304
rect 31754 19292 31760 19304
rect 31352 19264 31760 19292
rect 31352 19252 31358 19264
rect 31754 19252 31760 19264
rect 31812 19252 31818 19304
rect 32600 19292 32628 19320
rect 33318 19292 33324 19304
rect 32600 19264 33324 19292
rect 33318 19252 33324 19264
rect 33376 19292 33382 19304
rect 33413 19295 33471 19301
rect 33413 19292 33425 19295
rect 33376 19264 33425 19292
rect 33376 19252 33382 19264
rect 33413 19261 33425 19264
rect 33459 19261 33471 19295
rect 34698 19292 34704 19304
rect 34659 19264 34704 19292
rect 33413 19255 33471 19261
rect 34698 19252 34704 19264
rect 34756 19252 34762 19304
rect 40696 19301 40724 19332
rect 40773 19329 40785 19363
rect 40819 19329 40831 19363
rect 40773 19323 40831 19329
rect 40681 19295 40739 19301
rect 40681 19261 40693 19295
rect 40727 19292 40739 19295
rect 41601 19295 41659 19301
rect 41601 19292 41613 19295
rect 40727 19264 41613 19292
rect 40727 19261 40739 19264
rect 40681 19255 40739 19261
rect 41601 19261 41613 19264
rect 41647 19261 41659 19295
rect 41601 19255 41659 19261
rect 27065 19227 27123 19233
rect 20496 19196 23244 19224
rect 23308 19196 26740 19224
rect 20496 19184 20502 19196
rect 20530 19156 20536 19168
rect 17696 19128 20536 19156
rect 17589 19119 17647 19125
rect 20530 19116 20536 19128
rect 20588 19116 20594 19168
rect 22554 19116 22560 19168
rect 22612 19156 22618 19168
rect 23308 19156 23336 19196
rect 22612 19128 23336 19156
rect 26145 19159 26203 19165
rect 22612 19116 22618 19128
rect 26145 19125 26157 19159
rect 26191 19156 26203 19159
rect 26418 19156 26424 19168
rect 26191 19128 26424 19156
rect 26191 19125 26203 19128
rect 26145 19119 26203 19125
rect 26418 19116 26424 19128
rect 26476 19116 26482 19168
rect 26712 19156 26740 19196
rect 27065 19193 27077 19227
rect 27111 19224 27123 19227
rect 27111 19196 28120 19224
rect 27111 19193 27123 19196
rect 27065 19187 27123 19193
rect 27338 19156 27344 19168
rect 26712 19128 27344 19156
rect 27338 19116 27344 19128
rect 27396 19116 27402 19168
rect 27617 19159 27675 19165
rect 27617 19125 27629 19159
rect 27663 19156 27675 19159
rect 27798 19156 27804 19168
rect 27663 19128 27804 19156
rect 27663 19125 27675 19128
rect 27617 19119 27675 19125
rect 27798 19116 27804 19128
rect 27856 19116 27862 19168
rect 28092 19156 28120 19196
rect 30098 19184 30104 19236
rect 30156 19224 30162 19236
rect 38194 19224 38200 19236
rect 30156 19196 38200 19224
rect 30156 19184 30162 19196
rect 38194 19184 38200 19196
rect 38252 19184 38258 19236
rect 30116 19156 30144 19184
rect 28092 19128 30144 19156
rect 32030 19116 32036 19168
rect 32088 19156 32094 19168
rect 32490 19156 32496 19168
rect 32088 19128 32496 19156
rect 32088 19116 32094 19128
rect 32490 19116 32496 19128
rect 32548 19156 32554 19168
rect 32677 19159 32735 19165
rect 32677 19156 32689 19159
rect 32548 19128 32689 19156
rect 32548 19116 32554 19128
rect 32677 19125 32689 19128
rect 32723 19125 32735 19159
rect 32677 19119 32735 19125
rect 34698 19116 34704 19168
rect 34756 19156 34762 19168
rect 36262 19156 36268 19168
rect 34756 19128 36268 19156
rect 34756 19116 34762 19128
rect 36262 19116 36268 19128
rect 36320 19116 36326 19168
rect 36998 19116 37004 19168
rect 37056 19156 37062 19168
rect 38473 19159 38531 19165
rect 38473 19156 38485 19159
rect 37056 19128 38485 19156
rect 37056 19116 37062 19128
rect 38473 19125 38485 19128
rect 38519 19125 38531 19159
rect 38473 19119 38531 19125
rect 41049 19159 41107 19165
rect 41049 19125 41061 19159
rect 41095 19156 41107 19159
rect 41322 19156 41328 19168
rect 41095 19128 41328 19156
rect 41095 19125 41107 19128
rect 41049 19119 41107 19125
rect 41322 19116 41328 19128
rect 41380 19116 41386 19168
rect 1104 19066 68816 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 65654 19066
rect 65706 19014 65718 19066
rect 65770 19014 65782 19066
rect 65834 19014 65846 19066
rect 65898 19014 65910 19066
rect 65962 19014 68816 19066
rect 1104 18992 68816 19014
rect 7282 18952 7288 18964
rect 7195 18924 7288 18952
rect 7282 18912 7288 18924
rect 7340 18952 7346 18964
rect 13906 18952 13912 18964
rect 7340 18924 13912 18952
rect 7340 18912 7346 18924
rect 13906 18912 13912 18924
rect 13964 18912 13970 18964
rect 14090 18952 14096 18964
rect 14051 18924 14096 18952
rect 14090 18912 14096 18924
rect 14148 18912 14154 18964
rect 15565 18955 15623 18961
rect 15565 18921 15577 18955
rect 15611 18952 15623 18955
rect 15654 18952 15660 18964
rect 15611 18924 15660 18952
rect 15611 18921 15623 18924
rect 15565 18915 15623 18921
rect 15654 18912 15660 18924
rect 15712 18912 15718 18964
rect 24765 18955 24823 18961
rect 17236 18924 22094 18952
rect 15378 18844 15384 18896
rect 15436 18884 15442 18896
rect 15746 18884 15752 18896
rect 15436 18856 15752 18884
rect 15436 18844 15442 18856
rect 15746 18844 15752 18856
rect 15804 18844 15810 18896
rect 1486 18816 1492 18828
rect 1447 18788 1492 18816
rect 1486 18776 1492 18788
rect 1544 18776 1550 18828
rect 8662 18776 8668 18828
rect 8720 18816 8726 18828
rect 10321 18819 10379 18825
rect 10321 18816 10333 18819
rect 8720 18788 10333 18816
rect 8720 18776 8726 18788
rect 10321 18785 10333 18788
rect 10367 18785 10379 18819
rect 17236 18816 17264 18924
rect 18874 18844 18880 18896
rect 18932 18884 18938 18896
rect 19337 18887 19395 18893
rect 19337 18884 19349 18887
rect 18932 18856 19349 18884
rect 18932 18844 18938 18856
rect 19337 18853 19349 18856
rect 19383 18853 19395 18887
rect 22066 18884 22094 18924
rect 24765 18921 24777 18955
rect 24811 18952 24823 18955
rect 25498 18952 25504 18964
rect 24811 18924 25504 18952
rect 24811 18921 24823 18924
rect 24765 18915 24823 18921
rect 25498 18912 25504 18924
rect 25556 18912 25562 18964
rect 25593 18955 25651 18961
rect 25593 18921 25605 18955
rect 25639 18952 25651 18955
rect 25682 18952 25688 18964
rect 25639 18924 25688 18952
rect 25639 18921 25651 18924
rect 25593 18915 25651 18921
rect 25682 18912 25688 18924
rect 25740 18912 25746 18964
rect 29638 18952 29644 18964
rect 26344 18924 29644 18952
rect 22741 18887 22799 18893
rect 22741 18884 22753 18887
rect 22066 18856 22753 18884
rect 19337 18847 19395 18853
rect 22741 18853 22753 18856
rect 22787 18884 22799 18887
rect 23845 18887 23903 18893
rect 23845 18884 23857 18887
rect 22787 18856 23857 18884
rect 22787 18853 22799 18856
rect 22741 18847 22799 18853
rect 23845 18853 23857 18856
rect 23891 18884 23903 18887
rect 24946 18884 24952 18896
rect 23891 18856 24952 18884
rect 23891 18853 23903 18856
rect 23845 18847 23903 18853
rect 24946 18844 24952 18856
rect 25004 18884 25010 18896
rect 26050 18884 26056 18896
rect 25004 18856 26056 18884
rect 25004 18844 25010 18856
rect 26050 18844 26056 18856
rect 26108 18844 26114 18896
rect 10321 18779 10379 18785
rect 12406 18788 17264 18816
rect 18601 18819 18659 18825
rect 1762 18748 1768 18760
rect 1723 18720 1768 18748
rect 1762 18708 1768 18720
rect 1820 18708 1826 18760
rect 5077 18751 5135 18757
rect 5077 18717 5089 18751
rect 5123 18748 5135 18751
rect 5629 18751 5687 18757
rect 5629 18748 5641 18751
rect 5123 18720 5641 18748
rect 5123 18717 5135 18720
rect 5077 18711 5135 18717
rect 5629 18717 5641 18720
rect 5675 18748 5687 18751
rect 5810 18748 5816 18760
rect 5675 18720 5816 18748
rect 5675 18717 5687 18720
rect 5629 18711 5687 18717
rect 5810 18708 5816 18720
rect 5868 18748 5874 18760
rect 12406 18748 12434 18788
rect 18601 18785 18613 18819
rect 18647 18816 18659 18819
rect 19978 18816 19984 18828
rect 18647 18788 19984 18816
rect 18647 18785 18659 18788
rect 18601 18779 18659 18785
rect 19978 18776 19984 18788
rect 20036 18776 20042 18828
rect 20438 18776 20444 18828
rect 20496 18816 20502 18828
rect 20533 18819 20591 18825
rect 20533 18816 20545 18819
rect 20496 18788 20545 18816
rect 20496 18776 20502 18788
rect 20533 18785 20545 18788
rect 20579 18785 20591 18819
rect 22370 18816 22376 18828
rect 20533 18779 20591 18785
rect 21560 18788 22376 18816
rect 5868 18720 12434 18748
rect 5868 18708 5874 18720
rect 13446 18708 13452 18760
rect 13504 18748 13510 18760
rect 13541 18751 13599 18757
rect 13541 18748 13553 18751
rect 13504 18720 13553 18748
rect 13504 18708 13510 18720
rect 13541 18717 13553 18720
rect 13587 18748 13599 18751
rect 14182 18748 14188 18760
rect 13587 18720 14188 18748
rect 13587 18717 13599 18720
rect 13541 18711 13599 18717
rect 14182 18708 14188 18720
rect 14240 18748 14246 18760
rect 14323 18751 14381 18757
rect 14323 18748 14335 18751
rect 14240 18720 14335 18748
rect 14240 18708 14246 18720
rect 14323 18717 14335 18720
rect 14369 18717 14381 18751
rect 14458 18748 14464 18760
rect 14419 18720 14464 18748
rect 14323 18711 14381 18717
rect 14458 18708 14464 18720
rect 14516 18708 14522 18760
rect 14550 18708 14556 18760
rect 14608 18748 14614 18760
rect 14737 18751 14795 18757
rect 14608 18720 14653 18748
rect 14608 18708 14614 18720
rect 14737 18717 14749 18751
rect 14783 18717 14795 18751
rect 14737 18711 14795 18717
rect 10318 18640 10324 18692
rect 10376 18680 10382 18692
rect 10566 18683 10624 18689
rect 10566 18680 10578 18683
rect 10376 18652 10578 18680
rect 10376 18640 10382 18652
rect 10566 18649 10578 18652
rect 10612 18649 10624 18683
rect 14752 18680 14780 18711
rect 14918 18708 14924 18760
rect 14976 18748 14982 18760
rect 15197 18751 15255 18757
rect 15197 18748 15209 18751
rect 14976 18720 15209 18748
rect 14976 18708 14982 18720
rect 15197 18717 15209 18720
rect 15243 18717 15255 18751
rect 15378 18748 15384 18760
rect 15339 18720 15384 18748
rect 15197 18711 15255 18717
rect 15378 18708 15384 18720
rect 15436 18708 15442 18760
rect 15654 18708 15660 18760
rect 15712 18748 15718 18760
rect 16025 18751 16083 18757
rect 16025 18748 16037 18751
rect 15712 18720 16037 18748
rect 15712 18708 15718 18720
rect 16025 18717 16037 18720
rect 16071 18717 16083 18751
rect 16025 18711 16083 18717
rect 17310 18708 17316 18760
rect 17368 18748 17374 18760
rect 19521 18751 19579 18757
rect 17368 18720 18460 18748
rect 17368 18708 17374 18720
rect 16114 18680 16120 18692
rect 14752 18652 16120 18680
rect 10566 18643 10624 18649
rect 16114 18640 16120 18652
rect 16172 18640 16178 18692
rect 17586 18640 17592 18692
rect 17644 18680 17650 18692
rect 18334 18683 18392 18689
rect 18334 18680 18346 18683
rect 17644 18652 18346 18680
rect 17644 18640 17650 18652
rect 18334 18649 18346 18652
rect 18380 18649 18392 18683
rect 18432 18680 18460 18720
rect 19521 18717 19533 18751
rect 19567 18748 19579 18751
rect 20162 18748 20168 18760
rect 19567 18720 20168 18748
rect 19567 18717 19579 18720
rect 19521 18711 19579 18717
rect 20162 18708 20168 18720
rect 20220 18708 20226 18760
rect 20622 18708 20628 18760
rect 20680 18748 20686 18760
rect 21560 18757 21588 18788
rect 22370 18776 22376 18788
rect 22428 18776 22434 18828
rect 25406 18816 25412 18828
rect 25240 18788 25412 18816
rect 20809 18751 20867 18757
rect 20809 18748 20821 18751
rect 20680 18720 20821 18748
rect 20680 18708 20686 18720
rect 20809 18717 20821 18720
rect 20855 18717 20867 18751
rect 20809 18711 20867 18717
rect 21545 18751 21603 18757
rect 21545 18717 21557 18751
rect 21591 18717 21603 18751
rect 21910 18748 21916 18760
rect 21871 18720 21916 18748
rect 21545 18711 21603 18717
rect 21910 18708 21916 18720
rect 21968 18708 21974 18760
rect 22465 18751 22523 18757
rect 22465 18717 22477 18751
rect 22511 18748 22523 18751
rect 22554 18748 22560 18760
rect 22511 18720 22560 18748
rect 22511 18717 22523 18720
rect 22465 18711 22523 18717
rect 22554 18708 22560 18720
rect 22612 18708 22618 18760
rect 25240 18757 25268 18788
rect 25406 18776 25412 18788
rect 25464 18776 25470 18828
rect 25498 18776 25504 18828
rect 25556 18816 25562 18828
rect 25958 18816 25964 18828
rect 25556 18788 25964 18816
rect 25556 18776 25562 18788
rect 25958 18776 25964 18788
rect 26016 18816 26022 18828
rect 26344 18816 26372 18924
rect 29638 18912 29644 18924
rect 29696 18912 29702 18964
rect 30282 18952 30288 18964
rect 30243 18924 30288 18952
rect 30282 18912 30288 18924
rect 30340 18912 30346 18964
rect 30374 18912 30380 18964
rect 30432 18952 30438 18964
rect 37642 18952 37648 18964
rect 30432 18924 37648 18952
rect 30432 18912 30438 18924
rect 37642 18912 37648 18924
rect 37700 18952 37706 18964
rect 38286 18952 38292 18964
rect 37700 18924 38292 18952
rect 37700 18912 37706 18924
rect 38286 18912 38292 18924
rect 38344 18952 38350 18964
rect 39301 18955 39359 18961
rect 39301 18952 39313 18955
rect 38344 18924 39313 18952
rect 38344 18912 38350 18924
rect 39301 18921 39313 18924
rect 39347 18921 39359 18955
rect 40218 18952 40224 18964
rect 40179 18924 40224 18952
rect 39301 18915 39359 18921
rect 40218 18912 40224 18924
rect 40276 18912 40282 18964
rect 27338 18844 27344 18896
rect 27396 18884 27402 18896
rect 30558 18884 30564 18896
rect 27396 18856 30564 18884
rect 27396 18844 27402 18856
rect 30558 18844 30564 18856
rect 30616 18844 30622 18896
rect 34790 18844 34796 18896
rect 34848 18884 34854 18896
rect 34848 18856 35020 18884
rect 34848 18844 34854 18856
rect 30006 18816 30012 18828
rect 26016 18788 26372 18816
rect 29967 18788 30012 18816
rect 26016 18776 26022 18788
rect 30006 18776 30012 18788
rect 30064 18776 30070 18828
rect 34149 18819 34207 18825
rect 34149 18785 34161 18819
rect 34195 18816 34207 18819
rect 34992 18816 35020 18856
rect 36262 18844 36268 18896
rect 36320 18884 36326 18896
rect 41782 18884 41788 18896
rect 36320 18856 37228 18884
rect 41743 18856 41788 18884
rect 36320 18844 36326 18856
rect 34195 18788 34928 18816
rect 34195 18785 34207 18788
rect 34149 18779 34207 18785
rect 25225 18751 25283 18757
rect 25225 18717 25237 18751
rect 25271 18717 25283 18751
rect 25225 18711 25283 18717
rect 26329 18751 26387 18757
rect 26329 18717 26341 18751
rect 26375 18717 26387 18751
rect 26329 18711 26387 18717
rect 21637 18683 21695 18689
rect 21637 18680 21649 18683
rect 18432 18652 21649 18680
rect 18334 18643 18392 18649
rect 21637 18649 21649 18652
rect 21683 18649 21695 18683
rect 21637 18643 21695 18649
rect 21729 18683 21787 18689
rect 21729 18649 21741 18683
rect 21775 18680 21787 18683
rect 22094 18680 22100 18692
rect 21775 18652 22100 18680
rect 21775 18649 21787 18652
rect 21729 18643 21787 18649
rect 22094 18640 22100 18652
rect 22152 18640 22158 18692
rect 25130 18640 25136 18692
rect 25188 18680 25194 18692
rect 25409 18683 25467 18689
rect 25409 18680 25421 18683
rect 25188 18652 25421 18680
rect 25188 18640 25194 18652
rect 25409 18649 25421 18652
rect 25455 18649 25467 18683
rect 26344 18680 26372 18711
rect 26418 18708 26424 18760
rect 26476 18748 26482 18760
rect 26596 18751 26654 18757
rect 26596 18748 26608 18751
rect 26476 18720 26608 18748
rect 26476 18708 26482 18720
rect 26596 18717 26608 18720
rect 26642 18717 26654 18751
rect 28442 18748 28448 18760
rect 26596 18711 26654 18717
rect 26712 18720 28448 18748
rect 26712 18680 26740 18720
rect 28442 18708 28448 18720
rect 28500 18708 28506 18760
rect 29822 18708 29828 18760
rect 29880 18748 29886 18760
rect 29917 18751 29975 18757
rect 29917 18748 29929 18751
rect 29880 18720 29929 18748
rect 29880 18708 29886 18720
rect 29917 18717 29929 18720
rect 29963 18717 29975 18751
rect 32398 18748 32404 18760
rect 29917 18711 29975 18717
rect 31726 18720 32404 18748
rect 26344 18652 26740 18680
rect 25409 18643 25467 18649
rect 2501 18615 2559 18621
rect 2501 18581 2513 18615
rect 2547 18612 2559 18615
rect 4338 18612 4344 18624
rect 2547 18584 4344 18612
rect 2547 18581 2559 18584
rect 2501 18575 2559 18581
rect 4338 18572 4344 18584
rect 4396 18572 4402 18624
rect 4982 18612 4988 18624
rect 4943 18584 4988 18612
rect 4982 18572 4988 18584
rect 5040 18572 5046 18624
rect 11698 18612 11704 18624
rect 11659 18584 11704 18612
rect 11698 18572 11704 18584
rect 11756 18572 11762 18624
rect 15378 18572 15384 18624
rect 15436 18612 15442 18624
rect 15930 18612 15936 18624
rect 15436 18584 15936 18612
rect 15436 18572 15442 18584
rect 15930 18572 15936 18584
rect 15988 18612 15994 18624
rect 16209 18615 16267 18621
rect 16209 18612 16221 18615
rect 15988 18584 16221 18612
rect 15988 18572 15994 18584
rect 16209 18581 16221 18584
rect 16255 18581 16267 18615
rect 16758 18612 16764 18624
rect 16719 18584 16764 18612
rect 16209 18575 16267 18581
rect 16758 18572 16764 18584
rect 16816 18572 16822 18624
rect 17034 18572 17040 18624
rect 17092 18612 17098 18624
rect 17218 18612 17224 18624
rect 17092 18584 17224 18612
rect 17092 18572 17098 18584
rect 17218 18572 17224 18584
rect 17276 18572 17282 18624
rect 20622 18572 20628 18624
rect 20680 18612 20686 18624
rect 21361 18615 21419 18621
rect 21361 18612 21373 18615
rect 20680 18584 21373 18612
rect 20680 18572 20686 18584
rect 21361 18581 21373 18584
rect 21407 18581 21419 18615
rect 25424 18612 25452 18643
rect 27614 18640 27620 18692
rect 27672 18680 27678 18692
rect 31726 18680 31754 18720
rect 32398 18708 32404 18720
rect 32456 18748 32462 18760
rect 33042 18748 33048 18760
rect 32456 18720 33048 18748
rect 32456 18708 32462 18720
rect 33042 18708 33048 18720
rect 33100 18708 33106 18760
rect 33137 18751 33195 18757
rect 33137 18717 33149 18751
rect 33183 18748 33195 18751
rect 33502 18748 33508 18760
rect 33183 18720 33508 18748
rect 33183 18717 33195 18720
rect 33137 18711 33195 18717
rect 33502 18708 33508 18720
rect 33560 18708 33566 18760
rect 33778 18748 33784 18760
rect 33739 18720 33784 18748
rect 33778 18708 33784 18720
rect 33836 18708 33842 18760
rect 34606 18708 34612 18760
rect 34664 18748 34670 18760
rect 34900 18757 34928 18788
rect 34992 18788 37139 18816
rect 34992 18757 35020 18788
rect 34701 18751 34759 18757
rect 34701 18748 34713 18751
rect 34664 18720 34713 18748
rect 34664 18708 34670 18720
rect 34701 18717 34713 18720
rect 34747 18717 34759 18751
rect 34701 18711 34759 18717
rect 34885 18751 34943 18757
rect 34885 18717 34897 18751
rect 34931 18717 34943 18751
rect 34885 18711 34943 18717
rect 34977 18751 35035 18757
rect 34977 18717 34989 18751
rect 35023 18717 35035 18751
rect 34977 18711 35035 18717
rect 27672 18652 31754 18680
rect 27672 18640 27678 18652
rect 32674 18640 32680 18692
rect 32732 18680 32738 18692
rect 32870 18683 32928 18689
rect 32870 18680 32882 18683
rect 32732 18652 32882 18680
rect 32732 18640 32738 18652
rect 32870 18649 32882 18652
rect 32916 18649 32928 18683
rect 33962 18680 33968 18692
rect 33923 18652 33968 18680
rect 32870 18643 32928 18649
rect 33962 18640 33968 18652
rect 34020 18640 34026 18692
rect 34716 18680 34744 18711
rect 35066 18708 35072 18760
rect 35124 18748 35130 18760
rect 36722 18748 36728 18760
rect 35124 18720 35169 18748
rect 35866 18720 36728 18748
rect 35124 18708 35130 18720
rect 35866 18680 35894 18720
rect 36722 18708 36728 18720
rect 36780 18748 36786 18760
rect 36817 18751 36875 18757
rect 36817 18748 36829 18751
rect 36780 18720 36829 18748
rect 36780 18708 36786 18720
rect 36817 18717 36829 18720
rect 36863 18717 36875 18751
rect 36998 18748 37004 18760
rect 36959 18720 37004 18748
rect 36817 18711 36875 18717
rect 36998 18708 37004 18720
rect 37056 18708 37062 18760
rect 37111 18757 37139 18788
rect 37200 18757 37228 18856
rect 41782 18844 41788 18856
rect 41840 18844 41846 18896
rect 41322 18816 41328 18828
rect 41283 18788 41328 18816
rect 41322 18776 41328 18788
rect 41380 18776 41386 18828
rect 37093 18751 37151 18757
rect 37093 18717 37105 18751
rect 37139 18717 37151 18751
rect 37093 18711 37151 18717
rect 37185 18751 37243 18757
rect 37185 18717 37197 18751
rect 37231 18717 37243 18751
rect 37550 18748 37556 18760
rect 37185 18711 37243 18717
rect 37384 18720 37556 18748
rect 35986 18680 35992 18692
rect 34716 18652 35894 18680
rect 35947 18652 35992 18680
rect 35986 18640 35992 18652
rect 36044 18640 36050 18692
rect 36173 18683 36231 18689
rect 36173 18649 36185 18683
rect 36219 18680 36231 18683
rect 36446 18680 36452 18692
rect 36219 18652 36452 18680
rect 36219 18649 36231 18652
rect 36173 18643 36231 18649
rect 36446 18640 36452 18652
rect 36504 18640 36510 18692
rect 37111 18680 37139 18711
rect 37384 18680 37412 18720
rect 37550 18708 37556 18720
rect 37608 18708 37614 18760
rect 37921 18751 37979 18757
rect 37921 18717 37933 18751
rect 37967 18748 37979 18751
rect 38746 18748 38752 18760
rect 37967 18720 38752 18748
rect 37967 18717 37979 18720
rect 37921 18711 37979 18717
rect 38746 18708 38752 18720
rect 38804 18708 38810 18760
rect 41414 18748 41420 18760
rect 41375 18720 41420 18748
rect 41414 18708 41420 18720
rect 41472 18708 41478 18760
rect 68094 18748 68100 18760
rect 68055 18720 68100 18748
rect 68094 18708 68100 18720
rect 68152 18708 68158 18760
rect 37111 18652 37412 18680
rect 37461 18683 37519 18689
rect 37461 18649 37473 18683
rect 37507 18680 37519 18683
rect 38166 18683 38224 18689
rect 38166 18680 38178 18683
rect 37507 18652 38178 18680
rect 37507 18649 37519 18652
rect 37461 18643 37519 18649
rect 38166 18649 38178 18652
rect 38212 18649 38224 18683
rect 38166 18643 38224 18649
rect 27706 18612 27712 18624
rect 25424 18584 27712 18612
rect 21361 18575 21419 18581
rect 27706 18572 27712 18584
rect 27764 18572 27770 18624
rect 28074 18572 28080 18624
rect 28132 18612 28138 18624
rect 29546 18612 29552 18624
rect 28132 18584 29552 18612
rect 28132 18572 28138 18584
rect 29546 18572 29552 18584
rect 29604 18572 29610 18624
rect 31757 18615 31815 18621
rect 31757 18581 31769 18615
rect 31803 18612 31815 18615
rect 31846 18612 31852 18624
rect 31803 18584 31852 18612
rect 31803 18581 31815 18584
rect 31757 18575 31815 18581
rect 31846 18572 31852 18584
rect 31904 18612 31910 18624
rect 33318 18612 33324 18624
rect 31904 18584 33324 18612
rect 31904 18572 31910 18584
rect 33318 18572 33324 18584
rect 33376 18572 33382 18624
rect 34606 18572 34612 18624
rect 34664 18612 34670 18624
rect 35066 18612 35072 18624
rect 34664 18584 35072 18612
rect 34664 18572 34670 18584
rect 35066 18572 35072 18584
rect 35124 18572 35130 18624
rect 35342 18612 35348 18624
rect 35303 18584 35348 18612
rect 35342 18572 35348 18584
rect 35400 18572 35406 18624
rect 36357 18615 36415 18621
rect 36357 18581 36369 18615
rect 36403 18612 36415 18615
rect 37642 18612 37648 18624
rect 36403 18584 37648 18612
rect 36403 18581 36415 18584
rect 36357 18575 36415 18581
rect 37642 18572 37648 18584
rect 37700 18572 37706 18624
rect 1104 18522 68816 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 50294 18522
rect 50346 18470 50358 18522
rect 50410 18470 50422 18522
rect 50474 18470 50486 18522
rect 50538 18470 50550 18522
rect 50602 18470 68816 18522
rect 1104 18448 68816 18470
rect 2866 18408 2872 18420
rect 2827 18380 2872 18408
rect 2866 18368 2872 18380
rect 2924 18368 2930 18420
rect 8478 18368 8484 18420
rect 8536 18408 8542 18420
rect 8754 18408 8760 18420
rect 8536 18380 8760 18408
rect 8536 18368 8542 18380
rect 8754 18368 8760 18380
rect 8812 18368 8818 18420
rect 9858 18368 9864 18420
rect 9916 18368 9922 18420
rect 10318 18408 10324 18420
rect 10279 18380 10324 18408
rect 10318 18368 10324 18380
rect 10376 18368 10382 18420
rect 10873 18411 10931 18417
rect 10873 18377 10885 18411
rect 10919 18408 10931 18411
rect 14826 18408 14832 18420
rect 10919 18380 14832 18408
rect 10919 18377 10931 18380
rect 10873 18371 10931 18377
rect 4982 18340 4988 18352
rect 3910 18312 4988 18340
rect 4982 18300 4988 18312
rect 5040 18300 5046 18352
rect 7282 18340 7288 18352
rect 6748 18312 7288 18340
rect 2409 18275 2467 18281
rect 2409 18241 2421 18275
rect 2455 18272 2467 18275
rect 2774 18272 2780 18284
rect 2455 18244 2780 18272
rect 2455 18241 2467 18244
rect 2409 18235 2467 18241
rect 2774 18232 2780 18244
rect 2832 18232 2838 18284
rect 6748 18281 6776 18312
rect 7282 18300 7288 18312
rect 7340 18300 7346 18352
rect 8662 18340 8668 18352
rect 7760 18312 8668 18340
rect 6733 18275 6791 18281
rect 6733 18241 6745 18275
rect 6779 18241 6791 18275
rect 6733 18235 6791 18241
rect 6825 18275 6883 18281
rect 6825 18241 6837 18275
rect 6871 18241 6883 18275
rect 6825 18235 6883 18241
rect 4338 18204 4344 18216
rect 4299 18176 4344 18204
rect 4338 18164 4344 18176
rect 4396 18164 4402 18216
rect 4614 18204 4620 18216
rect 4575 18176 4620 18204
rect 4614 18164 4620 18176
rect 4672 18164 4678 18216
rect 2314 18068 2320 18080
rect 2275 18040 2320 18068
rect 2314 18028 2320 18040
rect 2372 18028 2378 18080
rect 6454 18068 6460 18080
rect 6415 18040 6460 18068
rect 6454 18028 6460 18040
rect 6512 18028 6518 18080
rect 6840 18068 6868 18235
rect 6914 18232 6920 18284
rect 6972 18272 6978 18284
rect 6972 18244 7017 18272
rect 6972 18232 6978 18244
rect 7098 18232 7104 18284
rect 7156 18272 7162 18284
rect 7156 18244 7201 18272
rect 7156 18232 7162 18244
rect 7650 18164 7656 18216
rect 7708 18204 7714 18216
rect 7760 18213 7788 18312
rect 8662 18300 8668 18312
rect 8720 18300 8726 18352
rect 9876 18340 9904 18368
rect 9692 18312 9904 18340
rect 8018 18281 8024 18284
rect 8012 18235 8024 18281
rect 8076 18272 8082 18284
rect 9692 18281 9720 18312
rect 10226 18300 10232 18352
rect 10284 18340 10290 18352
rect 10888 18340 10916 18371
rect 14826 18368 14832 18380
rect 14884 18368 14890 18420
rect 17126 18408 17132 18420
rect 17052 18380 17132 18408
rect 10284 18312 10916 18340
rect 14645 18343 14703 18349
rect 10284 18300 10290 18312
rect 14645 18309 14657 18343
rect 14691 18340 14703 18343
rect 15194 18340 15200 18352
rect 14691 18312 15200 18340
rect 14691 18309 14703 18312
rect 14645 18303 14703 18309
rect 15194 18300 15200 18312
rect 15252 18300 15258 18352
rect 16206 18340 16212 18352
rect 16040 18312 16212 18340
rect 9677 18275 9735 18281
rect 8076 18244 8112 18272
rect 8018 18232 8024 18235
rect 8076 18232 8082 18244
rect 9677 18241 9689 18275
rect 9723 18241 9735 18275
rect 9858 18272 9864 18284
rect 9819 18244 9864 18272
rect 9677 18235 9735 18241
rect 9858 18232 9864 18244
rect 9916 18232 9922 18284
rect 9953 18275 10011 18281
rect 9953 18241 9965 18275
rect 9999 18241 10011 18275
rect 9953 18235 10011 18241
rect 10045 18275 10103 18281
rect 10045 18241 10057 18275
rect 10091 18272 10103 18275
rect 10244 18272 10272 18300
rect 10091 18244 10272 18272
rect 14829 18275 14887 18281
rect 10091 18241 10103 18244
rect 10045 18235 10103 18241
rect 14829 18241 14841 18275
rect 14875 18241 14887 18275
rect 14829 18235 14887 18241
rect 15013 18275 15071 18281
rect 15013 18241 15025 18275
rect 15059 18272 15071 18275
rect 15378 18272 15384 18284
rect 15059 18244 15384 18272
rect 15059 18241 15071 18244
rect 15013 18235 15071 18241
rect 7745 18207 7803 18213
rect 7745 18204 7757 18207
rect 7708 18176 7757 18204
rect 7708 18164 7714 18176
rect 7745 18173 7757 18176
rect 7791 18173 7803 18207
rect 7745 18167 7803 18173
rect 8754 18164 8760 18216
rect 8812 18204 8818 18216
rect 9968 18204 9996 18235
rect 11054 18204 11060 18216
rect 8812 18176 11060 18204
rect 8812 18164 8818 18176
rect 11054 18164 11060 18176
rect 11112 18164 11118 18216
rect 14090 18164 14096 18216
rect 14148 18204 14154 18216
rect 14642 18204 14648 18216
rect 14148 18176 14648 18204
rect 14148 18164 14154 18176
rect 14642 18164 14648 18176
rect 14700 18204 14706 18216
rect 14844 18204 14872 18235
rect 15378 18232 15384 18244
rect 15436 18232 15442 18284
rect 15654 18232 15660 18284
rect 15712 18281 15718 18284
rect 15712 18275 15761 18281
rect 15712 18241 15715 18275
rect 15749 18241 15761 18275
rect 15712 18235 15761 18241
rect 15841 18275 15899 18281
rect 15841 18241 15853 18275
rect 15887 18241 15899 18275
rect 15841 18235 15899 18241
rect 15938 18275 15996 18281
rect 15938 18241 15950 18275
rect 15984 18272 15996 18275
rect 16040 18272 16068 18312
rect 16206 18300 16212 18312
rect 16264 18300 16270 18352
rect 15984 18244 16068 18272
rect 15984 18241 15996 18244
rect 15938 18235 15996 18241
rect 15712 18232 15718 18235
rect 15470 18204 15476 18216
rect 14700 18176 15476 18204
rect 14700 18164 14706 18176
rect 15470 18164 15476 18176
rect 15528 18164 15534 18216
rect 15856 18204 15884 18235
rect 16114 18232 16120 18284
rect 16172 18272 16178 18284
rect 16945 18275 17003 18281
rect 16945 18272 16957 18275
rect 16172 18244 16957 18272
rect 16172 18232 16178 18244
rect 16945 18241 16957 18244
rect 16991 18241 17003 18275
rect 17052 18272 17080 18380
rect 17126 18368 17132 18380
rect 17184 18368 17190 18420
rect 17586 18408 17592 18420
rect 17547 18380 17592 18408
rect 17586 18368 17592 18380
rect 17644 18368 17650 18420
rect 18325 18411 18383 18417
rect 18325 18377 18337 18411
rect 18371 18408 18383 18411
rect 18690 18408 18696 18420
rect 18371 18380 18696 18408
rect 18371 18377 18383 18380
rect 18325 18371 18383 18377
rect 18690 18368 18696 18380
rect 18748 18408 18754 18420
rect 19242 18408 19248 18420
rect 18748 18380 19248 18408
rect 18748 18368 18754 18380
rect 19242 18368 19248 18380
rect 19300 18368 19306 18420
rect 21910 18368 21916 18420
rect 21968 18408 21974 18420
rect 30374 18408 30380 18420
rect 21968 18380 30380 18408
rect 21968 18368 21974 18380
rect 30374 18368 30380 18380
rect 30432 18368 30438 18420
rect 32125 18411 32183 18417
rect 32125 18408 32137 18411
rect 31726 18380 32137 18408
rect 19429 18343 19487 18349
rect 19429 18309 19441 18343
rect 19475 18340 19487 18343
rect 20134 18343 20192 18349
rect 20134 18340 20146 18343
rect 19475 18312 20146 18340
rect 19475 18309 19487 18312
rect 19429 18303 19487 18309
rect 20134 18309 20146 18312
rect 20180 18309 20192 18343
rect 23566 18340 23572 18352
rect 20134 18303 20192 18309
rect 22066 18312 23572 18340
rect 22066 18284 22094 18312
rect 23566 18300 23572 18312
rect 23624 18300 23630 18352
rect 23692 18343 23750 18349
rect 23692 18309 23704 18343
rect 23738 18340 23750 18343
rect 24397 18343 24455 18349
rect 24397 18340 24409 18343
rect 23738 18312 24409 18340
rect 23738 18309 23750 18312
rect 23692 18303 23750 18309
rect 24397 18309 24409 18312
rect 24443 18309 24455 18343
rect 25130 18340 25136 18352
rect 24397 18303 24455 18309
rect 24688 18312 25136 18340
rect 17108 18275 17166 18281
rect 17108 18272 17120 18275
rect 17052 18244 17120 18272
rect 16945 18235 17003 18241
rect 17108 18241 17120 18244
rect 17154 18241 17166 18275
rect 17108 18235 17166 18241
rect 17221 18275 17279 18281
rect 17221 18241 17233 18275
rect 17267 18241 17279 18275
rect 17221 18235 17279 18241
rect 17313 18275 17371 18281
rect 17402 18275 17408 18284
rect 17313 18241 17325 18275
rect 17359 18247 17408 18275
rect 17359 18241 17371 18247
rect 17313 18235 17371 18241
rect 16206 18204 16212 18216
rect 15856 18176 16212 18204
rect 16206 18164 16212 18176
rect 16264 18204 16270 18216
rect 17223 18204 17251 18235
rect 17402 18232 17408 18247
rect 17460 18232 17466 18284
rect 18782 18272 18788 18284
rect 18743 18244 18788 18272
rect 18782 18232 18788 18244
rect 18840 18232 18846 18284
rect 18969 18275 19027 18281
rect 18969 18241 18981 18275
rect 19015 18241 19027 18275
rect 18969 18235 19027 18241
rect 16264 18176 17251 18204
rect 16264 18164 16270 18176
rect 18984 18136 19012 18235
rect 19058 18232 19064 18284
rect 19116 18272 19122 18284
rect 19242 18281 19248 18284
rect 19199 18275 19248 18281
rect 19116 18244 19161 18272
rect 19116 18232 19122 18244
rect 19199 18241 19211 18275
rect 19245 18241 19248 18275
rect 19199 18235 19248 18241
rect 19242 18232 19248 18235
rect 19300 18232 19306 18284
rect 19889 18275 19947 18281
rect 19889 18241 19901 18275
rect 19935 18272 19947 18275
rect 19978 18272 19984 18284
rect 19935 18244 19984 18272
rect 19935 18241 19947 18244
rect 19889 18235 19947 18241
rect 19978 18232 19984 18244
rect 20036 18232 20042 18284
rect 21726 18232 21732 18284
rect 21784 18272 21790 18284
rect 21821 18275 21879 18281
rect 21821 18272 21833 18275
rect 21784 18244 21833 18272
rect 21784 18232 21790 18244
rect 21821 18241 21833 18244
rect 21867 18241 21879 18275
rect 21821 18235 21879 18241
rect 22002 18232 22008 18284
rect 22060 18244 22094 18284
rect 24688 18281 24716 18312
rect 25130 18300 25136 18312
rect 25188 18300 25194 18352
rect 25406 18300 25412 18352
rect 25464 18340 25470 18352
rect 25593 18343 25651 18349
rect 25593 18340 25605 18343
rect 25464 18312 25605 18340
rect 25464 18300 25470 18312
rect 25593 18309 25605 18312
rect 25639 18309 25651 18343
rect 27614 18340 27620 18352
rect 27575 18312 27620 18340
rect 25593 18303 25651 18309
rect 27614 18300 27620 18312
rect 27672 18300 27678 18352
rect 28804 18343 28862 18349
rect 27724 18312 28028 18340
rect 24673 18275 24731 18281
rect 22060 18232 22066 18244
rect 24673 18241 24685 18275
rect 24719 18241 24731 18275
rect 24673 18235 24731 18241
rect 24765 18275 24823 18281
rect 24765 18241 24777 18275
rect 24811 18241 24823 18275
rect 24765 18235 24823 18241
rect 23934 18204 23940 18216
rect 23895 18176 23940 18204
rect 23934 18164 23940 18176
rect 23992 18164 23998 18216
rect 24780 18204 24808 18235
rect 24854 18232 24860 18284
rect 24912 18272 24918 18284
rect 24912 18244 24957 18272
rect 24912 18232 24918 18244
rect 25038 18232 25044 18284
rect 25096 18272 25102 18284
rect 25096 18244 25141 18272
rect 25096 18232 25102 18244
rect 25682 18232 25688 18284
rect 25740 18272 25746 18284
rect 25777 18275 25835 18281
rect 25777 18272 25789 18275
rect 25740 18244 25789 18272
rect 25740 18232 25746 18244
rect 25777 18241 25789 18244
rect 25823 18272 25835 18275
rect 25823 18244 26004 18272
rect 25823 18241 25835 18244
rect 25777 18235 25835 18241
rect 25222 18204 25228 18216
rect 24780 18176 25228 18204
rect 25222 18164 25228 18176
rect 25280 18164 25286 18216
rect 25976 18204 26004 18244
rect 26050 18232 26056 18284
rect 26108 18272 26114 18284
rect 27724 18272 27752 18312
rect 26108 18244 27752 18272
rect 27893 18275 27951 18281
rect 26108 18232 26114 18244
rect 27893 18241 27905 18275
rect 27939 18241 27951 18275
rect 28000 18272 28028 18312
rect 28804 18309 28816 18343
rect 28850 18340 28862 18343
rect 28994 18340 29000 18352
rect 28850 18312 29000 18340
rect 28850 18309 28862 18312
rect 28804 18303 28862 18309
rect 28994 18300 29000 18312
rect 29052 18300 29058 18352
rect 29638 18300 29644 18352
rect 29696 18340 29702 18352
rect 30190 18340 30196 18352
rect 29696 18312 30196 18340
rect 29696 18300 29702 18312
rect 30190 18300 30196 18312
rect 30248 18300 30254 18352
rect 31726 18272 31754 18380
rect 32125 18377 32137 18380
rect 32171 18377 32183 18411
rect 32125 18371 32183 18377
rect 28000 18244 31754 18272
rect 32140 18272 32168 18371
rect 33962 18368 33968 18420
rect 34020 18408 34026 18420
rect 35894 18408 35900 18420
rect 34020 18380 35900 18408
rect 34020 18368 34026 18380
rect 35894 18368 35900 18380
rect 35952 18408 35958 18420
rect 36173 18411 36231 18417
rect 36173 18408 36185 18411
rect 35952 18380 36185 18408
rect 35952 18368 35958 18380
rect 36173 18377 36185 18380
rect 36219 18377 36231 18411
rect 36173 18371 36231 18377
rect 40218 18368 40224 18420
rect 40276 18408 40282 18420
rect 40405 18411 40463 18417
rect 40405 18408 40417 18411
rect 40276 18380 40417 18408
rect 40276 18368 40282 18380
rect 40405 18377 40417 18380
rect 40451 18377 40463 18411
rect 40405 18371 40463 18377
rect 33594 18300 33600 18352
rect 33652 18340 33658 18352
rect 35060 18343 35118 18349
rect 33652 18312 34514 18340
rect 33652 18300 33658 18312
rect 32677 18275 32735 18281
rect 32677 18272 32689 18275
rect 32140 18244 32689 18272
rect 27893 18235 27951 18241
rect 32677 18241 32689 18244
rect 32723 18241 32735 18275
rect 34486 18272 34514 18312
rect 35060 18309 35072 18343
rect 35106 18340 35118 18343
rect 35342 18340 35348 18352
rect 35106 18312 35348 18340
rect 35106 18309 35118 18312
rect 35060 18303 35118 18309
rect 35342 18300 35348 18312
rect 35400 18300 35406 18352
rect 37550 18300 37556 18352
rect 37608 18340 37614 18352
rect 38105 18343 38163 18349
rect 37608 18312 37780 18340
rect 37608 18300 37614 18312
rect 34793 18275 34851 18281
rect 34793 18272 34805 18275
rect 34486 18244 34805 18272
rect 32677 18235 32735 18241
rect 34793 18241 34805 18244
rect 34839 18272 34851 18275
rect 36078 18272 36084 18284
rect 34839 18244 36084 18272
rect 34839 18241 34851 18244
rect 34793 18235 34851 18241
rect 27614 18204 27620 18216
rect 25976 18176 27620 18204
rect 27614 18164 27620 18176
rect 27672 18204 27678 18216
rect 27709 18207 27767 18213
rect 27709 18204 27721 18207
rect 27672 18176 27721 18204
rect 27672 18164 27678 18176
rect 27709 18173 27721 18176
rect 27755 18173 27767 18207
rect 27709 18167 27767 18173
rect 19610 18136 19616 18148
rect 18984 18108 19616 18136
rect 19610 18096 19616 18108
rect 19668 18096 19674 18148
rect 22002 18136 22008 18148
rect 21963 18108 22008 18136
rect 22002 18096 22008 18108
rect 22060 18096 22066 18148
rect 24578 18096 24584 18148
rect 24636 18136 24642 18148
rect 27908 18136 27936 18235
rect 36078 18232 36084 18244
rect 36136 18232 36142 18284
rect 36722 18232 36728 18284
rect 36780 18272 36786 18284
rect 37461 18275 37519 18281
rect 37461 18272 37473 18275
rect 36780 18244 37473 18272
rect 36780 18232 36786 18244
rect 37461 18241 37473 18244
rect 37507 18241 37519 18275
rect 37642 18272 37648 18284
rect 37603 18244 37648 18272
rect 37461 18235 37519 18241
rect 37642 18232 37648 18244
rect 37700 18232 37706 18284
rect 37752 18281 37780 18312
rect 38105 18309 38117 18343
rect 38151 18340 38163 18343
rect 39270 18343 39328 18349
rect 39270 18340 39282 18343
rect 38151 18312 39282 18340
rect 38151 18309 38163 18312
rect 38105 18303 38163 18309
rect 39270 18309 39282 18312
rect 39316 18309 39328 18343
rect 39270 18303 39328 18309
rect 37737 18275 37795 18281
rect 37737 18241 37749 18275
rect 37783 18241 37795 18275
rect 37737 18235 37795 18241
rect 37826 18232 37832 18284
rect 37884 18272 37890 18284
rect 37884 18244 37929 18272
rect 37884 18232 37890 18244
rect 38838 18232 38844 18284
rect 38896 18272 38902 18284
rect 39025 18275 39083 18281
rect 39025 18272 39037 18275
rect 38896 18244 39037 18272
rect 38896 18232 38902 18244
rect 39025 18241 39037 18244
rect 39071 18241 39083 18275
rect 39025 18235 39083 18241
rect 28442 18164 28448 18216
rect 28500 18204 28506 18216
rect 28537 18207 28595 18213
rect 28537 18204 28549 18207
rect 28500 18176 28549 18204
rect 28500 18164 28506 18176
rect 28537 18173 28549 18176
rect 28583 18173 28595 18207
rect 28537 18167 28595 18173
rect 29546 18164 29552 18216
rect 29604 18204 29610 18216
rect 33962 18204 33968 18216
rect 29604 18176 33968 18204
rect 29604 18164 29610 18176
rect 33962 18164 33968 18176
rect 34020 18204 34026 18216
rect 34333 18207 34391 18213
rect 34333 18204 34345 18207
rect 34020 18176 34345 18204
rect 34020 18164 34026 18176
rect 34333 18173 34345 18176
rect 34379 18173 34391 18207
rect 34333 18167 34391 18173
rect 30742 18136 30748 18148
rect 24636 18108 27936 18136
rect 29472 18108 30748 18136
rect 24636 18096 24642 18108
rect 8754 18068 8760 18080
rect 6840 18040 8760 18068
rect 8754 18028 8760 18040
rect 8812 18028 8818 18080
rect 9122 18068 9128 18080
rect 9083 18040 9128 18068
rect 9122 18028 9128 18040
rect 9180 18028 9186 18080
rect 13998 18028 14004 18080
rect 14056 18068 14062 18080
rect 14093 18071 14151 18077
rect 14093 18068 14105 18071
rect 14056 18040 14105 18068
rect 14056 18028 14062 18040
rect 14093 18037 14105 18040
rect 14139 18068 14151 18071
rect 14918 18068 14924 18080
rect 14139 18040 14924 18068
rect 14139 18037 14151 18040
rect 14093 18031 14151 18037
rect 14918 18028 14924 18040
rect 14976 18028 14982 18080
rect 15378 18028 15384 18080
rect 15436 18068 15442 18080
rect 15473 18071 15531 18077
rect 15473 18068 15485 18071
rect 15436 18040 15485 18068
rect 15436 18028 15442 18040
rect 15473 18037 15485 18040
rect 15519 18037 15531 18071
rect 21266 18068 21272 18080
rect 21227 18040 21272 18068
rect 15473 18031 15531 18037
rect 21266 18028 21272 18040
rect 21324 18028 21330 18080
rect 22557 18071 22615 18077
rect 22557 18037 22569 18071
rect 22603 18068 22615 18071
rect 23658 18068 23664 18080
rect 22603 18040 23664 18068
rect 22603 18037 22615 18040
rect 22557 18031 22615 18037
rect 23658 18028 23664 18040
rect 23716 18068 23722 18080
rect 24596 18068 24624 18096
rect 23716 18040 24624 18068
rect 25961 18071 26019 18077
rect 23716 18028 23722 18040
rect 25961 18037 25973 18071
rect 26007 18068 26019 18071
rect 26050 18068 26056 18080
rect 26007 18040 26056 18068
rect 26007 18037 26019 18040
rect 25961 18031 26019 18037
rect 26050 18028 26056 18040
rect 26108 18028 26114 18080
rect 27706 18068 27712 18080
rect 27667 18040 27712 18068
rect 27706 18028 27712 18040
rect 27764 18028 27770 18080
rect 28077 18071 28135 18077
rect 28077 18037 28089 18071
rect 28123 18068 28135 18071
rect 29472 18068 29500 18108
rect 30742 18096 30748 18108
rect 30800 18096 30806 18148
rect 33413 18139 33471 18145
rect 33413 18136 33425 18139
rect 32554 18108 33425 18136
rect 28123 18040 29500 18068
rect 28123 18037 28135 18040
rect 28077 18031 28135 18037
rect 29822 18028 29828 18080
rect 29880 18068 29886 18080
rect 29917 18071 29975 18077
rect 29917 18068 29929 18071
rect 29880 18040 29929 18068
rect 29880 18028 29886 18040
rect 29917 18037 29929 18040
rect 29963 18037 29975 18071
rect 29917 18031 29975 18037
rect 30190 18028 30196 18080
rect 30248 18068 30254 18080
rect 32554 18068 32582 18108
rect 33413 18105 33425 18108
rect 33459 18136 33471 18139
rect 33870 18136 33876 18148
rect 33459 18108 33876 18136
rect 33459 18105 33471 18108
rect 33413 18099 33471 18105
rect 33870 18096 33876 18108
rect 33928 18096 33934 18148
rect 30248 18040 32582 18068
rect 32861 18071 32919 18077
rect 30248 18028 30254 18040
rect 32861 18037 32873 18071
rect 32907 18068 32919 18071
rect 34698 18068 34704 18080
rect 32907 18040 34704 18068
rect 32907 18037 32919 18040
rect 32861 18031 32919 18037
rect 34698 18028 34704 18040
rect 34756 18028 34762 18080
rect 36446 18028 36452 18080
rect 36504 18068 36510 18080
rect 36633 18071 36691 18077
rect 36633 18068 36645 18071
rect 36504 18040 36645 18068
rect 36504 18028 36510 18040
rect 36633 18037 36645 18040
rect 36679 18068 36691 18071
rect 37734 18068 37740 18080
rect 36679 18040 37740 18068
rect 36679 18037 36691 18040
rect 36633 18031 36691 18037
rect 37734 18028 37740 18040
rect 37792 18028 37798 18080
rect 1104 17978 68816 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 65654 17978
rect 65706 17926 65718 17978
rect 65770 17926 65782 17978
rect 65834 17926 65846 17978
rect 65898 17926 65910 17978
rect 65962 17926 68816 17978
rect 1104 17904 68816 17926
rect 1854 17824 1860 17876
rect 1912 17864 1918 17876
rect 1949 17867 2007 17873
rect 1949 17864 1961 17867
rect 1912 17836 1961 17864
rect 1912 17824 1918 17836
rect 1949 17833 1961 17836
rect 1995 17833 2007 17867
rect 1949 17827 2007 17833
rect 4614 17824 4620 17876
rect 4672 17864 4678 17876
rect 7650 17864 7656 17876
rect 4672 17836 7656 17864
rect 4672 17824 4678 17836
rect 2866 17728 2872 17740
rect 1964 17700 2872 17728
rect 1964 17669 1992 17700
rect 2866 17688 2872 17700
rect 2924 17688 2930 17740
rect 1949 17663 2007 17669
rect 1949 17629 1961 17663
rect 1995 17629 2007 17663
rect 1949 17623 2007 17629
rect 2133 17663 2191 17669
rect 2133 17629 2145 17663
rect 2179 17660 2191 17663
rect 2314 17660 2320 17672
rect 2179 17632 2320 17660
rect 2179 17629 2191 17632
rect 2133 17623 2191 17629
rect 2314 17620 2320 17632
rect 2372 17620 2378 17672
rect 6656 17669 6684 17836
rect 7650 17824 7656 17836
rect 7708 17824 7714 17876
rect 8018 17864 8024 17876
rect 7979 17836 8024 17864
rect 8018 17824 8024 17836
rect 8076 17824 8082 17876
rect 9858 17824 9864 17876
rect 9916 17864 9922 17876
rect 10321 17867 10379 17873
rect 10321 17864 10333 17867
rect 9916 17836 10333 17864
rect 9916 17824 9922 17836
rect 10321 17833 10333 17836
rect 10367 17833 10379 17867
rect 14090 17864 14096 17876
rect 14051 17836 14096 17864
rect 10321 17827 10379 17833
rect 14090 17824 14096 17836
rect 14148 17824 14154 17876
rect 14826 17824 14832 17876
rect 14884 17864 14890 17876
rect 18782 17864 18788 17876
rect 14884 17836 18788 17864
rect 14884 17824 14890 17836
rect 18782 17824 18788 17836
rect 18840 17824 18846 17876
rect 19610 17864 19616 17876
rect 19571 17836 19616 17864
rect 19610 17824 19616 17836
rect 19668 17824 19674 17876
rect 21450 17864 21456 17876
rect 21411 17836 21456 17864
rect 21450 17824 21456 17836
rect 21508 17824 21514 17876
rect 22554 17824 22560 17876
rect 22612 17864 22618 17876
rect 22833 17867 22891 17873
rect 22833 17864 22845 17867
rect 22612 17836 22845 17864
rect 22612 17824 22618 17836
rect 22833 17833 22845 17836
rect 22879 17864 22891 17867
rect 23106 17864 23112 17876
rect 22879 17836 23112 17864
rect 22879 17833 22891 17836
rect 22833 17827 22891 17833
rect 23106 17824 23112 17836
rect 23164 17824 23170 17876
rect 23566 17824 23572 17876
rect 23624 17864 23630 17876
rect 23753 17867 23811 17873
rect 23753 17864 23765 17867
rect 23624 17836 23765 17864
rect 23624 17824 23630 17836
rect 23753 17833 23765 17836
rect 23799 17833 23811 17867
rect 23753 17827 23811 17833
rect 24765 17867 24823 17873
rect 24765 17833 24777 17867
rect 24811 17864 24823 17867
rect 24854 17864 24860 17876
rect 24811 17836 24860 17864
rect 24811 17833 24823 17836
rect 24765 17827 24823 17833
rect 24854 17824 24860 17836
rect 24912 17824 24918 17876
rect 27614 17824 27620 17876
rect 27672 17864 27678 17876
rect 27985 17867 28043 17873
rect 27985 17864 27997 17867
rect 27672 17836 27997 17864
rect 27672 17824 27678 17836
rect 27985 17833 27997 17836
rect 28031 17833 28043 17867
rect 32674 17864 32680 17876
rect 32635 17836 32680 17864
rect 27985 17827 28043 17833
rect 32674 17824 32680 17836
rect 32732 17824 32738 17876
rect 32968 17836 33364 17864
rect 9950 17796 9956 17808
rect 7392 17768 9956 17796
rect 7392 17669 7420 17768
rect 9950 17756 9956 17768
rect 10008 17756 10014 17808
rect 15654 17756 15660 17808
rect 15712 17796 15718 17808
rect 16666 17796 16672 17808
rect 15712 17768 16672 17796
rect 15712 17756 15718 17768
rect 16666 17756 16672 17768
rect 16724 17796 16730 17808
rect 17773 17799 17831 17805
rect 17773 17796 17785 17799
rect 16724 17768 17785 17796
rect 16724 17756 16730 17768
rect 17773 17765 17785 17768
rect 17819 17796 17831 17799
rect 20898 17796 20904 17808
rect 17819 17768 20904 17796
rect 17819 17765 17831 17768
rect 17773 17759 17831 17765
rect 20898 17756 20904 17768
rect 20956 17756 20962 17808
rect 20993 17799 21051 17805
rect 20993 17765 21005 17799
rect 21039 17796 21051 17799
rect 21910 17796 21916 17808
rect 21039 17768 21916 17796
rect 21039 17765 21051 17768
rect 20993 17759 21051 17765
rect 21910 17756 21916 17768
rect 21968 17756 21974 17808
rect 23934 17756 23940 17808
rect 23992 17796 23998 17808
rect 25682 17796 25688 17808
rect 23992 17768 25688 17796
rect 23992 17756 23998 17768
rect 25682 17756 25688 17768
rect 25740 17796 25746 17808
rect 31389 17799 31447 17805
rect 25740 17768 26648 17796
rect 25740 17756 25746 17768
rect 8754 17728 8760 17740
rect 7668 17700 8760 17728
rect 7668 17669 7696 17700
rect 8754 17688 8760 17700
rect 8812 17688 8818 17740
rect 12158 17728 12164 17740
rect 12119 17700 12164 17728
rect 12158 17688 12164 17700
rect 12216 17688 12222 17740
rect 16206 17728 16212 17740
rect 16119 17700 16212 17728
rect 16206 17688 16212 17700
rect 16264 17728 16270 17740
rect 19058 17728 19064 17740
rect 16264 17700 19064 17728
rect 16264 17688 16270 17700
rect 19058 17688 19064 17700
rect 19116 17688 19122 17740
rect 25222 17688 25228 17740
rect 25280 17728 25286 17740
rect 26326 17728 26332 17740
rect 25280 17700 25820 17728
rect 25280 17688 25286 17700
rect 6374 17663 6432 17669
rect 6374 17629 6386 17663
rect 6420 17629 6432 17663
rect 6374 17623 6432 17629
rect 6641 17663 6699 17669
rect 6641 17629 6653 17663
rect 6687 17629 6699 17663
rect 6641 17623 6699 17629
rect 7377 17663 7435 17669
rect 7377 17629 7389 17663
rect 7423 17629 7435 17663
rect 7377 17623 7435 17629
rect 7561 17663 7619 17669
rect 7561 17629 7573 17663
rect 7607 17629 7619 17663
rect 7561 17623 7619 17629
rect 7653 17663 7711 17669
rect 7653 17629 7665 17663
rect 7699 17629 7711 17663
rect 7653 17623 7711 17629
rect 1854 17552 1860 17604
rect 1912 17592 1918 17604
rect 6380 17592 6408 17623
rect 6454 17592 6460 17604
rect 1912 17564 5396 17592
rect 6380 17564 6460 17592
rect 1912 17552 1918 17564
rect 5258 17524 5264 17536
rect 5219 17496 5264 17524
rect 5258 17484 5264 17496
rect 5316 17484 5322 17536
rect 5368 17524 5396 17564
rect 6454 17552 6460 17564
rect 6512 17552 6518 17604
rect 7576 17592 7604 17623
rect 7742 17620 7748 17672
rect 7800 17660 7806 17672
rect 7800 17632 7845 17660
rect 7800 17620 7806 17632
rect 9214 17620 9220 17672
rect 9272 17660 9278 17672
rect 9309 17663 9367 17669
rect 9309 17660 9321 17663
rect 9272 17632 9321 17660
rect 9272 17620 9278 17632
rect 9309 17629 9321 17632
rect 9355 17660 9367 17663
rect 9953 17663 10011 17669
rect 9953 17660 9965 17663
rect 9355 17632 9965 17660
rect 9355 17629 9367 17632
rect 9309 17623 9367 17629
rect 9953 17629 9965 17632
rect 9999 17629 10011 17663
rect 9953 17623 10011 17629
rect 10137 17663 10195 17669
rect 10137 17629 10149 17663
rect 10183 17660 10195 17663
rect 11698 17660 11704 17672
rect 10183 17632 11704 17660
rect 10183 17629 10195 17632
rect 10137 17623 10195 17629
rect 8941 17595 8999 17601
rect 8941 17592 8953 17595
rect 7576 17564 8953 17592
rect 8941 17561 8953 17564
rect 8987 17561 8999 17595
rect 8941 17555 8999 17561
rect 9122 17552 9128 17604
rect 9180 17592 9186 17604
rect 9968 17592 9996 17623
rect 11698 17620 11704 17632
rect 11756 17620 11762 17672
rect 15217 17663 15275 17669
rect 15217 17629 15229 17663
rect 15263 17660 15275 17663
rect 15378 17660 15384 17672
rect 15263 17632 15384 17660
rect 15263 17629 15275 17632
rect 15217 17623 15275 17629
rect 15378 17620 15384 17632
rect 15436 17620 15442 17672
rect 15470 17620 15476 17672
rect 15528 17660 15534 17672
rect 15933 17663 15991 17669
rect 15528 17632 15573 17660
rect 15528 17620 15534 17632
rect 15933 17629 15945 17663
rect 15979 17660 15991 17663
rect 16298 17660 16304 17672
rect 15979 17632 16304 17660
rect 15979 17629 15991 17632
rect 15933 17623 15991 17629
rect 16298 17620 16304 17632
rect 16356 17660 16362 17672
rect 16942 17660 16948 17672
rect 16356 17632 16948 17660
rect 16356 17620 16362 17632
rect 16942 17620 16948 17632
rect 17000 17620 17006 17672
rect 17770 17620 17776 17672
rect 17828 17660 17834 17672
rect 19429 17663 19487 17669
rect 19429 17660 19441 17663
rect 17828 17632 19441 17660
rect 17828 17620 17834 17632
rect 19429 17629 19441 17632
rect 19475 17660 19487 17663
rect 21266 17660 21272 17672
rect 19475 17632 21272 17660
rect 19475 17629 19487 17632
rect 19429 17623 19487 17629
rect 21266 17620 21272 17632
rect 21324 17620 21330 17672
rect 21637 17663 21695 17669
rect 21637 17629 21649 17663
rect 21683 17629 21695 17663
rect 21637 17623 21695 17629
rect 11333 17595 11391 17601
rect 11333 17592 11345 17595
rect 9180 17564 9273 17592
rect 9968 17564 11345 17592
rect 9180 17552 9186 17564
rect 11333 17561 11345 17564
rect 11379 17561 11391 17595
rect 11333 17555 11391 17561
rect 11517 17595 11575 17601
rect 11517 17561 11529 17595
rect 11563 17592 11575 17595
rect 11606 17592 11612 17604
rect 11563 17564 11612 17592
rect 11563 17561 11575 17564
rect 11517 17555 11575 17561
rect 11606 17552 11612 17564
rect 11664 17592 11670 17604
rect 11664 17564 11928 17592
rect 11664 17552 11670 17564
rect 7006 17524 7012 17536
rect 5368 17496 7012 17524
rect 7006 17484 7012 17496
rect 7064 17484 7070 17536
rect 9140 17524 9168 17552
rect 11238 17524 11244 17536
rect 9140 17496 11244 17524
rect 11238 17484 11244 17496
rect 11296 17484 11302 17536
rect 11701 17527 11759 17533
rect 11701 17493 11713 17527
rect 11747 17524 11759 17527
rect 11790 17524 11796 17536
rect 11747 17496 11796 17524
rect 11747 17493 11759 17496
rect 11701 17487 11759 17493
rect 11790 17484 11796 17496
rect 11848 17484 11854 17536
rect 11900 17524 11928 17564
rect 12250 17552 12256 17604
rect 12308 17592 12314 17604
rect 12406 17595 12464 17601
rect 12406 17592 12418 17595
rect 12308 17564 12418 17592
rect 12308 17552 12314 17564
rect 12406 17561 12418 17564
rect 12452 17561 12464 17595
rect 12406 17555 12464 17561
rect 14918 17552 14924 17604
rect 14976 17592 14982 17604
rect 18601 17595 18659 17601
rect 18601 17592 18613 17595
rect 14976 17564 18613 17592
rect 14976 17552 14982 17564
rect 18601 17561 18613 17564
rect 18647 17561 18659 17595
rect 18601 17555 18659 17561
rect 13541 17527 13599 17533
rect 13541 17524 13553 17527
rect 11900 17496 13553 17524
rect 13541 17493 13553 17496
rect 13587 17524 13599 17527
rect 16574 17524 16580 17536
rect 13587 17496 16580 17524
rect 13587 17493 13599 17496
rect 13541 17487 13599 17493
rect 16574 17484 16580 17496
rect 16632 17484 16638 17536
rect 17218 17524 17224 17536
rect 17179 17496 17224 17524
rect 17218 17484 17224 17496
rect 17276 17484 17282 17536
rect 18616 17524 18644 17555
rect 19150 17552 19156 17604
rect 19208 17592 19214 17604
rect 19245 17595 19303 17601
rect 19245 17592 19257 17595
rect 19208 17564 19257 17592
rect 19208 17552 19214 17564
rect 19245 17561 19257 17564
rect 19291 17561 19303 17595
rect 21652 17592 21680 17623
rect 21726 17620 21732 17672
rect 21784 17660 21790 17672
rect 24397 17663 24455 17669
rect 21784 17632 22508 17660
rect 21784 17620 21790 17632
rect 22370 17592 22376 17604
rect 21652 17564 22376 17592
rect 19245 17555 19303 17561
rect 22370 17552 22376 17564
rect 22428 17552 22434 17604
rect 20349 17527 20407 17533
rect 20349 17524 20361 17527
rect 18616 17496 20361 17524
rect 20349 17493 20361 17496
rect 20395 17524 20407 17527
rect 21726 17524 21732 17536
rect 20395 17496 21732 17524
rect 20395 17493 20407 17496
rect 20349 17487 20407 17493
rect 21726 17484 21732 17496
rect 21784 17484 21790 17536
rect 22281 17527 22339 17533
rect 22281 17493 22293 17527
rect 22327 17524 22339 17527
rect 22480 17524 22508 17632
rect 24397 17629 24409 17663
rect 24443 17660 24455 17663
rect 24854 17660 24860 17672
rect 24443 17632 24860 17660
rect 24443 17629 24455 17632
rect 24397 17623 24455 17629
rect 24854 17620 24860 17632
rect 24912 17660 24918 17672
rect 25314 17660 25320 17672
rect 24912 17632 25320 17660
rect 24912 17620 24918 17632
rect 25314 17620 25320 17632
rect 25372 17620 25378 17672
rect 25498 17620 25504 17672
rect 25556 17669 25562 17672
rect 25792 17669 25820 17700
rect 25884 17700 26332 17728
rect 25884 17669 25912 17700
rect 26326 17688 26332 17700
rect 26384 17688 26390 17740
rect 26620 17737 26648 17768
rect 31389 17765 31401 17799
rect 31435 17796 31447 17799
rect 32968 17796 32996 17836
rect 33226 17796 33232 17808
rect 31435 17768 32996 17796
rect 33060 17768 33232 17796
rect 31435 17765 31447 17768
rect 31389 17759 31447 17765
rect 26605 17731 26663 17737
rect 26605 17697 26617 17731
rect 26651 17697 26663 17731
rect 26605 17691 26663 17697
rect 25556 17660 25565 17669
rect 25685 17663 25743 17669
rect 25556 17632 25601 17660
rect 25556 17623 25565 17632
rect 25685 17629 25697 17663
rect 25731 17629 25743 17663
rect 25685 17623 25743 17629
rect 25777 17663 25835 17669
rect 25777 17629 25789 17663
rect 25823 17629 25835 17663
rect 25777 17623 25835 17629
rect 25869 17663 25927 17669
rect 25869 17629 25881 17663
rect 25915 17629 25927 17663
rect 26620 17660 26648 17691
rect 32214 17688 32220 17740
rect 32272 17728 32278 17740
rect 32272 17700 32950 17728
rect 32272 17688 32278 17700
rect 28442 17660 28448 17672
rect 26620 17632 28448 17660
rect 25869 17623 25927 17629
rect 25556 17620 25562 17623
rect 24578 17592 24584 17604
rect 24539 17564 24584 17592
rect 24578 17552 24584 17564
rect 24636 17552 24642 17604
rect 25700 17592 25728 17623
rect 28442 17620 28448 17632
rect 28500 17620 28506 17672
rect 31110 17620 31116 17672
rect 31168 17660 31174 17672
rect 31297 17663 31355 17669
rect 31297 17660 31309 17663
rect 31168 17632 31309 17660
rect 31168 17620 31174 17632
rect 31297 17629 31309 17632
rect 31343 17629 31355 17663
rect 31478 17660 31484 17672
rect 31439 17632 31484 17660
rect 31297 17623 31355 17629
rect 31478 17620 31484 17632
rect 31536 17620 31542 17672
rect 32922 17669 32950 17700
rect 33060 17669 33088 17768
rect 33226 17756 33232 17768
rect 33284 17756 33290 17808
rect 33336 17728 33364 17836
rect 40034 17728 40040 17740
rect 33244 17700 33364 17728
rect 36740 17700 40040 17728
rect 32922 17663 32991 17669
rect 32922 17632 32945 17663
rect 32933 17629 32945 17632
rect 32979 17629 32991 17663
rect 32933 17623 32991 17629
rect 33045 17663 33103 17669
rect 33045 17629 33057 17663
rect 33091 17629 33103 17663
rect 33045 17623 33103 17629
rect 33158 17660 33216 17666
rect 33158 17626 33170 17660
rect 33204 17657 33216 17660
rect 33244 17657 33272 17700
rect 33204 17629 33272 17657
rect 33321 17663 33379 17669
rect 33321 17629 33333 17663
rect 33367 17660 33379 17663
rect 33410 17660 33416 17672
rect 33367 17632 33416 17660
rect 33367 17629 33379 17632
rect 33204 17626 33216 17629
rect 33158 17620 33216 17626
rect 33321 17623 33379 17629
rect 33410 17620 33416 17632
rect 33468 17620 33474 17672
rect 26050 17592 26056 17604
rect 25700 17564 26056 17592
rect 26050 17552 26056 17564
rect 26108 17552 26114 17604
rect 26145 17595 26203 17601
rect 26145 17561 26157 17595
rect 26191 17592 26203 17595
rect 26850 17595 26908 17601
rect 26850 17592 26862 17595
rect 26191 17564 26862 17592
rect 26191 17561 26203 17564
rect 26145 17555 26203 17561
rect 26850 17561 26862 17564
rect 26896 17561 26908 17595
rect 36740 17592 36768 17700
rect 40034 17688 40040 17700
rect 40092 17688 40098 17740
rect 36817 17663 36875 17669
rect 36817 17629 36829 17663
rect 36863 17660 36875 17663
rect 36863 17632 37688 17660
rect 36863 17629 36875 17632
rect 36817 17623 36875 17629
rect 37660 17604 37688 17632
rect 37734 17620 37740 17672
rect 37792 17660 37798 17672
rect 38473 17663 38531 17669
rect 38473 17660 38485 17663
rect 37792 17632 38485 17660
rect 37792 17620 37798 17632
rect 38473 17629 38485 17632
rect 38519 17629 38531 17663
rect 68094 17660 68100 17672
rect 68055 17632 68100 17660
rect 38473 17623 38531 17629
rect 68094 17620 68100 17632
rect 68152 17620 68158 17672
rect 37001 17595 37059 17601
rect 37001 17592 37013 17595
rect 26850 17555 26908 17561
rect 34624 17564 37013 17592
rect 26234 17524 26240 17536
rect 22327 17496 26240 17524
rect 22327 17493 22339 17496
rect 22281 17487 22339 17493
rect 26234 17484 26240 17496
rect 26292 17484 26298 17536
rect 32214 17524 32220 17536
rect 32175 17496 32220 17524
rect 32214 17484 32220 17496
rect 32272 17484 32278 17536
rect 32858 17484 32864 17536
rect 32916 17524 32922 17536
rect 34624 17524 34652 17564
rect 37001 17561 37013 17564
rect 37047 17561 37059 17595
rect 37642 17592 37648 17604
rect 37603 17564 37648 17592
rect 37001 17555 37059 17561
rect 37642 17552 37648 17564
rect 37700 17552 37706 17604
rect 37826 17592 37832 17604
rect 37787 17564 37832 17592
rect 37826 17552 37832 17564
rect 37884 17552 37890 17604
rect 32916 17496 34652 17524
rect 34793 17527 34851 17533
rect 32916 17484 32922 17496
rect 34793 17493 34805 17527
rect 34839 17524 34851 17527
rect 35434 17524 35440 17536
rect 34839 17496 35440 17524
rect 34839 17493 34851 17496
rect 34793 17487 34851 17493
rect 35434 17484 35440 17496
rect 35492 17524 35498 17536
rect 35618 17524 35624 17536
rect 35492 17496 35624 17524
rect 35492 17484 35498 17496
rect 35618 17484 35624 17496
rect 35676 17484 35682 17536
rect 35710 17484 35716 17536
rect 35768 17524 35774 17536
rect 36262 17524 36268 17536
rect 35768 17496 36268 17524
rect 35768 17484 35774 17496
rect 36262 17484 36268 17496
rect 36320 17484 36326 17536
rect 37182 17524 37188 17536
rect 37143 17496 37188 17524
rect 37182 17484 37188 17496
rect 37240 17484 37246 17536
rect 37458 17484 37464 17536
rect 37516 17524 37522 17536
rect 38013 17527 38071 17533
rect 38013 17524 38025 17527
rect 37516 17496 38025 17524
rect 37516 17484 37522 17496
rect 38013 17493 38025 17496
rect 38059 17493 38071 17527
rect 38013 17487 38071 17493
rect 1104 17434 68816 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 50294 17434
rect 50346 17382 50358 17434
rect 50410 17382 50422 17434
rect 50474 17382 50486 17434
rect 50538 17382 50550 17434
rect 50602 17382 68816 17434
rect 1104 17360 68816 17382
rect 1394 17320 1400 17332
rect 1355 17292 1400 17320
rect 1394 17280 1400 17292
rect 1452 17280 1458 17332
rect 1581 17323 1639 17329
rect 1581 17289 1593 17323
rect 1627 17320 1639 17323
rect 2866 17320 2872 17332
rect 1627 17292 2872 17320
rect 1627 17289 1639 17292
rect 1581 17283 1639 17289
rect 2866 17280 2872 17292
rect 2924 17280 2930 17332
rect 5813 17323 5871 17329
rect 5813 17289 5825 17323
rect 5859 17320 5871 17323
rect 6914 17320 6920 17332
rect 5859 17292 6920 17320
rect 5859 17289 5871 17292
rect 5813 17283 5871 17289
rect 6914 17280 6920 17292
rect 6972 17280 6978 17332
rect 12250 17320 12256 17332
rect 7116 17292 9812 17320
rect 12211 17292 12256 17320
rect 3234 17252 3240 17264
rect 2884 17224 3240 17252
rect 1578 17187 1636 17193
rect 1578 17153 1590 17187
rect 1624 17184 1636 17187
rect 2314 17184 2320 17196
rect 1624 17156 2320 17184
rect 1624 17153 1636 17156
rect 1578 17147 1636 17153
rect 2314 17144 2320 17156
rect 2372 17144 2378 17196
rect 2590 17144 2596 17196
rect 2648 17184 2654 17196
rect 2884 17193 2912 17224
rect 3234 17212 3240 17224
rect 3292 17212 3298 17264
rect 4614 17252 4620 17264
rect 3620 17224 4620 17252
rect 2731 17187 2789 17193
rect 2731 17184 2743 17187
rect 2648 17156 2743 17184
rect 2648 17144 2654 17156
rect 2731 17153 2743 17156
rect 2777 17153 2789 17187
rect 2731 17147 2789 17153
rect 2869 17187 2927 17193
rect 2869 17153 2881 17187
rect 2915 17153 2927 17187
rect 2869 17147 2927 17153
rect 2958 17144 2964 17196
rect 3016 17184 3022 17196
rect 3016 17156 3061 17184
rect 3016 17144 3022 17156
rect 3142 17144 3148 17196
rect 3200 17184 3206 17196
rect 3620 17193 3648 17224
rect 4614 17212 4620 17224
rect 4672 17212 4678 17264
rect 5258 17212 5264 17264
rect 5316 17252 5322 17264
rect 5629 17255 5687 17261
rect 5629 17252 5641 17255
rect 5316 17224 5641 17252
rect 5316 17212 5322 17224
rect 5629 17221 5641 17224
rect 5675 17252 5687 17255
rect 7116 17252 7144 17292
rect 8754 17252 8760 17264
rect 5675 17224 7144 17252
rect 7392 17224 8760 17252
rect 5675 17221 5687 17224
rect 5629 17215 5687 17221
rect 3605 17187 3663 17193
rect 3200 17156 3245 17184
rect 3200 17144 3206 17156
rect 3605 17153 3617 17187
rect 3651 17153 3663 17187
rect 3861 17187 3919 17193
rect 3861 17184 3873 17187
rect 3605 17147 3663 17153
rect 3712 17156 3873 17184
rect 2041 17119 2099 17125
rect 2041 17085 2053 17119
rect 2087 17116 2099 17119
rect 2406 17116 2412 17128
rect 2087 17088 2412 17116
rect 2087 17085 2099 17088
rect 2041 17079 2099 17085
rect 2406 17076 2412 17088
rect 2464 17076 2470 17128
rect 2501 17119 2559 17125
rect 2501 17085 2513 17119
rect 2547 17116 2559 17119
rect 3712 17116 3740 17156
rect 3861 17153 3873 17156
rect 3907 17153 3919 17187
rect 3861 17147 3919 17153
rect 4706 17144 4712 17196
rect 4764 17184 4770 17196
rect 7392 17193 7420 17224
rect 5445 17187 5503 17193
rect 5445 17184 5457 17187
rect 4764 17156 5457 17184
rect 4764 17144 4770 17156
rect 5445 17153 5457 17156
rect 5491 17153 5503 17187
rect 5445 17147 5503 17153
rect 7377 17187 7435 17193
rect 7377 17153 7389 17187
rect 7423 17153 7435 17187
rect 8113 17187 8171 17193
rect 8113 17184 8125 17187
rect 7377 17147 7435 17153
rect 7760 17156 8125 17184
rect 2547 17088 2774 17116
rect 2547 17085 2559 17088
rect 2501 17079 2559 17085
rect 1946 16980 1952 16992
rect 1907 16952 1952 16980
rect 1946 16940 1952 16952
rect 2004 16940 2010 16992
rect 2746 16980 2774 17088
rect 2976 17088 3740 17116
rect 2976 16980 3004 17088
rect 7466 17076 7472 17128
rect 7524 17116 7530 17128
rect 7653 17119 7711 17125
rect 7653 17116 7665 17119
rect 7524 17088 7665 17116
rect 7524 17076 7530 17088
rect 7653 17085 7665 17088
rect 7699 17085 7711 17119
rect 7653 17079 7711 17085
rect 7098 17048 7104 17060
rect 4908 17020 7104 17048
rect 2746 16952 3004 16980
rect 3142 16940 3148 16992
rect 3200 16980 3206 16992
rect 4908 16980 4936 17020
rect 7098 17008 7104 17020
rect 7156 17048 7162 17060
rect 7760 17048 7788 17156
rect 8113 17153 8125 17156
rect 8159 17153 8171 17187
rect 8113 17147 8171 17153
rect 8202 17144 8208 17196
rect 8260 17184 8266 17196
rect 8404 17193 8432 17224
rect 8754 17212 8760 17224
rect 8812 17212 8818 17264
rect 8297 17187 8355 17193
rect 8297 17184 8309 17187
rect 8260 17156 8309 17184
rect 8260 17144 8266 17156
rect 8297 17153 8309 17156
rect 8343 17153 8355 17187
rect 8297 17147 8355 17153
rect 8389 17187 8447 17193
rect 8389 17153 8401 17187
rect 8435 17153 8447 17187
rect 8389 17147 8447 17153
rect 8478 17144 8484 17196
rect 8536 17184 8542 17196
rect 9217 17187 9275 17193
rect 9217 17184 9229 17187
rect 8536 17156 9229 17184
rect 8536 17144 8542 17156
rect 9217 17153 9229 17156
rect 9263 17184 9275 17187
rect 9582 17184 9588 17196
rect 9263 17156 9588 17184
rect 9263 17153 9275 17156
rect 9217 17147 9275 17153
rect 9582 17144 9588 17156
rect 9640 17144 9646 17196
rect 9784 17048 9812 17292
rect 12250 17280 12256 17292
rect 12308 17280 12314 17332
rect 16114 17320 16120 17332
rect 15488 17292 16120 17320
rect 9950 17212 9956 17264
rect 10008 17252 10014 17264
rect 10686 17252 10692 17264
rect 10008 17224 10692 17252
rect 10008 17212 10014 17224
rect 10686 17212 10692 17224
rect 10744 17212 10750 17264
rect 11054 17212 11060 17264
rect 11112 17252 11118 17264
rect 11112 17224 11928 17252
rect 11112 17212 11118 17224
rect 10873 17187 10931 17193
rect 10873 17153 10885 17187
rect 10919 17184 10931 17187
rect 11514 17184 11520 17196
rect 10919 17156 11520 17184
rect 10919 17153 10931 17156
rect 10873 17147 10931 17153
rect 11514 17144 11520 17156
rect 11572 17144 11578 17196
rect 11609 17187 11667 17193
rect 11609 17153 11621 17187
rect 11655 17153 11667 17187
rect 11790 17184 11796 17196
rect 11751 17156 11796 17184
rect 11609 17147 11667 17153
rect 11422 17076 11428 17128
rect 11480 17116 11486 17128
rect 11624 17116 11652 17147
rect 11790 17144 11796 17156
rect 11848 17144 11854 17196
rect 11900 17193 11928 17224
rect 11885 17187 11943 17193
rect 11885 17153 11897 17187
rect 11931 17153 11943 17187
rect 11885 17147 11943 17153
rect 11974 17144 11980 17196
rect 12032 17184 12038 17196
rect 15488 17193 15516 17292
rect 16114 17280 16120 17292
rect 16172 17280 16178 17332
rect 16206 17280 16212 17332
rect 16264 17280 16270 17332
rect 18690 17280 18696 17332
rect 18748 17320 18754 17332
rect 21913 17323 21971 17329
rect 21913 17320 21925 17323
rect 18748 17292 21925 17320
rect 18748 17280 18754 17292
rect 21913 17289 21925 17292
rect 21959 17289 21971 17323
rect 23842 17320 23848 17332
rect 21913 17283 21971 17289
rect 22066 17292 23848 17320
rect 16224 17252 16252 17280
rect 15764 17224 16252 17252
rect 12713 17187 12771 17193
rect 12713 17184 12725 17187
rect 12032 17156 12725 17184
rect 12032 17144 12038 17156
rect 12713 17153 12725 17156
rect 12759 17153 12771 17187
rect 12713 17147 12771 17153
rect 15473 17187 15531 17193
rect 15473 17153 15485 17187
rect 15519 17153 15531 17187
rect 15654 17184 15660 17196
rect 15615 17156 15660 17184
rect 15473 17147 15531 17153
rect 15654 17144 15660 17156
rect 15712 17144 15718 17196
rect 15764 17193 15792 17224
rect 16390 17212 16396 17264
rect 16448 17252 16454 17264
rect 19978 17252 19984 17264
rect 16448 17224 19984 17252
rect 16448 17212 16454 17224
rect 15749 17187 15807 17193
rect 15749 17153 15761 17187
rect 15795 17153 15807 17187
rect 15749 17147 15807 17153
rect 15887 17187 15945 17193
rect 15887 17153 15899 17187
rect 15933 17184 15945 17187
rect 16206 17184 16212 17196
rect 15933 17156 16212 17184
rect 15933 17153 15945 17156
rect 15887 17147 15945 17153
rect 16206 17144 16212 17156
rect 16264 17144 16270 17196
rect 16592 17184 16620 17224
rect 19978 17212 19984 17224
rect 20036 17212 20042 17264
rect 20898 17212 20904 17264
rect 20956 17252 20962 17264
rect 22066 17252 22094 17292
rect 23842 17280 23848 17292
rect 23900 17280 23906 17332
rect 25222 17280 25228 17332
rect 25280 17280 25286 17332
rect 25314 17280 25320 17332
rect 25372 17280 25378 17332
rect 25498 17280 25504 17332
rect 25556 17280 25562 17332
rect 28534 17320 28540 17332
rect 28460 17292 28540 17320
rect 20956 17224 22094 17252
rect 23692 17255 23750 17261
rect 20956 17212 20962 17224
rect 23692 17221 23704 17255
rect 23738 17252 23750 17255
rect 24857 17255 24915 17261
rect 24857 17252 24869 17255
rect 23738 17224 24869 17252
rect 23738 17221 23750 17224
rect 23692 17215 23750 17221
rect 24857 17221 24869 17224
rect 24903 17221 24915 17255
rect 24857 17215 24915 17221
rect 16658 17187 16716 17193
rect 16658 17184 16670 17187
rect 16592 17156 16670 17184
rect 16658 17153 16670 17156
rect 16704 17153 16716 17187
rect 16925 17187 16983 17193
rect 16925 17184 16937 17187
rect 16658 17147 16716 17153
rect 16776 17156 16937 17184
rect 12066 17116 12072 17128
rect 11480 17088 12072 17116
rect 11480 17076 11486 17088
rect 12066 17076 12072 17088
rect 12124 17076 12130 17128
rect 16117 17119 16175 17125
rect 16117 17085 16129 17119
rect 16163 17116 16175 17119
rect 16776 17116 16804 17156
rect 16925 17153 16937 17156
rect 16971 17153 16983 17187
rect 19242 17184 19248 17196
rect 19203 17156 19248 17184
rect 16925 17147 16983 17153
rect 19242 17144 19248 17156
rect 19300 17144 19306 17196
rect 19426 17184 19432 17196
rect 19387 17156 19432 17184
rect 19426 17144 19432 17156
rect 19484 17144 19490 17196
rect 19521 17187 19579 17193
rect 19521 17153 19533 17187
rect 19567 17153 19579 17187
rect 19521 17147 19579 17153
rect 19613 17187 19671 17193
rect 19613 17153 19625 17187
rect 19659 17153 19671 17187
rect 19613 17147 19671 17153
rect 16163 17088 16804 17116
rect 16163 17085 16175 17088
rect 16117 17079 16175 17085
rect 19058 17076 19064 17128
rect 19116 17116 19122 17128
rect 19536 17116 19564 17147
rect 19116 17088 19564 17116
rect 19628 17116 19656 17147
rect 19702 17144 19708 17196
rect 19760 17184 19766 17196
rect 20254 17184 20260 17196
rect 19760 17156 20260 17184
rect 19760 17144 19766 17156
rect 20254 17144 20260 17156
rect 20312 17144 20318 17196
rect 21266 17184 21272 17196
rect 21227 17156 21272 17184
rect 21266 17144 21272 17156
rect 21324 17144 21330 17196
rect 22097 17187 22155 17193
rect 22097 17153 22109 17187
rect 22143 17184 22155 17187
rect 22830 17184 22836 17196
rect 22143 17156 22836 17184
rect 22143 17153 22155 17156
rect 22097 17147 22155 17153
rect 22830 17144 22836 17156
rect 22888 17144 22894 17196
rect 23934 17184 23940 17196
rect 23895 17156 23940 17184
rect 23934 17144 23940 17156
rect 23992 17144 23998 17196
rect 25240 17193 25268 17280
rect 25329 17199 25357 17280
rect 25516 17252 25544 17280
rect 25516 17224 25636 17252
rect 25317 17193 25375 17199
rect 25113 17187 25171 17193
rect 25113 17153 25125 17187
rect 25159 17184 25171 17187
rect 25225 17187 25283 17193
rect 25159 17153 25176 17184
rect 25113 17147 25176 17153
rect 25225 17153 25237 17187
rect 25271 17153 25283 17187
rect 25317 17159 25329 17193
rect 25363 17159 25375 17193
rect 25317 17153 25375 17159
rect 25501 17187 25559 17193
rect 25501 17153 25513 17187
rect 25547 17184 25559 17187
rect 25608 17184 25636 17224
rect 28350 17184 28356 17196
rect 25547 17156 25636 17184
rect 28311 17156 28356 17184
rect 25547 17153 25559 17156
rect 25225 17147 25283 17153
rect 25501 17147 25559 17153
rect 22186 17116 22192 17128
rect 19628 17088 22192 17116
rect 19116 17076 19122 17088
rect 13630 17048 13636 17060
rect 7156 17020 9628 17048
rect 9784 17020 13636 17048
rect 7156 17008 7162 17020
rect 3200 16952 4936 16980
rect 3200 16940 3206 16952
rect 4982 16940 4988 16992
rect 5040 16980 5046 16992
rect 8754 16980 8760 16992
rect 5040 16952 5085 16980
rect 8715 16952 8760 16980
rect 5040 16940 5046 16952
rect 8754 16940 8760 16952
rect 8812 16940 8818 16992
rect 9600 16980 9628 17020
rect 13630 17008 13636 17020
rect 13688 17008 13694 17060
rect 18782 17048 18788 17060
rect 18695 17020 18788 17048
rect 18782 17008 18788 17020
rect 18840 17048 18846 17060
rect 19628 17048 19656 17088
rect 22186 17076 22192 17088
rect 22244 17076 22250 17128
rect 25148 17116 25176 17147
rect 28350 17144 28356 17156
rect 28408 17144 28414 17196
rect 28460 17184 28488 17292
rect 28534 17280 28540 17292
rect 28592 17280 28598 17332
rect 28626 17280 28632 17332
rect 28684 17280 28690 17332
rect 28994 17320 29000 17332
rect 28955 17292 29000 17320
rect 28994 17280 29000 17292
rect 29052 17280 29058 17332
rect 37734 17320 37740 17332
rect 29104 17292 37740 17320
rect 28644 17193 28672 17280
rect 28902 17212 28908 17264
rect 28960 17252 28966 17264
rect 29104 17252 29132 17292
rect 37734 17280 37740 17292
rect 37792 17280 37798 17332
rect 37826 17280 37832 17332
rect 37884 17320 37890 17332
rect 40405 17323 40463 17329
rect 40405 17320 40417 17323
rect 37884 17292 40417 17320
rect 37884 17280 37890 17292
rect 40405 17289 40417 17292
rect 40451 17289 40463 17323
rect 40405 17283 40463 17289
rect 35710 17252 35716 17264
rect 28960 17224 29132 17252
rect 29196 17224 35716 17252
rect 28960 17212 28966 17224
rect 28516 17187 28574 17193
rect 28516 17184 28528 17187
rect 28460 17156 28528 17184
rect 28516 17153 28528 17156
rect 28562 17153 28574 17187
rect 28516 17147 28574 17153
rect 28629 17187 28687 17193
rect 28629 17153 28641 17187
rect 28675 17153 28687 17187
rect 28629 17147 28687 17153
rect 28721 17187 28779 17193
rect 28721 17153 28733 17187
rect 28767 17184 28779 17187
rect 29196 17184 29224 17224
rect 35710 17212 35716 17224
rect 35768 17212 35774 17264
rect 37921 17255 37979 17261
rect 37921 17221 37933 17255
rect 37967 17252 37979 17255
rect 39270 17255 39328 17261
rect 39270 17252 39282 17255
rect 37967 17224 39282 17252
rect 37967 17221 37979 17224
rect 37921 17215 37979 17221
rect 39270 17221 39282 17224
rect 39316 17221 39328 17255
rect 39270 17215 39328 17221
rect 28767 17156 28801 17184
rect 28966 17156 29224 17184
rect 28767 17153 28779 17156
rect 28721 17147 28779 17153
rect 26510 17116 26516 17128
rect 25148 17088 26516 17116
rect 26510 17076 26516 17088
rect 26568 17116 26574 17128
rect 27893 17119 27951 17125
rect 27893 17116 27905 17119
rect 26568 17088 27905 17116
rect 26568 17076 26574 17088
rect 27893 17085 27905 17088
rect 27939 17116 27951 17119
rect 28736 17116 28764 17147
rect 28966 17116 28994 17156
rect 29914 17144 29920 17196
rect 29972 17184 29978 17196
rect 30449 17187 30507 17193
rect 30449 17184 30461 17187
rect 29972 17156 30461 17184
rect 29972 17144 29978 17156
rect 30449 17153 30461 17156
rect 30495 17153 30507 17187
rect 33226 17184 33232 17196
rect 33187 17156 33232 17184
rect 30449 17147 30507 17153
rect 33226 17144 33232 17156
rect 33284 17144 33290 17196
rect 35342 17144 35348 17196
rect 35400 17184 35406 17196
rect 35814 17187 35872 17193
rect 35814 17184 35826 17187
rect 35400 17156 35826 17184
rect 35400 17144 35406 17156
rect 35814 17153 35826 17156
rect 35860 17153 35872 17187
rect 36078 17184 36084 17196
rect 36039 17156 36084 17184
rect 35814 17147 35872 17153
rect 36078 17144 36084 17156
rect 36136 17144 36142 17196
rect 37274 17184 37280 17196
rect 37235 17156 37280 17184
rect 37274 17144 37280 17156
rect 37332 17144 37338 17196
rect 37458 17184 37464 17196
rect 37419 17156 37464 17184
rect 37458 17144 37464 17156
rect 37516 17144 37522 17196
rect 37550 17144 37556 17196
rect 37608 17184 37614 17196
rect 37691 17187 37749 17193
rect 37608 17156 37653 17184
rect 37608 17144 37614 17156
rect 37691 17153 37703 17187
rect 37737 17184 37749 17187
rect 37737 17156 37872 17184
rect 37737 17153 37749 17156
rect 37691 17147 37749 17153
rect 27939 17088 28994 17116
rect 30193 17119 30251 17125
rect 27939 17085 27951 17088
rect 27893 17079 27951 17085
rect 30193 17085 30205 17119
rect 30239 17085 30251 17119
rect 30193 17079 30251 17085
rect 18840 17020 19656 17048
rect 18840 17008 18846 17020
rect 20898 17008 20904 17060
rect 20956 17048 20962 17060
rect 21085 17051 21143 17057
rect 21085 17048 21097 17051
rect 20956 17020 21097 17048
rect 20956 17008 20962 17020
rect 21085 17017 21097 17020
rect 21131 17017 21143 17051
rect 21085 17011 21143 17017
rect 11422 16980 11428 16992
rect 9600 16952 11428 16980
rect 11422 16940 11428 16952
rect 11480 16940 11486 16992
rect 17954 16940 17960 16992
rect 18012 16980 18018 16992
rect 18049 16983 18107 16989
rect 18049 16980 18061 16983
rect 18012 16952 18061 16980
rect 18012 16940 18018 16952
rect 18049 16949 18061 16952
rect 18095 16949 18107 16983
rect 18049 16943 18107 16949
rect 19889 16983 19947 16989
rect 19889 16949 19901 16983
rect 19935 16980 19947 16983
rect 20254 16980 20260 16992
rect 19935 16952 20260 16980
rect 19935 16949 19947 16952
rect 19889 16943 19947 16949
rect 20254 16940 20260 16952
rect 20312 16940 20318 16992
rect 20438 16980 20444 16992
rect 20399 16952 20444 16980
rect 20438 16940 20444 16952
rect 20496 16940 20502 16992
rect 22094 16940 22100 16992
rect 22152 16980 22158 16992
rect 22557 16983 22615 16989
rect 22557 16980 22569 16983
rect 22152 16952 22569 16980
rect 22152 16940 22158 16952
rect 22557 16949 22569 16952
rect 22603 16980 22615 16983
rect 25038 16980 25044 16992
rect 22603 16952 25044 16980
rect 22603 16949 22615 16952
rect 22557 16943 22615 16949
rect 25038 16940 25044 16952
rect 25096 16940 25102 16992
rect 26326 16980 26332 16992
rect 26239 16952 26332 16980
rect 26326 16940 26332 16952
rect 26384 16980 26390 16992
rect 27982 16980 27988 16992
rect 26384 16952 27988 16980
rect 26384 16940 26390 16952
rect 27982 16940 27988 16952
rect 28040 16940 28046 16992
rect 28442 16940 28448 16992
rect 28500 16980 28506 16992
rect 30208 16980 30236 17079
rect 31478 17076 31484 17128
rect 31536 17116 31542 17128
rect 32953 17119 33011 17125
rect 32953 17116 32965 17119
rect 31536 17088 32965 17116
rect 31536 17076 31542 17088
rect 32953 17085 32965 17088
rect 32999 17085 33011 17119
rect 32953 17079 33011 17085
rect 28500 16952 30236 16980
rect 28500 16940 28506 16952
rect 31202 16940 31208 16992
rect 31260 16980 31266 16992
rect 31573 16983 31631 16989
rect 31573 16980 31585 16983
rect 31260 16952 31585 16980
rect 31260 16940 31266 16952
rect 31573 16949 31585 16952
rect 31619 16949 31631 16983
rect 31573 16943 31631 16949
rect 34514 16940 34520 16992
rect 34572 16980 34578 16992
rect 34701 16983 34759 16989
rect 34701 16980 34713 16983
rect 34572 16952 34713 16980
rect 34572 16940 34578 16952
rect 34701 16949 34713 16952
rect 34747 16949 34759 16983
rect 34701 16943 34759 16949
rect 36078 16940 36084 16992
rect 36136 16980 36142 16992
rect 36725 16983 36783 16989
rect 36725 16980 36737 16983
rect 36136 16952 36737 16980
rect 36136 16940 36142 16952
rect 36725 16949 36737 16952
rect 36771 16980 36783 16983
rect 37844 16980 37872 17156
rect 38838 17144 38844 17196
rect 38896 17184 38902 17196
rect 39025 17187 39083 17193
rect 39025 17184 39037 17187
rect 38896 17156 39037 17184
rect 38896 17144 38902 17156
rect 39025 17153 39037 17156
rect 39071 17153 39083 17187
rect 39025 17147 39083 17153
rect 36771 16952 37872 16980
rect 36771 16949 36783 16952
rect 36725 16943 36783 16949
rect 1104 16890 68816 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 65654 16890
rect 65706 16838 65718 16890
rect 65770 16838 65782 16890
rect 65834 16838 65846 16890
rect 65898 16838 65910 16890
rect 65962 16838 68816 16890
rect 1104 16816 68816 16838
rect 1946 16736 1952 16788
rect 2004 16776 2010 16788
rect 2041 16779 2099 16785
rect 2041 16776 2053 16779
rect 2004 16748 2053 16776
rect 2004 16736 2010 16748
rect 2041 16745 2053 16748
rect 2087 16745 2099 16779
rect 2041 16739 2099 16745
rect 2501 16779 2559 16785
rect 2501 16745 2513 16779
rect 2547 16776 2559 16779
rect 2866 16776 2872 16788
rect 2547 16748 2872 16776
rect 2547 16745 2559 16748
rect 2501 16739 2559 16745
rect 2866 16736 2872 16748
rect 2924 16736 2930 16788
rect 2958 16736 2964 16788
rect 3016 16776 3022 16788
rect 4341 16779 4399 16785
rect 4341 16776 4353 16779
rect 3016 16748 4353 16776
rect 3016 16736 3022 16748
rect 4341 16745 4353 16748
rect 4387 16745 4399 16779
rect 4341 16739 4399 16745
rect 7561 16779 7619 16785
rect 7561 16745 7573 16779
rect 7607 16776 7619 16779
rect 8202 16776 8208 16788
rect 7607 16748 8208 16776
rect 7607 16745 7619 16748
rect 7561 16739 7619 16745
rect 8202 16736 8208 16748
rect 8260 16736 8266 16788
rect 15654 16776 15660 16788
rect 8312 16748 15516 16776
rect 15615 16748 15660 16776
rect 2590 16668 2596 16720
rect 2648 16708 2654 16720
rect 3881 16711 3939 16717
rect 3881 16708 3893 16711
rect 2648 16680 3893 16708
rect 2648 16668 2654 16680
rect 3881 16677 3893 16680
rect 3927 16708 3939 16711
rect 5074 16708 5080 16720
rect 3927 16680 5080 16708
rect 3927 16677 3939 16680
rect 3881 16671 3939 16677
rect 5074 16668 5080 16680
rect 5132 16668 5138 16720
rect 7742 16668 7748 16720
rect 7800 16708 7806 16720
rect 8113 16711 8171 16717
rect 8113 16708 8125 16711
rect 7800 16680 8125 16708
rect 7800 16668 7806 16680
rect 8113 16677 8125 16680
rect 8159 16708 8171 16711
rect 8312 16708 8340 16748
rect 8159 16680 8340 16708
rect 15488 16708 15516 16748
rect 15654 16736 15660 16748
rect 15712 16736 15718 16788
rect 19242 16736 19248 16788
rect 19300 16776 19306 16788
rect 23474 16776 23480 16788
rect 19300 16748 23480 16776
rect 19300 16736 19306 16748
rect 16206 16708 16212 16720
rect 15488 16680 16212 16708
rect 8159 16677 8171 16680
rect 8113 16671 8171 16677
rect 16206 16668 16212 16680
rect 16264 16708 16270 16720
rect 16485 16711 16543 16717
rect 16485 16708 16497 16711
rect 16264 16680 16497 16708
rect 16264 16668 16270 16680
rect 16485 16677 16497 16680
rect 16531 16708 16543 16711
rect 16850 16708 16856 16720
rect 16531 16680 16856 16708
rect 16531 16677 16543 16680
rect 16485 16671 16543 16677
rect 16850 16668 16856 16680
rect 16908 16668 16914 16720
rect 2409 16643 2467 16649
rect 2409 16609 2421 16643
rect 2455 16640 2467 16643
rect 2958 16640 2964 16652
rect 2455 16612 2964 16640
rect 2455 16609 2467 16612
rect 2409 16603 2467 16609
rect 2958 16600 2964 16612
rect 3016 16600 3022 16652
rect 3234 16600 3240 16652
rect 3292 16640 3298 16652
rect 5905 16643 5963 16649
rect 5905 16640 5917 16643
rect 3292 16612 5917 16640
rect 3292 16600 3298 16612
rect 5905 16609 5917 16612
rect 5951 16609 5963 16643
rect 5905 16603 5963 16609
rect 6012 16612 7512 16640
rect 2225 16575 2283 16581
rect 2225 16541 2237 16575
rect 2271 16572 2283 16575
rect 2314 16572 2320 16584
rect 2271 16544 2320 16572
rect 2271 16541 2283 16544
rect 2225 16535 2283 16541
rect 2314 16532 2320 16544
rect 2372 16532 2378 16584
rect 4525 16575 4583 16581
rect 4525 16541 4537 16575
rect 4571 16572 4583 16575
rect 4982 16572 4988 16584
rect 4571 16544 4988 16572
rect 4571 16541 4583 16544
rect 4525 16535 4583 16541
rect 4982 16532 4988 16544
rect 5040 16572 5046 16584
rect 5442 16572 5448 16584
rect 5040 16544 5448 16572
rect 5040 16532 5046 16544
rect 5442 16532 5448 16544
rect 5500 16532 5506 16584
rect 5629 16575 5687 16581
rect 5629 16541 5641 16575
rect 5675 16572 5687 16575
rect 6012 16572 6040 16612
rect 7484 16584 7512 16612
rect 8662 16600 8668 16652
rect 8720 16640 8726 16652
rect 8941 16643 8999 16649
rect 8941 16640 8953 16643
rect 8720 16612 8953 16640
rect 8720 16600 8726 16612
rect 8941 16609 8953 16612
rect 8987 16609 8999 16643
rect 8941 16603 8999 16609
rect 10686 16600 10692 16652
rect 10744 16640 10750 16652
rect 12158 16640 12164 16652
rect 10744 16612 11100 16640
rect 12119 16612 12164 16640
rect 10744 16600 10750 16612
rect 7466 16572 7472 16584
rect 5675 16544 6040 16572
rect 7427 16544 7472 16572
rect 5675 16541 5687 16544
rect 5629 16535 5687 16541
rect 7466 16532 7472 16544
rect 7524 16532 7530 16584
rect 7650 16572 7656 16584
rect 7611 16544 7656 16572
rect 7650 16532 7656 16544
rect 7708 16532 7714 16584
rect 8754 16532 8760 16584
rect 8812 16572 8818 16584
rect 11072 16581 11100 16612
rect 12158 16600 12164 16612
rect 12216 16600 12222 16652
rect 14918 16600 14924 16652
rect 14976 16640 14982 16652
rect 16298 16640 16304 16652
rect 14976 16612 16304 16640
rect 14976 16600 14982 16612
rect 16298 16600 16304 16612
rect 16356 16640 16362 16652
rect 16356 16612 18092 16640
rect 16356 16600 16362 16612
rect 9197 16575 9255 16581
rect 9197 16572 9209 16575
rect 8812 16544 9209 16572
rect 8812 16532 8818 16544
rect 9197 16541 9209 16544
rect 9243 16541 9255 16575
rect 9197 16535 9255 16541
rect 11057 16575 11115 16581
rect 11057 16541 11069 16575
rect 11103 16541 11115 16575
rect 11238 16572 11244 16584
rect 11199 16544 11244 16572
rect 11057 16535 11115 16541
rect 11238 16532 11244 16544
rect 11296 16532 11302 16584
rect 11333 16575 11391 16581
rect 11333 16541 11345 16575
rect 11379 16541 11391 16575
rect 11333 16535 11391 16541
rect 2501 16507 2559 16513
rect 2501 16473 2513 16507
rect 2547 16473 2559 16507
rect 4706 16504 4712 16516
rect 4667 16476 4712 16504
rect 2501 16467 2559 16473
rect 2516 16436 2544 16467
rect 4706 16464 4712 16476
rect 4764 16464 4770 16516
rect 10962 16464 10968 16516
rect 11020 16504 11026 16516
rect 11348 16504 11376 16535
rect 11422 16532 11428 16584
rect 11480 16572 11486 16584
rect 14090 16572 14096 16584
rect 11480 16544 11525 16572
rect 11624 16544 14096 16572
rect 11480 16532 11486 16544
rect 11020 16476 11376 16504
rect 11020 16464 11026 16476
rect 5350 16436 5356 16448
rect 2516 16408 5356 16436
rect 5350 16396 5356 16408
rect 5408 16396 5414 16448
rect 7006 16436 7012 16448
rect 6967 16408 7012 16436
rect 7006 16396 7012 16408
rect 7064 16396 7070 16448
rect 9490 16396 9496 16448
rect 9548 16436 9554 16448
rect 10321 16439 10379 16445
rect 10321 16436 10333 16439
rect 9548 16408 10333 16436
rect 9548 16396 9554 16408
rect 10321 16405 10333 16408
rect 10367 16436 10379 16439
rect 11624 16436 11652 16544
rect 14090 16532 14096 16544
rect 14148 16532 14154 16584
rect 17954 16572 17960 16584
rect 15856 16544 17960 16572
rect 11701 16507 11759 16513
rect 11701 16473 11713 16507
rect 11747 16504 11759 16507
rect 12406 16507 12464 16513
rect 12406 16504 12418 16507
rect 11747 16476 12418 16504
rect 11747 16473 11759 16476
rect 11701 16467 11759 16473
rect 12406 16473 12418 16476
rect 12452 16473 12464 16507
rect 12406 16467 12464 16473
rect 13078 16464 13084 16516
rect 13136 16504 13142 16516
rect 15856 16513 15884 16544
rect 17954 16532 17960 16544
rect 18012 16532 18018 16584
rect 18064 16572 18092 16612
rect 19444 16612 19656 16640
rect 19444 16572 19472 16612
rect 19628 16581 19656 16612
rect 19904 16581 19932 16748
rect 23474 16736 23480 16748
rect 23532 16736 23538 16788
rect 25225 16779 25283 16785
rect 25225 16745 25237 16779
rect 25271 16776 25283 16779
rect 25314 16776 25320 16788
rect 25271 16748 25320 16776
rect 25271 16745 25283 16748
rect 25225 16739 25283 16745
rect 25314 16736 25320 16748
rect 25372 16736 25378 16788
rect 26510 16776 26516 16788
rect 26471 16748 26516 16776
rect 26510 16736 26516 16748
rect 26568 16736 26574 16788
rect 28534 16736 28540 16788
rect 28592 16776 28598 16788
rect 28629 16779 28687 16785
rect 28629 16776 28641 16779
rect 28592 16748 28641 16776
rect 28592 16736 28598 16748
rect 28629 16745 28641 16748
rect 28675 16745 28687 16779
rect 29914 16776 29920 16788
rect 29875 16748 29920 16776
rect 28629 16739 28687 16745
rect 29914 16736 29920 16748
rect 29972 16736 29978 16788
rect 31386 16776 31392 16788
rect 30116 16748 31392 16776
rect 22186 16708 22192 16720
rect 22147 16680 22192 16708
rect 22186 16668 22192 16680
rect 22244 16668 22250 16720
rect 23566 16668 23572 16720
rect 23624 16708 23630 16720
rect 30116 16708 30144 16748
rect 31386 16736 31392 16748
rect 31444 16736 31450 16788
rect 31938 16736 31944 16788
rect 31996 16776 32002 16788
rect 32858 16776 32864 16788
rect 31996 16748 32864 16776
rect 31996 16736 32002 16748
rect 32858 16736 32864 16748
rect 32916 16736 32922 16788
rect 34698 16776 34704 16788
rect 32968 16748 34704 16776
rect 23624 16680 30144 16708
rect 23624 16668 23630 16680
rect 30190 16668 30196 16720
rect 30248 16708 30254 16720
rect 32968 16708 32996 16748
rect 34698 16736 34704 16748
rect 34756 16736 34762 16788
rect 35342 16776 35348 16788
rect 35303 16748 35348 16776
rect 35342 16736 35348 16748
rect 35400 16736 35406 16788
rect 35710 16736 35716 16788
rect 35768 16776 35774 16788
rect 35805 16779 35863 16785
rect 35805 16776 35817 16779
rect 35768 16748 35817 16776
rect 35768 16736 35774 16748
rect 35805 16745 35817 16748
rect 35851 16776 35863 16779
rect 35986 16776 35992 16788
rect 35851 16748 35992 16776
rect 35851 16745 35863 16748
rect 35805 16739 35863 16745
rect 35986 16736 35992 16748
rect 36044 16736 36050 16788
rect 36817 16779 36875 16785
rect 36817 16745 36829 16779
rect 36863 16776 36875 16779
rect 38286 16776 38292 16788
rect 36863 16748 38292 16776
rect 36863 16745 36875 16748
rect 36817 16739 36875 16745
rect 37826 16708 37832 16720
rect 30248 16680 32996 16708
rect 33060 16680 37832 16708
rect 30248 16668 30254 16680
rect 19978 16600 19984 16652
rect 20036 16640 20042 16652
rect 20349 16643 20407 16649
rect 20349 16640 20361 16643
rect 20036 16612 20361 16640
rect 20036 16600 20042 16612
rect 20349 16609 20361 16612
rect 20395 16609 20407 16643
rect 20349 16603 20407 16609
rect 23385 16643 23443 16649
rect 23385 16609 23397 16643
rect 23431 16640 23443 16643
rect 23750 16640 23756 16652
rect 23431 16612 23756 16640
rect 23431 16609 23443 16612
rect 23385 16603 23443 16609
rect 23750 16600 23756 16612
rect 23808 16600 23814 16652
rect 26973 16643 27031 16649
rect 26973 16640 26985 16643
rect 26252 16612 26985 16640
rect 18064 16544 19472 16572
rect 19521 16575 19579 16581
rect 19521 16541 19533 16575
rect 19567 16541 19579 16575
rect 19521 16535 19579 16541
rect 19613 16575 19671 16581
rect 19613 16541 19625 16575
rect 19659 16541 19671 16575
rect 19613 16535 19671 16541
rect 19705 16575 19763 16581
rect 19705 16541 19717 16575
rect 19751 16541 19763 16575
rect 19705 16535 19763 16541
rect 19889 16575 19947 16581
rect 19889 16541 19901 16575
rect 19935 16541 19947 16575
rect 19889 16535 19947 16541
rect 15841 16507 15899 16513
rect 15841 16504 15853 16507
rect 13136 16476 15853 16504
rect 13136 16464 13142 16476
rect 15841 16473 15853 16476
rect 15887 16473 15899 16507
rect 15841 16467 15899 16473
rect 15930 16464 15936 16516
rect 15988 16504 15994 16516
rect 16025 16507 16083 16513
rect 16025 16504 16037 16507
rect 15988 16476 16037 16504
rect 15988 16464 15994 16476
rect 16025 16473 16037 16476
rect 16071 16504 16083 16507
rect 18966 16504 18972 16516
rect 16071 16476 18972 16504
rect 16071 16473 16083 16476
rect 16025 16467 16083 16473
rect 18966 16464 18972 16476
rect 19024 16504 19030 16516
rect 19150 16504 19156 16516
rect 19024 16476 19156 16504
rect 19024 16464 19030 16476
rect 19150 16464 19156 16476
rect 19208 16464 19214 16516
rect 10367 16408 11652 16436
rect 10367 16405 10379 16408
rect 10321 16399 10379 16405
rect 11790 16396 11796 16448
rect 11848 16436 11854 16448
rect 13541 16439 13599 16445
rect 13541 16436 13553 16439
rect 11848 16408 13553 16436
rect 11848 16396 11854 16408
rect 13541 16405 13553 16408
rect 13587 16436 13599 16439
rect 17126 16436 17132 16448
rect 13587 16408 17132 16436
rect 13587 16405 13599 16408
rect 13541 16399 13599 16405
rect 17126 16396 17132 16408
rect 17184 16396 17190 16448
rect 19242 16436 19248 16448
rect 19203 16408 19248 16436
rect 19242 16396 19248 16408
rect 19300 16396 19306 16448
rect 19536 16436 19564 16535
rect 19720 16504 19748 16535
rect 20254 16532 20260 16584
rect 20312 16572 20318 16584
rect 20605 16575 20663 16581
rect 20605 16572 20617 16575
rect 20312 16544 20617 16572
rect 20312 16532 20318 16544
rect 20605 16541 20617 16544
rect 20651 16541 20663 16575
rect 20605 16535 20663 16541
rect 22002 16532 22008 16584
rect 22060 16572 22066 16584
rect 22094 16572 22100 16584
rect 22060 16544 22100 16572
rect 22060 16532 22066 16544
rect 22094 16532 22100 16544
rect 22152 16532 22158 16584
rect 24854 16572 24860 16584
rect 24815 16544 24860 16572
rect 24854 16532 24860 16544
rect 24912 16532 24918 16584
rect 25038 16572 25044 16584
rect 24999 16544 25044 16572
rect 25038 16532 25044 16544
rect 25096 16532 25102 16584
rect 25314 16532 25320 16584
rect 25372 16572 25378 16584
rect 25685 16575 25743 16581
rect 25685 16572 25697 16575
rect 25372 16544 25697 16572
rect 25372 16532 25378 16544
rect 25685 16541 25697 16544
rect 25731 16572 25743 16575
rect 26252 16572 26280 16612
rect 26973 16609 26985 16612
rect 27019 16609 27031 16643
rect 26973 16603 27031 16609
rect 27801 16643 27859 16649
rect 27801 16609 27813 16643
rect 27847 16640 27859 16643
rect 27982 16640 27988 16652
rect 27847 16612 27988 16640
rect 27847 16609 27859 16612
rect 27801 16603 27859 16609
rect 27982 16600 27988 16612
rect 28040 16640 28046 16652
rect 28902 16640 28908 16652
rect 28040 16612 28908 16640
rect 28040 16600 28046 16612
rect 28902 16600 28908 16612
rect 28960 16600 28966 16652
rect 25731 16544 26280 16572
rect 25731 16541 25743 16544
rect 25685 16535 25743 16541
rect 28350 16532 28356 16584
rect 28408 16572 28414 16584
rect 28810 16572 28816 16584
rect 28408 16544 28816 16572
rect 28408 16532 28414 16544
rect 28810 16532 28816 16544
rect 28868 16532 28874 16584
rect 30098 16532 30104 16584
rect 30156 16581 30162 16584
rect 30156 16575 30205 16581
rect 30156 16541 30159 16575
rect 30193 16541 30205 16575
rect 30156 16535 30205 16541
rect 30156 16532 30162 16535
rect 30287 16532 30293 16584
rect 30345 16575 30351 16584
rect 30576 16581 30604 16680
rect 31570 16600 31576 16652
rect 31628 16640 31634 16652
rect 33060 16649 33088 16680
rect 37826 16668 37832 16680
rect 37884 16668 37890 16720
rect 33045 16643 33103 16649
rect 33045 16640 33057 16643
rect 31628 16612 33057 16640
rect 31628 16600 31634 16612
rect 33045 16609 33057 16612
rect 33091 16609 33103 16643
rect 33045 16603 33103 16609
rect 34149 16643 34207 16649
rect 34149 16609 34161 16643
rect 34195 16640 34207 16643
rect 35618 16640 35624 16652
rect 34195 16612 34928 16640
rect 34195 16609 34207 16612
rect 34149 16603 34207 16609
rect 30398 16575 30456 16581
rect 30345 16532 30356 16575
rect 30398 16541 30410 16575
rect 30444 16572 30456 16575
rect 30561 16575 30619 16581
rect 30444 16544 30512 16572
rect 30444 16541 30456 16544
rect 30398 16535 30456 16541
rect 30298 16529 30356 16532
rect 19978 16504 19984 16516
rect 19720 16476 19984 16504
rect 19978 16464 19984 16476
rect 20036 16464 20042 16516
rect 22370 16504 22376 16516
rect 22283 16476 22376 16504
rect 22370 16464 22376 16476
rect 22428 16504 22434 16516
rect 25222 16504 25228 16516
rect 22428 16476 25228 16504
rect 22428 16464 22434 16476
rect 25222 16464 25228 16476
rect 25280 16464 25286 16516
rect 28258 16504 28264 16516
rect 28219 16476 28264 16504
rect 28258 16464 28264 16476
rect 28316 16464 28322 16516
rect 28445 16507 28503 16513
rect 28445 16473 28457 16507
rect 28491 16504 28503 16507
rect 29914 16504 29920 16516
rect 28491 16476 29920 16504
rect 28491 16473 28503 16476
rect 28445 16467 28503 16473
rect 29914 16464 29920 16476
rect 29972 16464 29978 16516
rect 19610 16436 19616 16448
rect 19536 16408 19616 16436
rect 19610 16396 19616 16408
rect 19668 16396 19674 16448
rect 21726 16436 21732 16448
rect 21687 16408 21732 16436
rect 21726 16396 21732 16408
rect 21784 16396 21790 16448
rect 25866 16436 25872 16448
rect 25827 16408 25872 16436
rect 25866 16396 25872 16408
rect 25924 16396 25930 16448
rect 30484 16436 30512 16544
rect 30561 16541 30573 16575
rect 30607 16541 30619 16575
rect 31202 16572 31208 16584
rect 31163 16544 31208 16572
rect 30561 16535 30619 16541
rect 31202 16532 31208 16544
rect 31260 16532 31266 16584
rect 32861 16575 32919 16581
rect 32861 16541 32873 16575
rect 32907 16572 32919 16575
rect 33594 16572 33600 16584
rect 32907 16544 33600 16572
rect 32907 16541 32919 16544
rect 32861 16535 32919 16541
rect 33594 16532 33600 16544
rect 33652 16532 33658 16584
rect 34698 16572 34704 16584
rect 34659 16544 34704 16572
rect 34698 16532 34704 16544
rect 34756 16532 34762 16584
rect 34900 16581 34928 16612
rect 35084 16612 35624 16640
rect 35084 16581 35112 16612
rect 35618 16600 35624 16612
rect 35676 16600 35682 16652
rect 34885 16575 34943 16581
rect 34885 16541 34897 16575
rect 34931 16541 34943 16575
rect 34977 16575 35035 16581
rect 34977 16572 34989 16575
rect 34885 16535 34943 16541
rect 34972 16541 34989 16572
rect 35023 16541 35035 16575
rect 34972 16535 35035 16541
rect 35069 16575 35127 16581
rect 35069 16541 35081 16575
rect 35115 16541 35127 16575
rect 35069 16535 35127 16541
rect 30834 16464 30840 16516
rect 30892 16504 30898 16516
rect 31021 16507 31079 16513
rect 31021 16504 31033 16507
rect 30892 16476 31033 16504
rect 30892 16464 30898 16476
rect 31021 16473 31033 16476
rect 31067 16473 31079 16507
rect 31021 16467 31079 16473
rect 33137 16507 33195 16513
rect 33137 16473 33149 16507
rect 33183 16504 33195 16507
rect 33318 16504 33324 16516
rect 33183 16476 33324 16504
rect 33183 16473 33195 16476
rect 33137 16467 33195 16473
rect 33318 16464 33324 16476
rect 33376 16464 33382 16516
rect 33778 16504 33784 16516
rect 33739 16476 33784 16504
rect 33778 16464 33784 16476
rect 33836 16464 33842 16516
rect 33965 16507 34023 16513
rect 33965 16473 33977 16507
rect 34011 16504 34023 16507
rect 34514 16504 34520 16516
rect 34011 16476 34520 16504
rect 34011 16473 34023 16476
rect 33965 16467 34023 16473
rect 34514 16464 34520 16476
rect 34572 16464 34578 16516
rect 31389 16439 31447 16445
rect 31389 16436 31401 16439
rect 30484 16408 31401 16436
rect 31389 16405 31401 16408
rect 31435 16405 31447 16439
rect 31389 16399 31447 16405
rect 32398 16396 32404 16448
rect 32456 16436 32462 16448
rect 32677 16439 32735 16445
rect 32677 16436 32689 16439
rect 32456 16408 32689 16436
rect 32456 16396 32462 16408
rect 32677 16405 32689 16408
rect 32723 16405 32735 16439
rect 32677 16399 32735 16405
rect 33226 16396 33232 16448
rect 33284 16436 33290 16448
rect 34972 16436 35000 16535
rect 35526 16532 35532 16584
rect 35584 16572 35590 16584
rect 37274 16572 37280 16584
rect 35584 16544 37280 16572
rect 35584 16532 35590 16544
rect 37274 16532 37280 16544
rect 37332 16532 37338 16584
rect 37440 16572 37498 16578
rect 37440 16538 37452 16572
rect 37486 16538 37498 16572
rect 37440 16532 37498 16538
rect 37540 16575 37598 16581
rect 37540 16541 37552 16575
rect 37586 16541 37598 16575
rect 37540 16535 37598 16541
rect 37691 16575 37749 16581
rect 37691 16541 37703 16575
rect 37737 16572 37749 16575
rect 37923 16572 37951 16748
rect 38286 16736 38292 16748
rect 38344 16736 38350 16788
rect 37737 16544 37951 16572
rect 37737 16541 37749 16544
rect 37691 16535 37749 16541
rect 37182 16464 37188 16516
rect 37240 16504 37246 16516
rect 37455 16504 37483 16532
rect 37240 16476 37483 16504
rect 37240 16464 37246 16476
rect 37568 16448 37596 16535
rect 37366 16436 37372 16448
rect 33284 16408 37372 16436
rect 33284 16396 33290 16408
rect 37366 16396 37372 16408
rect 37424 16436 37430 16448
rect 37550 16436 37556 16448
rect 37424 16408 37556 16436
rect 37424 16396 37430 16408
rect 37550 16396 37556 16408
rect 37608 16396 37614 16448
rect 37918 16436 37924 16448
rect 37879 16408 37924 16436
rect 37918 16396 37924 16408
rect 37976 16396 37982 16448
rect 1104 16346 68816 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 50294 16346
rect 50346 16294 50358 16346
rect 50410 16294 50422 16346
rect 50474 16294 50486 16346
rect 50538 16294 50550 16346
rect 50602 16294 68816 16346
rect 1104 16272 68816 16294
rect 3142 16232 3148 16244
rect 2976 16204 3148 16232
rect 2976 16105 3004 16204
rect 3142 16192 3148 16204
rect 3200 16192 3206 16244
rect 7650 16192 7656 16244
rect 7708 16232 7714 16244
rect 9401 16235 9459 16241
rect 9401 16232 9413 16235
rect 7708 16204 9413 16232
rect 7708 16192 7714 16204
rect 9401 16201 9413 16204
rect 9447 16201 9459 16235
rect 9401 16195 9459 16201
rect 10965 16235 11023 16241
rect 10965 16201 10977 16235
rect 11011 16232 11023 16235
rect 11238 16232 11244 16244
rect 11011 16204 11244 16232
rect 11011 16201 11023 16204
rect 10965 16195 11023 16201
rect 11238 16192 11244 16204
rect 11296 16192 11302 16244
rect 18230 16232 18236 16244
rect 18191 16204 18236 16232
rect 18230 16192 18236 16204
rect 18288 16192 18294 16244
rect 19337 16235 19395 16241
rect 19337 16201 19349 16235
rect 19383 16232 19395 16235
rect 19426 16232 19432 16244
rect 19383 16204 19432 16232
rect 19383 16201 19395 16204
rect 19337 16195 19395 16201
rect 19426 16192 19432 16204
rect 19484 16192 19490 16244
rect 20533 16235 20591 16241
rect 20533 16201 20545 16235
rect 20579 16232 20591 16235
rect 22370 16232 22376 16244
rect 20579 16204 22376 16232
rect 20579 16201 20591 16204
rect 20533 16195 20591 16201
rect 22370 16192 22376 16204
rect 22428 16192 22434 16244
rect 22925 16235 22983 16241
rect 22925 16201 22937 16235
rect 22971 16201 22983 16235
rect 22925 16195 22983 16201
rect 23569 16235 23627 16241
rect 23569 16201 23581 16235
rect 23615 16232 23627 16235
rect 24118 16232 24124 16244
rect 23615 16204 24124 16232
rect 23615 16201 23627 16204
rect 23569 16195 23627 16201
rect 9214 16164 9220 16176
rect 5828 16136 9220 16164
rect 2961 16099 3019 16105
rect 2961 16065 2973 16099
rect 3007 16065 3019 16099
rect 2961 16059 3019 16065
rect 3145 16102 3203 16108
rect 3145 16068 3157 16102
rect 3191 16068 3203 16102
rect 3145 16062 3203 16068
rect 3160 15972 3188 16062
rect 3234 16056 3240 16108
rect 3292 16096 3298 16108
rect 3418 16105 3424 16108
rect 3375 16099 3424 16105
rect 3292 16068 3337 16096
rect 3292 16056 3298 16068
rect 3375 16065 3387 16099
rect 3421 16065 3424 16099
rect 3375 16059 3424 16065
rect 3418 16056 3424 16059
rect 3476 16096 3482 16108
rect 5828 16105 5856 16136
rect 9214 16124 9220 16136
rect 9272 16164 9278 16176
rect 10597 16167 10655 16173
rect 10597 16164 10609 16167
rect 9272 16136 10609 16164
rect 9272 16124 9278 16136
rect 10597 16133 10609 16136
rect 10643 16133 10655 16167
rect 10597 16127 10655 16133
rect 10781 16167 10839 16173
rect 10781 16133 10793 16167
rect 10827 16164 10839 16167
rect 11790 16164 11796 16176
rect 10827 16136 11796 16164
rect 10827 16133 10839 16136
rect 10781 16127 10839 16133
rect 4065 16099 4123 16105
rect 4065 16096 4077 16099
rect 3476 16068 4077 16096
rect 3476 16056 3482 16068
rect 4065 16065 4077 16068
rect 4111 16065 4123 16099
rect 4065 16059 4123 16065
rect 5813 16099 5871 16105
rect 5813 16065 5825 16099
rect 5859 16065 5871 16099
rect 5813 16059 5871 16065
rect 6733 16099 6791 16105
rect 6733 16065 6745 16099
rect 6779 16065 6791 16099
rect 6733 16059 6791 16065
rect 6825 16099 6883 16105
rect 6825 16065 6837 16099
rect 6871 16065 6883 16099
rect 6825 16059 6883 16065
rect 3142 15920 3148 15972
rect 3200 15920 3206 15972
rect 6748 15960 6776 16059
rect 6840 16028 6868 16059
rect 6914 16056 6920 16108
rect 6972 16096 6978 16108
rect 7009 16099 7067 16105
rect 7009 16096 7021 16099
rect 6972 16068 7021 16096
rect 6972 16056 6978 16068
rect 7009 16065 7021 16068
rect 7055 16065 7067 16099
rect 7009 16059 7067 16065
rect 7101 16099 7159 16105
rect 7101 16065 7113 16099
rect 7147 16096 7159 16099
rect 9306 16096 9312 16108
rect 7147 16068 9312 16096
rect 7147 16065 7159 16068
rect 7101 16059 7159 16065
rect 9306 16056 9312 16068
rect 9364 16056 9370 16108
rect 9490 16096 9496 16108
rect 9451 16068 9496 16096
rect 9490 16056 9496 16068
rect 9548 16056 9554 16108
rect 7190 16028 7196 16040
rect 6840 16000 7196 16028
rect 7190 15988 7196 16000
rect 7248 15988 7254 16040
rect 7006 15960 7012 15972
rect 6748 15932 7012 15960
rect 7006 15920 7012 15932
rect 7064 15920 7070 15972
rect 10612 15960 10640 16127
rect 11790 16124 11796 16136
rect 11848 16124 11854 16176
rect 13630 16124 13636 16176
rect 13688 16164 13694 16176
rect 14921 16167 14979 16173
rect 14921 16164 14933 16167
rect 13688 16136 14933 16164
rect 13688 16124 13694 16136
rect 14921 16133 14933 16136
rect 14967 16133 14979 16167
rect 17770 16164 17776 16176
rect 17731 16136 17776 16164
rect 14921 16127 14979 16133
rect 17770 16124 17776 16136
rect 17828 16124 17834 16176
rect 18966 16164 18972 16176
rect 18927 16136 18972 16164
rect 18966 16124 18972 16136
rect 19024 16124 19030 16176
rect 19153 16167 19211 16173
rect 19153 16133 19165 16167
rect 19199 16164 19211 16167
rect 21726 16164 21732 16176
rect 19199 16136 21732 16164
rect 19199 16133 19211 16136
rect 19153 16127 19211 16133
rect 11514 16096 11520 16108
rect 11475 16068 11520 16096
rect 11514 16056 11520 16068
rect 11572 16056 11578 16108
rect 11698 16056 11704 16108
rect 11756 16096 11762 16108
rect 14553 16099 14611 16105
rect 14553 16096 14565 16099
rect 11756 16068 14565 16096
rect 11756 16056 11762 16068
rect 14553 16065 14565 16068
rect 14599 16065 14611 16099
rect 14553 16059 14611 16065
rect 14642 16056 14648 16108
rect 14700 16096 14706 16108
rect 14700 16068 14745 16096
rect 14700 16056 14706 16068
rect 14826 16056 14832 16108
rect 14884 16096 14890 16108
rect 14884 16068 14929 16096
rect 14884 16056 14890 16068
rect 15010 16056 15016 16108
rect 15068 16105 15074 16108
rect 15068 16096 15076 16105
rect 17954 16096 17960 16108
rect 15068 16068 15113 16096
rect 17915 16068 17960 16096
rect 15068 16059 15076 16068
rect 15068 16056 15074 16059
rect 17954 16056 17960 16068
rect 18012 16056 18018 16108
rect 18046 16056 18052 16108
rect 18104 16096 18110 16108
rect 18104 16068 18149 16096
rect 18104 16056 18110 16068
rect 11793 16031 11851 16037
rect 11793 15997 11805 16031
rect 11839 16028 11851 16031
rect 12066 16028 12072 16040
rect 11839 16000 12072 16028
rect 11839 15997 11851 16000
rect 11793 15991 11851 15997
rect 12066 15988 12072 16000
rect 12124 15988 12130 16040
rect 19168 16028 19196 16127
rect 21726 16124 21732 16136
rect 21784 16124 21790 16176
rect 22940 16164 22968 16195
rect 24118 16192 24124 16204
rect 24176 16192 24182 16244
rect 36446 16232 36452 16244
rect 25332 16204 36452 16232
rect 23198 16164 23204 16176
rect 22940 16136 23204 16164
rect 23198 16124 23204 16136
rect 23256 16164 23262 16176
rect 25332 16164 25360 16204
rect 36446 16192 36452 16204
rect 36504 16192 36510 16244
rect 40034 16232 40040 16244
rect 39995 16204 40040 16232
rect 40034 16192 40040 16204
rect 40092 16192 40098 16244
rect 23256 16136 25360 16164
rect 25440 16167 25498 16173
rect 23256 16124 23262 16136
rect 25440 16133 25452 16167
rect 25486 16164 25498 16167
rect 28169 16167 28227 16173
rect 28169 16164 28181 16167
rect 25486 16136 28181 16164
rect 25486 16133 25498 16136
rect 25440 16127 25498 16133
rect 28169 16133 28181 16136
rect 28215 16133 28227 16167
rect 35066 16164 35072 16176
rect 28169 16127 28227 16133
rect 31036 16136 35072 16164
rect 21085 16099 21143 16105
rect 21085 16065 21097 16099
rect 21131 16096 21143 16099
rect 22370 16096 22376 16108
rect 21131 16068 22376 16096
rect 21131 16065 21143 16068
rect 21085 16059 21143 16065
rect 22370 16056 22376 16068
rect 22428 16056 22434 16108
rect 22554 16096 22560 16108
rect 22515 16068 22560 16096
rect 22554 16056 22560 16068
rect 22612 16056 22618 16108
rect 23017 16099 23075 16105
rect 23017 16065 23029 16099
rect 23063 16065 23075 16099
rect 23750 16096 23756 16108
rect 23663 16068 23756 16096
rect 23017 16059 23075 16065
rect 18064 16000 19196 16028
rect 21269 16031 21327 16037
rect 11974 15960 11980 15972
rect 10612 15932 11980 15960
rect 11974 15920 11980 15932
rect 12032 15920 12038 15972
rect 3605 15895 3663 15901
rect 3605 15861 3617 15895
rect 3651 15892 3663 15895
rect 3878 15892 3884 15904
rect 3651 15864 3884 15892
rect 3651 15861 3663 15864
rect 3605 15855 3663 15861
rect 3878 15852 3884 15864
rect 3936 15852 3942 15904
rect 4706 15852 4712 15904
rect 4764 15892 4770 15904
rect 5629 15895 5687 15901
rect 5629 15892 5641 15895
rect 4764 15864 5641 15892
rect 4764 15852 4770 15864
rect 5629 15861 5641 15864
rect 5675 15861 5687 15895
rect 6546 15892 6552 15904
rect 6507 15864 6552 15892
rect 5629 15855 5687 15861
rect 6546 15852 6552 15864
rect 6604 15852 6610 15904
rect 15197 15895 15255 15901
rect 15197 15861 15209 15895
rect 15243 15892 15255 15895
rect 15562 15892 15568 15904
rect 15243 15864 15568 15892
rect 15243 15861 15255 15864
rect 15197 15855 15255 15861
rect 15562 15852 15568 15864
rect 15620 15852 15626 15904
rect 17034 15852 17040 15904
rect 17092 15892 17098 15904
rect 18064 15901 18092 16000
rect 21269 15997 21281 16031
rect 21315 16028 21327 16031
rect 22094 16028 22100 16040
rect 21315 16000 22100 16028
rect 21315 15997 21327 16000
rect 21269 15991 21327 15997
rect 22094 15988 22100 16000
rect 22152 16028 22158 16040
rect 23032 16028 23060 16059
rect 23750 16056 23756 16068
rect 23808 16096 23814 16108
rect 24578 16096 24584 16108
rect 23808 16068 24584 16096
rect 23808 16056 23814 16068
rect 24578 16056 24584 16068
rect 24636 16096 24642 16108
rect 24636 16068 25636 16096
rect 24636 16056 24642 16068
rect 22152 16000 23060 16028
rect 25608 16028 25636 16068
rect 25682 16056 25688 16108
rect 25740 16096 25746 16108
rect 26973 16099 27031 16105
rect 26973 16096 26985 16099
rect 25740 16068 25785 16096
rect 26344 16068 26985 16096
rect 25740 16056 25746 16068
rect 26344 16037 26372 16068
rect 26973 16065 26985 16068
rect 27019 16065 27031 16099
rect 26973 16059 27031 16065
rect 27706 16056 27712 16108
rect 27764 16096 27770 16108
rect 27982 16096 27988 16108
rect 27764 16068 27988 16096
rect 27764 16056 27770 16068
rect 27982 16056 27988 16068
rect 28040 16096 28046 16108
rect 28399 16099 28457 16105
rect 28399 16096 28411 16099
rect 28040 16068 28411 16096
rect 28040 16056 28046 16068
rect 28399 16065 28411 16068
rect 28445 16065 28457 16099
rect 28534 16096 28540 16108
rect 28495 16068 28540 16096
rect 28399 16059 28457 16065
rect 28534 16056 28540 16068
rect 28592 16056 28598 16108
rect 28629 16099 28687 16105
rect 28629 16065 28641 16099
rect 28675 16096 28687 16099
rect 28718 16096 28724 16108
rect 28675 16068 28724 16096
rect 28675 16065 28687 16068
rect 28629 16059 28687 16065
rect 28718 16056 28724 16068
rect 28776 16056 28782 16108
rect 28810 16056 28816 16108
rect 28868 16096 28874 16108
rect 30745 16099 30803 16105
rect 30745 16096 30757 16099
rect 28868 16068 30757 16096
rect 28868 16056 28874 16068
rect 30745 16065 30757 16068
rect 30791 16065 30803 16099
rect 30745 16059 30803 16065
rect 26329 16031 26387 16037
rect 26329 16028 26341 16031
rect 25608 16000 26341 16028
rect 22152 15988 22158 16000
rect 26329 15997 26341 16000
rect 26375 15997 26387 16031
rect 26329 15991 26387 15997
rect 30466 15988 30472 16040
rect 30524 16028 30530 16040
rect 31036 16037 31064 16136
rect 35066 16124 35072 16136
rect 35124 16124 35130 16176
rect 37918 16124 37924 16176
rect 37976 16164 37982 16176
rect 38902 16167 38960 16173
rect 38902 16164 38914 16167
rect 37976 16136 38914 16164
rect 37976 16124 37982 16136
rect 38902 16133 38914 16136
rect 38948 16133 38960 16167
rect 38902 16127 38960 16133
rect 32858 16056 32864 16108
rect 32916 16096 32922 16108
rect 33238 16099 33296 16105
rect 33238 16096 33250 16099
rect 32916 16068 33250 16096
rect 32916 16056 32922 16068
rect 33238 16065 33250 16068
rect 33284 16065 33296 16099
rect 33502 16096 33508 16108
rect 33463 16068 33508 16096
rect 33238 16059 33296 16065
rect 33502 16056 33508 16068
rect 33560 16056 33566 16108
rect 34882 16056 34888 16108
rect 34940 16096 34946 16108
rect 35526 16096 35532 16108
rect 34940 16068 35532 16096
rect 34940 16056 34946 16068
rect 35526 16056 35532 16068
rect 35584 16056 35590 16108
rect 35692 16099 35750 16105
rect 35692 16096 35704 16099
rect 35627 16068 35704 16096
rect 31021 16031 31079 16037
rect 31021 16028 31033 16031
rect 30524 16000 31033 16028
rect 30524 15988 30530 16000
rect 31021 15997 31033 16000
rect 31067 15997 31079 16031
rect 31021 15991 31079 15997
rect 33686 15988 33692 16040
rect 33744 16028 33750 16040
rect 34698 16028 34704 16040
rect 33744 16000 34704 16028
rect 33744 15988 33750 16000
rect 34698 15988 34704 16000
rect 34756 16028 34762 16040
rect 34793 16031 34851 16037
rect 34793 16028 34805 16031
rect 34756 16000 34805 16028
rect 34756 15988 34762 16000
rect 34793 15997 34805 16000
rect 34839 15997 34851 16031
rect 35066 16028 35072 16040
rect 35027 16000 35072 16028
rect 34793 15991 34851 15997
rect 35066 15988 35072 16000
rect 35124 16028 35130 16040
rect 35342 16028 35348 16040
rect 35124 16000 35348 16028
rect 35124 15988 35130 16000
rect 35342 15988 35348 16000
rect 35400 15988 35406 16040
rect 35434 15988 35440 16040
rect 35492 16028 35498 16040
rect 35627 16028 35655 16068
rect 35692 16065 35704 16068
rect 35738 16065 35750 16099
rect 35692 16059 35750 16065
rect 35802 16056 35808 16108
rect 35860 16096 35866 16108
rect 35986 16105 35992 16108
rect 35943 16099 35992 16105
rect 35860 16068 35905 16096
rect 35860 16056 35866 16068
rect 35943 16065 35955 16099
rect 35989 16065 35992 16099
rect 35943 16059 35992 16065
rect 35986 16056 35992 16059
rect 36044 16056 36050 16108
rect 37461 16099 37519 16105
rect 37461 16065 37473 16099
rect 37507 16065 37519 16099
rect 37642 16096 37648 16108
rect 37603 16068 37648 16096
rect 37461 16059 37519 16065
rect 35492 16000 35655 16028
rect 37476 16028 37504 16059
rect 37642 16056 37648 16068
rect 37700 16056 37706 16108
rect 38657 16099 38715 16105
rect 38657 16065 38669 16099
rect 38703 16096 38715 16099
rect 38746 16096 38752 16108
rect 38703 16068 38752 16096
rect 38703 16065 38715 16068
rect 38657 16059 38715 16065
rect 38746 16056 38752 16068
rect 38804 16056 38810 16108
rect 37918 16028 37924 16040
rect 37476 16000 37924 16028
rect 35492 15988 35498 16000
rect 37918 15988 37924 16000
rect 37976 15988 37982 16040
rect 18138 15920 18144 15972
rect 18196 15960 18202 15972
rect 22281 15963 22339 15969
rect 22281 15960 22293 15963
rect 18196 15932 22293 15960
rect 18196 15920 18202 15932
rect 22281 15929 22293 15932
rect 22327 15929 22339 15963
rect 22281 15923 22339 15929
rect 22649 15963 22707 15969
rect 22649 15929 22661 15963
rect 22695 15960 22707 15963
rect 24670 15960 24676 15972
rect 22695 15932 24676 15960
rect 22695 15929 22707 15932
rect 22649 15923 22707 15929
rect 24670 15920 24676 15932
rect 24728 15920 24734 15972
rect 28994 15960 29000 15972
rect 26252 15932 29000 15960
rect 18049 15895 18107 15901
rect 18049 15892 18061 15895
rect 17092 15864 18061 15892
rect 17092 15852 17098 15864
rect 18049 15861 18061 15864
rect 18095 15861 18107 15895
rect 18049 15855 18107 15861
rect 22738 15852 22744 15904
rect 22796 15892 22802 15904
rect 22796 15864 22841 15892
rect 22796 15852 22802 15864
rect 23474 15852 23480 15904
rect 23532 15892 23538 15904
rect 24305 15895 24363 15901
rect 24305 15892 24317 15895
rect 23532 15864 24317 15892
rect 23532 15852 23538 15864
rect 24305 15861 24317 15864
rect 24351 15892 24363 15895
rect 26252 15892 26280 15932
rect 28994 15920 29000 15932
rect 29052 15920 29058 15972
rect 27154 15892 27160 15904
rect 24351 15864 26280 15892
rect 27115 15864 27160 15892
rect 24351 15861 24363 15864
rect 24305 15855 24363 15861
rect 27154 15852 27160 15864
rect 27212 15852 27218 15904
rect 28350 15852 28356 15904
rect 28408 15892 28414 15904
rect 29641 15895 29699 15901
rect 29641 15892 29653 15895
rect 28408 15864 29653 15892
rect 28408 15852 28414 15864
rect 29641 15861 29653 15864
rect 29687 15892 29699 15895
rect 30006 15892 30012 15904
rect 29687 15864 30012 15892
rect 29687 15861 29699 15864
rect 29641 15855 29699 15861
rect 30006 15852 30012 15864
rect 30064 15852 30070 15904
rect 30098 15852 30104 15904
rect 30156 15892 30162 15904
rect 32125 15895 32183 15901
rect 32125 15892 32137 15895
rect 30156 15864 32137 15892
rect 30156 15852 30162 15864
rect 32125 15861 32137 15864
rect 32171 15892 32183 15895
rect 33594 15892 33600 15904
rect 32171 15864 33600 15892
rect 32171 15861 32183 15864
rect 32125 15855 32183 15861
rect 33594 15852 33600 15864
rect 33652 15852 33658 15904
rect 36170 15892 36176 15904
rect 36131 15864 36176 15892
rect 36170 15852 36176 15864
rect 36228 15852 36234 15904
rect 37277 15895 37335 15901
rect 37277 15861 37289 15895
rect 37323 15892 37335 15895
rect 37458 15892 37464 15904
rect 37323 15864 37464 15892
rect 37323 15861 37335 15864
rect 37277 15855 37335 15861
rect 37458 15852 37464 15864
rect 37516 15852 37522 15904
rect 67634 15892 67640 15904
rect 67595 15864 67640 15892
rect 67634 15852 67640 15864
rect 67692 15852 67698 15904
rect 1104 15802 68816 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 65654 15802
rect 65706 15750 65718 15802
rect 65770 15750 65782 15802
rect 65834 15750 65846 15802
rect 65898 15750 65910 15802
rect 65962 15750 68816 15802
rect 1104 15728 68816 15750
rect 1489 15691 1547 15697
rect 1489 15657 1501 15691
rect 1535 15688 1547 15691
rect 1762 15688 1768 15700
rect 1535 15660 1768 15688
rect 1535 15657 1547 15660
rect 1489 15651 1547 15657
rect 1762 15648 1768 15660
rect 1820 15648 1826 15700
rect 2774 15648 2780 15700
rect 2832 15688 2838 15700
rect 2832 15660 2877 15688
rect 2832 15648 2838 15660
rect 6454 15648 6460 15700
rect 6512 15688 6518 15700
rect 7193 15691 7251 15697
rect 7193 15688 7205 15691
rect 6512 15660 7205 15688
rect 6512 15648 6518 15660
rect 7193 15657 7205 15660
rect 7239 15657 7251 15691
rect 7193 15651 7251 15657
rect 9306 15648 9312 15700
rect 9364 15688 9370 15700
rect 11057 15691 11115 15697
rect 11057 15688 11069 15691
rect 9364 15660 11069 15688
rect 9364 15648 9370 15660
rect 11057 15657 11069 15660
rect 11103 15657 11115 15691
rect 11057 15651 11115 15657
rect 11517 15691 11575 15697
rect 11517 15657 11529 15691
rect 11563 15688 11575 15691
rect 11882 15688 11888 15700
rect 11563 15660 11888 15688
rect 11563 15657 11575 15660
rect 11517 15651 11575 15657
rect 11882 15648 11888 15660
rect 11940 15648 11946 15700
rect 11974 15648 11980 15700
rect 12032 15688 12038 15700
rect 14829 15691 14887 15697
rect 12032 15660 12077 15688
rect 12032 15648 12038 15660
rect 14829 15657 14841 15691
rect 14875 15688 14887 15691
rect 14918 15688 14924 15700
rect 14875 15660 14924 15688
rect 14875 15657 14887 15660
rect 14829 15651 14887 15657
rect 14918 15648 14924 15660
rect 14976 15648 14982 15700
rect 18322 15648 18328 15700
rect 18380 15688 18386 15700
rect 18509 15691 18567 15697
rect 18509 15688 18521 15691
rect 18380 15660 18521 15688
rect 18380 15648 18386 15660
rect 18509 15657 18521 15660
rect 18555 15657 18567 15691
rect 18509 15651 18567 15657
rect 19613 15691 19671 15697
rect 19613 15657 19625 15691
rect 19659 15688 19671 15691
rect 19978 15688 19984 15700
rect 19659 15660 19984 15688
rect 19659 15657 19671 15660
rect 19613 15651 19671 15657
rect 19978 15648 19984 15660
rect 20036 15648 20042 15700
rect 24581 15691 24639 15697
rect 24581 15657 24593 15691
rect 24627 15688 24639 15691
rect 27798 15688 27804 15700
rect 24627 15660 27804 15688
rect 24627 15657 24639 15660
rect 24581 15651 24639 15657
rect 27798 15648 27804 15660
rect 27856 15648 27862 15700
rect 28629 15691 28687 15697
rect 28629 15657 28641 15691
rect 28675 15688 28687 15691
rect 28718 15688 28724 15700
rect 28675 15660 28724 15688
rect 28675 15657 28687 15660
rect 28629 15651 28687 15657
rect 28718 15648 28724 15660
rect 28776 15648 28782 15700
rect 32858 15688 32864 15700
rect 32819 15660 32864 15688
rect 32858 15648 32864 15660
rect 32916 15648 32922 15700
rect 36906 15688 36912 15700
rect 36819 15660 36912 15688
rect 36906 15648 36912 15660
rect 36964 15688 36970 15700
rect 38102 15688 38108 15700
rect 36964 15660 38108 15688
rect 36964 15648 36970 15660
rect 38102 15648 38108 15660
rect 38160 15648 38166 15700
rect 9493 15623 9551 15629
rect 6196 15592 7328 15620
rect 2958 15552 2964 15564
rect 2792 15524 2964 15552
rect 1394 15444 1400 15496
rect 1452 15484 1458 15496
rect 1673 15487 1731 15493
rect 1673 15484 1685 15487
rect 1452 15456 1685 15484
rect 1452 15444 1458 15456
rect 1673 15453 1685 15456
rect 1719 15453 1731 15487
rect 1673 15447 1731 15453
rect 1949 15487 2007 15493
rect 1949 15453 1961 15487
rect 1995 15453 2007 15487
rect 2130 15484 2136 15496
rect 2091 15456 2136 15484
rect 1949 15447 2007 15453
rect 1964 15416 1992 15447
rect 2130 15444 2136 15456
rect 2188 15444 2194 15496
rect 2792 15493 2820 15524
rect 2958 15512 2964 15524
rect 3016 15552 3022 15564
rect 3418 15552 3424 15564
rect 3016 15524 3424 15552
rect 3016 15512 3022 15524
rect 3418 15512 3424 15524
rect 3476 15512 3482 15564
rect 2777 15487 2835 15493
rect 2777 15453 2789 15487
rect 2823 15453 2835 15487
rect 2777 15447 2835 15453
rect 2869 15487 2927 15493
rect 2869 15453 2881 15487
rect 2915 15453 2927 15487
rect 2869 15447 2927 15453
rect 1964 15388 2636 15416
rect 2608 15357 2636 15388
rect 2593 15351 2651 15357
rect 2593 15317 2605 15351
rect 2639 15317 2651 15351
rect 2884 15348 2912 15447
rect 3602 15444 3608 15496
rect 3660 15484 3666 15496
rect 3789 15487 3847 15493
rect 3789 15484 3801 15487
rect 3660 15456 3801 15484
rect 3660 15444 3666 15456
rect 3789 15453 3801 15456
rect 3835 15453 3847 15487
rect 3789 15447 3847 15453
rect 3878 15444 3884 15496
rect 3936 15484 3942 15496
rect 6196 15493 6224 15592
rect 7190 15552 7196 15564
rect 7151 15524 7196 15552
rect 7190 15512 7196 15524
rect 7248 15512 7254 15564
rect 7300 15561 7328 15592
rect 9493 15589 9505 15623
rect 9539 15620 9551 15623
rect 9539 15592 12940 15620
rect 9539 15589 9551 15592
rect 9493 15583 9551 15589
rect 7285 15555 7343 15561
rect 7285 15521 7297 15555
rect 7331 15552 7343 15555
rect 7926 15552 7932 15564
rect 7331 15524 7932 15552
rect 7331 15521 7343 15524
rect 7285 15515 7343 15521
rect 7926 15512 7932 15524
rect 7984 15512 7990 15564
rect 9582 15552 9588 15564
rect 8036 15524 9588 15552
rect 4045 15487 4103 15493
rect 4045 15484 4057 15487
rect 3936 15456 4057 15484
rect 3936 15444 3942 15456
rect 4045 15453 4057 15456
rect 4091 15453 4103 15487
rect 4045 15447 4103 15453
rect 6181 15487 6239 15493
rect 6181 15453 6193 15487
rect 6227 15453 6239 15487
rect 6181 15447 6239 15453
rect 6273 15487 6331 15493
rect 6273 15453 6285 15487
rect 6319 15453 6331 15487
rect 6454 15484 6460 15496
rect 6415 15456 6460 15484
rect 6273 15447 6331 15453
rect 3053 15419 3111 15425
rect 3053 15385 3065 15419
rect 3099 15416 3111 15419
rect 5997 15419 6055 15425
rect 5997 15416 6009 15419
rect 3099 15388 6009 15416
rect 3099 15385 3111 15388
rect 3053 15379 3111 15385
rect 5997 15385 6009 15388
rect 6043 15385 6055 15419
rect 6288 15416 6316 15447
rect 6454 15444 6460 15456
rect 6512 15444 6518 15496
rect 6546 15444 6552 15496
rect 6604 15484 6610 15496
rect 7377 15487 7435 15493
rect 7377 15484 7389 15487
rect 6604 15456 6649 15484
rect 6748 15456 7389 15484
rect 6604 15444 6610 15456
rect 6748 15416 6776 15456
rect 7377 15453 7389 15456
rect 7423 15484 7435 15487
rect 7650 15484 7656 15496
rect 7423 15456 7656 15484
rect 7423 15453 7435 15456
rect 7377 15447 7435 15453
rect 7650 15444 7656 15456
rect 7708 15444 7714 15496
rect 8036 15493 8064 15524
rect 7837 15487 7895 15493
rect 7837 15453 7849 15487
rect 7883 15453 7895 15487
rect 7837 15447 7895 15453
rect 8021 15487 8079 15493
rect 8021 15453 8033 15487
rect 8067 15453 8079 15487
rect 8021 15447 8079 15453
rect 8205 15487 8263 15493
rect 8205 15453 8217 15487
rect 8251 15484 8263 15487
rect 8386 15484 8392 15496
rect 8251 15456 8392 15484
rect 8251 15453 8263 15456
rect 8205 15447 8263 15453
rect 7006 15416 7012 15428
rect 6288 15388 6776 15416
rect 6967 15388 7012 15416
rect 5997 15379 6055 15385
rect 7006 15376 7012 15388
rect 7064 15376 7070 15428
rect 4890 15348 4896 15360
rect 2884 15320 4896 15348
rect 2593 15311 2651 15317
rect 4890 15308 4896 15320
rect 4948 15308 4954 15360
rect 5169 15351 5227 15357
rect 5169 15317 5181 15351
rect 5215 15348 5227 15351
rect 5258 15348 5264 15360
rect 5215 15320 5264 15348
rect 5215 15317 5227 15320
rect 5169 15311 5227 15317
rect 5258 15308 5264 15320
rect 5316 15308 5322 15360
rect 6638 15308 6644 15360
rect 6696 15348 6702 15360
rect 7852 15348 7880 15447
rect 8386 15444 8392 15456
rect 8444 15444 8450 15496
rect 8478 15444 8484 15496
rect 8536 15484 8542 15496
rect 9140 15493 9168 15524
rect 9582 15512 9588 15524
rect 9640 15512 9646 15564
rect 11790 15552 11796 15564
rect 9692 15524 10456 15552
rect 8941 15487 8999 15493
rect 8941 15484 8953 15487
rect 8536 15456 8953 15484
rect 8536 15444 8542 15456
rect 8941 15453 8953 15456
rect 8987 15453 8999 15487
rect 8941 15447 8999 15453
rect 9125 15487 9183 15493
rect 9125 15453 9137 15487
rect 9171 15484 9183 15487
rect 9309 15487 9367 15493
rect 9171 15456 9205 15484
rect 9171 15453 9183 15456
rect 9125 15447 9183 15453
rect 9309 15453 9321 15487
rect 9355 15484 9367 15487
rect 9692 15484 9720 15524
rect 9355 15456 9720 15484
rect 9355 15453 9367 15456
rect 9309 15447 9367 15453
rect 9766 15444 9772 15496
rect 9824 15484 9830 15496
rect 10045 15487 10103 15493
rect 10045 15484 10057 15487
rect 9824 15456 10057 15484
rect 9824 15444 9830 15456
rect 10045 15453 10057 15456
rect 10091 15453 10103 15487
rect 10318 15484 10324 15496
rect 10279 15456 10324 15484
rect 10045 15447 10103 15453
rect 10318 15444 10324 15456
rect 10376 15444 10382 15496
rect 10428 15493 10456 15524
rect 11256 15524 11796 15552
rect 10413 15487 10471 15493
rect 10413 15453 10425 15487
rect 10459 15484 10471 15487
rect 10686 15484 10692 15496
rect 10459 15456 10692 15484
rect 10459 15453 10471 15456
rect 10413 15447 10471 15453
rect 10686 15444 10692 15456
rect 10744 15444 10750 15496
rect 11256 15493 11284 15524
rect 11790 15512 11796 15524
rect 11848 15512 11854 15564
rect 11241 15487 11299 15493
rect 11241 15453 11253 15487
rect 11287 15453 11299 15487
rect 11241 15447 11299 15453
rect 11330 15444 11336 15496
rect 11388 15484 11394 15496
rect 11517 15487 11575 15493
rect 11388 15456 11433 15484
rect 11388 15444 11394 15456
rect 11517 15453 11529 15487
rect 11563 15484 11575 15487
rect 11606 15484 11612 15496
rect 11563 15456 11612 15484
rect 11563 15453 11575 15456
rect 11517 15447 11575 15453
rect 11606 15444 11612 15456
rect 11664 15444 11670 15496
rect 12161 15487 12219 15493
rect 12161 15453 12173 15487
rect 12207 15453 12219 15487
rect 12161 15447 12219 15453
rect 12345 15487 12403 15493
rect 12345 15453 12357 15487
rect 12391 15484 12403 15487
rect 12618 15484 12624 15496
rect 12391 15456 12624 15484
rect 12391 15453 12403 15456
rect 12345 15447 12403 15453
rect 8110 15416 8116 15428
rect 8071 15388 8116 15416
rect 8110 15376 8116 15388
rect 8168 15376 8174 15428
rect 8846 15376 8852 15428
rect 8904 15416 8910 15428
rect 9217 15419 9275 15425
rect 9217 15416 9229 15419
rect 8904 15388 9229 15416
rect 8904 15376 8910 15388
rect 9217 15385 9229 15388
rect 9263 15385 9275 15419
rect 9217 15379 9275 15385
rect 9582 15376 9588 15428
rect 9640 15416 9646 15428
rect 10229 15419 10287 15425
rect 10229 15416 10241 15419
rect 9640 15388 10241 15416
rect 9640 15376 9646 15388
rect 10229 15385 10241 15388
rect 10275 15385 10287 15419
rect 11698 15416 11704 15428
rect 10229 15379 10287 15385
rect 10428 15388 11704 15416
rect 6696 15320 7880 15348
rect 8389 15351 8447 15357
rect 6696 15308 6702 15320
rect 8389 15317 8401 15351
rect 8435 15348 8447 15351
rect 10428 15348 10456 15388
rect 11698 15376 11704 15388
rect 11756 15376 11762 15428
rect 12176 15416 12204 15447
rect 12618 15444 12624 15456
rect 12676 15444 12682 15496
rect 12912 15493 12940 15592
rect 12986 15580 12992 15632
rect 13044 15620 13050 15632
rect 17862 15620 17868 15632
rect 13044 15592 13446 15620
rect 13044 15580 13050 15592
rect 13418 15552 13446 15592
rect 15120 15592 17868 15620
rect 15010 15552 15016 15564
rect 13418 15524 15016 15552
rect 13078 15493 13084 15496
rect 12897 15487 12955 15493
rect 12897 15453 12909 15487
rect 12943 15453 12955 15487
rect 12897 15447 12955 15453
rect 13045 15487 13084 15493
rect 13045 15453 13057 15487
rect 13045 15447 13084 15453
rect 13078 15444 13084 15447
rect 13136 15444 13142 15496
rect 13418 15493 13446 15524
rect 15010 15512 15016 15524
rect 15068 15512 15074 15564
rect 13403 15487 13461 15493
rect 13403 15453 13415 15487
rect 13449 15453 13461 15487
rect 13403 15447 13461 15453
rect 14274 15444 14280 15496
rect 14332 15484 14338 15496
rect 14737 15487 14795 15493
rect 14737 15484 14749 15487
rect 14332 15456 14749 15484
rect 14332 15444 14338 15456
rect 14737 15453 14749 15456
rect 14783 15484 14795 15487
rect 14826 15484 14832 15496
rect 14783 15456 14832 15484
rect 14783 15453 14795 15456
rect 14737 15447 14795 15453
rect 14826 15444 14832 15456
rect 14884 15444 14890 15496
rect 14918 15444 14924 15496
rect 14976 15484 14982 15496
rect 15120 15484 15148 15592
rect 17862 15580 17868 15592
rect 17920 15580 17926 15632
rect 23293 15623 23351 15629
rect 23293 15589 23305 15623
rect 23339 15589 23351 15623
rect 23293 15583 23351 15589
rect 25409 15623 25467 15629
rect 25409 15589 25421 15623
rect 25455 15620 25467 15623
rect 25958 15620 25964 15632
rect 25455 15592 25964 15620
rect 25455 15589 25467 15592
rect 25409 15583 25467 15589
rect 15194 15512 15200 15564
rect 15252 15552 15258 15564
rect 23308 15552 23336 15583
rect 25958 15580 25964 15592
rect 26016 15580 26022 15632
rect 29730 15580 29736 15632
rect 29788 15620 29794 15632
rect 34057 15623 34115 15629
rect 34057 15620 34069 15623
rect 29788 15592 34069 15620
rect 29788 15580 29794 15592
rect 34057 15589 34069 15592
rect 34103 15620 34115 15623
rect 34514 15620 34520 15632
rect 34103 15592 34520 15620
rect 34103 15589 34115 15592
rect 34057 15583 34115 15589
rect 34514 15580 34520 15592
rect 34572 15580 34578 15632
rect 27522 15552 27528 15564
rect 15252 15524 26464 15552
rect 15252 15512 15258 15524
rect 14976 15456 15148 15484
rect 15565 15487 15623 15493
rect 14976 15444 14982 15456
rect 15565 15453 15577 15487
rect 15611 15484 15623 15487
rect 15746 15484 15752 15496
rect 15611 15456 15752 15484
rect 15611 15453 15623 15456
rect 15565 15447 15623 15453
rect 15746 15444 15752 15456
rect 15804 15444 15810 15496
rect 15841 15487 15899 15493
rect 15841 15453 15853 15487
rect 15887 15453 15899 15487
rect 16850 15484 16856 15496
rect 16811 15456 16856 15484
rect 15841 15447 15899 15453
rect 12802 15416 12808 15428
rect 11808 15388 12112 15416
rect 12176 15388 12808 15416
rect 10594 15348 10600 15360
rect 8435 15320 10456 15348
rect 10555 15320 10600 15348
rect 8435 15317 8447 15320
rect 8389 15311 8447 15317
rect 10594 15308 10600 15320
rect 10652 15308 10658 15360
rect 11330 15308 11336 15360
rect 11388 15348 11394 15360
rect 11808 15348 11836 15388
rect 11388 15320 11836 15348
rect 12084 15348 12112 15388
rect 12802 15376 12808 15388
rect 12860 15376 12866 15428
rect 13170 15416 13176 15428
rect 13131 15388 13176 15416
rect 13170 15376 13176 15388
rect 13228 15376 13234 15428
rect 13265 15419 13323 15425
rect 13265 15385 13277 15419
rect 13311 15385 13323 15419
rect 14844 15416 14872 15444
rect 15856 15416 15884 15447
rect 16850 15444 16856 15456
rect 16908 15444 16914 15496
rect 17034 15493 17040 15496
rect 17001 15487 17040 15493
rect 17001 15453 17013 15487
rect 17001 15447 17040 15453
rect 17034 15444 17040 15447
rect 17092 15444 17098 15496
rect 17218 15484 17224 15496
rect 17179 15456 17224 15484
rect 17218 15444 17224 15456
rect 17276 15444 17282 15496
rect 17310 15444 17316 15496
rect 17368 15493 17374 15496
rect 17368 15484 17376 15493
rect 17368 15456 17413 15484
rect 17368 15447 17376 15456
rect 17368 15444 17374 15447
rect 18046 15444 18052 15496
rect 18104 15484 18110 15496
rect 19429 15487 19487 15493
rect 19429 15484 19441 15487
rect 18104 15456 19441 15484
rect 18104 15444 18110 15456
rect 19429 15453 19441 15456
rect 19475 15484 19487 15487
rect 20254 15484 20260 15496
rect 19475 15456 20260 15484
rect 19475 15453 19487 15456
rect 19429 15447 19487 15453
rect 20254 15444 20260 15456
rect 20312 15444 20318 15496
rect 24394 15484 24400 15496
rect 24355 15456 24400 15484
rect 24394 15444 24400 15456
rect 24452 15444 24458 15496
rect 25222 15484 25228 15496
rect 25183 15456 25228 15484
rect 25222 15444 25228 15456
rect 25280 15444 25286 15496
rect 26436 15484 26464 15524
rect 27356 15524 27528 15552
rect 26878 15484 26884 15496
rect 26436 15456 26884 15484
rect 26878 15444 26884 15456
rect 26936 15484 26942 15496
rect 27356 15484 27384 15524
rect 27522 15512 27528 15524
rect 27580 15512 27586 15564
rect 27798 15512 27804 15564
rect 27856 15552 27862 15564
rect 30558 15552 30564 15564
rect 27856 15524 30564 15552
rect 27856 15512 27862 15524
rect 30558 15512 30564 15524
rect 30616 15552 30622 15564
rect 30929 15555 30987 15561
rect 30929 15552 30941 15555
rect 30616 15524 30941 15552
rect 30616 15512 30622 15524
rect 30929 15521 30941 15524
rect 30975 15552 30987 15555
rect 31110 15552 31116 15564
rect 30975 15524 31116 15552
rect 30975 15521 30987 15524
rect 30929 15515 30987 15521
rect 31110 15512 31116 15524
rect 31168 15512 31174 15564
rect 31478 15552 31484 15564
rect 31439 15524 31484 15552
rect 31478 15512 31484 15524
rect 31536 15552 31542 15564
rect 34701 15555 34759 15561
rect 34701 15552 34713 15555
rect 31536 15524 33272 15552
rect 31536 15512 31542 15524
rect 26936 15456 27384 15484
rect 27433 15487 27491 15493
rect 26936 15444 26942 15456
rect 27433 15453 27445 15487
rect 27479 15484 27491 15487
rect 27614 15484 27620 15496
rect 27479 15456 27620 15484
rect 27479 15453 27491 15456
rect 27433 15447 27491 15453
rect 27614 15444 27620 15456
rect 27672 15444 27678 15496
rect 28534 15444 28540 15496
rect 28592 15484 28598 15496
rect 28592 15456 29132 15484
rect 28592 15444 28598 15456
rect 14844 15388 15884 15416
rect 13265 15379 13323 15385
rect 13280 15348 13308 15379
rect 15930 15376 15936 15428
rect 15988 15416 15994 15428
rect 17129 15419 17187 15425
rect 17129 15416 17141 15419
rect 15988 15388 17141 15416
rect 15988 15376 15994 15388
rect 17129 15385 17141 15388
rect 17175 15385 17187 15419
rect 17129 15379 17187 15385
rect 18414 15376 18420 15428
rect 18472 15416 18478 15428
rect 18601 15419 18659 15425
rect 18601 15416 18613 15419
rect 18472 15388 18613 15416
rect 18472 15376 18478 15388
rect 18601 15385 18613 15388
rect 18647 15385 18659 15419
rect 18601 15379 18659 15385
rect 18966 15376 18972 15428
rect 19024 15416 19030 15428
rect 19245 15419 19303 15425
rect 19245 15416 19257 15419
rect 19024 15388 19257 15416
rect 19024 15376 19030 15388
rect 19245 15385 19257 15388
rect 19291 15385 19303 15419
rect 19245 15379 19303 15385
rect 20901 15419 20959 15425
rect 20901 15385 20913 15419
rect 20947 15416 20959 15419
rect 21266 15416 21272 15428
rect 20947 15388 21272 15416
rect 20947 15385 20959 15388
rect 20901 15379 20959 15385
rect 21266 15376 21272 15388
rect 21324 15416 21330 15428
rect 21818 15416 21824 15428
rect 21324 15388 21824 15416
rect 21324 15376 21330 15388
rect 21818 15376 21824 15388
rect 21876 15376 21882 15428
rect 22002 15416 22008 15428
rect 21963 15388 22008 15416
rect 22002 15376 22008 15388
rect 22060 15376 22066 15428
rect 25314 15416 25320 15428
rect 24412 15388 25320 15416
rect 13538 15348 13544 15360
rect 12084 15320 13308 15348
rect 13499 15320 13544 15348
rect 11388 15308 11394 15320
rect 13538 15308 13544 15320
rect 13596 15308 13602 15360
rect 14277 15351 14335 15357
rect 14277 15317 14289 15351
rect 14323 15348 14335 15351
rect 14366 15348 14372 15360
rect 14323 15320 14372 15348
rect 14323 15317 14335 15320
rect 14277 15311 14335 15317
rect 14366 15308 14372 15320
rect 14424 15348 14430 15360
rect 14918 15348 14924 15360
rect 14424 15320 14924 15348
rect 14424 15308 14430 15320
rect 14918 15308 14924 15320
rect 14976 15308 14982 15360
rect 17497 15351 17555 15357
rect 17497 15317 17509 15351
rect 17543 15348 17555 15351
rect 18230 15348 18236 15360
rect 17543 15320 18236 15348
rect 17543 15317 17555 15320
rect 17497 15311 17555 15317
rect 18230 15308 18236 15320
rect 18288 15308 18294 15360
rect 21545 15351 21603 15357
rect 21545 15317 21557 15351
rect 21591 15348 21603 15351
rect 22830 15348 22836 15360
rect 21591 15320 22836 15348
rect 21591 15317 21603 15320
rect 21545 15311 21603 15317
rect 22830 15308 22836 15320
rect 22888 15348 22894 15360
rect 24412 15348 24440 15388
rect 25314 15376 25320 15388
rect 25372 15376 25378 15428
rect 27188 15419 27246 15425
rect 27188 15385 27200 15419
rect 27234 15416 27246 15419
rect 27234 15388 28212 15416
rect 27234 15385 27246 15388
rect 27188 15379 27246 15385
rect 22888 15320 24440 15348
rect 22888 15308 22894 15320
rect 25682 15308 25688 15360
rect 25740 15348 25746 15360
rect 26053 15351 26111 15357
rect 26053 15348 26065 15351
rect 25740 15320 26065 15348
rect 25740 15308 25746 15320
rect 26053 15317 26065 15320
rect 26099 15317 26111 15351
rect 28184 15348 28212 15388
rect 28258 15376 28264 15428
rect 28316 15416 28322 15428
rect 28445 15419 28503 15425
rect 28316 15388 28361 15416
rect 28316 15376 28322 15388
rect 28445 15385 28457 15419
rect 28491 15416 28503 15419
rect 28994 15416 29000 15428
rect 28491 15388 29000 15416
rect 28491 15385 28503 15388
rect 28445 15379 28503 15385
rect 28994 15376 29000 15388
rect 29052 15376 29058 15428
rect 29104 15416 29132 15456
rect 29638 15444 29644 15496
rect 29696 15484 29702 15496
rect 29822 15484 29828 15496
rect 29696 15456 29828 15484
rect 29696 15444 29702 15456
rect 29822 15444 29828 15456
rect 29880 15444 29886 15496
rect 29917 15487 29975 15493
rect 29917 15453 29929 15487
rect 29963 15453 29975 15487
rect 29917 15447 29975 15453
rect 29932 15416 29960 15447
rect 30006 15444 30012 15496
rect 30064 15484 30070 15496
rect 30064 15456 30109 15484
rect 30064 15444 30070 15456
rect 30190 15444 30196 15496
rect 30248 15484 30254 15496
rect 31754 15484 31760 15496
rect 30248 15456 30293 15484
rect 31036 15456 31760 15484
rect 30248 15444 30254 15456
rect 30282 15416 30288 15428
rect 29104 15388 30288 15416
rect 30282 15376 30288 15388
rect 30340 15416 30346 15428
rect 31036 15416 31064 15456
rect 31754 15444 31760 15456
rect 31812 15444 31818 15496
rect 33244 15493 33272 15524
rect 33336 15524 34713 15552
rect 33336 15493 33364 15524
rect 34701 15521 34713 15524
rect 34747 15521 34759 15555
rect 34701 15515 34759 15521
rect 33137 15487 33195 15493
rect 33137 15453 33149 15487
rect 33183 15453 33195 15487
rect 33137 15447 33195 15453
rect 33229 15487 33287 15493
rect 33229 15453 33241 15487
rect 33275 15453 33287 15487
rect 33229 15447 33287 15453
rect 33321 15487 33379 15493
rect 33321 15453 33333 15487
rect 33367 15453 33379 15487
rect 33321 15447 33379 15453
rect 30340 15388 31064 15416
rect 30340 15376 30346 15388
rect 31110 15376 31116 15428
rect 31168 15416 31174 15428
rect 33152 15416 33180 15447
rect 33410 15444 33416 15496
rect 33468 15484 33474 15496
rect 33505 15487 33563 15493
rect 33505 15484 33517 15487
rect 33468 15456 33517 15484
rect 33468 15444 33474 15456
rect 33505 15453 33517 15456
rect 33551 15453 33563 15487
rect 33505 15447 33563 15453
rect 31168 15388 33180 15416
rect 33520 15416 33548 15447
rect 33594 15444 33600 15496
rect 33652 15484 33658 15496
rect 34885 15487 34943 15493
rect 34885 15484 34897 15487
rect 33652 15456 34897 15484
rect 33652 15444 33658 15456
rect 34885 15453 34897 15456
rect 34931 15453 34943 15487
rect 34885 15447 34943 15453
rect 35342 15444 35348 15496
rect 35400 15484 35406 15496
rect 35529 15487 35587 15493
rect 35529 15484 35541 15487
rect 35400 15456 35541 15484
rect 35400 15444 35406 15456
rect 35529 15453 35541 15456
rect 35575 15453 35587 15487
rect 35529 15447 35587 15453
rect 35796 15487 35854 15493
rect 35796 15453 35808 15487
rect 35842 15484 35854 15487
rect 36170 15484 36176 15496
rect 35842 15456 36176 15484
rect 35842 15453 35854 15456
rect 35796 15447 35854 15453
rect 36170 15444 36176 15456
rect 36228 15444 36234 15496
rect 39298 15484 39304 15496
rect 39259 15456 39304 15484
rect 39298 15444 39304 15456
rect 39356 15444 39362 15496
rect 34790 15416 34796 15428
rect 33520 15388 34796 15416
rect 31168 15376 31174 15388
rect 34790 15376 34796 15388
rect 34848 15376 34854 15428
rect 35069 15419 35127 15425
rect 35069 15385 35081 15419
rect 35115 15416 35127 15419
rect 37642 15416 37648 15428
rect 35115 15388 37648 15416
rect 35115 15385 35127 15388
rect 35069 15379 35127 15385
rect 29549 15351 29607 15357
rect 29549 15348 29561 15351
rect 28184 15320 29561 15348
rect 26053 15311 26111 15317
rect 29549 15317 29561 15320
rect 29595 15317 29607 15351
rect 29549 15311 29607 15317
rect 30374 15308 30380 15360
rect 30432 15348 30438 15360
rect 30834 15348 30840 15360
rect 30432 15320 30840 15348
rect 30432 15308 30438 15320
rect 30834 15308 30840 15320
rect 30892 15308 30898 15360
rect 32122 15308 32128 15360
rect 32180 15348 32186 15360
rect 33686 15348 33692 15360
rect 32180 15320 33692 15348
rect 32180 15308 32186 15320
rect 33686 15308 33692 15320
rect 33744 15308 33750 15360
rect 33778 15308 33784 15360
rect 33836 15348 33842 15360
rect 35084 15348 35112 15379
rect 37642 15376 37648 15388
rect 37700 15376 37706 15428
rect 38654 15376 38660 15428
rect 38712 15416 38718 15428
rect 39034 15419 39092 15425
rect 39034 15416 39046 15419
rect 38712 15388 39046 15416
rect 38712 15376 38718 15388
rect 39034 15385 39046 15388
rect 39080 15385 39092 15419
rect 39034 15379 39092 15385
rect 37918 15348 37924 15360
rect 33836 15320 35112 15348
rect 37879 15320 37924 15348
rect 33836 15308 33842 15320
rect 37918 15308 37924 15320
rect 37976 15308 37982 15360
rect 1104 15258 68816 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 50294 15258
rect 50346 15206 50358 15258
rect 50410 15206 50422 15258
rect 50474 15206 50486 15258
rect 50538 15206 50550 15258
rect 50602 15206 68816 15258
rect 1104 15184 68816 15206
rect 3142 15104 3148 15156
rect 3200 15144 3206 15156
rect 3329 15147 3387 15153
rect 3329 15144 3341 15147
rect 3200 15116 3341 15144
rect 3200 15104 3206 15116
rect 3329 15113 3341 15116
rect 3375 15113 3387 15147
rect 4890 15144 4896 15156
rect 4851 15116 4896 15144
rect 3329 15107 3387 15113
rect 4890 15104 4896 15116
rect 4948 15104 4954 15156
rect 7834 15104 7840 15156
rect 7892 15144 7898 15156
rect 8205 15147 8263 15153
rect 8205 15144 8217 15147
rect 7892 15116 8217 15144
rect 7892 15104 7898 15116
rect 8205 15113 8217 15116
rect 8251 15113 8263 15147
rect 8205 15107 8263 15113
rect 8938 15104 8944 15156
rect 8996 15144 9002 15156
rect 9493 15147 9551 15153
rect 9493 15144 9505 15147
rect 8996 15116 9505 15144
rect 8996 15104 9002 15116
rect 9493 15113 9505 15116
rect 9539 15113 9551 15147
rect 11054 15144 11060 15156
rect 9493 15107 9551 15113
rect 9600 15116 11060 15144
rect 4706 15076 4712 15088
rect 2976 15048 4712 15076
rect 2590 14968 2596 15020
rect 2648 15008 2654 15020
rect 2976 15017 3004 15048
rect 4706 15036 4712 15048
rect 4764 15036 4770 15088
rect 7466 15036 7472 15088
rect 7524 15076 7530 15088
rect 9600 15076 9628 15116
rect 11054 15104 11060 15116
rect 11112 15144 11118 15156
rect 11793 15147 11851 15153
rect 11793 15144 11805 15147
rect 11112 15116 11805 15144
rect 11112 15104 11118 15116
rect 11793 15113 11805 15116
rect 11839 15113 11851 15147
rect 11793 15107 11851 15113
rect 12618 15104 12624 15156
rect 12676 15104 12682 15156
rect 16942 15144 16948 15156
rect 14108 15116 16948 15144
rect 7524 15048 9628 15076
rect 7524 15036 7530 15048
rect 11698 15036 11704 15088
rect 11756 15076 11762 15088
rect 12636 15076 12664 15104
rect 11756 15048 12664 15076
rect 12805 15079 12863 15085
rect 11756 15036 11762 15048
rect 12805 15045 12817 15079
rect 12851 15076 12863 15079
rect 13170 15076 13176 15088
rect 12851 15048 13176 15076
rect 12851 15045 12863 15048
rect 12805 15039 12863 15045
rect 13170 15036 13176 15048
rect 13228 15036 13234 15088
rect 2961 15011 3019 15017
rect 2961 15008 2973 15011
rect 2648 14980 2973 15008
rect 2648 14968 2654 14980
rect 2961 14977 2973 14980
rect 3007 14977 3019 15011
rect 2961 14971 3019 14977
rect 3145 15011 3203 15017
rect 3145 14977 3157 15011
rect 3191 15008 3203 15011
rect 5077 15011 5135 15017
rect 3191 14980 3924 15008
rect 3191 14977 3203 14980
rect 3145 14971 3203 14977
rect 3896 14949 3924 14980
rect 5077 14977 5089 15011
rect 5123 15008 5135 15011
rect 5166 15008 5172 15020
rect 5123 14980 5172 15008
rect 5123 14977 5135 14980
rect 5077 14971 5135 14977
rect 5166 14968 5172 14980
rect 5224 14968 5230 15020
rect 5350 14968 5356 15020
rect 5408 15008 5414 15020
rect 7558 15008 7564 15020
rect 5408 14980 7564 15008
rect 5408 14968 5414 14980
rect 7558 14968 7564 14980
rect 7616 14968 7622 15020
rect 8386 15008 8392 15020
rect 8347 14980 8392 15008
rect 8386 14968 8392 14980
rect 8444 15008 8450 15020
rect 8846 15008 8852 15020
rect 8444 14980 8852 15008
rect 8444 14968 8450 14980
rect 8846 14968 8852 14980
rect 8904 15008 8910 15020
rect 9401 15011 9459 15017
rect 9401 15008 9413 15011
rect 8904 14980 9413 15008
rect 8904 14968 8910 14980
rect 9401 14977 9413 14980
rect 9447 14977 9459 15011
rect 9401 14971 9459 14977
rect 9585 15011 9643 15017
rect 9585 14977 9597 15011
rect 9631 15008 9643 15011
rect 10226 15008 10232 15020
rect 9631 14980 10232 15008
rect 9631 14977 9643 14980
rect 9585 14971 9643 14977
rect 10226 14968 10232 14980
rect 10284 15008 10290 15020
rect 11790 15008 11796 15020
rect 10284 14980 11796 15008
rect 10284 14968 10290 14980
rect 11790 14968 11796 14980
rect 11848 14968 11854 15020
rect 11974 14968 11980 15020
rect 12032 15008 12038 15020
rect 12526 15008 12532 15020
rect 12032 14980 12077 15008
rect 12487 14980 12532 15008
rect 12032 14968 12038 14980
rect 12526 14968 12532 14980
rect 12584 14968 12590 15020
rect 12710 15017 12716 15020
rect 12677 15011 12716 15017
rect 12677 14977 12689 15011
rect 12677 14971 12716 14977
rect 12710 14968 12716 14971
rect 12768 14968 12774 15020
rect 12897 15011 12955 15017
rect 12897 14977 12909 15011
rect 12943 14977 12955 15011
rect 12897 14971 12955 14977
rect 3881 14943 3939 14949
rect 3881 14909 3893 14943
rect 3927 14940 3939 14943
rect 5258 14940 5264 14952
rect 3927 14912 5264 14940
rect 3927 14909 3939 14912
rect 3881 14903 3939 14909
rect 5258 14900 5264 14912
rect 5316 14900 5322 14952
rect 8573 14943 8631 14949
rect 8573 14909 8585 14943
rect 8619 14940 8631 14943
rect 11698 14940 11704 14952
rect 8619 14912 11704 14940
rect 8619 14909 8631 14912
rect 8573 14903 8631 14909
rect 8386 14832 8392 14884
rect 8444 14872 8450 14884
rect 8588 14872 8616 14903
rect 11698 14900 11704 14912
rect 11756 14900 11762 14952
rect 12912 14940 12940 14971
rect 12986 14968 12992 15020
rect 13044 15017 13050 15020
rect 13044 15008 13052 15017
rect 13044 14980 13089 15008
rect 13044 14971 13052 14980
rect 13044 14968 13050 14971
rect 11946 14912 12940 14940
rect 13188 14940 13216 15036
rect 13722 14968 13728 15020
rect 13780 15008 13786 15020
rect 14108 15017 14136 15116
rect 16942 15104 16948 15116
rect 17000 15104 17006 15156
rect 17218 15104 17224 15156
rect 17276 15144 17282 15156
rect 18046 15144 18052 15156
rect 17276 15116 18052 15144
rect 17276 15104 17282 15116
rect 18046 15104 18052 15116
rect 18104 15104 18110 15156
rect 19058 15104 19064 15156
rect 19116 15104 19122 15156
rect 20254 15144 20260 15156
rect 20215 15116 20260 15144
rect 20254 15104 20260 15116
rect 20312 15104 20318 15156
rect 21821 15147 21879 15153
rect 21821 15113 21833 15147
rect 21867 15144 21879 15147
rect 22738 15144 22744 15156
rect 21867 15116 22744 15144
rect 21867 15113 21879 15116
rect 21821 15107 21879 15113
rect 22738 15104 22744 15116
rect 22796 15104 22802 15156
rect 22833 15147 22891 15153
rect 22833 15113 22845 15147
rect 22879 15144 22891 15147
rect 27985 15147 28043 15153
rect 22879 15116 24808 15144
rect 22879 15113 22891 15116
rect 22833 15107 22891 15113
rect 14182 15036 14188 15088
rect 14240 15076 14246 15088
rect 14369 15079 14427 15085
rect 14369 15076 14381 15079
rect 14240 15048 14381 15076
rect 14240 15036 14246 15048
rect 14369 15045 14381 15048
rect 14415 15045 14427 15079
rect 14369 15039 14427 15045
rect 14642 15036 14648 15088
rect 14700 15076 14706 15088
rect 15841 15079 15899 15085
rect 15841 15076 15853 15079
rect 14700 15048 15853 15076
rect 14700 15036 14706 15048
rect 15841 15045 15853 15048
rect 15887 15045 15899 15079
rect 15841 15039 15899 15045
rect 16574 15036 16580 15088
rect 16632 15076 16638 15088
rect 17589 15079 17647 15085
rect 17589 15076 17601 15079
rect 16632 15048 17601 15076
rect 16632 15036 16638 15048
rect 17589 15045 17601 15048
rect 17635 15045 17647 15079
rect 17589 15039 17647 15045
rect 17678 15036 17684 15088
rect 17736 15076 17742 15088
rect 18414 15076 18420 15088
rect 17736 15048 17781 15076
rect 18375 15048 18420 15076
rect 17736 15036 17742 15048
rect 18414 15036 18420 15048
rect 18472 15036 18478 15088
rect 14001 15011 14059 15017
rect 14001 15008 14013 15011
rect 13780 14980 14013 15008
rect 13780 14968 13786 14980
rect 14001 14977 14013 14980
rect 14047 14977 14059 15011
rect 14001 14971 14059 14977
rect 14093 15011 14151 15017
rect 14093 14977 14105 15011
rect 14139 14977 14151 15011
rect 14274 15008 14280 15020
rect 14187 14980 14280 15008
rect 14093 14971 14151 14977
rect 14274 14968 14280 14980
rect 14332 14968 14338 15020
rect 14461 15011 14519 15017
rect 14461 14977 14473 15011
rect 14507 15008 14519 15011
rect 15010 15008 15016 15020
rect 14507 14980 15016 15008
rect 14507 14977 14519 14980
rect 14461 14971 14519 14977
rect 15010 14968 15016 14980
rect 15068 14968 15074 15020
rect 15286 14968 15292 15020
rect 15344 15008 15350 15020
rect 15565 15011 15623 15017
rect 15565 15008 15577 15011
rect 15344 14980 15577 15008
rect 15344 14968 15350 14980
rect 15565 14977 15577 14980
rect 15611 14977 15623 15011
rect 15746 15008 15752 15020
rect 15707 14980 15752 15008
rect 15565 14971 15623 14977
rect 15746 14968 15752 14980
rect 15804 14968 15810 15020
rect 15933 15011 15991 15017
rect 15933 14977 15945 15011
rect 15979 15008 15991 15011
rect 17497 15011 17555 15017
rect 17497 15008 17509 15011
rect 15979 14980 17509 15008
rect 15979 14977 15991 14980
rect 15933 14971 15991 14977
rect 17497 14977 17509 14980
rect 17543 14977 17555 15011
rect 17497 14971 17555 14977
rect 14292 14940 14320 14968
rect 13188 14912 14320 14940
rect 14553 14943 14611 14949
rect 11946 14872 11974 14912
rect 14553 14909 14565 14943
rect 14599 14940 14611 14943
rect 17402 14940 17408 14952
rect 14599 14912 17408 14940
rect 14599 14909 14611 14912
rect 14553 14903 14611 14909
rect 17402 14900 17408 14912
rect 17460 14900 17466 14952
rect 17512 14940 17540 14971
rect 17770 14968 17776 15020
rect 17828 15008 17834 15020
rect 17865 15011 17923 15017
rect 17865 15008 17877 15011
rect 17828 14980 17877 15008
rect 17828 14968 17834 14980
rect 17865 14977 17877 14980
rect 17911 14977 17923 15011
rect 19076 15008 19104 15104
rect 24780 15088 24808 15116
rect 27985 15113 27997 15147
rect 28031 15144 28043 15147
rect 28258 15144 28264 15156
rect 28031 15116 28264 15144
rect 28031 15113 28043 15116
rect 27985 15107 28043 15113
rect 28258 15104 28264 15116
rect 28316 15144 28322 15156
rect 29641 15147 29699 15153
rect 28316 15116 29316 15144
rect 28316 15104 28322 15116
rect 19144 15079 19202 15085
rect 19144 15045 19156 15079
rect 19190 15076 19202 15079
rect 19242 15076 19248 15088
rect 19190 15048 19248 15076
rect 19190 15045 19202 15048
rect 19144 15039 19202 15045
rect 19242 15036 19248 15048
rect 19300 15036 19306 15088
rect 22189 15079 22247 15085
rect 22189 15045 22201 15079
rect 22235 15076 22247 15079
rect 22922 15076 22928 15088
rect 22235 15048 22928 15076
rect 22235 15045 22247 15048
rect 22189 15039 22247 15045
rect 22922 15036 22928 15048
rect 22980 15036 22986 15088
rect 24762 15036 24768 15088
rect 24820 15076 24826 15088
rect 25225 15079 25283 15085
rect 25225 15076 25237 15079
rect 24820 15048 25237 15076
rect 24820 15036 24826 15048
rect 25225 15045 25237 15048
rect 25271 15045 25283 15079
rect 25225 15039 25283 15045
rect 26234 15036 26240 15088
rect 26292 15076 26298 15088
rect 29288 15085 29316 15116
rect 29641 15113 29653 15147
rect 29687 15144 29699 15147
rect 30006 15144 30012 15156
rect 29687 15116 30012 15144
rect 29687 15113 29699 15116
rect 29641 15107 29699 15113
rect 30006 15104 30012 15116
rect 30064 15104 30070 15156
rect 30650 15144 30656 15156
rect 30611 15116 30656 15144
rect 30650 15104 30656 15116
rect 30708 15104 30714 15156
rect 31389 15147 31447 15153
rect 31389 15113 31401 15147
rect 31435 15144 31447 15147
rect 31478 15144 31484 15156
rect 31435 15116 31484 15144
rect 31435 15113 31447 15116
rect 31389 15107 31447 15113
rect 31478 15104 31484 15116
rect 31536 15104 31542 15156
rect 31754 15104 31760 15156
rect 31812 15144 31818 15156
rect 33873 15147 33931 15153
rect 31812 15116 32444 15144
rect 31812 15104 31818 15116
rect 27249 15079 27307 15085
rect 27249 15076 27261 15079
rect 26292 15048 27261 15076
rect 26292 15036 26298 15048
rect 27249 15045 27261 15048
rect 27295 15076 27307 15079
rect 29273 15079 29331 15085
rect 27295 15048 28488 15076
rect 27295 15045 27307 15048
rect 27249 15039 27307 15045
rect 20717 15011 20775 15017
rect 20717 15008 20729 15011
rect 19076 14980 20729 15008
rect 17865 14971 17923 14977
rect 20717 14977 20729 14980
rect 20763 14977 20775 15011
rect 20898 15008 20904 15020
rect 20859 14980 20904 15008
rect 20717 14971 20775 14977
rect 20898 14968 20904 14980
rect 20956 14968 20962 15020
rect 20993 15011 21051 15017
rect 20993 14977 21005 15011
rect 21039 14977 21051 15011
rect 20993 14971 21051 14977
rect 21085 15011 21143 15017
rect 21085 14977 21097 15011
rect 21131 15008 21143 15011
rect 22005 15011 22063 15017
rect 22005 15008 22017 15011
rect 21131 14980 22017 15008
rect 21131 14977 21143 14980
rect 21085 14971 21143 14977
rect 22005 14977 22017 14980
rect 22051 14977 22063 15011
rect 22005 14971 22063 14977
rect 22097 15011 22155 15017
rect 22097 14977 22109 15011
rect 22143 15008 22155 15011
rect 22278 15008 22284 15020
rect 22143 14980 22284 15008
rect 22143 14977 22155 14980
rect 22097 14971 22155 14977
rect 18874 14940 18880 14952
rect 17512 14912 17908 14940
rect 18835 14912 18880 14940
rect 8444 14844 8616 14872
rect 8680 14844 11974 14872
rect 8444 14832 8450 14844
rect 5353 14807 5411 14813
rect 5353 14773 5365 14807
rect 5399 14804 5411 14807
rect 5442 14804 5448 14816
rect 5399 14776 5448 14804
rect 5399 14773 5411 14776
rect 5353 14767 5411 14773
rect 5442 14764 5448 14776
rect 5500 14764 5506 14816
rect 6178 14764 6184 14816
rect 6236 14804 6242 14816
rect 6917 14807 6975 14813
rect 6917 14804 6929 14807
rect 6236 14776 6929 14804
rect 6236 14764 6242 14776
rect 6917 14773 6929 14776
rect 6963 14804 6975 14807
rect 7006 14804 7012 14816
rect 6963 14776 7012 14804
rect 6963 14773 6975 14776
rect 6917 14767 6975 14773
rect 7006 14764 7012 14776
rect 7064 14764 7070 14816
rect 7098 14764 7104 14816
rect 7156 14804 7162 14816
rect 8680 14804 8708 14844
rect 15746 14832 15752 14884
rect 15804 14872 15810 14884
rect 16298 14872 16304 14884
rect 15804 14844 16304 14872
rect 15804 14832 15810 14844
rect 16298 14832 16304 14844
rect 16356 14872 16362 14884
rect 17678 14872 17684 14884
rect 16356 14844 17684 14872
rect 16356 14832 16362 14844
rect 17678 14832 17684 14844
rect 17736 14832 17742 14884
rect 7156 14776 8708 14804
rect 7156 14764 7162 14776
rect 11974 14764 11980 14816
rect 12032 14804 12038 14816
rect 12986 14804 12992 14816
rect 12032 14776 12992 14804
rect 12032 14764 12038 14776
rect 12986 14764 12992 14776
rect 13044 14764 13050 14816
rect 13173 14807 13231 14813
rect 13173 14773 13185 14807
rect 13219 14804 13231 14807
rect 15286 14804 15292 14816
rect 13219 14776 15292 14804
rect 13219 14773 13231 14776
rect 13173 14767 13231 14773
rect 15286 14764 15292 14776
rect 15344 14764 15350 14816
rect 15930 14764 15936 14816
rect 15988 14804 15994 14816
rect 16117 14807 16175 14813
rect 16117 14804 16129 14807
rect 15988 14776 16129 14804
rect 15988 14764 15994 14776
rect 16117 14773 16129 14776
rect 16163 14773 16175 14807
rect 16117 14767 16175 14773
rect 17313 14807 17371 14813
rect 17313 14773 17325 14807
rect 17359 14804 17371 14807
rect 17770 14804 17776 14816
rect 17359 14776 17776 14804
rect 17359 14773 17371 14776
rect 17313 14767 17371 14773
rect 17770 14764 17776 14776
rect 17828 14764 17834 14816
rect 17880 14804 17908 14912
rect 18874 14900 18880 14912
rect 18932 14900 18938 14952
rect 20806 14900 20812 14952
rect 20864 14940 20870 14952
rect 21008 14940 21036 14971
rect 20864 14912 21036 14940
rect 20864 14900 20870 14912
rect 19978 14832 19984 14884
rect 20036 14872 20042 14884
rect 21100 14872 21128 14971
rect 22278 14968 22284 14980
rect 22336 14968 22342 15020
rect 22373 15011 22431 15017
rect 22373 14977 22385 15011
rect 22419 15008 22431 15011
rect 23474 15008 23480 15020
rect 22419 14980 23480 15008
rect 22419 14977 22431 14980
rect 22373 14971 22431 14977
rect 23474 14968 23480 14980
rect 23532 14968 23538 15020
rect 23957 15011 24015 15017
rect 23957 14977 23969 15011
rect 24003 15008 24015 15011
rect 24946 15008 24952 15020
rect 24003 14980 24952 15008
rect 24003 14977 24015 14980
rect 23957 14971 24015 14977
rect 24946 14968 24952 14980
rect 25004 14968 25010 15020
rect 25038 14968 25044 15020
rect 25096 15008 25102 15020
rect 25096 14980 25141 15008
rect 25096 14968 25102 14980
rect 25682 14968 25688 15020
rect 25740 15008 25746 15020
rect 27801 15011 27859 15017
rect 25740 14980 26234 15008
rect 25740 14968 25746 14980
rect 24210 14940 24216 14952
rect 24171 14912 24216 14940
rect 24210 14900 24216 14912
rect 24268 14900 24274 14952
rect 26206 14940 26234 14980
rect 27801 14977 27813 15011
rect 27847 15008 27859 15011
rect 28166 15008 28172 15020
rect 27847 14980 28172 15008
rect 27847 14977 27859 14980
rect 27801 14971 27859 14977
rect 28166 14968 28172 14980
rect 28224 14968 28230 15020
rect 28460 15017 28488 15048
rect 29273 15045 29285 15079
rect 29319 15076 29331 15079
rect 30190 15076 30196 15088
rect 29319 15048 30196 15076
rect 29319 15045 29331 15048
rect 29273 15039 29331 15045
rect 30190 15036 30196 15048
rect 30248 15036 30254 15088
rect 28445 15011 28503 15017
rect 28445 14977 28457 15011
rect 28491 14977 28503 15011
rect 28445 14971 28503 14977
rect 28626 14968 28632 15020
rect 28684 15008 28690 15020
rect 29457 15011 29515 15017
rect 28684 14980 28729 15008
rect 28684 14968 28690 14980
rect 29457 14977 29469 15011
rect 29503 14977 29515 15011
rect 29457 14971 29515 14977
rect 29472 14940 29500 14971
rect 30282 14968 30288 15020
rect 30340 15008 30346 15020
rect 30469 15011 30527 15017
rect 30340 14980 30385 15008
rect 30340 14968 30346 14980
rect 30469 14977 30481 15011
rect 30515 15008 30527 15011
rect 30650 15008 30656 15020
rect 30515 14980 30656 15008
rect 30515 14977 30527 14980
rect 30469 14971 30527 14977
rect 24320 14912 26004 14940
rect 26206 14912 29500 14940
rect 20036 14844 21128 14872
rect 20036 14832 20042 14844
rect 17954 14804 17960 14816
rect 17880 14776 17960 14804
rect 17954 14764 17960 14776
rect 18012 14804 18018 14816
rect 19996 14804 20024 14832
rect 21266 14804 21272 14816
rect 18012 14776 20024 14804
rect 21227 14776 21272 14804
rect 18012 14764 18018 14776
rect 21266 14764 21272 14776
rect 21324 14764 21330 14816
rect 22554 14764 22560 14816
rect 22612 14804 22618 14816
rect 24320 14804 24348 14912
rect 24854 14832 24860 14884
rect 24912 14872 24918 14884
rect 25222 14872 25228 14884
rect 24912 14844 25228 14872
rect 24912 14832 24918 14844
rect 25222 14832 25228 14844
rect 25280 14872 25286 14884
rect 25869 14875 25927 14881
rect 25869 14872 25881 14875
rect 25280 14844 25881 14872
rect 25280 14832 25286 14844
rect 25869 14841 25881 14844
rect 25915 14841 25927 14875
rect 25869 14835 25927 14841
rect 25406 14804 25412 14816
rect 22612 14776 24348 14804
rect 25367 14776 25412 14804
rect 22612 14764 22618 14776
rect 25406 14764 25412 14776
rect 25464 14764 25470 14816
rect 25976 14804 26004 14912
rect 28074 14804 28080 14816
rect 25976 14776 28080 14804
rect 28074 14764 28080 14776
rect 28132 14764 28138 14816
rect 28166 14764 28172 14816
rect 28224 14804 28230 14816
rect 28810 14804 28816 14816
rect 28224 14776 28816 14804
rect 28224 14764 28230 14776
rect 28810 14764 28816 14776
rect 28868 14764 28874 14816
rect 29472 14804 29500 14912
rect 30006 14900 30012 14952
rect 30064 14940 30070 14952
rect 30484 14940 30512 14971
rect 30650 14968 30656 14980
rect 30708 14968 30714 15020
rect 31018 14968 31024 15020
rect 31076 15008 31082 15020
rect 31205 15011 31263 15017
rect 31205 15008 31217 15011
rect 31076 14980 31217 15008
rect 31076 14968 31082 14980
rect 31205 14977 31217 14980
rect 31251 14977 31263 15011
rect 31386 15008 31392 15020
rect 31347 14980 31392 15008
rect 31205 14971 31263 14977
rect 31386 14968 31392 14980
rect 31444 14968 31450 15020
rect 32122 15008 32128 15020
rect 32083 14980 32128 15008
rect 32122 14968 32128 14980
rect 32180 14968 32186 15020
rect 32306 15008 32312 15020
rect 32267 14980 32312 15008
rect 32306 14968 32312 14980
rect 32364 14968 32370 15020
rect 32416 15017 32444 15116
rect 33873 15113 33885 15147
rect 33919 15144 33931 15147
rect 35434 15144 35440 15156
rect 33919 15116 35440 15144
rect 33919 15113 33931 15116
rect 33873 15107 33931 15113
rect 35434 15104 35440 15116
rect 35492 15104 35498 15156
rect 36630 15144 36636 15156
rect 36591 15116 36636 15144
rect 36630 15104 36636 15116
rect 36688 15144 36694 15156
rect 37921 15147 37979 15153
rect 36688 15116 37734 15144
rect 36688 15104 36694 15116
rect 33502 15076 33508 15088
rect 33463 15048 33508 15076
rect 33502 15036 33508 15048
rect 33560 15036 33566 15088
rect 33689 15079 33747 15085
rect 33689 15045 33701 15079
rect 33735 15076 33747 15079
rect 33962 15076 33968 15088
rect 33735 15048 33968 15076
rect 33735 15045 33747 15048
rect 33689 15039 33747 15045
rect 33962 15036 33968 15048
rect 34020 15076 34026 15088
rect 36906 15076 36912 15088
rect 34020 15048 36912 15076
rect 34020 15036 34026 15048
rect 36906 15036 36912 15048
rect 36964 15036 36970 15088
rect 37366 15036 37372 15088
rect 37424 15076 37430 15088
rect 37424 15048 37596 15076
rect 37424 15036 37430 15048
rect 32416 15011 32478 15017
rect 32416 14980 32432 15011
rect 32420 14977 32432 14980
rect 32466 14977 32478 15011
rect 32420 14971 32478 14977
rect 32539 15011 32597 15017
rect 32539 14977 32551 15011
rect 32585 15008 32597 15011
rect 32858 15008 32864 15020
rect 32585 14980 32864 15008
rect 32585 14977 32597 14980
rect 32539 14971 32597 14977
rect 32858 14968 32864 14980
rect 32916 14968 32922 15020
rect 34790 14968 34796 15020
rect 34848 15008 34854 15020
rect 34885 15011 34943 15017
rect 34885 15008 34897 15011
rect 34848 14980 34897 15008
rect 34848 14968 34854 14980
rect 34885 14977 34897 14980
rect 34931 14977 34943 15011
rect 37277 15011 37335 15017
rect 37277 15008 37289 15011
rect 34885 14971 34943 14977
rect 34972 14980 37289 15008
rect 30064 14912 30512 14940
rect 30064 14900 30070 14912
rect 34698 14900 34704 14952
rect 34756 14940 34762 14952
rect 34972 14940 35000 14980
rect 37277 14977 37289 14980
rect 37323 14977 37335 15011
rect 37458 15008 37464 15020
rect 37419 14980 37464 15008
rect 37277 14971 37335 14977
rect 37458 14968 37464 14980
rect 37516 14968 37522 15020
rect 37568 15017 37596 15048
rect 37706 15017 37734 15116
rect 37921 15113 37933 15147
rect 37967 15144 37979 15147
rect 38654 15144 38660 15156
rect 37967 15116 38660 15144
rect 37967 15113 37979 15116
rect 37921 15107 37979 15113
rect 38654 15104 38660 15116
rect 38712 15104 38718 15156
rect 40497 15147 40555 15153
rect 40497 15113 40509 15147
rect 40543 15144 40555 15147
rect 41414 15144 41420 15156
rect 40543 15116 41420 15144
rect 40543 15113 40555 15116
rect 40497 15107 40555 15113
rect 40512 15076 40540 15107
rect 41414 15104 41420 15116
rect 41472 15104 41478 15156
rect 38028 15048 40540 15076
rect 37553 15011 37611 15017
rect 37553 14977 37565 15011
rect 37599 14977 37611 15011
rect 37553 14971 37611 14977
rect 37691 15011 37749 15017
rect 37691 14977 37703 15011
rect 37737 14977 37749 15011
rect 37691 14971 37749 14977
rect 34756 14912 35000 14940
rect 35161 14943 35219 14949
rect 34756 14900 34762 14912
rect 35161 14909 35173 14943
rect 35207 14940 35219 14943
rect 35250 14940 35256 14952
rect 35207 14912 35256 14940
rect 35207 14909 35219 14912
rect 35161 14903 35219 14909
rect 35250 14900 35256 14912
rect 35308 14940 35314 14952
rect 35526 14940 35532 14952
rect 35308 14912 35532 14940
rect 35308 14900 35314 14912
rect 35526 14900 35532 14912
rect 35584 14900 35590 14952
rect 30190 14832 30196 14884
rect 30248 14872 30254 14884
rect 31202 14872 31208 14884
rect 30248 14844 31208 14872
rect 30248 14832 30254 14844
rect 31202 14832 31208 14844
rect 31260 14832 31266 14884
rect 32674 14832 32680 14884
rect 32732 14872 32738 14884
rect 37918 14872 37924 14884
rect 32732 14844 37924 14872
rect 32732 14832 32738 14844
rect 37918 14832 37924 14844
rect 37976 14832 37982 14884
rect 30285 14807 30343 14813
rect 30285 14804 30297 14807
rect 29472 14776 30297 14804
rect 30285 14773 30297 14776
rect 30331 14773 30343 14807
rect 32766 14804 32772 14816
rect 32727 14776 32772 14804
rect 30285 14767 30343 14773
rect 32766 14764 32772 14776
rect 32824 14764 32830 14816
rect 37090 14764 37096 14816
rect 37148 14804 37154 14816
rect 38028 14804 38056 15048
rect 38378 14968 38384 15020
rect 38436 15008 38442 15020
rect 39373 15011 39431 15017
rect 39373 15008 39385 15011
rect 38436 14980 39385 15008
rect 38436 14968 38442 14980
rect 39373 14977 39385 14980
rect 39419 14977 39431 15011
rect 39373 14971 39431 14977
rect 39117 14943 39175 14949
rect 39117 14909 39129 14943
rect 39163 14909 39175 14943
rect 39117 14903 39175 14909
rect 37148 14776 38056 14804
rect 39132 14804 39160 14903
rect 39298 14804 39304 14816
rect 39132 14776 39304 14804
rect 37148 14764 37154 14776
rect 39298 14764 39304 14776
rect 39356 14804 39362 14816
rect 39850 14804 39856 14816
rect 39356 14776 39856 14804
rect 39356 14764 39362 14776
rect 39850 14764 39856 14776
rect 39908 14764 39914 14816
rect 1104 14714 68816 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 65654 14714
rect 65706 14662 65718 14714
rect 65770 14662 65782 14714
rect 65834 14662 65846 14714
rect 65898 14662 65910 14714
rect 65962 14662 68816 14714
rect 1104 14640 68816 14662
rect 2685 14603 2743 14609
rect 2685 14569 2697 14603
rect 2731 14600 2743 14603
rect 2866 14600 2872 14612
rect 2731 14572 2872 14600
rect 2731 14569 2743 14572
rect 2685 14563 2743 14569
rect 2866 14560 2872 14572
rect 2924 14600 2930 14612
rect 3326 14600 3332 14612
rect 2924 14572 3332 14600
rect 2924 14560 2930 14572
rect 3326 14560 3332 14572
rect 3384 14560 3390 14612
rect 8389 14603 8447 14609
rect 8389 14569 8401 14603
rect 8435 14600 8447 14603
rect 8570 14600 8576 14612
rect 8435 14572 8576 14600
rect 8435 14569 8447 14572
rect 8389 14563 8447 14569
rect 8570 14560 8576 14572
rect 8628 14600 8634 14612
rect 8754 14600 8760 14612
rect 8628 14572 8760 14600
rect 8628 14560 8634 14572
rect 8754 14560 8760 14572
rect 8812 14560 8818 14612
rect 9030 14560 9036 14612
rect 9088 14600 9094 14612
rect 12526 14600 12532 14612
rect 9088 14572 12532 14600
rect 9088 14560 9094 14572
rect 12526 14560 12532 14572
rect 12584 14560 12590 14612
rect 13998 14600 14004 14612
rect 12636 14572 14004 14600
rect 11425 14535 11483 14541
rect 11425 14501 11437 14535
rect 11471 14501 11483 14535
rect 11425 14495 11483 14501
rect 12253 14535 12311 14541
rect 12253 14501 12265 14535
rect 12299 14532 12311 14535
rect 12636 14532 12664 14572
rect 13998 14560 14004 14572
rect 14056 14560 14062 14612
rect 14642 14560 14648 14612
rect 14700 14600 14706 14612
rect 15838 14600 15844 14612
rect 14700 14572 15844 14600
rect 14700 14560 14706 14572
rect 15838 14560 15844 14572
rect 15896 14560 15902 14612
rect 16684 14572 17816 14600
rect 16022 14532 16028 14544
rect 12299 14504 12664 14532
rect 14532 14504 16028 14532
rect 12299 14501 12311 14504
rect 12253 14495 12311 14501
rect 7466 14464 7472 14476
rect 5644 14436 7472 14464
rect 5644 14405 5672 14436
rect 7466 14424 7472 14436
rect 7524 14424 7530 14476
rect 10962 14464 10968 14476
rect 9876 14436 10968 14464
rect 2501 14399 2559 14405
rect 2501 14396 2513 14399
rect 2332 14368 2513 14396
rect 2332 14272 2360 14368
rect 2501 14365 2513 14368
rect 2547 14365 2559 14399
rect 2501 14359 2559 14365
rect 5629 14399 5687 14405
rect 5629 14365 5641 14399
rect 5675 14365 5687 14399
rect 5629 14359 5687 14365
rect 5813 14399 5871 14405
rect 5813 14365 5825 14399
rect 5859 14396 5871 14399
rect 7190 14396 7196 14408
rect 5859 14368 7196 14396
rect 5859 14365 5871 14368
rect 5813 14359 5871 14365
rect 7190 14356 7196 14368
rect 7248 14356 7254 14408
rect 7285 14399 7343 14405
rect 7285 14365 7297 14399
rect 7331 14396 7343 14399
rect 7742 14396 7748 14408
rect 7331 14368 7748 14396
rect 7331 14365 7343 14368
rect 7285 14359 7343 14365
rect 7742 14356 7748 14368
rect 7800 14356 7806 14408
rect 9876 14405 9904 14436
rect 10962 14424 10968 14436
rect 11020 14424 11026 14476
rect 11440 14464 11468 14495
rect 11440 14436 14412 14464
rect 9861 14399 9919 14405
rect 9861 14365 9873 14399
rect 9907 14365 9919 14399
rect 10229 14399 10287 14405
rect 9861 14359 9919 14365
rect 9968 14368 10180 14396
rect 5258 14288 5264 14340
rect 5316 14328 5322 14340
rect 5316 14300 6408 14328
rect 5316 14288 5322 14300
rect 2041 14263 2099 14269
rect 2041 14229 2053 14263
rect 2087 14260 2099 14263
rect 2314 14260 2320 14272
rect 2087 14232 2320 14260
rect 2087 14229 2099 14232
rect 2041 14223 2099 14229
rect 2314 14220 2320 14232
rect 2372 14220 2378 14272
rect 5626 14220 5632 14272
rect 5684 14260 5690 14272
rect 6380 14269 6408 14300
rect 9398 14288 9404 14340
rect 9456 14328 9462 14340
rect 9968 14328 9996 14368
rect 10152 14337 10180 14368
rect 10229 14365 10241 14399
rect 10275 14396 10287 14399
rect 10410 14396 10416 14408
rect 10275 14368 10416 14396
rect 10275 14365 10287 14368
rect 10229 14359 10287 14365
rect 10410 14356 10416 14368
rect 10468 14356 10474 14408
rect 10502 14356 10508 14408
rect 10560 14396 10566 14408
rect 10873 14399 10931 14405
rect 10873 14396 10885 14399
rect 10560 14368 10885 14396
rect 10560 14356 10566 14368
rect 10873 14365 10885 14368
rect 10919 14365 10931 14399
rect 11146 14396 11152 14408
rect 11107 14368 11152 14396
rect 10873 14359 10931 14365
rect 11146 14356 11152 14368
rect 11204 14356 11210 14408
rect 11238 14356 11244 14408
rect 11296 14396 11302 14408
rect 12069 14399 12127 14405
rect 11296 14368 11341 14396
rect 11296 14356 11302 14368
rect 12069 14365 12081 14399
rect 12115 14396 12127 14399
rect 12342 14396 12348 14408
rect 12115 14368 12348 14396
rect 12115 14365 12127 14368
rect 12069 14359 12127 14365
rect 12342 14356 12348 14368
rect 12400 14356 12406 14408
rect 12710 14396 12716 14408
rect 12671 14368 12716 14396
rect 12710 14356 12716 14368
rect 12768 14356 12774 14408
rect 14384 14405 14412 14436
rect 14532 14405 14560 14504
rect 16022 14492 16028 14504
rect 16080 14492 16086 14544
rect 16574 14532 16580 14544
rect 16132 14504 16580 14532
rect 16132 14464 16160 14504
rect 16574 14492 16580 14504
rect 16632 14492 16638 14544
rect 16298 14464 16304 14476
rect 14936 14436 16160 14464
rect 16259 14436 16304 14464
rect 14369 14399 14427 14405
rect 14369 14365 14381 14399
rect 14415 14365 14427 14399
rect 14369 14359 14427 14365
rect 14517 14399 14575 14405
rect 14517 14365 14529 14399
rect 14563 14365 14575 14399
rect 14517 14359 14575 14365
rect 14834 14399 14892 14405
rect 14834 14365 14846 14399
rect 14880 14396 14892 14399
rect 14936 14396 14964 14436
rect 16298 14424 16304 14436
rect 16356 14424 16362 14476
rect 16684 14464 16712 14572
rect 17788 14532 17816 14572
rect 17862 14560 17868 14612
rect 17920 14600 17926 14612
rect 20438 14600 20444 14612
rect 17920 14572 20444 14600
rect 17920 14560 17926 14572
rect 20438 14560 20444 14572
rect 20496 14560 20502 14612
rect 23198 14600 23204 14612
rect 23159 14572 23204 14600
rect 23198 14560 23204 14572
rect 23256 14560 23262 14612
rect 24394 14600 24400 14612
rect 24355 14572 24400 14600
rect 24394 14560 24400 14572
rect 24452 14560 24458 14612
rect 28350 14600 28356 14612
rect 25884 14572 28356 14600
rect 19150 14532 19156 14544
rect 17788 14504 19156 14532
rect 19150 14492 19156 14504
rect 19208 14492 19214 14544
rect 19334 14532 19340 14544
rect 19295 14504 19340 14532
rect 19334 14492 19340 14504
rect 19392 14492 19398 14544
rect 23014 14532 23020 14544
rect 19536 14504 23020 14532
rect 16408 14436 16712 14464
rect 16761 14467 16819 14473
rect 14880 14368 14964 14396
rect 14880 14365 14892 14368
rect 14834 14359 14892 14365
rect 9456 14300 9996 14328
rect 10045 14331 10103 14337
rect 9456 14288 9462 14300
rect 10045 14297 10057 14331
rect 10091 14297 10103 14331
rect 10045 14291 10103 14297
rect 10137 14331 10195 14337
rect 10137 14297 10149 14331
rect 10183 14297 10195 14331
rect 11057 14331 11115 14337
rect 11057 14328 11069 14331
rect 10137 14291 10195 14297
rect 10244 14300 11069 14328
rect 5721 14263 5779 14269
rect 5721 14260 5733 14263
rect 5684 14232 5733 14260
rect 5684 14220 5690 14232
rect 5721 14229 5733 14232
rect 5767 14229 5779 14263
rect 5721 14223 5779 14229
rect 6365 14263 6423 14269
rect 6365 14229 6377 14263
rect 6411 14260 6423 14263
rect 9122 14260 9128 14272
rect 6411 14232 9128 14260
rect 6411 14229 6423 14232
rect 6365 14223 6423 14229
rect 9122 14220 9128 14232
rect 9180 14220 9186 14272
rect 10060 14260 10088 14291
rect 10244 14260 10272 14300
rect 11057 14297 11069 14300
rect 11103 14328 11115 14331
rect 11422 14328 11428 14340
rect 11103 14300 11428 14328
rect 11103 14297 11115 14300
rect 11057 14291 11115 14297
rect 11422 14288 11428 14300
rect 11480 14288 11486 14340
rect 14642 14328 14648 14340
rect 14603 14300 14648 14328
rect 14642 14288 14648 14300
rect 14700 14288 14706 14340
rect 14734 14288 14740 14340
rect 14792 14328 14798 14340
rect 14792 14300 14837 14328
rect 14792 14288 14798 14300
rect 10410 14260 10416 14272
rect 10060 14232 10272 14260
rect 10371 14232 10416 14260
rect 10410 14220 10416 14232
rect 10468 14220 10474 14272
rect 11790 14220 11796 14272
rect 11848 14260 11854 14272
rect 12943 14263 13001 14269
rect 12943 14260 12955 14263
rect 11848 14232 12955 14260
rect 11848 14220 11854 14232
rect 12943 14229 12955 14232
rect 12989 14260 13001 14263
rect 13446 14260 13452 14272
rect 12989 14232 13452 14260
rect 12989 14229 13001 14232
rect 12943 14223 13001 14229
rect 13446 14220 13452 14232
rect 13504 14220 13510 14272
rect 13630 14220 13636 14272
rect 13688 14260 13694 14272
rect 14936 14260 14964 14368
rect 15838 14356 15844 14408
rect 15896 14396 15902 14408
rect 16025 14399 16083 14405
rect 16025 14396 16037 14399
rect 15896 14368 16037 14396
rect 15896 14356 15902 14368
rect 16025 14365 16037 14368
rect 16071 14365 16083 14399
rect 16025 14359 16083 14365
rect 13688 14232 14964 14260
rect 15013 14263 15071 14269
rect 13688 14220 13694 14232
rect 15013 14229 15025 14263
rect 15059 14260 15071 14263
rect 16408 14260 16436 14436
rect 16761 14433 16773 14467
rect 16807 14464 16819 14467
rect 17954 14464 17960 14476
rect 16807 14436 17960 14464
rect 16807 14433 16819 14436
rect 16761 14427 16819 14433
rect 17954 14424 17960 14436
rect 18012 14424 18018 14476
rect 16574 14356 16580 14408
rect 16632 14396 16638 14408
rect 17037 14399 17095 14405
rect 17037 14396 17049 14399
rect 16632 14368 17049 14396
rect 16632 14356 16638 14368
rect 17037 14365 17049 14368
rect 17083 14396 17095 14399
rect 17310 14396 17316 14408
rect 17083 14368 17316 14396
rect 17083 14365 17095 14368
rect 17037 14359 17095 14365
rect 17310 14356 17316 14368
rect 17368 14356 17374 14408
rect 19536 14405 19564 14504
rect 23014 14492 23020 14504
rect 23072 14492 23078 14544
rect 20622 14424 20628 14476
rect 20680 14464 20686 14476
rect 21821 14467 21879 14473
rect 21821 14464 21833 14467
rect 20680 14436 21833 14464
rect 20680 14424 20686 14436
rect 21821 14433 21833 14436
rect 21867 14464 21879 14467
rect 22002 14464 22008 14476
rect 21867 14436 22008 14464
rect 21867 14433 21879 14436
rect 21821 14427 21879 14433
rect 22002 14424 22008 14436
rect 22060 14424 22066 14476
rect 25774 14464 25780 14476
rect 25424 14436 25780 14464
rect 18693 14399 18751 14405
rect 18693 14365 18705 14399
rect 18739 14396 18751 14399
rect 19521 14399 19579 14405
rect 19521 14396 19533 14399
rect 18739 14368 19533 14396
rect 18739 14365 18751 14368
rect 18693 14359 18751 14365
rect 19521 14365 19533 14368
rect 19567 14365 19579 14399
rect 19521 14359 19579 14365
rect 20438 14356 20444 14408
rect 20496 14396 20502 14408
rect 20993 14399 21051 14405
rect 20993 14396 21005 14399
rect 20496 14368 21005 14396
rect 20496 14356 20502 14368
rect 20993 14365 21005 14368
rect 21039 14365 21051 14399
rect 20993 14359 21051 14365
rect 21269 14399 21327 14405
rect 21269 14365 21281 14399
rect 21315 14396 21327 14399
rect 21910 14396 21916 14408
rect 21315 14368 21916 14396
rect 21315 14365 21327 14368
rect 21269 14359 21327 14365
rect 21910 14356 21916 14368
rect 21968 14356 21974 14408
rect 25133 14399 25191 14405
rect 25133 14365 25145 14399
rect 25179 14365 25191 14399
rect 25314 14396 25320 14408
rect 25275 14368 25320 14396
rect 25133 14359 25191 14365
rect 17586 14288 17592 14340
rect 17644 14328 17650 14340
rect 20533 14331 20591 14337
rect 20533 14328 20545 14331
rect 17644 14300 20545 14328
rect 17644 14288 17650 14300
rect 20533 14297 20545 14300
rect 20579 14328 20591 14331
rect 20806 14328 20812 14340
rect 20579 14300 20812 14328
rect 20579 14297 20591 14300
rect 20533 14291 20591 14297
rect 20806 14288 20812 14300
rect 20864 14288 20870 14340
rect 21177 14331 21235 14337
rect 21177 14297 21189 14331
rect 21223 14328 21235 14331
rect 22186 14328 22192 14340
rect 21223 14300 22192 14328
rect 21223 14297 21235 14300
rect 21177 14291 21235 14297
rect 22186 14288 22192 14300
rect 22244 14288 22250 14340
rect 25148 14328 25176 14359
rect 25314 14356 25320 14368
rect 25372 14356 25378 14408
rect 25424 14405 25452 14436
rect 25774 14424 25780 14436
rect 25832 14424 25838 14476
rect 25409 14399 25467 14405
rect 25409 14365 25421 14399
rect 25455 14365 25467 14399
rect 25409 14359 25467 14365
rect 25501 14399 25559 14405
rect 25501 14365 25513 14399
rect 25547 14396 25559 14399
rect 25884 14396 25912 14572
rect 28350 14560 28356 14572
rect 28408 14560 28414 14612
rect 30190 14600 30196 14612
rect 30151 14572 30196 14600
rect 30190 14560 30196 14572
rect 30248 14560 30254 14612
rect 30282 14560 30288 14612
rect 30340 14600 30346 14612
rect 30377 14603 30435 14609
rect 30377 14600 30389 14603
rect 30340 14572 30389 14600
rect 30340 14560 30346 14572
rect 30377 14569 30389 14572
rect 30423 14569 30435 14603
rect 30377 14563 30435 14569
rect 31205 14603 31263 14609
rect 31205 14569 31217 14603
rect 31251 14600 31263 14603
rect 32306 14600 32312 14612
rect 31251 14572 32312 14600
rect 31251 14569 31263 14572
rect 31205 14563 31263 14569
rect 32306 14560 32312 14572
rect 32364 14560 32370 14612
rect 33137 14603 33195 14609
rect 33137 14569 33149 14603
rect 33183 14600 33195 14603
rect 33778 14600 33784 14612
rect 33183 14572 33784 14600
rect 33183 14569 33195 14572
rect 33137 14563 33195 14569
rect 33778 14560 33784 14572
rect 33836 14560 33842 14612
rect 38378 14600 38384 14612
rect 38339 14572 38384 14600
rect 38378 14560 38384 14572
rect 38436 14560 38442 14612
rect 28810 14492 28816 14544
rect 28868 14532 28874 14544
rect 28868 14504 32996 14532
rect 28868 14492 28874 14504
rect 28994 14424 29000 14476
rect 29052 14464 29058 14476
rect 30009 14467 30067 14473
rect 30009 14464 30021 14467
rect 29052 14436 30021 14464
rect 29052 14424 29058 14436
rect 30009 14433 30021 14436
rect 30055 14433 30067 14467
rect 30009 14427 30067 14433
rect 30116 14436 31156 14464
rect 26050 14396 26056 14408
rect 25547 14368 26056 14396
rect 25547 14365 25559 14368
rect 25501 14359 25559 14365
rect 26050 14356 26056 14368
rect 26108 14356 26114 14408
rect 26234 14396 26240 14408
rect 26195 14368 26240 14396
rect 26234 14356 26240 14368
rect 26292 14356 26298 14408
rect 30116 14396 30144 14436
rect 26620 14368 30144 14396
rect 30193 14399 30251 14405
rect 25777 14331 25835 14337
rect 25148 14300 25268 14328
rect 21082 14260 21088 14272
rect 15059 14232 16436 14260
rect 21043 14232 21088 14260
rect 15059 14229 15071 14232
rect 15013 14223 15071 14229
rect 21082 14220 21088 14232
rect 21140 14220 21146 14272
rect 22370 14260 22376 14272
rect 22331 14232 22376 14260
rect 22370 14220 22376 14232
rect 22428 14220 22434 14272
rect 25240 14260 25268 14300
rect 25777 14297 25789 14331
rect 25823 14328 25835 14331
rect 26482 14331 26540 14337
rect 26482 14328 26494 14331
rect 25823 14300 26494 14328
rect 25823 14297 25835 14300
rect 25777 14291 25835 14297
rect 26482 14297 26494 14300
rect 26528 14297 26540 14331
rect 26482 14291 26540 14297
rect 25590 14260 25596 14272
rect 25240 14232 25596 14260
rect 25590 14220 25596 14232
rect 25648 14260 25654 14272
rect 26326 14260 26332 14272
rect 25648 14232 26332 14260
rect 25648 14220 25654 14232
rect 26326 14220 26332 14232
rect 26384 14260 26390 14272
rect 26620 14260 26648 14368
rect 30193 14365 30205 14399
rect 30239 14396 30251 14399
rect 31018 14396 31024 14408
rect 30239 14368 31024 14396
rect 30239 14365 30251 14368
rect 30193 14359 30251 14365
rect 31018 14356 31024 14368
rect 31076 14356 31082 14408
rect 31128 14396 31156 14436
rect 31386 14424 31392 14476
rect 31444 14464 31450 14476
rect 31665 14467 31723 14473
rect 31665 14464 31677 14467
rect 31444 14436 31677 14464
rect 31444 14424 31450 14436
rect 31665 14433 31677 14436
rect 31711 14464 31723 14467
rect 32674 14464 32680 14476
rect 31711 14436 32680 14464
rect 31711 14433 31723 14436
rect 31665 14427 31723 14433
rect 32674 14424 32680 14436
rect 32732 14424 32738 14476
rect 32490 14396 32496 14408
rect 31128 14368 32496 14396
rect 32490 14356 32496 14368
rect 32548 14356 32554 14408
rect 32968 14405 32996 14504
rect 37734 14492 37740 14544
rect 37792 14492 37798 14544
rect 35253 14467 35311 14473
rect 35253 14433 35265 14467
rect 35299 14464 35311 14467
rect 35434 14464 35440 14476
rect 35299 14436 35440 14464
rect 35299 14433 35311 14436
rect 35253 14427 35311 14433
rect 35434 14424 35440 14436
rect 35492 14464 35498 14476
rect 37752 14464 37780 14492
rect 38841 14467 38899 14473
rect 38841 14464 38853 14467
rect 35492 14436 37688 14464
rect 37752 14436 38853 14464
rect 35492 14424 35498 14436
rect 37660 14408 37688 14436
rect 32953 14399 33011 14405
rect 32953 14365 32965 14399
rect 32999 14365 33011 14399
rect 35526 14396 35532 14408
rect 35487 14368 35532 14396
rect 32953 14359 33011 14365
rect 35526 14356 35532 14368
rect 35584 14356 35590 14408
rect 37642 14356 37648 14408
rect 37700 14396 37706 14408
rect 38120 14405 38148 14436
rect 38841 14433 38853 14436
rect 38887 14433 38899 14467
rect 38841 14427 38899 14433
rect 37737 14399 37795 14405
rect 37737 14396 37749 14399
rect 37700 14368 37749 14396
rect 37700 14356 37706 14368
rect 37737 14365 37749 14368
rect 37783 14365 37795 14399
rect 37737 14359 37795 14365
rect 37921 14399 37979 14405
rect 37921 14365 37933 14399
rect 37967 14365 37979 14399
rect 37921 14359 37979 14365
rect 38013 14399 38071 14405
rect 38013 14365 38025 14399
rect 38059 14365 38071 14399
rect 38013 14359 38071 14365
rect 38105 14399 38163 14405
rect 38105 14365 38117 14399
rect 38151 14365 38163 14399
rect 68094 14396 68100 14408
rect 68055 14368 68100 14396
rect 38105 14359 38163 14365
rect 27798 14288 27804 14340
rect 27856 14328 27862 14340
rect 28261 14331 28319 14337
rect 28261 14328 28273 14331
rect 27856 14300 28273 14328
rect 27856 14288 27862 14300
rect 28261 14297 28273 14300
rect 28307 14297 28319 14331
rect 29914 14328 29920 14340
rect 29875 14300 29920 14328
rect 28261 14291 28319 14297
rect 29914 14288 29920 14300
rect 29972 14288 29978 14340
rect 30834 14328 30840 14340
rect 30795 14300 30840 14328
rect 30834 14288 30840 14300
rect 30892 14288 30898 14340
rect 33134 14288 33140 14340
rect 33192 14328 33198 14340
rect 33318 14328 33324 14340
rect 33192 14300 33324 14328
rect 33192 14288 33198 14300
rect 33318 14288 33324 14300
rect 33376 14288 33382 14340
rect 34514 14288 34520 14340
rect 34572 14328 34578 14340
rect 36906 14328 36912 14340
rect 34572 14300 36912 14328
rect 34572 14288 34578 14300
rect 36906 14288 36912 14300
rect 36964 14288 36970 14340
rect 37090 14328 37096 14340
rect 37051 14300 37096 14328
rect 37090 14288 37096 14300
rect 37148 14288 37154 14340
rect 37277 14331 37335 14337
rect 37277 14297 37289 14331
rect 37323 14328 37335 14331
rect 37936 14328 37964 14359
rect 37323 14300 37964 14328
rect 37323 14297 37335 14300
rect 37277 14291 37335 14297
rect 26384 14232 26648 14260
rect 26384 14220 26390 14232
rect 27522 14220 27528 14272
rect 27580 14260 27586 14272
rect 27617 14263 27675 14269
rect 27617 14260 27629 14263
rect 27580 14232 27629 14260
rect 27580 14220 27586 14232
rect 27617 14229 27629 14232
rect 27663 14229 27675 14263
rect 28902 14260 28908 14272
rect 28863 14232 28908 14260
rect 27617 14223 27675 14229
rect 28902 14220 28908 14232
rect 28960 14220 28966 14272
rect 37826 14220 37832 14272
rect 37884 14260 37890 14272
rect 38028 14260 38056 14359
rect 68094 14356 68100 14368
rect 68152 14356 68158 14408
rect 37884 14232 38056 14260
rect 37884 14220 37890 14232
rect 1104 14170 68816 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 50294 14170
rect 50346 14118 50358 14170
rect 50410 14118 50422 14170
rect 50474 14118 50486 14170
rect 50538 14118 50550 14170
rect 50602 14118 68816 14170
rect 1104 14096 68816 14118
rect 2682 14056 2688 14068
rect 1596 14028 2688 14056
rect 1596 13929 1624 14028
rect 2682 14016 2688 14028
rect 2740 14056 2746 14068
rect 4985 14059 5043 14065
rect 4985 14056 4997 14059
rect 2740 14028 4997 14056
rect 2740 14016 2746 14028
rect 4985 14025 4997 14028
rect 5031 14056 5043 14059
rect 7098 14056 7104 14068
rect 5031 14028 7104 14056
rect 5031 14025 5043 14028
rect 4985 14019 5043 14025
rect 7098 14016 7104 14028
rect 7156 14016 7162 14068
rect 7742 14056 7748 14068
rect 7703 14028 7748 14056
rect 7742 14016 7748 14028
rect 7800 14016 7806 14068
rect 9030 14056 9036 14068
rect 8991 14028 9036 14056
rect 9030 14016 9036 14028
rect 9088 14016 9094 14068
rect 9122 14016 9128 14068
rect 9180 14056 9186 14068
rect 17586 14056 17592 14068
rect 9180 14028 17592 14056
rect 9180 14016 9186 14028
rect 17586 14016 17592 14028
rect 17644 14016 17650 14068
rect 17681 14059 17739 14065
rect 17681 14025 17693 14059
rect 17727 14056 17739 14059
rect 18322 14056 18328 14068
rect 17727 14028 18328 14056
rect 17727 14025 17739 14028
rect 17681 14019 17739 14025
rect 18322 14016 18328 14028
rect 18380 14016 18386 14068
rect 19886 14056 19892 14068
rect 19847 14028 19892 14056
rect 19886 14016 19892 14028
rect 19944 14016 19950 14068
rect 22186 14016 22192 14068
rect 22244 14056 22250 14068
rect 22373 14059 22431 14065
rect 22373 14056 22385 14059
rect 22244 14028 22385 14056
rect 22244 14016 22250 14028
rect 22373 14025 22385 14028
rect 22419 14056 22431 14059
rect 22554 14056 22560 14068
rect 22419 14028 22560 14056
rect 22419 14025 22431 14028
rect 22373 14019 22431 14025
rect 22554 14016 22560 14028
rect 22612 14016 22618 14068
rect 24946 14056 24952 14068
rect 24907 14028 24952 14056
rect 24946 14016 24952 14028
rect 25004 14016 25010 14068
rect 25314 14016 25320 14068
rect 25372 14056 25378 14068
rect 27433 14059 27491 14065
rect 27433 14056 27445 14059
rect 25372 14028 27445 14056
rect 25372 14016 25378 14028
rect 27433 14025 27445 14028
rect 27479 14025 27491 14059
rect 27433 14019 27491 14025
rect 28997 14059 29055 14065
rect 28997 14025 29009 14059
rect 29043 14056 29055 14059
rect 29086 14056 29092 14068
rect 29043 14028 29092 14056
rect 29043 14025 29055 14028
rect 28997 14019 29055 14025
rect 29086 14016 29092 14028
rect 29144 14016 29150 14068
rect 31018 14016 31024 14068
rect 31076 14056 31082 14068
rect 31662 14056 31668 14068
rect 31076 14028 31668 14056
rect 31076 14016 31082 14028
rect 31662 14016 31668 14028
rect 31720 14056 31726 14068
rect 32125 14059 32183 14065
rect 32125 14056 32137 14059
rect 31720 14028 32137 14056
rect 31720 14016 31726 14028
rect 32125 14025 32137 14028
rect 32171 14025 32183 14059
rect 36725 14059 36783 14065
rect 36725 14056 36737 14059
rect 32125 14019 32183 14025
rect 34716 14028 36737 14056
rect 3050 13988 3056 14000
rect 2792 13960 3056 13988
rect 1581 13923 1639 13929
rect 1581 13889 1593 13923
rect 1627 13889 1639 13923
rect 2498 13920 2504 13932
rect 2459 13892 2504 13920
rect 1581 13883 1639 13889
rect 2498 13880 2504 13892
rect 2556 13880 2562 13932
rect 2792 13929 2820 13960
rect 3050 13948 3056 13960
rect 3108 13948 3114 14000
rect 3145 13991 3203 13997
rect 3145 13957 3157 13991
rect 3191 13988 3203 13991
rect 3850 13991 3908 13997
rect 3850 13988 3862 13991
rect 3191 13960 3862 13988
rect 3191 13957 3203 13960
rect 3145 13951 3203 13957
rect 3850 13957 3862 13960
rect 3896 13957 3908 13991
rect 3850 13951 3908 13957
rect 8754 13948 8760 14000
rect 8812 13988 8818 14000
rect 8812 13960 8857 13988
rect 8812 13948 8818 13960
rect 9582 13948 9588 14000
rect 9640 13988 9646 14000
rect 9640 13960 11836 13988
rect 9640 13948 9646 13960
rect 2685 13923 2743 13929
rect 2685 13889 2697 13923
rect 2731 13889 2743 13923
rect 2685 13883 2743 13889
rect 2777 13923 2835 13929
rect 2777 13889 2789 13923
rect 2823 13889 2835 13923
rect 2777 13883 2835 13889
rect 1486 13852 1492 13864
rect 1447 13824 1492 13852
rect 1486 13812 1492 13824
rect 1544 13812 1550 13864
rect 2700 13852 2728 13883
rect 2866 13880 2872 13932
rect 2924 13920 2930 13932
rect 3602 13920 3608 13932
rect 2924 13892 2969 13920
rect 3563 13892 3608 13920
rect 2924 13880 2930 13892
rect 3602 13880 3608 13892
rect 3660 13880 3666 13932
rect 6086 13880 6092 13932
rect 6144 13920 6150 13932
rect 6621 13923 6679 13929
rect 6621 13920 6633 13923
rect 6144 13892 6633 13920
rect 6144 13880 6150 13892
rect 6621 13889 6633 13892
rect 6667 13889 6679 13923
rect 6621 13883 6679 13889
rect 8294 13880 8300 13932
rect 8352 13920 8358 13932
rect 8662 13929 8668 13932
rect 8481 13923 8539 13929
rect 8481 13920 8493 13923
rect 8352 13892 8493 13920
rect 8352 13880 8358 13892
rect 8481 13889 8493 13892
rect 8527 13889 8539 13923
rect 8481 13883 8539 13889
rect 8619 13923 8668 13929
rect 8619 13889 8631 13923
rect 8665 13889 8668 13923
rect 8619 13883 8668 13889
rect 8662 13880 8668 13883
rect 8720 13880 8726 13932
rect 8846 13920 8852 13932
rect 8807 13892 8852 13920
rect 8846 13880 8852 13892
rect 8904 13920 8910 13932
rect 9398 13920 9404 13932
rect 8904 13892 9404 13920
rect 8904 13880 8910 13892
rect 9398 13880 9404 13892
rect 9456 13920 9462 13932
rect 11808 13929 11836 13960
rect 15838 13948 15844 14000
rect 15896 13988 15902 14000
rect 17313 13991 17371 13997
rect 17313 13988 17325 13991
rect 15896 13960 17325 13988
rect 15896 13948 15902 13960
rect 17313 13957 17325 13960
rect 17359 13957 17371 13991
rect 17313 13951 17371 13957
rect 19150 13948 19156 14000
rect 19208 13988 19214 14000
rect 19429 13991 19487 13997
rect 19429 13988 19441 13991
rect 19208 13960 19441 13988
rect 19208 13948 19214 13960
rect 19429 13957 19441 13960
rect 19475 13957 19487 13991
rect 20898 13988 20904 14000
rect 19429 13951 19487 13957
rect 19536 13960 20904 13988
rect 10045 13923 10103 13929
rect 10045 13920 10057 13923
rect 9456 13892 10057 13920
rect 9456 13880 9462 13892
rect 10045 13889 10057 13892
rect 10091 13889 10103 13923
rect 10045 13883 10103 13889
rect 11793 13923 11851 13929
rect 11793 13889 11805 13923
rect 11839 13889 11851 13923
rect 11793 13883 11851 13889
rect 12986 13880 12992 13932
rect 13044 13920 13050 13932
rect 13357 13923 13415 13929
rect 13357 13920 13369 13923
rect 13044 13892 13369 13920
rect 13044 13880 13050 13892
rect 13357 13889 13369 13892
rect 13403 13889 13415 13923
rect 13357 13883 13415 13889
rect 13446 13880 13452 13932
rect 13504 13920 13510 13932
rect 14093 13923 14151 13929
rect 14093 13920 14105 13923
rect 13504 13892 14105 13920
rect 13504 13880 13510 13892
rect 14093 13889 14105 13892
rect 14139 13889 14151 13923
rect 15470 13920 15476 13932
rect 15431 13892 15476 13920
rect 14093 13883 14151 13889
rect 15470 13880 15476 13892
rect 15528 13880 15534 13932
rect 15657 13923 15715 13929
rect 15657 13889 15669 13923
rect 15703 13920 15715 13923
rect 17034 13920 17040 13932
rect 15703 13892 16896 13920
rect 16995 13892 17040 13920
rect 15703 13889 15715 13892
rect 15657 13883 15715 13889
rect 6362 13852 6368 13864
rect 2700 13824 2820 13852
rect 6323 13824 6368 13852
rect 2792 13784 2820 13824
rect 6362 13812 6368 13824
rect 6420 13812 6426 13864
rect 10318 13852 10324 13864
rect 10231 13824 10324 13852
rect 10318 13812 10324 13824
rect 10376 13852 10382 13864
rect 11238 13852 11244 13864
rect 10376 13824 11244 13852
rect 10376 13812 10382 13824
rect 11238 13812 11244 13824
rect 11296 13812 11302 13864
rect 11514 13852 11520 13864
rect 11475 13824 11520 13852
rect 11514 13812 11520 13824
rect 11572 13812 11578 13864
rect 12802 13812 12808 13864
rect 12860 13852 12866 13864
rect 13630 13852 13636 13864
rect 12860 13824 13636 13852
rect 12860 13812 12866 13824
rect 13630 13812 13636 13824
rect 13688 13812 13694 13864
rect 15289 13855 15347 13861
rect 15289 13821 15301 13855
rect 15335 13852 15347 13855
rect 16390 13852 16396 13864
rect 15335 13824 16396 13852
rect 15335 13821 15347 13824
rect 15289 13815 15347 13821
rect 16390 13812 16396 13824
rect 16448 13812 16454 13864
rect 16868 13852 16896 13892
rect 17034 13880 17040 13892
rect 17092 13880 17098 13932
rect 17218 13929 17224 13932
rect 17185 13923 17224 13929
rect 17185 13889 17197 13923
rect 17185 13883 17224 13889
rect 17218 13880 17224 13883
rect 17276 13880 17282 13932
rect 17402 13920 17408 13932
rect 17363 13892 17408 13920
rect 17402 13880 17408 13892
rect 17460 13880 17466 13932
rect 17494 13880 17500 13932
rect 17552 13929 17558 13932
rect 17552 13920 17560 13929
rect 17552 13892 17597 13920
rect 17552 13883 17560 13892
rect 17552 13880 17558 13883
rect 17678 13880 17684 13932
rect 17736 13920 17742 13932
rect 18141 13923 18199 13929
rect 18141 13920 18153 13923
rect 17736 13892 18153 13920
rect 17736 13880 17742 13892
rect 18141 13889 18153 13892
rect 18187 13889 18199 13923
rect 18141 13883 18199 13889
rect 18325 13923 18383 13929
rect 18325 13889 18337 13923
rect 18371 13920 18383 13923
rect 19536 13920 19564 13960
rect 20898 13948 20904 13960
rect 20956 13948 20962 14000
rect 25774 13988 25780 14000
rect 25332 13960 25780 13988
rect 19702 13920 19708 13932
rect 18371 13892 19564 13920
rect 19663 13892 19708 13920
rect 18371 13889 18383 13892
rect 18325 13883 18383 13889
rect 19702 13880 19708 13892
rect 19760 13880 19766 13932
rect 20254 13880 20260 13932
rect 20312 13920 20318 13932
rect 20349 13923 20407 13929
rect 20349 13920 20361 13923
rect 20312 13892 20361 13920
rect 20312 13880 20318 13892
rect 20349 13889 20361 13892
rect 20395 13920 20407 13923
rect 20714 13920 20720 13932
rect 20395 13892 20720 13920
rect 20395 13889 20407 13892
rect 20349 13883 20407 13889
rect 20714 13880 20720 13892
rect 20772 13880 20778 13932
rect 23753 13923 23811 13929
rect 23753 13920 23765 13923
rect 23124 13892 23765 13920
rect 18509 13855 18567 13861
rect 16868 13824 18460 13852
rect 2866 13784 2872 13796
rect 2792 13756 2872 13784
rect 2866 13744 2872 13756
rect 2924 13744 2930 13796
rect 13262 13744 13268 13796
rect 13320 13784 13326 13796
rect 18046 13784 18052 13796
rect 13320 13756 18052 13784
rect 13320 13744 13326 13756
rect 18046 13744 18052 13756
rect 18104 13744 18110 13796
rect 1857 13719 1915 13725
rect 1857 13685 1869 13719
rect 1903 13716 1915 13719
rect 2774 13716 2780 13728
rect 1903 13688 2780 13716
rect 1903 13685 1915 13688
rect 1857 13679 1915 13685
rect 2774 13676 2780 13688
rect 2832 13676 2838 13728
rect 3602 13676 3608 13728
rect 3660 13716 3666 13728
rect 3786 13716 3792 13728
rect 3660 13688 3792 13716
rect 3660 13676 3666 13688
rect 3786 13676 3792 13688
rect 3844 13676 3850 13728
rect 10686 13676 10692 13728
rect 10744 13716 10750 13728
rect 13814 13716 13820 13728
rect 10744 13688 13820 13716
rect 10744 13676 10750 13688
rect 13814 13676 13820 13688
rect 13872 13676 13878 13728
rect 14277 13719 14335 13725
rect 14277 13685 14289 13719
rect 14323 13716 14335 13719
rect 14366 13716 14372 13728
rect 14323 13688 14372 13716
rect 14323 13685 14335 13688
rect 14277 13679 14335 13685
rect 14366 13676 14372 13688
rect 14424 13676 14430 13728
rect 18432 13716 18460 13824
rect 18509 13821 18521 13855
rect 18555 13852 18567 13855
rect 19426 13852 19432 13864
rect 18555 13824 19432 13852
rect 18555 13821 18567 13824
rect 18509 13815 18567 13821
rect 19426 13812 19432 13824
rect 19484 13812 19490 13864
rect 19613 13855 19671 13861
rect 19613 13821 19625 13855
rect 19659 13852 19671 13855
rect 20530 13852 20536 13864
rect 19659 13824 20536 13852
rect 19659 13821 19671 13824
rect 19613 13815 19671 13821
rect 20530 13812 20536 13824
rect 20588 13812 20594 13864
rect 22830 13852 22836 13864
rect 20640 13824 22836 13852
rect 18966 13744 18972 13796
rect 19024 13784 19030 13796
rect 20640 13784 20668 13824
rect 22830 13812 22836 13824
rect 22888 13852 22894 13864
rect 23124 13861 23152 13892
rect 23753 13889 23765 13892
rect 23799 13889 23811 13923
rect 23753 13883 23811 13889
rect 23937 13923 23995 13929
rect 23937 13889 23949 13923
rect 23983 13920 23995 13923
rect 25130 13920 25136 13932
rect 23983 13892 25136 13920
rect 23983 13889 23995 13892
rect 23937 13883 23995 13889
rect 25130 13880 25136 13892
rect 25188 13929 25194 13932
rect 25332 13929 25360 13960
rect 25774 13948 25780 13960
rect 25832 13948 25838 14000
rect 26050 13988 26056 14000
rect 26011 13960 26056 13988
rect 26050 13948 26056 13960
rect 26108 13948 26114 14000
rect 29270 13988 29276 14000
rect 29231 13960 29276 13988
rect 29270 13948 29276 13960
rect 29328 13948 29334 14000
rect 32766 13948 32772 14000
rect 32824 13988 32830 14000
rect 33238 13991 33296 13997
rect 33238 13988 33250 13991
rect 32824 13960 33250 13988
rect 32824 13948 32830 13960
rect 33238 13957 33250 13960
rect 33284 13957 33296 13991
rect 33238 13951 33296 13957
rect 33502 13948 33508 14000
rect 33560 13988 33566 14000
rect 34514 13988 34520 14000
rect 33560 13960 34520 13988
rect 33560 13948 33566 13960
rect 34514 13948 34520 13960
rect 34572 13948 34578 14000
rect 34716 13932 34744 14028
rect 36725 14025 36737 14028
rect 36771 14056 36783 14059
rect 37366 14056 37372 14068
rect 36771 14028 37372 14056
rect 36771 14025 36783 14028
rect 36725 14019 36783 14025
rect 37366 14016 37372 14028
rect 37424 14016 37430 14068
rect 25188 13923 25237 13929
rect 25188 13889 25191 13923
rect 25225 13889 25237 13923
rect 25188 13883 25237 13889
rect 25314 13923 25372 13929
rect 25314 13889 25326 13923
rect 25360 13889 25372 13923
rect 25314 13883 25372 13889
rect 25188 13880 25194 13883
rect 25406 13880 25412 13932
rect 25464 13929 25470 13932
rect 25464 13920 25472 13929
rect 25464 13892 25509 13920
rect 25464 13883 25472 13892
rect 25464 13880 25470 13883
rect 25590 13880 25596 13932
rect 25648 13920 25654 13932
rect 25648 13892 25693 13920
rect 25648 13880 25654 13892
rect 26142 13880 26148 13932
rect 26200 13920 26206 13932
rect 27065 13923 27123 13929
rect 27065 13920 27077 13923
rect 26200 13892 27077 13920
rect 26200 13880 26206 13892
rect 27065 13889 27077 13892
rect 27111 13889 27123 13923
rect 27065 13883 27123 13889
rect 27249 13923 27307 13929
rect 27249 13889 27261 13923
rect 27295 13920 27307 13923
rect 27522 13920 27528 13932
rect 27295 13892 27528 13920
rect 27295 13889 27307 13892
rect 27249 13883 27307 13889
rect 27522 13880 27528 13892
rect 27580 13880 27586 13932
rect 27798 13880 27804 13932
rect 27856 13920 27862 13932
rect 27985 13923 28043 13929
rect 27985 13920 27997 13923
rect 27856 13892 27997 13920
rect 27856 13880 27862 13892
rect 27985 13889 27997 13892
rect 28031 13889 28043 13923
rect 29178 13920 29184 13932
rect 29139 13892 29184 13920
rect 27985 13883 28043 13889
rect 29178 13880 29184 13892
rect 29236 13880 29242 13932
rect 29365 13923 29423 13929
rect 29365 13889 29377 13923
rect 29411 13889 29423 13923
rect 29546 13920 29552 13932
rect 29507 13892 29552 13920
rect 29365 13883 29423 13889
rect 23109 13855 23167 13861
rect 23109 13852 23121 13855
rect 22888 13824 23121 13852
rect 22888 13812 22894 13824
rect 23109 13821 23121 13824
rect 23155 13821 23167 13855
rect 23109 13815 23167 13821
rect 25774 13812 25780 13864
rect 25832 13852 25838 13864
rect 26786 13852 26792 13864
rect 25832 13824 26792 13852
rect 25832 13812 25838 13824
rect 26786 13812 26792 13824
rect 26844 13812 26850 13864
rect 27614 13852 27620 13864
rect 27527 13824 27620 13852
rect 27586 13812 27620 13824
rect 27672 13852 27678 13864
rect 28166 13852 28172 13864
rect 27672 13824 28172 13852
rect 27672 13812 27678 13824
rect 28166 13812 28172 13824
rect 28224 13812 28230 13864
rect 28534 13812 28540 13864
rect 28592 13852 28598 13864
rect 29380 13852 29408 13883
rect 29546 13880 29552 13892
rect 29604 13880 29610 13932
rect 34698 13920 34704 13932
rect 34659 13892 34704 13920
rect 34698 13880 34704 13892
rect 34756 13880 34762 13932
rect 35342 13920 35348 13932
rect 35303 13892 35348 13920
rect 35342 13880 35348 13892
rect 35400 13880 35406 13932
rect 35618 13929 35624 13932
rect 35612 13883 35624 13929
rect 35676 13920 35682 13932
rect 37642 13920 37648 13932
rect 35676 13892 35712 13920
rect 37603 13892 37648 13920
rect 35618 13880 35624 13883
rect 35676 13880 35682 13892
rect 37642 13880 37648 13892
rect 37700 13880 37706 13932
rect 37808 13926 37866 13932
rect 37808 13923 37820 13926
rect 37798 13892 37820 13923
rect 37854 13892 37866 13926
rect 37798 13886 37866 13892
rect 28592 13824 29408 13852
rect 33505 13855 33563 13861
rect 28592 13812 28598 13824
rect 33505 13821 33517 13855
rect 33551 13852 33563 13855
rect 35360 13852 35388 13880
rect 33551 13824 35388 13852
rect 33551 13821 33563 13824
rect 33505 13815 33563 13821
rect 19024 13756 20668 13784
rect 19024 13744 19030 13756
rect 26234 13744 26240 13796
rect 26292 13784 26298 13796
rect 27246 13784 27252 13796
rect 26292 13756 27252 13784
rect 26292 13744 26298 13756
rect 27246 13744 27252 13756
rect 27304 13784 27310 13796
rect 27586 13784 27614 13812
rect 37798 13796 37826 13886
rect 37918 13880 37924 13932
rect 37976 13920 37982 13932
rect 38059 13923 38117 13929
rect 37976 13892 38021 13920
rect 37976 13880 37982 13892
rect 38059 13889 38071 13923
rect 38105 13920 38117 13923
rect 38194 13920 38200 13932
rect 38105 13892 38200 13920
rect 38105 13889 38117 13892
rect 38059 13883 38117 13889
rect 38194 13880 38200 13892
rect 38252 13880 38258 13932
rect 38289 13855 38347 13861
rect 38289 13821 38301 13855
rect 38335 13852 38347 13855
rect 39942 13852 39948 13864
rect 38335 13824 39948 13852
rect 38335 13821 38347 13824
rect 38289 13815 38347 13821
rect 39942 13812 39948 13824
rect 40000 13812 40006 13864
rect 27304 13756 27614 13784
rect 27304 13744 27310 13756
rect 29086 13744 29092 13796
rect 29144 13784 29150 13796
rect 29822 13784 29828 13796
rect 29144 13756 29828 13784
rect 29144 13744 29150 13756
rect 29822 13744 29828 13756
rect 29880 13744 29886 13796
rect 37734 13744 37740 13796
rect 37792 13756 37826 13796
rect 37792 13744 37798 13756
rect 19610 13716 19616 13728
rect 18432 13688 19616 13716
rect 19610 13676 19616 13688
rect 19668 13676 19674 13728
rect 19705 13719 19763 13725
rect 19705 13685 19717 13719
rect 19751 13716 19763 13719
rect 20254 13716 20260 13728
rect 19751 13688 20260 13716
rect 19751 13685 19763 13688
rect 19705 13679 19763 13685
rect 20254 13676 20260 13688
rect 20312 13676 20318 13728
rect 27522 13676 27528 13728
rect 27580 13716 27586 13728
rect 29638 13716 29644 13728
rect 27580 13688 29644 13716
rect 27580 13676 27586 13688
rect 29638 13676 29644 13688
rect 29696 13676 29702 13728
rect 34790 13676 34796 13728
rect 34848 13716 34854 13728
rect 34885 13719 34943 13725
rect 34885 13716 34897 13719
rect 34848 13688 34897 13716
rect 34848 13676 34854 13688
rect 34885 13685 34897 13688
rect 34931 13685 34943 13719
rect 34885 13679 34943 13685
rect 1104 13626 68816 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 65654 13626
rect 65706 13574 65718 13626
rect 65770 13574 65782 13626
rect 65834 13574 65846 13626
rect 65898 13574 65910 13626
rect 65962 13574 68816 13626
rect 1104 13552 68816 13574
rect 2866 13512 2872 13524
rect 2827 13484 2872 13512
rect 2866 13472 2872 13484
rect 2924 13472 2930 13524
rect 2958 13472 2964 13524
rect 3016 13512 3022 13524
rect 3789 13515 3847 13521
rect 3789 13512 3801 13515
rect 3016 13484 3801 13512
rect 3016 13472 3022 13484
rect 3789 13481 3801 13484
rect 3835 13481 3847 13515
rect 6086 13512 6092 13524
rect 6047 13484 6092 13512
rect 3789 13475 3847 13481
rect 6086 13472 6092 13484
rect 6144 13472 6150 13524
rect 9493 13515 9551 13521
rect 9493 13481 9505 13515
rect 9539 13512 9551 13515
rect 13722 13512 13728 13524
rect 9539 13484 13728 13512
rect 9539 13481 9551 13484
rect 9493 13475 9551 13481
rect 13722 13472 13728 13484
rect 13780 13472 13786 13524
rect 13814 13472 13820 13524
rect 13872 13512 13878 13524
rect 14550 13512 14556 13524
rect 13872 13484 14556 13512
rect 13872 13472 13878 13484
rect 14550 13472 14556 13484
rect 14608 13472 14614 13524
rect 15289 13515 15347 13521
rect 15289 13481 15301 13515
rect 15335 13512 15347 13515
rect 15470 13512 15476 13524
rect 15335 13484 15476 13512
rect 15335 13481 15347 13484
rect 15289 13475 15347 13481
rect 15470 13472 15476 13484
rect 15528 13472 15534 13524
rect 15838 13472 15844 13524
rect 15896 13512 15902 13524
rect 16482 13512 16488 13524
rect 15896 13484 16488 13512
rect 15896 13472 15902 13484
rect 16482 13472 16488 13484
rect 16540 13472 16546 13524
rect 19245 13515 19303 13521
rect 16592 13484 17540 13512
rect 11330 13444 11336 13456
rect 5460 13416 11336 13444
rect 2498 13336 2504 13388
rect 2556 13376 2562 13388
rect 5460 13376 5488 13416
rect 11330 13404 11336 13416
rect 11388 13404 11394 13456
rect 16592 13444 16620 13484
rect 11716 13416 16620 13444
rect 17405 13447 17463 13453
rect 8662 13376 8668 13388
rect 2556 13348 5488 13376
rect 2556 13336 2562 13348
rect 2682 13308 2688 13320
rect 2643 13280 2688 13308
rect 2682 13268 2688 13280
rect 2740 13268 2746 13320
rect 5460 13317 5488 13348
rect 8036 13348 8668 13376
rect 5445 13311 5503 13317
rect 5445 13277 5457 13311
rect 5491 13277 5503 13311
rect 5626 13308 5632 13320
rect 5587 13280 5632 13308
rect 5445 13271 5503 13277
rect 5626 13268 5632 13280
rect 5684 13268 5690 13320
rect 5721 13311 5779 13317
rect 5721 13277 5733 13311
rect 5767 13277 5779 13311
rect 5721 13271 5779 13277
rect 5813 13311 5871 13317
rect 5813 13277 5825 13311
rect 5859 13308 5871 13311
rect 6546 13308 6552 13320
rect 5859 13280 6552 13308
rect 5859 13277 5871 13280
rect 5813 13271 5871 13277
rect 2501 13243 2559 13249
rect 2501 13209 2513 13243
rect 2547 13240 2559 13243
rect 2590 13240 2596 13252
rect 2547 13212 2596 13240
rect 2547 13209 2559 13212
rect 2501 13203 2559 13209
rect 2590 13200 2596 13212
rect 2648 13200 2654 13252
rect 3050 13200 3056 13252
rect 3108 13240 3114 13252
rect 5736 13240 5764 13271
rect 6546 13268 6552 13280
rect 6604 13268 6610 13320
rect 8036 13317 8064 13348
rect 8662 13336 8668 13348
rect 8720 13376 8726 13388
rect 9582 13376 9588 13388
rect 8720 13348 9588 13376
rect 8720 13336 8726 13348
rect 9582 13336 9588 13348
rect 9640 13336 9646 13388
rect 11514 13336 11520 13388
rect 11572 13376 11578 13388
rect 11716 13385 11744 13416
rect 17405 13413 17417 13447
rect 17451 13413 17463 13447
rect 17512 13444 17540 13484
rect 19245 13481 19257 13515
rect 19291 13512 19303 13515
rect 19978 13512 19984 13524
rect 19291 13484 19984 13512
rect 19291 13481 19303 13484
rect 19245 13475 19303 13481
rect 19978 13472 19984 13484
rect 20036 13472 20042 13524
rect 20441 13515 20499 13521
rect 20441 13481 20453 13515
rect 20487 13512 20499 13515
rect 21637 13515 21695 13521
rect 21637 13512 21649 13515
rect 20487 13484 21649 13512
rect 20487 13481 20499 13484
rect 20441 13475 20499 13481
rect 21637 13481 21649 13484
rect 21683 13481 21695 13515
rect 21637 13475 21695 13481
rect 22462 13472 22468 13524
rect 22520 13512 22526 13524
rect 22741 13515 22799 13521
rect 22741 13512 22753 13515
rect 22520 13484 22753 13512
rect 22520 13472 22526 13484
rect 22741 13481 22753 13484
rect 22787 13481 22799 13515
rect 22741 13475 22799 13481
rect 24026 13472 24032 13524
rect 24084 13512 24090 13524
rect 28534 13512 28540 13524
rect 24084 13484 28540 13512
rect 24084 13472 24090 13484
rect 28534 13472 28540 13484
rect 28592 13472 28598 13524
rect 28718 13512 28724 13524
rect 28679 13484 28724 13512
rect 28718 13472 28724 13484
rect 28776 13472 28782 13524
rect 29822 13472 29828 13524
rect 29880 13512 29886 13524
rect 34057 13515 34115 13521
rect 34057 13512 34069 13515
rect 29880 13484 34069 13512
rect 29880 13472 29886 13484
rect 34057 13481 34069 13484
rect 34103 13481 34115 13515
rect 34057 13475 34115 13481
rect 18325 13447 18383 13453
rect 18325 13444 18337 13447
rect 17512 13416 18337 13444
rect 17405 13407 17463 13413
rect 18325 13413 18337 13416
rect 18371 13413 18383 13447
rect 24302 13444 24308 13456
rect 18325 13407 18383 13413
rect 21008 13416 24308 13444
rect 11701 13379 11759 13385
rect 11701 13376 11713 13379
rect 11572 13348 11713 13376
rect 11572 13336 11578 13348
rect 11701 13345 11713 13348
rect 11747 13345 11759 13379
rect 11701 13339 11759 13345
rect 12434 13336 12440 13388
rect 12492 13376 12498 13388
rect 12621 13379 12679 13385
rect 12621 13376 12633 13379
rect 12492 13348 12633 13376
rect 12492 13336 12498 13348
rect 12621 13345 12633 13348
rect 12667 13376 12679 13379
rect 13446 13376 13452 13388
rect 12667 13348 13452 13376
rect 12667 13345 12679 13348
rect 12621 13339 12679 13345
rect 13446 13336 13452 13348
rect 13504 13336 13510 13388
rect 15654 13376 15660 13388
rect 15488 13348 15660 13376
rect 8021 13311 8079 13317
rect 8021 13277 8033 13311
rect 8067 13277 8079 13311
rect 8021 13271 8079 13277
rect 8205 13311 8263 13317
rect 8205 13277 8217 13311
rect 8251 13308 8263 13311
rect 8386 13308 8392 13320
rect 8251 13280 8392 13308
rect 8251 13277 8263 13280
rect 8205 13271 8263 13277
rect 8386 13268 8392 13280
rect 8444 13268 8450 13320
rect 8938 13308 8944 13320
rect 8899 13280 8944 13308
rect 8938 13268 8944 13280
rect 8996 13268 9002 13320
rect 9309 13311 9367 13317
rect 9048 13280 9260 13308
rect 3108 13212 5764 13240
rect 3108 13200 3114 13212
rect 7374 13200 7380 13252
rect 7432 13240 7438 13252
rect 9048 13240 9076 13280
rect 9232 13249 9260 13280
rect 9309 13277 9321 13311
rect 9355 13308 9367 13311
rect 9398 13308 9404 13320
rect 9355 13280 9404 13308
rect 9355 13277 9367 13280
rect 9309 13271 9367 13277
rect 9398 13268 9404 13280
rect 9456 13268 9462 13320
rect 11422 13308 11428 13320
rect 11383 13280 11428 13308
rect 11422 13268 11428 13280
rect 11480 13268 11486 13320
rect 12894 13308 12900 13320
rect 12855 13280 12900 13308
rect 12894 13268 12900 13280
rect 12952 13268 12958 13320
rect 15488 13317 15516 13348
rect 15654 13336 15660 13348
rect 15712 13336 15718 13388
rect 16482 13376 16488 13388
rect 15764 13348 16488 13376
rect 15764 13317 15792 13348
rect 16482 13336 16488 13348
rect 16540 13336 16546 13388
rect 16574 13336 16580 13388
rect 16632 13376 16638 13388
rect 17420 13376 17448 13407
rect 18966 13376 18972 13388
rect 16632 13348 17448 13376
rect 17604 13348 18972 13376
rect 16632 13336 16638 13348
rect 15473 13311 15531 13317
rect 15473 13277 15485 13311
rect 15519 13277 15531 13311
rect 15473 13271 15531 13277
rect 15565 13311 15623 13317
rect 15565 13277 15577 13311
rect 15611 13277 15623 13311
rect 15565 13271 15623 13277
rect 15749 13311 15807 13317
rect 15749 13277 15761 13311
rect 15795 13277 15807 13311
rect 15749 13271 15807 13277
rect 7432 13212 9076 13240
rect 9125 13243 9183 13249
rect 7432 13200 7438 13212
rect 9125 13209 9137 13243
rect 9171 13209 9183 13243
rect 9125 13203 9183 13209
rect 9217 13243 9275 13249
rect 9217 13209 9229 13243
rect 9263 13209 9275 13243
rect 9217 13203 9275 13209
rect 6822 13132 6828 13184
rect 6880 13172 6886 13184
rect 7837 13175 7895 13181
rect 7837 13172 7849 13175
rect 6880 13144 7849 13172
rect 6880 13132 6886 13144
rect 7837 13141 7849 13144
rect 7883 13141 7895 13175
rect 7837 13135 7895 13141
rect 8846 13132 8852 13184
rect 8904 13172 8910 13184
rect 9140 13172 9168 13203
rect 14642 13200 14648 13252
rect 14700 13240 14706 13252
rect 14700 13212 14745 13240
rect 14700 13200 14706 13212
rect 10870 13172 10876 13184
rect 8904 13144 10876 13172
rect 8904 13132 8910 13144
rect 10870 13132 10876 13144
rect 10928 13172 10934 13184
rect 15488 13172 15516 13271
rect 10928 13144 15516 13172
rect 15580 13172 15608 13271
rect 15838 13268 15844 13320
rect 15896 13308 15902 13320
rect 15896 13280 15941 13308
rect 15896 13268 15902 13280
rect 16022 13268 16028 13320
rect 16080 13308 16086 13320
rect 17604 13317 17632 13348
rect 18966 13336 18972 13348
rect 19024 13336 19030 13388
rect 19058 13336 19064 13388
rect 19116 13376 19122 13388
rect 20346 13376 20352 13388
rect 19116 13348 20352 13376
rect 19116 13336 19122 13348
rect 20346 13336 20352 13348
rect 20404 13376 20410 13388
rect 20404 13348 20668 13376
rect 20404 13336 20410 13348
rect 16393 13311 16451 13317
rect 16393 13308 16405 13311
rect 16080 13280 16405 13308
rect 16080 13268 16086 13280
rect 16393 13277 16405 13280
rect 16439 13277 16451 13311
rect 16393 13271 16451 13277
rect 17589 13311 17647 13317
rect 17589 13277 17601 13311
rect 17635 13277 17647 13311
rect 17589 13271 17647 13277
rect 18509 13311 18567 13317
rect 18509 13277 18521 13311
rect 18555 13277 18567 13311
rect 18509 13271 18567 13277
rect 18693 13311 18751 13317
rect 18693 13277 18705 13311
rect 18739 13308 18751 13311
rect 19334 13308 19340 13320
rect 18739 13280 19340 13308
rect 18739 13277 18751 13280
rect 18693 13271 18751 13277
rect 16577 13243 16635 13249
rect 16577 13209 16589 13243
rect 16623 13240 16635 13243
rect 16758 13240 16764 13252
rect 16623 13212 16764 13240
rect 16623 13209 16635 13212
rect 16577 13203 16635 13209
rect 16758 13200 16764 13212
rect 16816 13240 16822 13252
rect 17494 13240 17500 13252
rect 16816 13212 17500 13240
rect 16816 13200 16822 13212
rect 17494 13200 17500 13212
rect 17552 13200 17558 13252
rect 18524 13240 18552 13271
rect 19334 13268 19340 13280
rect 19392 13268 19398 13320
rect 19426 13268 19432 13320
rect 19484 13308 19490 13320
rect 19613 13311 19671 13317
rect 19484 13280 19529 13308
rect 19484 13268 19490 13280
rect 19613 13277 19625 13311
rect 19659 13308 19671 13311
rect 19978 13308 19984 13320
rect 19659 13280 19984 13308
rect 19659 13277 19671 13280
rect 19613 13271 19671 13277
rect 19978 13268 19984 13280
rect 20036 13268 20042 13320
rect 20640 13317 20668 13348
rect 20625 13311 20683 13317
rect 20625 13277 20637 13311
rect 20671 13277 20683 13311
rect 20625 13271 20683 13277
rect 20714 13268 20720 13320
rect 20772 13308 20778 13320
rect 21008 13317 21036 13416
rect 24302 13404 24308 13416
rect 24360 13404 24366 13456
rect 26510 13444 26516 13456
rect 26471 13416 26516 13444
rect 26510 13404 26516 13416
rect 26568 13404 26574 13456
rect 27617 13447 27675 13453
rect 27617 13413 27629 13447
rect 27663 13413 27675 13447
rect 31386 13444 31392 13456
rect 31347 13416 31392 13444
rect 27617 13407 27675 13413
rect 21266 13336 21272 13388
rect 21324 13376 21330 13388
rect 21729 13379 21787 13385
rect 21729 13376 21741 13379
rect 21324 13348 21741 13376
rect 21324 13336 21330 13348
rect 21729 13345 21741 13348
rect 21775 13345 21787 13379
rect 25130 13376 25136 13388
rect 21729 13339 21787 13345
rect 23584 13348 25136 13376
rect 20993 13311 21051 13317
rect 20772 13280 20817 13308
rect 20772 13268 20778 13280
rect 20993 13277 21005 13311
rect 21039 13277 21051 13311
rect 21634 13308 21640 13320
rect 21595 13280 21640 13308
rect 20993 13271 21051 13277
rect 21634 13268 21640 13280
rect 21692 13268 21698 13320
rect 22002 13268 22008 13320
rect 22060 13308 22066 13320
rect 22373 13311 22431 13317
rect 22373 13308 22385 13311
rect 22060 13280 22385 13308
rect 22060 13268 22066 13280
rect 22373 13277 22385 13280
rect 22419 13277 22431 13311
rect 22554 13308 22560 13320
rect 22515 13280 22560 13308
rect 22373 13271 22431 13277
rect 22554 13268 22560 13280
rect 22612 13268 22618 13320
rect 23382 13308 23388 13320
rect 23343 13280 23388 13308
rect 23382 13268 23388 13280
rect 23440 13268 23446 13320
rect 23584 13317 23612 13348
rect 25130 13336 25136 13348
rect 25188 13376 25194 13388
rect 25188 13348 27292 13376
rect 25188 13336 25194 13348
rect 23569 13311 23627 13317
rect 23569 13277 23581 13311
rect 23615 13277 23627 13311
rect 23750 13308 23756 13320
rect 23711 13280 23756 13308
rect 23569 13271 23627 13277
rect 23750 13268 23756 13280
rect 23808 13268 23814 13320
rect 25409 13311 25467 13317
rect 25409 13277 25421 13311
rect 25455 13308 25467 13311
rect 25590 13308 25596 13320
rect 25455 13280 25596 13308
rect 25455 13277 25467 13280
rect 25409 13271 25467 13277
rect 25590 13268 25596 13280
rect 25648 13308 25654 13320
rect 27264 13317 27292 13348
rect 27065 13311 27123 13317
rect 27065 13308 27077 13311
rect 25648 13280 27077 13308
rect 25648 13268 25654 13280
rect 27065 13277 27077 13280
rect 27111 13277 27123 13311
rect 27065 13271 27123 13277
rect 27249 13311 27307 13317
rect 27249 13277 27261 13311
rect 27295 13277 27307 13311
rect 27430 13308 27436 13320
rect 27391 13280 27436 13308
rect 27249 13271 27307 13277
rect 27430 13268 27436 13280
rect 27488 13268 27494 13320
rect 27632 13308 27660 13407
rect 31386 13404 31392 13416
rect 31444 13404 31450 13456
rect 34072 13444 34100 13475
rect 34974 13472 34980 13524
rect 35032 13512 35038 13524
rect 35434 13512 35440 13524
rect 35032 13484 35440 13512
rect 35032 13472 35038 13484
rect 35434 13472 35440 13484
rect 35492 13472 35498 13524
rect 35618 13512 35624 13524
rect 35579 13484 35624 13512
rect 35618 13472 35624 13484
rect 35676 13472 35682 13524
rect 36541 13515 36599 13521
rect 36541 13481 36553 13515
rect 36587 13512 36599 13515
rect 36630 13512 36636 13524
rect 36587 13484 36636 13512
rect 36587 13481 36599 13484
rect 36541 13475 36599 13481
rect 36630 13472 36636 13484
rect 36688 13512 36694 13524
rect 36998 13512 37004 13524
rect 36688 13484 37004 13512
rect 36688 13472 36694 13484
rect 36998 13472 37004 13484
rect 37056 13472 37062 13524
rect 37734 13512 37740 13524
rect 37695 13484 37740 13512
rect 37734 13472 37740 13484
rect 37792 13472 37798 13524
rect 38194 13512 38200 13524
rect 38155 13484 38200 13512
rect 38194 13472 38200 13484
rect 38252 13472 38258 13524
rect 35452 13444 35480 13472
rect 35802 13444 35808 13456
rect 34072 13416 35368 13444
rect 35452 13416 35808 13444
rect 30190 13336 30196 13388
rect 30248 13376 30254 13388
rect 30248 13348 30328 13376
rect 30248 13336 30254 13348
rect 28258 13317 28264 13320
rect 28077 13311 28135 13317
rect 28077 13308 28089 13311
rect 27632 13280 28089 13308
rect 28077 13277 28089 13280
rect 28123 13277 28135 13311
rect 28077 13271 28135 13277
rect 28225 13311 28264 13317
rect 28225 13277 28237 13311
rect 28225 13271 28264 13277
rect 28258 13268 28264 13271
rect 28316 13268 28322 13320
rect 28350 13268 28356 13320
rect 28408 13308 28414 13320
rect 28583 13311 28641 13317
rect 28408 13280 28453 13308
rect 28408 13268 28414 13280
rect 28583 13277 28595 13311
rect 28629 13308 28641 13311
rect 29454 13308 29460 13320
rect 28629 13280 29460 13308
rect 28629 13277 28641 13280
rect 28583 13271 28641 13277
rect 29454 13268 29460 13280
rect 29512 13268 29518 13320
rect 29638 13268 29644 13320
rect 29696 13308 29702 13320
rect 30300 13317 30328 13348
rect 34790 13336 34796 13388
rect 34848 13376 34854 13388
rect 35340 13376 35368 13416
rect 35802 13404 35808 13416
rect 35860 13404 35866 13456
rect 34848 13348 35204 13376
rect 35340 13348 35480 13376
rect 34848 13336 34854 13348
rect 30009 13311 30067 13317
rect 30009 13308 30021 13311
rect 29696 13280 30021 13308
rect 29696 13268 29702 13280
rect 30009 13277 30021 13280
rect 30055 13277 30067 13311
rect 30009 13271 30067 13277
rect 30285 13311 30343 13317
rect 30285 13277 30297 13311
rect 30331 13277 30343 13311
rect 30285 13271 30343 13277
rect 30377 13311 30435 13317
rect 30377 13277 30389 13311
rect 30423 13308 30435 13311
rect 31386 13308 31392 13320
rect 30423 13280 31392 13308
rect 30423 13277 30435 13280
rect 30377 13271 30435 13277
rect 31386 13268 31392 13280
rect 31444 13308 31450 13320
rect 31527 13311 31585 13317
rect 31527 13308 31539 13311
rect 31444 13280 31539 13308
rect 31444 13268 31450 13280
rect 31527 13277 31539 13280
rect 31573 13277 31585 13311
rect 31662 13308 31668 13320
rect 31623 13280 31668 13308
rect 31527 13271 31585 13277
rect 31662 13268 31668 13280
rect 31720 13268 31726 13320
rect 31941 13311 31999 13317
rect 31941 13277 31953 13311
rect 31987 13308 31999 13311
rect 33502 13308 33508 13320
rect 31987 13280 33508 13308
rect 31987 13277 31999 13280
rect 31941 13271 31999 13277
rect 33502 13268 33508 13280
rect 33560 13268 33566 13320
rect 34146 13268 34152 13320
rect 34204 13308 34210 13320
rect 34974 13308 34980 13320
rect 34204 13280 34980 13308
rect 34204 13268 34210 13280
rect 34974 13268 34980 13280
rect 35032 13268 35038 13320
rect 35176 13317 35204 13348
rect 35161 13311 35219 13317
rect 35365 13311 35423 13317
rect 35161 13277 35173 13311
rect 35207 13277 35219 13311
rect 35161 13271 35219 13277
rect 35256 13305 35314 13311
rect 35365 13308 35377 13311
rect 35256 13271 35268 13305
rect 35302 13271 35314 13305
rect 35360 13277 35377 13308
rect 35411 13305 35423 13311
rect 35452 13305 35480 13348
rect 35411 13277 35480 13305
rect 35365 13271 35423 13277
rect 35256 13265 35314 13271
rect 36906 13268 36912 13320
rect 36964 13308 36970 13320
rect 37369 13311 37427 13317
rect 37369 13308 37381 13311
rect 36964 13280 37381 13308
rect 36964 13268 36970 13280
rect 37369 13277 37381 13280
rect 37415 13277 37427 13311
rect 39850 13308 39856 13320
rect 39811 13280 39856 13308
rect 37369 13271 37427 13277
rect 39850 13268 39856 13280
rect 39908 13268 39914 13320
rect 39942 13268 39948 13320
rect 40000 13308 40006 13320
rect 40109 13311 40167 13317
rect 40109 13308 40121 13311
rect 40000 13280 40121 13308
rect 40000 13268 40006 13280
rect 40109 13277 40121 13280
rect 40155 13277 40167 13311
rect 40109 13271 40167 13277
rect 20438 13240 20444 13252
rect 18524 13212 20444 13240
rect 20438 13200 20444 13212
rect 20496 13200 20502 13252
rect 20806 13240 20812 13252
rect 20767 13212 20812 13240
rect 20806 13200 20812 13212
rect 20864 13200 20870 13252
rect 21913 13243 21971 13249
rect 21913 13209 21925 13243
rect 21959 13240 21971 13243
rect 23477 13243 23535 13249
rect 21959 13212 23244 13240
rect 21959 13209 21971 13212
rect 21913 13203 21971 13209
rect 15838 13172 15844 13184
rect 15580 13144 15844 13172
rect 10928 13132 10934 13144
rect 15838 13132 15844 13144
rect 15896 13132 15902 13184
rect 16298 13132 16304 13184
rect 16356 13172 16362 13184
rect 18138 13172 18144 13184
rect 16356 13144 18144 13172
rect 16356 13132 16362 13144
rect 18138 13132 18144 13144
rect 18196 13132 18202 13184
rect 19610 13132 19616 13184
rect 19668 13172 19674 13184
rect 23216 13181 23244 13212
rect 23477 13209 23489 13243
rect 23523 13240 23535 13243
rect 23658 13240 23664 13252
rect 23523 13212 23664 13240
rect 23523 13209 23535 13212
rect 23477 13203 23535 13209
rect 23658 13200 23664 13212
rect 23716 13200 23722 13252
rect 25038 13200 25044 13252
rect 25096 13240 25102 13252
rect 25225 13243 25283 13249
rect 25225 13240 25237 13243
rect 25096 13212 25237 13240
rect 25096 13200 25102 13212
rect 25225 13209 25237 13212
rect 25271 13240 25283 13243
rect 26142 13240 26148 13252
rect 25271 13212 26148 13240
rect 25271 13209 25283 13212
rect 25225 13203 25283 13209
rect 26142 13200 26148 13212
rect 26200 13200 26206 13252
rect 26326 13240 26332 13252
rect 26287 13212 26332 13240
rect 26326 13200 26332 13212
rect 26384 13200 26390 13252
rect 27341 13243 27399 13249
rect 27341 13209 27353 13243
rect 27387 13240 27399 13243
rect 28445 13243 28503 13249
rect 27387 13212 28396 13240
rect 27387 13209 27399 13212
rect 27341 13203 27399 13209
rect 21453 13175 21511 13181
rect 21453 13172 21465 13175
rect 19668 13144 21465 13172
rect 19668 13132 19674 13144
rect 21453 13141 21465 13144
rect 21499 13141 21511 13175
rect 21453 13135 21511 13141
rect 23201 13175 23259 13181
rect 23201 13141 23213 13175
rect 23247 13141 23259 13175
rect 24670 13172 24676 13184
rect 24631 13144 24676 13172
rect 23201 13135 23259 13141
rect 24670 13132 24676 13144
rect 24728 13132 24734 13184
rect 25593 13175 25651 13181
rect 25593 13141 25605 13175
rect 25639 13172 25651 13175
rect 25958 13172 25964 13184
rect 25639 13144 25964 13172
rect 25639 13141 25651 13144
rect 25593 13135 25651 13141
rect 25958 13132 25964 13144
rect 26016 13132 26022 13184
rect 27430 13132 27436 13184
rect 27488 13172 27494 13184
rect 27982 13172 27988 13184
rect 27488 13144 27988 13172
rect 27488 13132 27494 13144
rect 27982 13132 27988 13144
rect 28040 13132 28046 13184
rect 28368 13172 28396 13212
rect 28445 13209 28457 13243
rect 28491 13240 28503 13243
rect 28491 13212 30098 13240
rect 28491 13209 28503 13212
rect 28445 13203 28503 13209
rect 29914 13172 29920 13184
rect 28368 13144 29920 13172
rect 29914 13132 29920 13144
rect 29972 13132 29978 13184
rect 30070 13172 30098 13212
rect 30190 13200 30196 13252
rect 30248 13240 30254 13252
rect 31757 13243 31815 13249
rect 30248 13212 30293 13240
rect 30484 13212 31524 13240
rect 30248 13200 30254 13212
rect 30484 13172 30512 13212
rect 30070 13144 30512 13172
rect 30561 13175 30619 13181
rect 30561 13141 30573 13175
rect 30607 13172 30619 13175
rect 30650 13172 30656 13184
rect 30607 13144 30656 13172
rect 30607 13141 30619 13144
rect 30561 13135 30619 13141
rect 30650 13132 30656 13144
rect 30708 13132 30714 13184
rect 31496 13172 31524 13212
rect 31757 13209 31769 13243
rect 31803 13240 31815 13243
rect 33870 13240 33876 13252
rect 31803 13212 33876 13240
rect 31803 13209 31815 13212
rect 31757 13203 31815 13209
rect 33870 13200 33876 13212
rect 33928 13200 33934 13252
rect 35271 13184 35299 13265
rect 37553 13243 37611 13249
rect 37553 13209 37565 13243
rect 37599 13240 37611 13243
rect 37642 13240 37648 13252
rect 37599 13212 37648 13240
rect 37599 13209 37611 13212
rect 37553 13203 37611 13209
rect 37642 13200 37648 13212
rect 37700 13240 37706 13252
rect 37700 13212 41276 13240
rect 37700 13200 37706 13212
rect 33962 13172 33968 13184
rect 31496 13144 33968 13172
rect 33962 13132 33968 13144
rect 34020 13132 34026 13184
rect 35250 13132 35256 13184
rect 35308 13132 35314 13184
rect 41248 13181 41276 13212
rect 41233 13175 41291 13181
rect 41233 13141 41245 13175
rect 41279 13141 41291 13175
rect 41233 13135 41291 13141
rect 1104 13082 68816 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 50294 13082
rect 50346 13030 50358 13082
rect 50410 13030 50422 13082
rect 50474 13030 50486 13082
rect 50538 13030 50550 13082
rect 50602 13030 68816 13082
rect 1104 13008 68816 13030
rect 4614 12968 4620 12980
rect 2332 12940 4620 12968
rect 1673 12835 1731 12841
rect 1673 12801 1685 12835
rect 1719 12832 1731 12835
rect 2038 12832 2044 12844
rect 1719 12804 2044 12832
rect 1719 12801 1731 12804
rect 1673 12795 1731 12801
rect 2038 12792 2044 12804
rect 2096 12832 2102 12844
rect 2332 12841 2360 12940
rect 4614 12928 4620 12940
rect 4672 12928 4678 12980
rect 10042 12968 10048 12980
rect 9968 12940 10048 12968
rect 2501 12903 2559 12909
rect 2501 12869 2513 12903
rect 2547 12900 2559 12903
rect 2590 12900 2596 12912
rect 2547 12872 2596 12900
rect 2547 12869 2559 12872
rect 2501 12863 2559 12869
rect 2590 12860 2596 12872
rect 2648 12860 2654 12912
rect 3786 12900 3792 12912
rect 3068 12872 3792 12900
rect 3068 12841 3096 12872
rect 3786 12860 3792 12872
rect 3844 12860 3850 12912
rect 7561 12903 7619 12909
rect 7561 12869 7573 12903
rect 7607 12900 7619 12903
rect 8938 12900 8944 12912
rect 7607 12872 8944 12900
rect 7607 12869 7619 12872
rect 7561 12863 7619 12869
rect 8938 12860 8944 12872
rect 8996 12860 9002 12912
rect 9968 12909 9996 12940
rect 10042 12928 10048 12940
rect 10100 12928 10106 12980
rect 10870 12968 10876 12980
rect 10831 12940 10876 12968
rect 10870 12928 10876 12940
rect 10928 12928 10934 12980
rect 11330 12928 11336 12980
rect 11388 12968 11394 12980
rect 11698 12968 11704 12980
rect 11388 12940 11704 12968
rect 11388 12928 11394 12940
rect 11698 12928 11704 12940
rect 11756 12928 11762 12980
rect 12066 12928 12072 12980
rect 12124 12968 12130 12980
rect 13262 12968 13268 12980
rect 12124 12940 13268 12968
rect 12124 12928 12130 12940
rect 13262 12928 13268 12940
rect 13320 12928 13326 12980
rect 15657 12971 15715 12977
rect 15657 12937 15669 12971
rect 15703 12968 15715 12971
rect 17218 12968 17224 12980
rect 15703 12940 17224 12968
rect 15703 12937 15715 12940
rect 15657 12931 15715 12937
rect 17218 12928 17224 12940
rect 17276 12928 17282 12980
rect 18046 12928 18052 12980
rect 18104 12968 18110 12980
rect 18417 12971 18475 12977
rect 18417 12968 18429 12971
rect 18104 12940 18429 12968
rect 18104 12928 18110 12940
rect 18417 12937 18429 12940
rect 18463 12968 18475 12971
rect 18782 12968 18788 12980
rect 18463 12940 18788 12968
rect 18463 12937 18475 12940
rect 18417 12931 18475 12937
rect 18782 12928 18788 12940
rect 18840 12928 18846 12980
rect 18966 12968 18972 12980
rect 18927 12940 18972 12968
rect 18966 12928 18972 12940
rect 19024 12928 19030 12980
rect 20533 12971 20591 12977
rect 20533 12937 20545 12971
rect 20579 12968 20591 12971
rect 20990 12968 20996 12980
rect 20579 12940 20996 12968
rect 20579 12937 20591 12940
rect 20533 12931 20591 12937
rect 20990 12928 20996 12940
rect 21048 12928 21054 12980
rect 21634 12928 21640 12980
rect 21692 12968 21698 12980
rect 21821 12971 21879 12977
rect 21821 12968 21833 12971
rect 21692 12940 21833 12968
rect 21692 12928 21698 12940
rect 21821 12937 21833 12940
rect 21867 12937 21879 12971
rect 21821 12931 21879 12937
rect 21989 12971 22047 12977
rect 21989 12937 22001 12971
rect 22035 12968 22047 12971
rect 22278 12968 22284 12980
rect 22035 12940 22284 12968
rect 22035 12937 22047 12940
rect 21989 12931 22047 12937
rect 22278 12928 22284 12940
rect 22336 12968 22342 12980
rect 22554 12968 22560 12980
rect 22336 12940 22560 12968
rect 22336 12928 22342 12940
rect 22554 12928 22560 12940
rect 22612 12928 22618 12980
rect 25406 12968 25412 12980
rect 23400 12940 25412 12968
rect 9953 12903 10011 12909
rect 9953 12869 9965 12903
rect 9999 12869 10011 12903
rect 11606 12900 11612 12912
rect 11567 12872 11612 12900
rect 9953 12863 10011 12869
rect 11606 12860 11612 12872
rect 11664 12860 11670 12912
rect 18874 12900 18880 12912
rect 13096 12872 16252 12900
rect 2317 12835 2375 12841
rect 2317 12832 2329 12835
rect 2096 12804 2329 12832
rect 2096 12792 2102 12804
rect 2317 12801 2329 12804
rect 2363 12801 2375 12835
rect 2317 12795 2375 12801
rect 3053 12835 3111 12841
rect 3053 12801 3065 12835
rect 3099 12801 3111 12835
rect 3053 12795 3111 12801
rect 3142 12792 3148 12844
rect 3200 12832 3206 12844
rect 3309 12835 3367 12841
rect 3309 12832 3321 12835
rect 3200 12804 3321 12832
rect 3200 12792 3206 12804
rect 3309 12801 3321 12804
rect 3355 12801 3367 12835
rect 7742 12832 7748 12844
rect 7703 12804 7748 12832
rect 3309 12795 3367 12801
rect 7742 12792 7748 12804
rect 7800 12792 7806 12844
rect 9674 12832 9680 12844
rect 9635 12804 9680 12832
rect 9674 12792 9680 12804
rect 9732 12792 9738 12844
rect 9861 12835 9919 12841
rect 9861 12801 9873 12835
rect 9907 12801 9919 12835
rect 9861 12795 9919 12801
rect 10045 12835 10103 12841
rect 10045 12801 10057 12835
rect 10091 12832 10103 12835
rect 10686 12832 10692 12844
rect 10091 12804 10692 12832
rect 10091 12801 10103 12804
rect 10045 12795 10103 12801
rect 9876 12764 9904 12795
rect 10686 12792 10692 12804
rect 10744 12792 10750 12844
rect 10781 12835 10839 12841
rect 10781 12801 10793 12835
rect 10827 12832 10839 12835
rect 11422 12832 11428 12844
rect 10827 12804 11428 12832
rect 10827 12801 10839 12804
rect 10781 12795 10839 12801
rect 10796 12764 10824 12795
rect 11422 12792 11428 12804
rect 11480 12792 11486 12844
rect 12526 12832 12532 12844
rect 12487 12804 12532 12832
rect 12526 12792 12532 12804
rect 12584 12792 12590 12844
rect 13096 12841 13124 12872
rect 16224 12844 16252 12872
rect 17052 12872 18880 12900
rect 13354 12841 13360 12844
rect 13081 12835 13139 12841
rect 13081 12801 13093 12835
rect 13127 12801 13139 12835
rect 13081 12795 13139 12801
rect 13348 12795 13360 12841
rect 13412 12832 13418 12844
rect 15841 12835 15899 12841
rect 13412 12804 13448 12832
rect 13354 12792 13360 12795
rect 13412 12792 13418 12804
rect 15841 12801 15853 12835
rect 15887 12801 15899 12835
rect 16114 12832 16120 12844
rect 16075 12804 16120 12832
rect 15841 12795 15899 12801
rect 9876 12736 10824 12764
rect 10060 12708 10088 12736
rect 4433 12699 4491 12705
rect 4433 12665 4445 12699
rect 4479 12696 4491 12699
rect 4614 12696 4620 12708
rect 4479 12668 4620 12696
rect 4479 12665 4491 12668
rect 4433 12659 4491 12665
rect 4614 12656 4620 12668
rect 4672 12656 4678 12708
rect 6546 12656 6552 12708
rect 6604 12696 6610 12708
rect 6604 12668 9996 12696
rect 6604 12656 6610 12668
rect 2133 12631 2191 12637
rect 2133 12597 2145 12631
rect 2179 12628 2191 12631
rect 2682 12628 2688 12640
rect 2179 12600 2688 12628
rect 2179 12597 2191 12600
rect 2133 12591 2191 12597
rect 2682 12588 2688 12600
rect 2740 12588 2746 12640
rect 7377 12631 7435 12637
rect 7377 12597 7389 12631
rect 7423 12628 7435 12631
rect 7466 12628 7472 12640
rect 7423 12600 7472 12628
rect 7423 12597 7435 12600
rect 7377 12591 7435 12597
rect 7466 12588 7472 12600
rect 7524 12588 7530 12640
rect 8297 12631 8355 12637
rect 8297 12597 8309 12631
rect 8343 12628 8355 12631
rect 8386 12628 8392 12640
rect 8343 12600 8392 12628
rect 8343 12597 8355 12600
rect 8297 12591 8355 12597
rect 8386 12588 8392 12600
rect 8444 12588 8450 12640
rect 9968 12628 9996 12668
rect 10042 12656 10048 12708
rect 10100 12656 10106 12708
rect 10229 12699 10287 12705
rect 10229 12665 10241 12699
rect 10275 12696 10287 12699
rect 15856 12696 15884 12795
rect 16114 12792 16120 12804
rect 16172 12792 16178 12844
rect 16206 12792 16212 12844
rect 16264 12832 16270 12844
rect 17052 12841 17080 12872
rect 18874 12860 18880 12872
rect 18932 12860 18938 12912
rect 22186 12900 22192 12912
rect 22147 12872 22192 12900
rect 22186 12860 22192 12872
rect 22244 12860 22250 12912
rect 23400 12909 23428 12940
rect 25406 12928 25412 12940
rect 25464 12928 25470 12980
rect 25774 12928 25780 12980
rect 25832 12928 25838 12980
rect 26142 12928 26148 12980
rect 26200 12968 26206 12980
rect 34698 12968 34704 12980
rect 26200 12940 34704 12968
rect 26200 12928 26206 12940
rect 34698 12928 34704 12940
rect 34756 12928 34762 12980
rect 36495 12971 36553 12977
rect 36495 12968 36507 12971
rect 36372 12940 36507 12968
rect 23385 12903 23443 12909
rect 23385 12869 23397 12903
rect 23431 12869 23443 12903
rect 23385 12863 23443 12869
rect 23474 12860 23480 12912
rect 23532 12900 23538 12912
rect 23532 12872 23577 12900
rect 23532 12860 23538 12872
rect 17037 12835 17095 12841
rect 17037 12832 17049 12835
rect 16264 12804 17049 12832
rect 16264 12792 16270 12804
rect 17037 12801 17049 12804
rect 17083 12801 17095 12835
rect 17037 12795 17095 12801
rect 17126 12792 17132 12844
rect 17184 12832 17190 12844
rect 17293 12835 17351 12841
rect 17293 12832 17305 12835
rect 17184 12804 17305 12832
rect 17184 12792 17190 12804
rect 17293 12801 17305 12804
rect 17339 12801 17351 12835
rect 17293 12795 17351 12801
rect 19334 12792 19340 12844
rect 19392 12832 19398 12844
rect 20165 12835 20223 12841
rect 20165 12832 20177 12835
rect 19392 12804 20177 12832
rect 19392 12792 19398 12804
rect 20165 12801 20177 12804
rect 20211 12801 20223 12835
rect 20165 12795 20223 12801
rect 20349 12835 20407 12841
rect 20349 12801 20361 12835
rect 20395 12832 20407 12835
rect 20898 12832 20904 12844
rect 20395 12804 20904 12832
rect 20395 12801 20407 12804
rect 20349 12795 20407 12801
rect 20898 12792 20904 12804
rect 20956 12792 20962 12844
rect 23293 12835 23351 12841
rect 23293 12801 23305 12835
rect 23339 12801 23351 12835
rect 23293 12795 23351 12801
rect 16025 12767 16083 12773
rect 16025 12733 16037 12767
rect 16071 12733 16083 12767
rect 16025 12727 16083 12733
rect 10275 12668 13124 12696
rect 10275 12665 10287 12668
rect 10229 12659 10287 12665
rect 12250 12628 12256 12640
rect 9968 12600 12256 12628
rect 12250 12588 12256 12600
rect 12308 12628 12314 12640
rect 12345 12631 12403 12637
rect 12345 12628 12357 12631
rect 12308 12600 12357 12628
rect 12308 12588 12314 12600
rect 12345 12597 12357 12600
rect 12391 12597 12403 12631
rect 13096 12628 13124 12668
rect 14016 12668 15884 12696
rect 14016 12628 14044 12668
rect 14458 12628 14464 12640
rect 13096 12600 14044 12628
rect 14419 12600 14464 12628
rect 12345 12591 12403 12597
rect 14458 12588 14464 12600
rect 14516 12588 14522 12640
rect 14918 12588 14924 12640
rect 14976 12628 14982 12640
rect 15013 12631 15071 12637
rect 15013 12628 15025 12631
rect 14976 12600 15025 12628
rect 14976 12588 14982 12600
rect 15013 12597 15025 12600
rect 15059 12597 15071 12631
rect 15930 12628 15936 12640
rect 15891 12600 15936 12628
rect 15013 12591 15071 12597
rect 15930 12588 15936 12600
rect 15988 12588 15994 12640
rect 16040 12628 16068 12727
rect 23109 12699 23167 12705
rect 23109 12696 23121 12699
rect 18340 12668 23121 12696
rect 18340 12628 18368 12668
rect 23109 12665 23121 12668
rect 23155 12665 23167 12699
rect 23308 12696 23336 12795
rect 23492 12764 23520 12860
rect 25792 12847 25820 12928
rect 25958 12860 25964 12912
rect 26016 12860 26022 12912
rect 26973 12903 27031 12909
rect 26973 12869 26985 12903
rect 27019 12900 27031 12903
rect 27522 12900 27528 12912
rect 27019 12872 27528 12900
rect 27019 12869 27031 12872
rect 26973 12863 27031 12869
rect 27522 12860 27528 12872
rect 27580 12860 27586 12912
rect 29362 12860 29368 12912
rect 29420 12900 29426 12912
rect 30926 12900 30932 12912
rect 29420 12872 30932 12900
rect 29420 12860 29426 12872
rect 30926 12860 30932 12872
rect 30984 12860 30990 12912
rect 31021 12903 31079 12909
rect 31021 12869 31033 12903
rect 31067 12900 31079 12903
rect 33689 12903 33747 12909
rect 31067 12872 33456 12900
rect 31067 12869 31079 12872
rect 31021 12863 31079 12869
rect 23661 12835 23719 12841
rect 23661 12801 23673 12835
rect 23707 12832 23719 12835
rect 23750 12832 23756 12844
rect 23707 12804 23756 12832
rect 23707 12801 23719 12804
rect 23661 12795 23719 12801
rect 23750 12792 23756 12804
rect 23808 12792 23814 12844
rect 24026 12792 24032 12844
rect 24084 12832 24090 12844
rect 25774 12841 25832 12847
rect 24397 12835 24455 12841
rect 24397 12832 24409 12835
rect 24084 12804 24409 12832
rect 24084 12792 24090 12804
rect 24397 12801 24409 12804
rect 24443 12801 24455 12835
rect 24397 12795 24455 12801
rect 25685 12835 25743 12841
rect 25685 12801 25697 12835
rect 25731 12801 25743 12835
rect 25774 12807 25786 12841
rect 25820 12807 25832 12841
rect 25774 12801 25832 12807
rect 25869 12835 25927 12841
rect 25869 12801 25881 12835
rect 25915 12832 25927 12835
rect 25976 12832 26004 12860
rect 25915 12804 26004 12832
rect 26053 12835 26111 12841
rect 25915 12801 25927 12804
rect 25685 12795 25743 12801
rect 25869 12795 25927 12801
rect 26053 12801 26065 12835
rect 26099 12832 26111 12835
rect 26234 12832 26240 12844
rect 26099 12804 26240 12832
rect 26099 12801 26111 12804
rect 26053 12795 26111 12801
rect 24118 12764 24124 12776
rect 23492 12736 24124 12764
rect 24118 12724 24124 12736
rect 24176 12724 24182 12776
rect 25700 12764 25728 12795
rect 26234 12792 26240 12804
rect 26292 12832 26298 12844
rect 26418 12832 26424 12844
rect 26292 12804 26424 12832
rect 26292 12792 26298 12804
rect 26418 12792 26424 12804
rect 26476 12792 26482 12844
rect 27249 12835 27307 12841
rect 27249 12801 27261 12835
rect 27295 12801 27307 12835
rect 27982 12832 27988 12844
rect 27943 12804 27988 12832
rect 27249 12795 27307 12801
rect 26510 12764 26516 12776
rect 25700 12736 26516 12764
rect 26510 12724 26516 12736
rect 26568 12724 26574 12776
rect 27062 12764 27068 12776
rect 27023 12736 27068 12764
rect 27062 12724 27068 12736
rect 27120 12724 27126 12776
rect 27264 12764 27292 12795
rect 27982 12792 27988 12804
rect 28040 12792 28046 12844
rect 28261 12835 28319 12841
rect 28261 12801 28273 12835
rect 28307 12832 28319 12835
rect 28350 12832 28356 12844
rect 28307 12804 28356 12832
rect 28307 12801 28319 12804
rect 28261 12795 28319 12801
rect 28350 12792 28356 12804
rect 28408 12832 28414 12844
rect 28626 12832 28632 12844
rect 28408 12804 28632 12832
rect 28408 12792 28414 12804
rect 28626 12792 28632 12804
rect 28684 12792 28690 12844
rect 29178 12792 29184 12844
rect 29236 12832 29242 12844
rect 29273 12835 29331 12841
rect 29273 12832 29285 12835
rect 29236 12804 29285 12832
rect 29236 12792 29242 12804
rect 29273 12801 29285 12804
rect 29319 12801 29331 12835
rect 29273 12795 29331 12801
rect 29454 12792 29460 12844
rect 29512 12832 29518 12844
rect 29549 12835 29607 12841
rect 29549 12832 29561 12835
rect 29512 12804 29561 12832
rect 29512 12792 29518 12804
rect 29549 12801 29561 12804
rect 29595 12801 29607 12835
rect 30650 12832 30656 12844
rect 30611 12804 30656 12832
rect 29549 12795 29607 12801
rect 30650 12792 30656 12804
rect 30708 12792 30714 12844
rect 30742 12792 30748 12844
rect 30800 12832 30806 12844
rect 30800 12804 30845 12832
rect 30800 12792 30806 12804
rect 31110 12792 31116 12844
rect 31168 12841 31174 12844
rect 31168 12832 31176 12841
rect 33318 12832 33324 12844
rect 31168 12804 31213 12832
rect 33279 12804 33324 12832
rect 31168 12795 31176 12804
rect 31168 12792 31174 12795
rect 33318 12792 33324 12804
rect 33376 12792 33382 12844
rect 29638 12764 29644 12776
rect 27264 12736 29644 12764
rect 29638 12724 29644 12736
rect 29696 12724 29702 12776
rect 23934 12696 23940 12708
rect 23308 12668 23940 12696
rect 23109 12659 23167 12665
rect 23934 12656 23940 12668
rect 23992 12656 23998 12708
rect 33428 12696 33456 12872
rect 33689 12869 33701 12903
rect 33735 12900 33747 12903
rect 35250 12900 35256 12912
rect 33735 12872 34376 12900
rect 33735 12869 33747 12872
rect 33689 12863 33747 12869
rect 33502 12792 33508 12844
rect 33560 12832 33566 12844
rect 34146 12832 34152 12844
rect 33560 12804 33605 12832
rect 34107 12804 34152 12832
rect 33560 12792 33566 12804
rect 34146 12792 34152 12804
rect 34204 12792 34210 12844
rect 34348 12841 34376 12872
rect 34440 12872 35256 12900
rect 34440 12841 34468 12872
rect 35250 12860 35256 12872
rect 35308 12900 35314 12912
rect 35894 12900 35900 12912
rect 35308 12872 35900 12900
rect 35308 12860 35314 12872
rect 35894 12860 35900 12872
rect 35952 12900 35958 12912
rect 36372 12900 36400 12940
rect 36495 12937 36507 12940
rect 36541 12968 36553 12971
rect 37826 12968 37832 12980
rect 36541 12940 37832 12968
rect 36541 12937 36553 12940
rect 36495 12931 36553 12937
rect 37826 12928 37832 12940
rect 37884 12928 37890 12980
rect 37921 12971 37979 12977
rect 37921 12937 37933 12971
rect 37967 12968 37979 12971
rect 38010 12968 38016 12980
rect 37967 12940 38016 12968
rect 37967 12937 37979 12940
rect 37921 12931 37979 12937
rect 38010 12928 38016 12940
rect 38068 12928 38074 12980
rect 41325 12971 41383 12977
rect 41325 12937 41337 12971
rect 41371 12968 41383 12971
rect 41690 12968 41696 12980
rect 41371 12940 41696 12968
rect 41371 12937 41383 12940
rect 41325 12931 41383 12937
rect 41340 12900 41368 12931
rect 41690 12928 41696 12940
rect 41748 12928 41754 12980
rect 35952 12872 36400 12900
rect 36740 12872 40632 12900
rect 35952 12860 35958 12872
rect 36740 12844 36768 12872
rect 34333 12835 34391 12841
rect 34333 12801 34345 12835
rect 34379 12801 34391 12835
rect 34333 12795 34391 12801
rect 34425 12835 34483 12841
rect 34425 12801 34437 12835
rect 34471 12801 34483 12835
rect 34425 12795 34483 12801
rect 34517 12835 34575 12841
rect 34517 12801 34529 12835
rect 34563 12832 34575 12835
rect 34606 12832 34612 12844
rect 34563 12804 34612 12832
rect 34563 12801 34575 12804
rect 34517 12795 34575 12801
rect 34606 12792 34612 12804
rect 34664 12792 34670 12844
rect 36722 12832 36728 12844
rect 36635 12804 36728 12832
rect 36722 12792 36728 12804
rect 36780 12792 36786 12844
rect 37461 12835 37519 12841
rect 37461 12801 37473 12835
rect 37507 12832 37519 12835
rect 37642 12832 37648 12844
rect 37507 12804 37648 12832
rect 37507 12801 37519 12804
rect 37461 12795 37519 12801
rect 37642 12792 37648 12804
rect 37700 12792 37706 12844
rect 37737 12835 37795 12841
rect 37737 12801 37749 12835
rect 37783 12832 37795 12835
rect 37826 12832 37832 12844
rect 37783 12804 37832 12832
rect 37783 12801 37795 12804
rect 37737 12795 37795 12801
rect 37826 12792 37832 12804
rect 37884 12792 37890 12844
rect 40604 12841 40632 12872
rect 40788 12872 41368 12900
rect 40788 12841 40816 12872
rect 40589 12835 40647 12841
rect 40589 12801 40601 12835
rect 40635 12801 40647 12835
rect 40589 12795 40647 12801
rect 40773 12835 40831 12841
rect 40773 12801 40785 12835
rect 40819 12801 40831 12835
rect 41230 12832 41236 12844
rect 41191 12804 41236 12832
rect 40773 12795 40831 12801
rect 41230 12792 41236 12804
rect 41288 12792 41294 12844
rect 33520 12764 33548 12792
rect 36078 12764 36084 12776
rect 33520 12736 36084 12764
rect 36078 12724 36084 12736
rect 36136 12764 36142 12776
rect 37553 12767 37611 12773
rect 37553 12764 37565 12767
rect 36136 12736 37565 12764
rect 36136 12724 36142 12736
rect 37553 12733 37565 12736
rect 37599 12733 37611 12767
rect 37553 12727 37611 12733
rect 37660 12696 37688 12792
rect 67634 12696 67640 12708
rect 33428 12668 37688 12696
rect 67595 12668 67640 12696
rect 67634 12656 67640 12668
rect 67692 12656 67698 12708
rect 16040 12600 18368 12628
rect 19426 12588 19432 12640
rect 19484 12628 19490 12640
rect 20714 12628 20720 12640
rect 19484 12600 20720 12628
rect 19484 12588 19490 12600
rect 20714 12588 20720 12600
rect 20772 12628 20778 12640
rect 22002 12628 22008 12640
rect 20772 12600 22008 12628
rect 20772 12588 20778 12600
rect 22002 12588 22008 12600
rect 22060 12588 22066 12640
rect 24486 12588 24492 12640
rect 24544 12628 24550 12640
rect 25409 12631 25467 12637
rect 25409 12628 25421 12631
rect 24544 12600 25421 12628
rect 24544 12588 24550 12600
rect 25409 12597 25421 12600
rect 25455 12597 25467 12631
rect 25409 12591 25467 12597
rect 25958 12588 25964 12640
rect 26016 12628 26022 12640
rect 26973 12631 27031 12637
rect 26973 12628 26985 12631
rect 26016 12600 26985 12628
rect 26016 12588 26022 12600
rect 26973 12597 26985 12600
rect 27019 12597 27031 12631
rect 26973 12591 27031 12597
rect 27338 12588 27344 12640
rect 27396 12628 27402 12640
rect 27433 12631 27491 12637
rect 27433 12628 27445 12631
rect 27396 12600 27445 12628
rect 27396 12588 27402 12600
rect 27433 12597 27445 12600
rect 27479 12597 27491 12631
rect 27433 12591 27491 12597
rect 29454 12588 29460 12640
rect 29512 12628 29518 12640
rect 29730 12628 29736 12640
rect 29512 12600 29736 12628
rect 29512 12588 29518 12600
rect 29730 12588 29736 12600
rect 29788 12588 29794 12640
rect 31294 12628 31300 12640
rect 31255 12600 31300 12628
rect 31294 12588 31300 12600
rect 31352 12588 31358 12640
rect 34790 12628 34796 12640
rect 34751 12600 34796 12628
rect 34790 12588 34796 12600
rect 34848 12588 34854 12640
rect 37366 12588 37372 12640
rect 37424 12628 37430 12640
rect 37461 12631 37519 12637
rect 37461 12628 37473 12631
rect 37424 12600 37473 12628
rect 37424 12588 37430 12600
rect 37461 12597 37473 12600
rect 37507 12597 37519 12631
rect 38378 12628 38384 12640
rect 38339 12600 38384 12628
rect 37461 12591 37519 12597
rect 38378 12588 38384 12600
rect 38436 12588 38442 12640
rect 38654 12588 38660 12640
rect 38712 12628 38718 12640
rect 40681 12631 40739 12637
rect 40681 12628 40693 12631
rect 38712 12600 40693 12628
rect 38712 12588 38718 12600
rect 40681 12597 40693 12600
rect 40727 12597 40739 12631
rect 40681 12591 40739 12597
rect 1104 12538 68816 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 65654 12538
rect 65706 12486 65718 12538
rect 65770 12486 65782 12538
rect 65834 12486 65846 12538
rect 65898 12486 65910 12538
rect 65962 12486 68816 12538
rect 1104 12464 68816 12486
rect 3142 12424 3148 12436
rect 3103 12396 3148 12424
rect 3142 12384 3148 12396
rect 3200 12384 3206 12436
rect 3694 12384 3700 12436
rect 3752 12424 3758 12436
rect 3789 12427 3847 12433
rect 3789 12424 3801 12427
rect 3752 12396 3801 12424
rect 3752 12384 3758 12396
rect 3789 12393 3801 12396
rect 3835 12393 3847 12427
rect 3789 12387 3847 12393
rect 6362 12384 6368 12436
rect 6420 12424 6426 12436
rect 7098 12424 7104 12436
rect 6420 12396 7104 12424
rect 6420 12384 6426 12396
rect 7098 12384 7104 12396
rect 7156 12384 7162 12436
rect 13262 12424 13268 12436
rect 13223 12396 13268 12424
rect 13262 12384 13268 12396
rect 13320 12384 13326 12436
rect 16485 12427 16543 12433
rect 16485 12393 16497 12427
rect 16531 12424 16543 12427
rect 16666 12424 16672 12436
rect 16531 12396 16672 12424
rect 16531 12393 16543 12396
rect 16485 12387 16543 12393
rect 16666 12384 16672 12396
rect 16724 12384 16730 12436
rect 17770 12424 17776 12436
rect 17731 12396 17776 12424
rect 17770 12384 17776 12396
rect 17828 12384 17834 12436
rect 20806 12384 20812 12436
rect 20864 12424 20870 12436
rect 20901 12427 20959 12433
rect 20901 12424 20913 12427
rect 20864 12396 20913 12424
rect 20864 12384 20870 12396
rect 20901 12393 20913 12396
rect 20947 12393 20959 12427
rect 20901 12387 20959 12393
rect 20990 12384 20996 12436
rect 21048 12424 21054 12436
rect 23753 12427 23811 12433
rect 23753 12424 23765 12427
rect 21048 12396 23765 12424
rect 21048 12384 21054 12396
rect 23753 12393 23765 12396
rect 23799 12393 23811 12427
rect 23753 12387 23811 12393
rect 2041 12359 2099 12365
rect 2041 12325 2053 12359
rect 2087 12356 2099 12359
rect 2087 12328 3188 12356
rect 2087 12325 2099 12328
rect 2041 12319 2099 12325
rect 3050 12288 3056 12300
rect 2792 12260 3056 12288
rect 2498 12220 2504 12232
rect 2459 12192 2504 12220
rect 2498 12180 2504 12192
rect 2556 12180 2562 12232
rect 2682 12220 2688 12232
rect 2643 12192 2688 12220
rect 2682 12180 2688 12192
rect 2740 12180 2746 12232
rect 2792 12229 2820 12260
rect 3050 12248 3056 12260
rect 3108 12248 3114 12300
rect 2777 12223 2835 12229
rect 2777 12189 2789 12223
rect 2823 12189 2835 12223
rect 2777 12183 2835 12189
rect 2869 12223 2927 12229
rect 2869 12189 2881 12223
rect 2915 12220 2927 12223
rect 3160 12220 3188 12328
rect 5810 12316 5816 12368
rect 5868 12356 5874 12368
rect 6822 12356 6828 12368
rect 5868 12328 6828 12356
rect 5868 12316 5874 12328
rect 6822 12316 6828 12328
rect 6880 12316 6886 12368
rect 7650 12316 7656 12368
rect 7708 12356 7714 12368
rect 8386 12356 8392 12368
rect 7708 12328 8392 12356
rect 7708 12316 7714 12328
rect 8386 12316 8392 12328
rect 8444 12316 8450 12368
rect 10413 12359 10471 12365
rect 10413 12325 10425 12359
rect 10459 12356 10471 12359
rect 23768 12356 23796 12387
rect 24670 12384 24676 12436
rect 24728 12424 24734 12436
rect 25130 12424 25136 12436
rect 24728 12396 25136 12424
rect 24728 12384 24734 12396
rect 25130 12384 25136 12396
rect 25188 12424 25194 12436
rect 25866 12424 25872 12436
rect 25188 12396 25872 12424
rect 25188 12384 25194 12396
rect 25866 12384 25872 12396
rect 25924 12384 25930 12436
rect 26510 12424 26516 12436
rect 26471 12396 26516 12424
rect 26510 12384 26516 12396
rect 26568 12384 26574 12436
rect 26878 12384 26884 12436
rect 26936 12424 26942 12436
rect 26973 12427 27031 12433
rect 26973 12424 26985 12427
rect 26936 12396 26985 12424
rect 26936 12384 26942 12396
rect 26973 12393 26985 12396
rect 27019 12393 27031 12427
rect 31386 12424 31392 12436
rect 26973 12387 27031 12393
rect 27632 12396 31392 12424
rect 10459 12328 17632 12356
rect 10459 12325 10471 12328
rect 10413 12319 10471 12325
rect 6914 12288 6920 12300
rect 6564 12260 6920 12288
rect 3694 12220 3700 12232
rect 2915 12192 3700 12220
rect 2915 12189 2927 12192
rect 2869 12183 2927 12189
rect 3694 12180 3700 12192
rect 3752 12180 3758 12232
rect 3786 12180 3792 12232
rect 3844 12220 3850 12232
rect 4341 12223 4399 12229
rect 4341 12220 4353 12223
rect 3844 12192 4353 12220
rect 3844 12180 3850 12192
rect 4341 12189 4353 12192
rect 4387 12220 4399 12223
rect 6362 12220 6368 12232
rect 4387 12192 6368 12220
rect 4387 12189 4399 12192
rect 4341 12183 4399 12189
rect 6362 12180 6368 12192
rect 6420 12180 6426 12232
rect 6564 12229 6592 12260
rect 6914 12248 6920 12260
rect 6972 12288 6978 12300
rect 12345 12291 12403 12297
rect 6972 12260 7604 12288
rect 6972 12248 6978 12260
rect 6457 12223 6515 12229
rect 6457 12189 6469 12223
rect 6503 12189 6515 12223
rect 6457 12183 6515 12189
rect 6549 12223 6607 12229
rect 6549 12189 6561 12223
rect 6595 12189 6607 12223
rect 6549 12183 6607 12189
rect 6641 12223 6699 12229
rect 6641 12189 6653 12223
rect 6687 12220 6699 12223
rect 6730 12220 6736 12232
rect 6687 12192 6736 12220
rect 6687 12189 6699 12192
rect 6641 12183 6699 12189
rect 1857 12155 1915 12161
rect 1857 12121 1869 12155
rect 1903 12152 1915 12155
rect 4608 12155 4666 12161
rect 1903 12124 2360 12152
rect 1903 12121 1915 12124
rect 1857 12115 1915 12121
rect 2332 12084 2360 12124
rect 4608 12121 4620 12155
rect 4654 12152 4666 12155
rect 6181 12155 6239 12161
rect 6181 12152 6193 12155
rect 4654 12124 6193 12152
rect 4654 12121 4666 12124
rect 4608 12115 4666 12121
rect 6181 12121 6193 12124
rect 6227 12121 6239 12155
rect 6181 12115 6239 12121
rect 3142 12084 3148 12096
rect 2332 12056 3148 12084
rect 3142 12044 3148 12056
rect 3200 12044 3206 12096
rect 5718 12084 5724 12096
rect 5679 12056 5724 12084
rect 5718 12044 5724 12056
rect 5776 12044 5782 12096
rect 6472 12084 6500 12183
rect 6730 12180 6736 12192
rect 6788 12180 6794 12232
rect 6822 12180 6828 12232
rect 6880 12220 6886 12232
rect 7285 12223 7343 12229
rect 7285 12220 7297 12223
rect 6880 12192 7297 12220
rect 6880 12180 6886 12192
rect 7285 12189 7297 12192
rect 7331 12189 7343 12223
rect 7466 12220 7472 12232
rect 7427 12192 7472 12220
rect 7285 12183 7343 12189
rect 7466 12180 7472 12192
rect 7524 12180 7530 12232
rect 7576 12229 7604 12260
rect 12345 12257 12357 12291
rect 12391 12288 12403 12291
rect 17126 12288 17132 12300
rect 12391 12260 17132 12288
rect 12391 12257 12403 12260
rect 12345 12251 12403 12257
rect 17126 12248 17132 12260
rect 17184 12248 17190 12300
rect 7561 12223 7619 12229
rect 7561 12189 7573 12223
rect 7607 12189 7619 12223
rect 7561 12183 7619 12189
rect 7650 12180 7656 12232
rect 7708 12220 7714 12232
rect 9858 12220 9864 12232
rect 7708 12192 7753 12220
rect 9819 12192 9864 12220
rect 7708 12180 7714 12192
rect 9858 12180 9864 12192
rect 9916 12180 9922 12232
rect 10042 12220 10048 12232
rect 10003 12192 10048 12220
rect 10042 12180 10048 12192
rect 10100 12180 10106 12232
rect 10229 12223 10287 12229
rect 10229 12189 10241 12223
rect 10275 12220 10287 12223
rect 10318 12220 10324 12232
rect 10275 12192 10324 12220
rect 10275 12189 10287 12192
rect 10229 12183 10287 12189
rect 10318 12180 10324 12192
rect 10376 12180 10382 12232
rect 10873 12223 10931 12229
rect 10873 12189 10885 12223
rect 10919 12220 10931 12223
rect 11330 12220 11336 12232
rect 10919 12192 11336 12220
rect 10919 12189 10931 12192
rect 10873 12183 10931 12189
rect 11330 12180 11336 12192
rect 11388 12180 11394 12232
rect 11698 12220 11704 12232
rect 11659 12192 11704 12220
rect 11698 12180 11704 12192
rect 11756 12180 11762 12232
rect 11885 12223 11943 12229
rect 11885 12189 11897 12223
rect 11931 12189 11943 12223
rect 11885 12183 11943 12189
rect 11977 12223 12035 12229
rect 11977 12189 11989 12223
rect 12023 12189 12035 12223
rect 11977 12183 12035 12189
rect 10134 12152 10140 12164
rect 10095 12124 10140 12152
rect 10134 12112 10140 12124
rect 10192 12112 10198 12164
rect 11054 12152 11060 12164
rect 11015 12124 11060 12152
rect 11054 12112 11060 12124
rect 11112 12112 11118 12164
rect 11241 12155 11299 12161
rect 11241 12121 11253 12155
rect 11287 12152 11299 12155
rect 11900 12152 11928 12183
rect 11287 12124 11928 12152
rect 11992 12152 12020 12183
rect 12066 12180 12072 12232
rect 12124 12220 12130 12232
rect 12989 12223 13047 12229
rect 12124 12192 12169 12220
rect 12124 12180 12130 12192
rect 12989 12189 13001 12223
rect 13035 12189 13047 12223
rect 12989 12183 13047 12189
rect 13081 12223 13139 12229
rect 13081 12189 13093 12223
rect 13127 12220 13139 12223
rect 13814 12220 13820 12232
rect 13127 12192 13820 12220
rect 13127 12189 13139 12192
rect 13081 12183 13139 12189
rect 12250 12152 12256 12164
rect 11992 12124 12256 12152
rect 11287 12121 11299 12124
rect 11241 12115 11299 12121
rect 12250 12112 12256 12124
rect 12308 12112 12314 12164
rect 13004 12152 13032 12183
rect 13814 12180 13820 12192
rect 13872 12220 13878 12232
rect 14458 12220 14464 12232
rect 13872 12192 14464 12220
rect 13872 12180 13878 12192
rect 14458 12180 14464 12192
rect 14516 12180 14522 12232
rect 14645 12223 14703 12229
rect 14645 12189 14657 12223
rect 14691 12220 14703 12223
rect 14734 12220 14740 12232
rect 14691 12192 14740 12220
rect 14691 12189 14703 12192
rect 14645 12183 14703 12189
rect 14734 12180 14740 12192
rect 14792 12180 14798 12232
rect 14918 12220 14924 12232
rect 14879 12192 14924 12220
rect 14918 12180 14924 12192
rect 14976 12180 14982 12232
rect 15102 12180 15108 12232
rect 15160 12220 15166 12232
rect 15381 12223 15439 12229
rect 15381 12220 15393 12223
rect 15160 12192 15393 12220
rect 15160 12180 15166 12192
rect 15381 12189 15393 12192
rect 15427 12189 15439 12223
rect 15381 12183 15439 12189
rect 15470 12180 15476 12232
rect 15528 12220 15534 12232
rect 15654 12220 15660 12232
rect 15528 12192 15573 12220
rect 15615 12192 15660 12220
rect 15528 12180 15534 12192
rect 15654 12180 15660 12192
rect 15712 12180 15718 12232
rect 15746 12180 15752 12232
rect 15804 12220 15810 12232
rect 16669 12223 16727 12229
rect 15804 12192 15849 12220
rect 15804 12180 15810 12192
rect 16669 12189 16681 12223
rect 16715 12220 16727 12223
rect 16758 12220 16764 12232
rect 16715 12192 16764 12220
rect 16715 12189 16727 12192
rect 16669 12183 16727 12189
rect 16758 12180 16764 12192
rect 16816 12180 16822 12232
rect 17604 12229 17632 12328
rect 17880 12328 23612 12356
rect 23768 12328 23888 12356
rect 17589 12223 17647 12229
rect 17589 12189 17601 12223
rect 17635 12189 17647 12223
rect 17589 12183 17647 12189
rect 17678 12180 17684 12232
rect 17736 12220 17742 12232
rect 17880 12229 17908 12328
rect 19426 12248 19432 12300
rect 19484 12288 19490 12300
rect 19978 12288 19984 12300
rect 19484 12260 19984 12288
rect 19484 12248 19490 12260
rect 19978 12248 19984 12260
rect 20036 12248 20042 12300
rect 22922 12248 22928 12300
rect 22980 12288 22986 12300
rect 23017 12291 23075 12297
rect 23017 12288 23029 12291
rect 22980 12260 23029 12288
rect 22980 12248 22986 12260
rect 23017 12257 23029 12260
rect 23063 12288 23075 12291
rect 23474 12288 23480 12300
rect 23063 12260 23480 12288
rect 23063 12257 23075 12260
rect 23017 12251 23075 12257
rect 23474 12248 23480 12260
rect 23532 12248 23538 12300
rect 17865 12223 17923 12229
rect 17736 12192 17781 12220
rect 17736 12180 17742 12192
rect 17865 12189 17877 12223
rect 17911 12189 17923 12223
rect 17865 12183 17923 12189
rect 20254 12180 20260 12232
rect 20312 12220 20318 12232
rect 20533 12223 20591 12229
rect 20533 12220 20545 12223
rect 20312 12192 20545 12220
rect 20312 12180 20318 12192
rect 20533 12189 20545 12192
rect 20579 12189 20591 12223
rect 20533 12183 20591 12189
rect 20717 12223 20775 12229
rect 20717 12189 20729 12223
rect 20763 12220 20775 12223
rect 22186 12220 22192 12232
rect 20763 12192 22192 12220
rect 20763 12189 20775 12192
rect 20717 12183 20775 12189
rect 22186 12180 22192 12192
rect 22244 12180 22250 12232
rect 23584 12220 23612 12328
rect 23860 12220 23888 12328
rect 24578 12316 24584 12368
rect 24636 12356 24642 12368
rect 24762 12356 24768 12368
rect 24636 12328 24768 12356
rect 24636 12316 24642 12328
rect 24762 12316 24768 12328
rect 24820 12316 24826 12368
rect 25406 12356 25412 12368
rect 25367 12328 25412 12356
rect 25406 12316 25412 12328
rect 25464 12316 25470 12368
rect 26602 12316 26608 12368
rect 26660 12356 26666 12368
rect 27632 12356 27660 12396
rect 27982 12356 27988 12368
rect 26660 12328 27660 12356
rect 27724 12328 27988 12356
rect 26660 12316 26666 12328
rect 26234 12248 26240 12300
rect 26292 12288 26298 12300
rect 27724 12288 27752 12328
rect 27982 12316 27988 12328
rect 28040 12316 28046 12368
rect 29454 12288 29460 12300
rect 26292 12260 27752 12288
rect 26292 12248 26298 12260
rect 24397 12223 24455 12229
rect 24397 12220 24409 12223
rect 23584 12192 23704 12220
rect 23860 12192 24409 12220
rect 13265 12155 13323 12161
rect 12406 12124 13124 12152
rect 7190 12084 7196 12096
rect 6472 12056 7196 12084
rect 7190 12044 7196 12056
rect 7248 12044 7254 12096
rect 7929 12087 7987 12093
rect 7929 12053 7941 12087
rect 7975 12084 7987 12087
rect 8018 12084 8024 12096
rect 7975 12056 8024 12084
rect 7975 12053 7987 12056
rect 7929 12047 7987 12053
rect 8018 12044 8024 12056
rect 8076 12044 8082 12096
rect 8294 12044 8300 12096
rect 8352 12084 8358 12096
rect 8941 12087 8999 12093
rect 8941 12084 8953 12087
rect 8352 12056 8953 12084
rect 8352 12044 8358 12056
rect 8941 12053 8953 12056
rect 8987 12053 8999 12087
rect 8941 12047 8999 12053
rect 9950 12044 9956 12096
rect 10008 12084 10014 12096
rect 12406 12084 12434 12124
rect 12802 12084 12808 12096
rect 10008 12056 12434 12084
rect 12763 12056 12808 12084
rect 10008 12044 10014 12056
rect 12802 12044 12808 12056
rect 12860 12044 12866 12096
rect 13096 12084 13124 12124
rect 13265 12121 13277 12155
rect 13311 12152 13323 12155
rect 13630 12152 13636 12164
rect 13311 12124 13636 12152
rect 13311 12121 13323 12124
rect 13265 12115 13323 12121
rect 13630 12112 13636 12124
rect 13688 12112 13694 12164
rect 14550 12112 14556 12164
rect 14608 12152 14614 12164
rect 20990 12152 20996 12164
rect 14608 12124 20996 12152
rect 14608 12112 14614 12124
rect 20990 12112 20996 12124
rect 21048 12112 21054 12164
rect 22094 12112 22100 12164
rect 22152 12152 22158 12164
rect 22833 12155 22891 12161
rect 22833 12152 22845 12155
rect 22152 12124 22845 12152
rect 22152 12112 22158 12124
rect 22833 12121 22845 12124
rect 22879 12121 22891 12155
rect 23676 12152 23704 12192
rect 24397 12189 24409 12192
rect 24443 12189 24455 12223
rect 24578 12220 24584 12232
rect 24539 12192 24584 12220
rect 24397 12183 24455 12189
rect 24578 12180 24584 12192
rect 24636 12180 24642 12232
rect 25130 12180 25136 12232
rect 25188 12220 25194 12232
rect 25593 12223 25651 12229
rect 25593 12220 25605 12223
rect 25188 12192 25605 12220
rect 25188 12180 25194 12192
rect 25593 12189 25605 12192
rect 25639 12189 25651 12223
rect 25593 12183 25651 12189
rect 25682 12180 25688 12232
rect 25740 12220 25746 12232
rect 25961 12223 26019 12229
rect 25740 12192 25785 12220
rect 25740 12180 25746 12192
rect 25961 12189 25973 12223
rect 26007 12214 26019 12223
rect 26050 12214 26056 12232
rect 26007 12189 26056 12214
rect 25961 12186 26056 12189
rect 25961 12183 26019 12186
rect 26050 12180 26056 12186
rect 26108 12180 26114 12232
rect 27724 12229 27752 12260
rect 27816 12260 29460 12288
rect 27816 12229 27844 12260
rect 29454 12248 29460 12260
rect 29512 12248 29518 12300
rect 29822 12288 29828 12300
rect 29656 12260 29828 12288
rect 29656 12232 29684 12260
rect 29822 12248 29828 12260
rect 29880 12248 29886 12300
rect 29932 12288 29960 12396
rect 31386 12384 31392 12396
rect 31444 12384 31450 12436
rect 36078 12424 36084 12436
rect 34624 12396 35940 12424
rect 36039 12396 36084 12424
rect 31110 12316 31116 12368
rect 31168 12356 31174 12368
rect 31168 12328 33088 12356
rect 31168 12316 31174 12328
rect 29932 12260 30052 12288
rect 27709 12223 27767 12229
rect 27709 12189 27721 12223
rect 27755 12189 27767 12223
rect 27709 12183 27767 12189
rect 27801 12223 27859 12229
rect 27801 12189 27813 12223
rect 27847 12189 27859 12223
rect 27801 12183 27859 12189
rect 28077 12223 28135 12229
rect 28077 12189 28089 12223
rect 28123 12220 28135 12223
rect 29638 12220 29644 12232
rect 28123 12192 29500 12220
rect 29599 12192 29644 12220
rect 28123 12189 28135 12192
rect 28077 12183 28135 12189
rect 23676 12124 24624 12152
rect 22833 12115 22891 12121
rect 14826 12084 14832 12096
rect 13096 12056 14832 12084
rect 14826 12044 14832 12056
rect 14884 12044 14890 12096
rect 15746 12044 15752 12096
rect 15804 12084 15810 12096
rect 15933 12087 15991 12093
rect 15933 12084 15945 12087
rect 15804 12056 15945 12084
rect 15804 12044 15810 12056
rect 15933 12053 15945 12056
rect 15979 12053 15991 12087
rect 15933 12047 15991 12053
rect 16666 12044 16672 12096
rect 16724 12084 16730 12096
rect 17405 12087 17463 12093
rect 17405 12084 17417 12087
rect 16724 12056 17417 12084
rect 16724 12044 16730 12056
rect 17405 12053 17417 12056
rect 17451 12053 17463 12087
rect 17405 12047 17463 12053
rect 17862 12044 17868 12096
rect 17920 12084 17926 12096
rect 18325 12087 18383 12093
rect 18325 12084 18337 12087
rect 17920 12056 18337 12084
rect 17920 12044 17926 12056
rect 18325 12053 18337 12056
rect 18371 12053 18383 12087
rect 18325 12047 18383 12053
rect 20438 12044 20444 12096
rect 20496 12084 20502 12096
rect 20714 12084 20720 12096
rect 20496 12056 20720 12084
rect 20496 12044 20502 12056
rect 20714 12044 20720 12056
rect 20772 12044 20778 12096
rect 22189 12087 22247 12093
rect 22189 12053 22201 12087
rect 22235 12084 22247 12087
rect 22922 12084 22928 12096
rect 22235 12056 22928 12084
rect 22235 12053 22247 12056
rect 22189 12047 22247 12053
rect 22922 12044 22928 12056
rect 22980 12044 22986 12096
rect 24394 12084 24400 12096
rect 24355 12056 24400 12084
rect 24394 12044 24400 12056
rect 24452 12044 24458 12096
rect 24596 12084 24624 12124
rect 25406 12112 25412 12164
rect 25464 12152 25470 12164
rect 25777 12155 25835 12161
rect 25777 12152 25789 12155
rect 25464 12124 25789 12152
rect 25464 12112 25470 12124
rect 25777 12121 25789 12124
rect 25823 12121 25835 12155
rect 25777 12115 25835 12121
rect 25866 12112 25872 12164
rect 25924 12152 25930 12164
rect 27893 12155 27951 12161
rect 27893 12152 27905 12155
rect 25924 12124 27905 12152
rect 25924 12112 25930 12124
rect 27893 12121 27905 12124
rect 27939 12152 27951 12155
rect 27982 12152 27988 12164
rect 27939 12124 27988 12152
rect 27939 12121 27951 12124
rect 27893 12115 27951 12121
rect 27982 12112 27988 12124
rect 28040 12112 28046 12164
rect 28626 12152 28632 12164
rect 28587 12124 28632 12152
rect 28626 12112 28632 12124
rect 28684 12112 28690 12164
rect 29472 12152 29500 12192
rect 29638 12180 29644 12192
rect 29696 12180 29702 12232
rect 29914 12220 29920 12232
rect 29875 12192 29920 12220
rect 29914 12180 29920 12192
rect 29972 12180 29978 12232
rect 30024 12229 30052 12260
rect 30926 12248 30932 12300
rect 30984 12288 30990 12300
rect 32490 12288 32496 12300
rect 30984 12260 32496 12288
rect 30984 12248 30990 12260
rect 32490 12248 32496 12260
rect 32548 12288 32554 12300
rect 33060 12297 33088 12328
rect 33045 12291 33103 12297
rect 32548 12260 32812 12288
rect 32548 12248 32554 12260
rect 30009 12223 30067 12229
rect 30009 12189 30021 12223
rect 30055 12189 30067 12223
rect 30009 12183 30067 12189
rect 30190 12180 30196 12232
rect 30248 12180 30254 12232
rect 31294 12220 31300 12232
rect 31255 12192 31300 12220
rect 31294 12180 31300 12192
rect 31352 12180 31358 12232
rect 31386 12180 31392 12232
rect 31444 12220 31450 12232
rect 31665 12223 31723 12229
rect 31665 12222 31677 12223
rect 31588 12220 31677 12222
rect 31444 12194 31677 12220
rect 31444 12192 31616 12194
rect 31444 12180 31450 12192
rect 31665 12189 31677 12194
rect 31711 12189 31723 12223
rect 31665 12183 31723 12189
rect 32122 12180 32128 12232
rect 32180 12220 32186 12232
rect 32309 12223 32367 12229
rect 32309 12220 32321 12223
rect 32180 12192 32321 12220
rect 32180 12180 32186 12192
rect 32309 12189 32321 12192
rect 32355 12189 32367 12223
rect 32309 12183 32367 12189
rect 32585 12223 32643 12229
rect 32585 12189 32597 12223
rect 32631 12220 32643 12223
rect 32674 12220 32680 12232
rect 32631 12192 32680 12220
rect 32631 12189 32643 12192
rect 32585 12183 32643 12189
rect 32674 12180 32680 12192
rect 32732 12180 32738 12232
rect 32784 12229 32812 12260
rect 33045 12257 33057 12291
rect 33091 12288 33103 12291
rect 33594 12288 33600 12300
rect 33091 12260 33600 12288
rect 33091 12257 33103 12260
rect 33045 12251 33103 12257
rect 33594 12248 33600 12260
rect 33652 12288 33658 12300
rect 33781 12291 33839 12297
rect 33781 12288 33793 12291
rect 33652 12260 33793 12288
rect 33652 12248 33658 12260
rect 33781 12257 33793 12260
rect 33827 12257 33839 12291
rect 33781 12251 33839 12257
rect 32769 12223 32827 12229
rect 32769 12189 32781 12223
rect 32815 12189 32827 12223
rect 32769 12183 32827 12189
rect 33137 12223 33195 12229
rect 33137 12189 33149 12223
rect 33183 12220 33195 12223
rect 34624 12220 34652 12396
rect 35912 12356 35940 12396
rect 36078 12384 36084 12396
rect 36136 12384 36142 12436
rect 41230 12424 41236 12436
rect 38580 12396 41236 12424
rect 38580 12356 38608 12396
rect 41230 12384 41236 12396
rect 41288 12384 41294 12436
rect 35912 12328 38608 12356
rect 38654 12288 38660 12300
rect 38028 12260 38660 12288
rect 33183 12192 34652 12220
rect 34701 12223 34759 12229
rect 33183 12189 33195 12192
rect 33137 12183 33195 12189
rect 34701 12189 34713 12223
rect 34747 12220 34759 12223
rect 35342 12220 35348 12232
rect 34747 12192 35348 12220
rect 34747 12189 34759 12192
rect 34701 12183 34759 12189
rect 35342 12180 35348 12192
rect 35400 12180 35406 12232
rect 35802 12180 35808 12232
rect 35860 12220 35866 12232
rect 36633 12223 36691 12229
rect 36633 12220 36645 12223
rect 35860 12192 36645 12220
rect 35860 12180 35866 12192
rect 36633 12189 36645 12192
rect 36679 12189 36691 12223
rect 36814 12220 36820 12232
rect 36775 12192 36820 12220
rect 36633 12183 36691 12189
rect 36814 12180 36820 12192
rect 36872 12180 36878 12232
rect 36909 12223 36967 12229
rect 36909 12189 36921 12223
rect 36955 12189 36967 12223
rect 36909 12183 36967 12189
rect 29546 12152 29552 12164
rect 29472 12124 29552 12152
rect 29546 12112 29552 12124
rect 29604 12112 29610 12164
rect 29825 12155 29883 12161
rect 29825 12121 29837 12155
rect 29871 12152 29883 12155
rect 30208 12152 30236 12180
rect 31481 12155 31539 12161
rect 31481 12152 31493 12155
rect 29871 12124 31493 12152
rect 29871 12121 29883 12124
rect 29825 12115 29883 12121
rect 31481 12121 31493 12124
rect 31527 12121 31539 12155
rect 31481 12115 31539 12121
rect 27525 12087 27583 12093
rect 27525 12084 27537 12087
rect 24596 12056 27537 12084
rect 27525 12053 27537 12056
rect 27571 12053 27583 12087
rect 28718 12084 28724 12096
rect 28679 12056 28724 12084
rect 27525 12047 27583 12053
rect 28718 12044 28724 12056
rect 28776 12044 28782 12096
rect 28994 12044 29000 12096
rect 29052 12084 29058 12096
rect 29840 12084 29868 12115
rect 31570 12112 31576 12164
rect 31628 12152 31634 12164
rect 32398 12152 32404 12164
rect 31628 12124 31673 12152
rect 32359 12124 32404 12152
rect 31628 12112 31634 12124
rect 32398 12112 32404 12124
rect 32456 12112 32462 12164
rect 33502 12112 33508 12164
rect 33560 12152 33566 12164
rect 33870 12152 33876 12164
rect 33560 12124 33876 12152
rect 33560 12112 33566 12124
rect 33870 12112 33876 12124
rect 33928 12152 33934 12164
rect 33965 12155 34023 12161
rect 33965 12152 33977 12155
rect 33928 12124 33977 12152
rect 33928 12112 33934 12124
rect 33965 12121 33977 12124
rect 34011 12121 34023 12155
rect 33965 12115 34023 12121
rect 34790 12112 34796 12164
rect 34848 12152 34854 12164
rect 34946 12155 35004 12161
rect 34946 12152 34958 12155
rect 34848 12124 34958 12152
rect 34848 12112 34854 12124
rect 34946 12121 34958 12124
rect 34992 12121 35004 12155
rect 36924 12152 36952 12183
rect 36998 12180 37004 12232
rect 37056 12220 37062 12232
rect 37056 12192 37101 12220
rect 37056 12180 37062 12192
rect 37550 12180 37556 12232
rect 37608 12220 37614 12232
rect 38028 12229 38056 12260
rect 38654 12248 38660 12260
rect 38712 12248 38718 12300
rect 37829 12223 37887 12229
rect 37829 12220 37841 12223
rect 37608 12192 37841 12220
rect 37608 12180 37614 12192
rect 37829 12189 37841 12192
rect 37875 12189 37887 12223
rect 37829 12183 37887 12189
rect 38013 12223 38071 12229
rect 38013 12189 38025 12223
rect 38059 12189 38071 12223
rect 38013 12183 38071 12189
rect 38105 12223 38163 12229
rect 38105 12189 38117 12223
rect 38151 12189 38163 12223
rect 38105 12183 38163 12189
rect 38197 12223 38255 12229
rect 38197 12189 38209 12223
rect 38243 12220 38255 12223
rect 38378 12220 38384 12232
rect 38243 12192 38384 12220
rect 38243 12189 38255 12192
rect 38197 12183 38255 12189
rect 37918 12152 37924 12164
rect 36924 12124 37924 12152
rect 34946 12115 35004 12121
rect 37918 12112 37924 12124
rect 37976 12152 37982 12164
rect 38120 12152 38148 12183
rect 38378 12180 38384 12192
rect 38436 12180 38442 12232
rect 39022 12180 39028 12232
rect 39080 12220 39086 12232
rect 39850 12220 39856 12232
rect 39080 12192 39856 12220
rect 39080 12180 39086 12192
rect 39850 12180 39856 12192
rect 39908 12180 39914 12232
rect 37976 12124 38148 12152
rect 38473 12155 38531 12161
rect 37976 12112 37982 12124
rect 38473 12121 38485 12155
rect 38519 12152 38531 12155
rect 40098 12155 40156 12161
rect 40098 12152 40110 12155
rect 38519 12124 40110 12152
rect 38519 12121 38531 12124
rect 38473 12115 38531 12121
rect 40098 12121 40110 12124
rect 40144 12121 40156 12155
rect 40098 12115 40156 12121
rect 29052 12056 29868 12084
rect 30193 12087 30251 12093
rect 29052 12044 29058 12056
rect 30193 12053 30205 12087
rect 30239 12084 30251 12087
rect 30374 12084 30380 12096
rect 30239 12056 30380 12084
rect 30239 12053 30251 12056
rect 30193 12047 30251 12053
rect 30374 12044 30380 12056
rect 30432 12044 30438 12096
rect 31849 12087 31907 12093
rect 31849 12053 31861 12087
rect 31895 12084 31907 12087
rect 32214 12084 32220 12096
rect 31895 12056 32220 12084
rect 31895 12053 31907 12056
rect 31849 12047 31907 12053
rect 32214 12044 32220 12056
rect 32272 12044 32278 12096
rect 37274 12084 37280 12096
rect 37235 12056 37280 12084
rect 37274 12044 37280 12056
rect 37332 12044 37338 12096
rect 1104 11994 68816 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 50294 11994
rect 50346 11942 50358 11994
rect 50410 11942 50422 11994
rect 50474 11942 50486 11994
rect 50538 11942 50550 11994
rect 50602 11942 68816 11994
rect 1104 11920 68816 11942
rect 2130 11840 2136 11892
rect 2188 11880 2194 11892
rect 2225 11883 2283 11889
rect 2225 11880 2237 11883
rect 2188 11852 2237 11880
rect 2188 11840 2194 11852
rect 2225 11849 2237 11852
rect 2271 11849 2283 11883
rect 2225 11843 2283 11849
rect 2406 11840 2412 11892
rect 2464 11880 2470 11892
rect 2685 11883 2743 11889
rect 2685 11880 2697 11883
rect 2464 11852 2697 11880
rect 2464 11840 2470 11852
rect 2685 11849 2697 11852
rect 2731 11849 2743 11883
rect 2685 11843 2743 11849
rect 4157 11883 4215 11889
rect 4157 11849 4169 11883
rect 4203 11880 4215 11883
rect 4614 11880 4620 11892
rect 4203 11852 4620 11880
rect 4203 11849 4215 11852
rect 4157 11843 4215 11849
rect 4614 11840 4620 11852
rect 4672 11840 4678 11892
rect 6730 11880 6736 11892
rect 6691 11852 6736 11880
rect 6730 11840 6736 11852
rect 6788 11840 6794 11892
rect 7190 11880 7196 11892
rect 7151 11852 7196 11880
rect 7190 11840 7196 11852
rect 7248 11880 7254 11892
rect 7248 11852 8892 11880
rect 7248 11840 7254 11852
rect 1765 11815 1823 11821
rect 1765 11781 1777 11815
rect 1811 11812 1823 11815
rect 1946 11812 1952 11824
rect 1811 11784 1952 11812
rect 1811 11781 1823 11784
rect 1765 11775 1823 11781
rect 1946 11772 1952 11784
rect 2004 11812 2010 11824
rect 2004 11784 2774 11812
rect 2004 11772 2010 11784
rect 2038 11744 2044 11756
rect 1999 11716 2044 11744
rect 2038 11704 2044 11716
rect 2096 11704 2102 11756
rect 2746 11744 2774 11784
rect 5718 11772 5724 11824
rect 5776 11812 5782 11824
rect 6549 11815 6607 11821
rect 6549 11812 6561 11815
rect 5776 11784 6561 11812
rect 5776 11772 5782 11784
rect 6549 11781 6561 11784
rect 6595 11812 6607 11815
rect 8478 11812 8484 11824
rect 6595 11784 8484 11812
rect 6595 11781 6607 11784
rect 6549 11775 6607 11781
rect 8478 11772 8484 11784
rect 8536 11772 8542 11824
rect 3053 11747 3111 11753
rect 3053 11744 3065 11747
rect 2746 11716 3065 11744
rect 3053 11713 3065 11716
rect 3099 11713 3111 11747
rect 3053 11707 3111 11713
rect 5629 11747 5687 11753
rect 5629 11713 5641 11747
rect 5675 11744 5687 11747
rect 5810 11744 5816 11756
rect 5675 11716 5816 11744
rect 5675 11713 5687 11716
rect 5629 11707 5687 11713
rect 5810 11704 5816 11716
rect 5868 11704 5874 11756
rect 5994 11704 6000 11756
rect 6052 11744 6058 11756
rect 8018 11753 8024 11756
rect 6365 11747 6423 11753
rect 6365 11744 6377 11747
rect 6052 11716 6377 11744
rect 6052 11704 6058 11716
rect 6365 11713 6377 11716
rect 6411 11713 6423 11747
rect 8012 11744 8024 11753
rect 7979 11716 8024 11744
rect 6365 11707 6423 11713
rect 8012 11707 8024 11716
rect 8018 11704 8024 11707
rect 8076 11704 8082 11756
rect 1949 11679 2007 11685
rect 1949 11645 1961 11679
rect 1995 11676 2007 11679
rect 2498 11676 2504 11688
rect 1995 11648 2504 11676
rect 1995 11645 2007 11648
rect 1949 11639 2007 11645
rect 2498 11636 2504 11648
rect 2556 11636 2562 11688
rect 2961 11679 3019 11685
rect 2961 11645 2973 11679
rect 3007 11676 3019 11679
rect 3007 11648 3041 11676
rect 3007 11645 3019 11648
rect 2961 11639 3019 11645
rect 2976 11608 3004 11639
rect 7098 11636 7104 11688
rect 7156 11676 7162 11688
rect 7745 11679 7803 11685
rect 7745 11676 7757 11679
rect 7156 11648 7757 11676
rect 7156 11636 7162 11648
rect 7745 11645 7757 11648
rect 7791 11645 7803 11679
rect 7745 11639 7803 11645
rect 3234 11608 3240 11620
rect 2056 11580 3240 11608
rect 2056 11549 2084 11580
rect 3234 11568 3240 11580
rect 3292 11568 3298 11620
rect 8864 11608 8892 11852
rect 8938 11840 8944 11892
rect 8996 11880 9002 11892
rect 9125 11883 9183 11889
rect 9125 11880 9137 11883
rect 8996 11852 9137 11880
rect 8996 11840 9002 11852
rect 9125 11849 9137 11852
rect 9171 11849 9183 11883
rect 9125 11843 9183 11849
rect 17126 11840 17132 11892
rect 17184 11880 17190 11892
rect 17865 11883 17923 11889
rect 17865 11880 17877 11883
rect 17184 11852 17877 11880
rect 17184 11840 17190 11852
rect 17865 11849 17877 11852
rect 17911 11849 17923 11883
rect 18782 11880 18788 11892
rect 18743 11852 18788 11880
rect 17865 11843 17923 11849
rect 18782 11840 18788 11852
rect 18840 11840 18846 11892
rect 23290 11880 23296 11892
rect 23251 11852 23296 11880
rect 23290 11840 23296 11852
rect 23348 11840 23354 11892
rect 25498 11880 25504 11892
rect 23584 11852 25504 11880
rect 10042 11772 10048 11824
rect 10100 11812 10106 11824
rect 11701 11815 11759 11821
rect 11701 11812 11713 11815
rect 10100 11784 11713 11812
rect 10100 11772 10106 11784
rect 11701 11781 11713 11784
rect 11747 11812 11759 11815
rect 11747 11784 12434 11812
rect 11747 11781 11759 11784
rect 11701 11775 11759 11781
rect 11330 11704 11336 11756
rect 11388 11744 11394 11756
rect 11517 11747 11575 11753
rect 11517 11744 11529 11747
rect 11388 11716 11529 11744
rect 11388 11704 11394 11716
rect 11517 11713 11529 11716
rect 11563 11713 11575 11747
rect 12406 11744 12434 11784
rect 13170 11772 13176 11824
rect 13228 11812 13234 11824
rect 15013 11815 15071 11821
rect 15013 11812 15025 11815
rect 13228 11784 15025 11812
rect 13228 11772 13234 11784
rect 15013 11781 15025 11784
rect 15059 11812 15071 11815
rect 16206 11812 16212 11824
rect 15059 11784 16212 11812
rect 15059 11781 15071 11784
rect 15013 11775 15071 11781
rect 16206 11772 16212 11784
rect 16264 11772 16270 11824
rect 23198 11812 23204 11824
rect 17052 11784 23204 11812
rect 12897 11747 12955 11753
rect 12897 11744 12909 11747
rect 12406 11716 12909 11744
rect 11517 11707 11575 11713
rect 12897 11713 12909 11716
rect 12943 11713 12955 11747
rect 12897 11707 12955 11713
rect 14185 11747 14243 11753
rect 14185 11713 14197 11747
rect 14231 11744 14243 11747
rect 15194 11744 15200 11756
rect 14231 11716 15200 11744
rect 14231 11713 14243 11716
rect 14185 11707 14243 11713
rect 15194 11704 15200 11716
rect 15252 11704 15258 11756
rect 15746 11744 15752 11756
rect 15707 11716 15752 11744
rect 15746 11704 15752 11716
rect 15804 11704 15810 11756
rect 15933 11747 15991 11753
rect 15933 11713 15945 11747
rect 15979 11744 15991 11747
rect 16298 11744 16304 11756
rect 15979 11716 16304 11744
rect 15979 11713 15991 11716
rect 15933 11707 15991 11713
rect 16298 11704 16304 11716
rect 16356 11704 16362 11756
rect 17052 11753 17080 11784
rect 23198 11772 23204 11784
rect 23256 11772 23262 11824
rect 23584 11821 23612 11852
rect 25498 11840 25504 11852
rect 25556 11840 25562 11892
rect 28994 11880 29000 11892
rect 26068 11852 29000 11880
rect 23569 11815 23627 11821
rect 23569 11781 23581 11815
rect 23615 11781 23627 11815
rect 23569 11775 23627 11781
rect 23661 11815 23719 11821
rect 23661 11781 23673 11815
rect 23707 11812 23719 11815
rect 23934 11812 23940 11824
rect 23707 11784 23940 11812
rect 23707 11781 23719 11784
rect 23661 11775 23719 11781
rect 23934 11772 23940 11784
rect 23992 11772 23998 11824
rect 24118 11772 24124 11824
rect 24176 11812 24182 11824
rect 24397 11815 24455 11821
rect 24397 11812 24409 11815
rect 24176 11784 24409 11812
rect 24176 11772 24182 11784
rect 24397 11781 24409 11784
rect 24443 11812 24455 11815
rect 24762 11812 24768 11824
rect 24443 11784 24768 11812
rect 24443 11781 24455 11784
rect 24397 11775 24455 11781
rect 24762 11772 24768 11784
rect 24820 11772 24826 11824
rect 25130 11812 25136 11824
rect 25091 11784 25136 11812
rect 25130 11772 25136 11784
rect 25188 11772 25194 11824
rect 25406 11772 25412 11824
rect 25464 11812 25470 11824
rect 26068 11812 26096 11852
rect 28994 11840 29000 11852
rect 29052 11840 29058 11892
rect 29089 11883 29147 11889
rect 29089 11849 29101 11883
rect 29135 11880 29147 11883
rect 29454 11880 29460 11892
rect 29135 11852 29460 11880
rect 29135 11849 29147 11852
rect 29089 11843 29147 11849
rect 29454 11840 29460 11852
rect 29512 11840 29518 11892
rect 29638 11840 29644 11892
rect 29696 11880 29702 11892
rect 33042 11880 33048 11892
rect 29696 11852 33048 11880
rect 29696 11840 29702 11852
rect 33042 11840 33048 11852
rect 33100 11840 33106 11892
rect 34514 11840 34520 11892
rect 34572 11880 34578 11892
rect 35253 11883 35311 11889
rect 35253 11880 35265 11883
rect 34572 11852 35265 11880
rect 34572 11840 34578 11852
rect 35253 11849 35265 11852
rect 35299 11849 35311 11883
rect 35253 11843 35311 11849
rect 35618 11840 35624 11892
rect 35676 11880 35682 11892
rect 35676 11852 37320 11880
rect 35676 11840 35682 11852
rect 29270 11812 29276 11824
rect 25464 11784 26096 11812
rect 26160 11784 29276 11812
rect 25464 11772 25470 11784
rect 17037 11747 17095 11753
rect 17037 11713 17049 11747
rect 17083 11713 17095 11747
rect 17037 11707 17095 11713
rect 17126 11704 17132 11756
rect 17184 11744 17190 11756
rect 17221 11747 17279 11753
rect 17221 11744 17233 11747
rect 17184 11716 17233 11744
rect 17184 11704 17190 11716
rect 17221 11713 17233 11716
rect 17267 11713 17279 11747
rect 17221 11707 17279 11713
rect 17405 11747 17463 11753
rect 17405 11713 17417 11747
rect 17451 11744 17463 11747
rect 18506 11744 18512 11756
rect 17451 11716 18512 11744
rect 17451 11713 17463 11716
rect 17405 11707 17463 11713
rect 15286 11636 15292 11688
rect 15344 11676 15350 11688
rect 16945 11679 17003 11685
rect 16945 11676 16957 11679
rect 15344 11648 16957 11676
rect 15344 11636 15350 11648
rect 16945 11645 16957 11648
rect 16991 11645 17003 11679
rect 17420 11676 17448 11707
rect 18506 11704 18512 11716
rect 18564 11744 18570 11756
rect 18693 11747 18751 11753
rect 18693 11744 18705 11747
rect 18564 11716 18705 11744
rect 18564 11704 18570 11716
rect 18693 11713 18705 11716
rect 18739 11713 18751 11747
rect 18693 11707 18751 11713
rect 19061 11747 19119 11753
rect 19061 11713 19073 11747
rect 19107 11744 19119 11747
rect 20070 11744 20076 11756
rect 19107 11716 20076 11744
rect 19107 11713 19119 11716
rect 19061 11707 19119 11713
rect 20070 11704 20076 11716
rect 20128 11704 20134 11756
rect 20349 11747 20407 11753
rect 20349 11744 20361 11747
rect 20180 11716 20361 11744
rect 16945 11639 17003 11645
rect 17052 11648 17448 11676
rect 17052 11620 17080 11648
rect 18230 11636 18236 11688
rect 18288 11676 18294 11688
rect 19153 11679 19211 11685
rect 19153 11676 19165 11679
rect 18288 11648 19165 11676
rect 18288 11636 18294 11648
rect 19153 11645 19165 11648
rect 19199 11645 19211 11679
rect 19153 11639 19211 11645
rect 11514 11608 11520 11620
rect 8864 11580 11520 11608
rect 11514 11568 11520 11580
rect 11572 11568 11578 11620
rect 17034 11568 17040 11620
rect 17092 11568 17098 11620
rect 17129 11611 17187 11617
rect 17129 11577 17141 11611
rect 17175 11608 17187 11611
rect 17402 11608 17408 11620
rect 17175 11580 17408 11608
rect 17175 11577 17187 11580
rect 17129 11571 17187 11577
rect 17402 11568 17408 11580
rect 17460 11568 17466 11620
rect 19242 11568 19248 11620
rect 19300 11608 19306 11620
rect 19429 11611 19487 11617
rect 19429 11608 19441 11611
rect 19300 11580 19441 11608
rect 19300 11568 19306 11580
rect 19429 11577 19441 11580
rect 19475 11577 19487 11611
rect 19429 11571 19487 11577
rect 2041 11543 2099 11549
rect 2041 11509 2053 11543
rect 2087 11509 2099 11543
rect 2041 11503 2099 11509
rect 2498 11500 2504 11552
rect 2556 11540 2562 11552
rect 2869 11543 2927 11549
rect 2869 11540 2881 11543
rect 2556 11512 2881 11540
rect 2556 11500 2562 11512
rect 2869 11509 2881 11512
rect 2915 11540 2927 11543
rect 3513 11543 3571 11549
rect 3513 11540 3525 11543
rect 2915 11512 3525 11540
rect 2915 11509 2927 11512
rect 2869 11503 2927 11509
rect 3513 11509 3525 11512
rect 3559 11509 3571 11543
rect 3513 11503 3571 11509
rect 5813 11543 5871 11549
rect 5813 11509 5825 11543
rect 5859 11540 5871 11543
rect 5994 11540 6000 11552
rect 5859 11512 6000 11540
rect 5859 11509 5871 11512
rect 5813 11503 5871 11509
rect 5994 11500 6000 11512
rect 6052 11500 6058 11552
rect 10870 11500 10876 11552
rect 10928 11540 10934 11552
rect 10965 11543 11023 11549
rect 10965 11540 10977 11543
rect 10928 11512 10977 11540
rect 10928 11500 10934 11512
rect 10965 11509 10977 11512
rect 11011 11540 11023 11543
rect 11054 11540 11060 11552
rect 11011 11512 11060 11540
rect 11011 11509 11023 11512
rect 10965 11503 11023 11509
rect 11054 11500 11060 11512
rect 11112 11500 11118 11552
rect 11885 11543 11943 11549
rect 11885 11509 11897 11543
rect 11931 11540 11943 11543
rect 12066 11540 12072 11552
rect 11931 11512 12072 11540
rect 11931 11509 11943 11512
rect 11885 11503 11943 11509
rect 12066 11500 12072 11512
rect 12124 11500 12130 11552
rect 12437 11543 12495 11549
rect 12437 11509 12449 11543
rect 12483 11540 12495 11543
rect 12618 11540 12624 11552
rect 12483 11512 12624 11540
rect 12483 11509 12495 11512
rect 12437 11503 12495 11509
rect 12618 11500 12624 11512
rect 12676 11500 12682 11552
rect 15565 11543 15623 11549
rect 15565 11509 15577 11543
rect 15611 11540 15623 11543
rect 15930 11540 15936 11552
rect 15611 11512 15936 11540
rect 15611 11509 15623 11512
rect 15565 11503 15623 11509
rect 15930 11500 15936 11512
rect 15988 11500 15994 11552
rect 16574 11500 16580 11552
rect 16632 11540 16638 11552
rect 16669 11543 16727 11549
rect 16669 11540 16681 11543
rect 16632 11512 16681 11540
rect 16632 11500 16638 11512
rect 16669 11509 16681 11512
rect 16715 11509 16727 11543
rect 18966 11540 18972 11552
rect 18927 11512 18972 11540
rect 16669 11503 16727 11509
rect 18966 11500 18972 11512
rect 19024 11500 19030 11552
rect 19518 11500 19524 11552
rect 19576 11540 19582 11552
rect 20070 11540 20076 11552
rect 19576 11512 20076 11540
rect 19576 11500 19582 11512
rect 20070 11500 20076 11512
rect 20128 11500 20134 11552
rect 20180 11540 20208 11716
rect 20349 11713 20361 11716
rect 20395 11713 20407 11747
rect 20530 11744 20536 11756
rect 20491 11716 20536 11744
rect 20349 11707 20407 11713
rect 20530 11704 20536 11716
rect 20588 11704 20594 11756
rect 20625 11747 20683 11753
rect 20625 11713 20637 11747
rect 20671 11713 20683 11747
rect 20625 11707 20683 11713
rect 20717 11747 20775 11753
rect 20717 11713 20729 11747
rect 20763 11713 20775 11747
rect 20717 11707 20775 11713
rect 22189 11747 22247 11753
rect 22189 11713 22201 11747
rect 22235 11713 22247 11747
rect 22370 11744 22376 11756
rect 22331 11716 22376 11744
rect 22189 11707 22247 11713
rect 20254 11636 20260 11688
rect 20312 11676 20318 11688
rect 20640 11676 20668 11707
rect 20312 11648 20668 11676
rect 20312 11636 20318 11648
rect 20732 11608 20760 11707
rect 20990 11636 20996 11688
rect 21048 11676 21054 11688
rect 22005 11679 22063 11685
rect 22005 11676 22017 11679
rect 21048 11648 22017 11676
rect 21048 11636 21054 11648
rect 22005 11645 22017 11648
rect 22051 11645 22063 11679
rect 22204 11676 22232 11707
rect 22370 11704 22376 11716
rect 22428 11704 22434 11756
rect 22557 11747 22615 11753
rect 22557 11713 22569 11747
rect 22603 11744 22615 11747
rect 22833 11747 22891 11753
rect 22603 11716 22692 11744
rect 22603 11713 22615 11716
rect 22557 11707 22615 11713
rect 22204 11648 22416 11676
rect 22005 11639 22063 11645
rect 22278 11608 22284 11620
rect 20732 11580 22284 11608
rect 22278 11568 22284 11580
rect 22336 11568 22342 11620
rect 20714 11540 20720 11552
rect 20180 11512 20720 11540
rect 20714 11500 20720 11512
rect 20772 11500 20778 11552
rect 20901 11543 20959 11549
rect 20901 11509 20913 11543
rect 20947 11540 20959 11543
rect 22388 11540 22416 11648
rect 22664 11608 22692 11716
rect 22833 11713 22845 11747
rect 22879 11744 22891 11747
rect 22922 11744 22928 11756
rect 22879 11716 22928 11744
rect 22879 11713 22891 11716
rect 22833 11707 22891 11713
rect 22922 11704 22928 11716
rect 22980 11704 22986 11756
rect 23474 11744 23480 11756
rect 23435 11716 23480 11744
rect 23474 11704 23480 11716
rect 23532 11704 23538 11756
rect 23845 11747 23903 11753
rect 23845 11713 23857 11747
rect 23891 11744 23903 11747
rect 24578 11744 24584 11756
rect 23891 11716 24440 11744
rect 24539 11716 24584 11744
rect 23891 11713 23903 11716
rect 23845 11707 23903 11713
rect 24412 11676 24440 11716
rect 24578 11704 24584 11716
rect 24636 11744 24642 11756
rect 26160 11744 26188 11784
rect 29270 11772 29276 11784
rect 29328 11812 29334 11824
rect 30101 11815 30159 11821
rect 30101 11812 30113 11815
rect 29328 11784 30113 11812
rect 29328 11772 29334 11784
rect 30101 11781 30113 11784
rect 30147 11781 30159 11815
rect 30101 11775 30159 11781
rect 35342 11772 35348 11824
rect 35400 11812 35406 11824
rect 35802 11812 35808 11824
rect 35400 11784 35808 11812
rect 35400 11772 35406 11784
rect 35802 11772 35808 11784
rect 35860 11812 35866 11824
rect 36449 11815 36507 11821
rect 36449 11812 36461 11815
rect 35860 11784 36461 11812
rect 35860 11772 35866 11784
rect 36449 11781 36461 11784
rect 36495 11781 36507 11815
rect 36449 11775 36507 11781
rect 24636 11716 26188 11744
rect 24636 11704 24642 11716
rect 26234 11704 26240 11756
rect 26292 11744 26298 11756
rect 26292 11716 26385 11744
rect 26292 11704 26298 11716
rect 26418 11704 26424 11756
rect 26476 11744 26482 11756
rect 27341 11747 27399 11753
rect 27341 11744 27353 11747
rect 26476 11716 27353 11744
rect 26476 11704 26482 11716
rect 27341 11713 27353 11716
rect 27387 11713 27399 11747
rect 27341 11707 27399 11713
rect 27430 11704 27436 11756
rect 27488 11744 27494 11756
rect 27525 11747 27583 11753
rect 27525 11744 27537 11747
rect 27488 11716 27537 11744
rect 27488 11704 27494 11716
rect 27525 11713 27537 11716
rect 27571 11713 27583 11747
rect 27525 11707 27583 11713
rect 27617 11747 27675 11753
rect 27617 11713 27629 11747
rect 27663 11713 27675 11747
rect 27617 11707 27675 11713
rect 26252 11676 26280 11704
rect 26694 11676 26700 11688
rect 24412 11648 25636 11676
rect 26252 11648 26700 11676
rect 23750 11608 23756 11620
rect 22664 11580 23756 11608
rect 23750 11568 23756 11580
rect 23808 11568 23814 11620
rect 23934 11568 23940 11620
rect 23992 11608 23998 11620
rect 25406 11608 25412 11620
rect 23992 11580 25412 11608
rect 23992 11568 23998 11580
rect 25406 11568 25412 11580
rect 25464 11568 25470 11620
rect 20947 11512 22416 11540
rect 25608 11540 25636 11648
rect 26694 11636 26700 11648
rect 26752 11636 26758 11688
rect 26786 11636 26792 11688
rect 26844 11676 26850 11688
rect 27635 11676 27663 11707
rect 27706 11704 27712 11756
rect 27764 11744 27770 11756
rect 27764 11716 27809 11744
rect 27764 11704 27770 11716
rect 29822 11704 29828 11756
rect 29880 11753 29886 11756
rect 29880 11747 29929 11753
rect 29880 11713 29883 11747
rect 29917 11713 29929 11747
rect 29880 11707 29929 11713
rect 30012 11747 30070 11753
rect 30012 11713 30024 11747
rect 30058 11713 30070 11747
rect 30012 11707 30070 11713
rect 29880 11704 29886 11707
rect 26844 11648 27663 11676
rect 26844 11636 26850 11648
rect 25685 11611 25743 11617
rect 25685 11577 25697 11611
rect 25731 11608 25743 11611
rect 26421 11611 26479 11617
rect 26421 11608 26433 11611
rect 25731 11580 26433 11608
rect 25731 11577 25743 11580
rect 25685 11571 25743 11577
rect 26421 11577 26433 11580
rect 26467 11608 26479 11611
rect 27724 11608 27752 11704
rect 26467 11580 27752 11608
rect 30027 11608 30055 11707
rect 30190 11704 30196 11756
rect 30248 11753 30254 11756
rect 30248 11747 30287 11753
rect 30275 11713 30287 11747
rect 30248 11707 30287 11713
rect 30248 11704 30254 11707
rect 30374 11704 30380 11756
rect 30432 11744 30438 11756
rect 30432 11716 30477 11744
rect 30432 11704 30438 11716
rect 32858 11704 32864 11756
rect 32916 11744 32922 11756
rect 33413 11747 33471 11753
rect 33413 11744 33425 11747
rect 32916 11716 33425 11744
rect 32916 11704 32922 11716
rect 33413 11713 33425 11716
rect 33459 11713 33471 11747
rect 33594 11744 33600 11756
rect 33555 11716 33600 11744
rect 33413 11707 33471 11713
rect 33594 11704 33600 11716
rect 33652 11704 33658 11756
rect 34790 11704 34796 11756
rect 34848 11744 34854 11756
rect 37292 11753 37320 11852
rect 35069 11747 35127 11753
rect 35069 11744 35081 11747
rect 34848 11716 35081 11744
rect 34848 11704 34854 11716
rect 35069 11713 35081 11716
rect 35115 11713 35127 11747
rect 35069 11707 35127 11713
rect 35713 11747 35771 11753
rect 35713 11713 35725 11747
rect 35759 11713 35771 11747
rect 35713 11707 35771 11713
rect 37277 11747 37335 11753
rect 37277 11713 37289 11747
rect 37323 11713 37335 11747
rect 37550 11744 37556 11756
rect 37511 11716 37556 11744
rect 37277 11707 37335 11713
rect 34514 11676 34520 11688
rect 34475 11648 34520 11676
rect 34514 11636 34520 11648
rect 34572 11676 34578 11688
rect 35728 11676 35756 11707
rect 37550 11704 37556 11716
rect 37608 11704 37614 11756
rect 34572 11648 35756 11676
rect 34572 11636 34578 11648
rect 33505 11611 33563 11617
rect 30027 11580 32996 11608
rect 26467 11577 26479 11580
rect 26421 11571 26479 11577
rect 27706 11540 27712 11552
rect 25608 11512 27712 11540
rect 20947 11509 20959 11512
rect 20901 11503 20959 11509
rect 27706 11500 27712 11512
rect 27764 11500 27770 11552
rect 27798 11500 27804 11552
rect 27856 11540 27862 11552
rect 27985 11543 28043 11549
rect 27985 11540 27997 11543
rect 27856 11512 27997 11540
rect 27856 11500 27862 11512
rect 27985 11509 27997 11512
rect 28031 11509 28043 11543
rect 27985 11503 28043 11509
rect 28074 11500 28080 11552
rect 28132 11540 28138 11552
rect 28445 11543 28503 11549
rect 28445 11540 28457 11543
rect 28132 11512 28457 11540
rect 28132 11500 28138 11512
rect 28445 11509 28457 11512
rect 28491 11540 28503 11543
rect 28626 11540 28632 11552
rect 28491 11512 28632 11540
rect 28491 11509 28503 11512
rect 28445 11503 28503 11509
rect 28626 11500 28632 11512
rect 28684 11500 28690 11552
rect 29730 11540 29736 11552
rect 29691 11512 29736 11540
rect 29730 11500 29736 11512
rect 29788 11500 29794 11552
rect 30006 11500 30012 11552
rect 30064 11540 30070 11552
rect 30190 11540 30196 11552
rect 30064 11512 30196 11540
rect 30064 11500 30070 11512
rect 30190 11500 30196 11512
rect 30248 11500 30254 11552
rect 32858 11540 32864 11552
rect 32819 11512 32864 11540
rect 32858 11500 32864 11512
rect 32916 11500 32922 11552
rect 32968 11540 32996 11580
rect 33505 11577 33517 11611
rect 33551 11608 33563 11611
rect 36630 11608 36636 11620
rect 33551 11580 36636 11608
rect 33551 11577 33563 11580
rect 33505 11571 33563 11577
rect 36630 11568 36636 11580
rect 36688 11568 36694 11620
rect 36906 11540 36912 11552
rect 32968 11512 36912 11540
rect 36906 11500 36912 11512
rect 36964 11540 36970 11552
rect 37826 11540 37832 11552
rect 36964 11512 37832 11540
rect 36964 11500 36970 11512
rect 37826 11500 37832 11512
rect 37884 11500 37890 11552
rect 67634 11540 67640 11552
rect 67595 11512 67640 11540
rect 67634 11500 67640 11512
rect 67692 11500 67698 11552
rect 1104 11450 68816 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 65654 11450
rect 65706 11398 65718 11450
rect 65770 11398 65782 11450
rect 65834 11398 65846 11450
rect 65898 11398 65910 11450
rect 65962 11398 68816 11450
rect 1104 11376 68816 11398
rect 9217 11339 9275 11345
rect 9217 11305 9229 11339
rect 9263 11336 9275 11339
rect 9950 11336 9956 11348
rect 9263 11308 9956 11336
rect 9263 11305 9275 11308
rect 9217 11299 9275 11305
rect 9950 11296 9956 11308
rect 10008 11296 10014 11348
rect 12805 11339 12863 11345
rect 12805 11305 12817 11339
rect 12851 11336 12863 11339
rect 13354 11336 13360 11348
rect 12851 11308 13360 11336
rect 12851 11305 12863 11308
rect 12805 11299 12863 11305
rect 13354 11296 13360 11308
rect 13412 11296 13418 11348
rect 13538 11296 13544 11348
rect 13596 11336 13602 11348
rect 15013 11339 15071 11345
rect 15013 11336 15025 11339
rect 13596 11308 15025 11336
rect 13596 11296 13602 11308
rect 15013 11305 15025 11308
rect 15059 11305 15071 11339
rect 15013 11299 15071 11305
rect 15102 11296 15108 11348
rect 15160 11336 15166 11348
rect 15160 11308 15205 11336
rect 15160 11296 15166 11308
rect 15562 11296 15568 11348
rect 15620 11336 15626 11348
rect 16577 11339 16635 11345
rect 16577 11336 16589 11339
rect 15620 11308 16589 11336
rect 15620 11296 15626 11308
rect 16577 11305 16589 11308
rect 16623 11305 16635 11339
rect 16577 11299 16635 11305
rect 18325 11339 18383 11345
rect 18325 11305 18337 11339
rect 18371 11336 18383 11339
rect 18414 11336 18420 11348
rect 18371 11308 18420 11336
rect 18371 11305 18383 11308
rect 18325 11299 18383 11305
rect 18414 11296 18420 11308
rect 18472 11296 18478 11348
rect 19705 11339 19763 11345
rect 19705 11305 19717 11339
rect 19751 11336 19763 11339
rect 20162 11336 20168 11348
rect 19751 11308 20168 11336
rect 19751 11305 19763 11308
rect 19705 11299 19763 11305
rect 20162 11296 20168 11308
rect 20220 11296 20226 11348
rect 21085 11339 21143 11345
rect 21085 11305 21097 11339
rect 21131 11336 21143 11339
rect 22094 11336 22100 11348
rect 21131 11308 22100 11336
rect 21131 11305 21143 11308
rect 21085 11299 21143 11305
rect 22094 11296 22100 11308
rect 22152 11296 22158 11348
rect 22370 11336 22376 11348
rect 22331 11308 22376 11336
rect 22370 11296 22376 11308
rect 22428 11296 22434 11348
rect 23750 11336 23756 11348
rect 23663 11308 23756 11336
rect 23750 11296 23756 11308
rect 23808 11336 23814 11348
rect 24670 11336 24676 11348
rect 23808 11308 24676 11336
rect 23808 11296 23814 11308
rect 24670 11296 24676 11308
rect 24728 11296 24734 11348
rect 28718 11296 28724 11348
rect 28776 11336 28782 11348
rect 28776 11308 34192 11336
rect 28776 11296 28782 11308
rect 5169 11271 5227 11277
rect 5169 11237 5181 11271
rect 5215 11237 5227 11271
rect 5169 11231 5227 11237
rect 2225 11135 2283 11141
rect 2225 11101 2237 11135
rect 2271 11132 2283 11135
rect 3142 11132 3148 11144
rect 2271 11104 3148 11132
rect 2271 11101 2283 11104
rect 2225 11095 2283 11101
rect 3142 11092 3148 11104
rect 3200 11092 3206 11144
rect 3786 11132 3792 11144
rect 3747 11104 3792 11132
rect 3786 11092 3792 11104
rect 3844 11092 3850 11144
rect 5184 11132 5212 11231
rect 11422 11228 11428 11280
rect 11480 11268 11486 11280
rect 11606 11268 11612 11280
rect 11480 11240 11612 11268
rect 11480 11228 11486 11240
rect 11606 11228 11612 11240
rect 11664 11268 11670 11280
rect 14734 11268 14740 11280
rect 11664 11240 14740 11268
rect 11664 11228 11670 11240
rect 14734 11228 14740 11240
rect 14792 11228 14798 11280
rect 14826 11228 14832 11280
rect 14884 11268 14890 11280
rect 14884 11240 17448 11268
rect 14884 11228 14890 11240
rect 6086 11160 6092 11212
rect 6144 11200 6150 11212
rect 6457 11203 6515 11209
rect 6457 11200 6469 11203
rect 6144 11172 6469 11200
rect 6144 11160 6150 11172
rect 6457 11169 6469 11172
rect 6503 11169 6515 11203
rect 6457 11163 6515 11169
rect 7098 11160 7104 11212
rect 7156 11200 7162 11212
rect 7469 11203 7527 11209
rect 7469 11200 7481 11203
rect 7156 11172 7481 11200
rect 7156 11160 7162 11172
rect 7469 11169 7481 11172
rect 7515 11169 7527 11203
rect 7469 11163 7527 11169
rect 15197 11203 15255 11209
rect 15197 11169 15209 11203
rect 15243 11200 15255 11203
rect 16482 11200 16488 11212
rect 15243 11172 16488 11200
rect 15243 11169 15255 11172
rect 15197 11163 15255 11169
rect 16482 11160 16488 11172
rect 16540 11160 16546 11212
rect 16669 11203 16727 11209
rect 16669 11169 16681 11203
rect 16715 11200 16727 11203
rect 17310 11200 17316 11212
rect 16715 11172 17316 11200
rect 16715 11169 16727 11172
rect 16669 11163 16727 11169
rect 17310 11160 17316 11172
rect 17368 11160 17374 11212
rect 17420 11200 17448 11240
rect 17678 11228 17684 11280
rect 17736 11268 17742 11280
rect 24397 11271 24455 11277
rect 24397 11268 24409 11271
rect 17736 11240 24409 11268
rect 17736 11228 17742 11240
rect 24397 11237 24409 11240
rect 24443 11237 24455 11271
rect 29822 11268 29828 11280
rect 29783 11240 29828 11268
rect 24397 11231 24455 11237
rect 29822 11228 29828 11240
rect 29880 11228 29886 11280
rect 32858 11268 32864 11280
rect 29932 11240 31754 11268
rect 32819 11240 32864 11268
rect 17420 11172 18184 11200
rect 5813 11135 5871 11141
rect 5813 11132 5825 11135
rect 5184 11104 5825 11132
rect 5813 11101 5825 11104
rect 5859 11132 5871 11135
rect 9766 11132 9772 11144
rect 5859 11104 9772 11132
rect 5859 11101 5871 11104
rect 5813 11095 5871 11101
rect 9766 11092 9772 11104
rect 9824 11092 9830 11144
rect 10597 11135 10655 11141
rect 10597 11101 10609 11135
rect 10643 11132 10655 11135
rect 11606 11132 11612 11144
rect 10643 11104 11612 11132
rect 10643 11101 10655 11104
rect 10597 11095 10655 11101
rect 11606 11092 11612 11104
rect 11664 11092 11670 11144
rect 11882 11092 11888 11144
rect 11940 11132 11946 11144
rect 12161 11135 12219 11141
rect 12161 11132 12173 11135
rect 11940 11104 12173 11132
rect 11940 11092 11946 11104
rect 12161 11101 12173 11104
rect 12207 11101 12219 11135
rect 12161 11095 12219 11101
rect 12345 11135 12403 11141
rect 12345 11101 12357 11135
rect 12391 11101 12403 11135
rect 12345 11095 12403 11101
rect 4056 11067 4114 11073
rect 4056 11033 4068 11067
rect 4102 11064 4114 11067
rect 5074 11064 5080 11076
rect 4102 11036 5080 11064
rect 4102 11033 4114 11036
rect 4056 11027 4114 11033
rect 5074 11024 5080 11036
rect 5132 11024 5138 11076
rect 5994 11064 6000 11076
rect 5907 11036 6000 11064
rect 5994 11024 6000 11036
rect 6052 11024 6058 11076
rect 6638 11064 6644 11076
rect 6599 11036 6644 11064
rect 6638 11024 6644 11036
rect 6696 11024 6702 11076
rect 6825 11067 6883 11073
rect 6825 11033 6837 11067
rect 6871 11033 6883 11067
rect 8294 11064 8300 11076
rect 8255 11036 8300 11064
rect 6825 11027 6883 11033
rect 2498 10956 2504 11008
rect 2556 10996 2562 11008
rect 2685 10999 2743 11005
rect 2685 10996 2697 10999
rect 2556 10968 2697 10996
rect 2556 10956 2562 10968
rect 2685 10965 2697 10968
rect 2731 10965 2743 10999
rect 5626 10996 5632 11008
rect 5587 10968 5632 10996
rect 2685 10959 2743 10965
rect 5626 10956 5632 10968
rect 5684 10956 5690 11008
rect 6012 10996 6040 11024
rect 6840 10996 6868 11027
rect 8294 11024 8300 11036
rect 8352 11024 8358 11076
rect 10226 11024 10232 11076
rect 10284 11064 10290 11076
rect 10330 11067 10388 11073
rect 10330 11064 10342 11067
rect 10284 11036 10342 11064
rect 10284 11024 10290 11036
rect 10330 11033 10342 11036
rect 10376 11033 10388 11067
rect 10330 11027 10388 11033
rect 10502 11024 10508 11076
rect 10560 11064 10566 11076
rect 11330 11064 11336 11076
rect 10560 11036 11336 11064
rect 10560 11024 10566 11036
rect 11330 11024 11336 11036
rect 11388 11024 11394 11076
rect 11514 11064 11520 11076
rect 11475 11036 11520 11064
rect 11514 11024 11520 11036
rect 11572 11064 11578 11076
rect 11701 11067 11759 11073
rect 11572 11036 11652 11064
rect 11572 11024 11578 11036
rect 7742 10996 7748 11008
rect 6012 10968 7748 10996
rect 7742 10956 7748 10968
rect 7800 10996 7806 11008
rect 8938 10996 8944 11008
rect 7800 10968 8944 10996
rect 7800 10956 7806 10968
rect 8938 10956 8944 10968
rect 8996 10956 9002 11008
rect 11624 10996 11652 11036
rect 11701 11033 11713 11067
rect 11747 11064 11759 11067
rect 12360 11064 12388 11095
rect 12434 11092 12440 11144
rect 12492 11132 12498 11144
rect 12575 11135 12633 11141
rect 12492 11104 12537 11132
rect 12492 11092 12498 11104
rect 12575 11101 12587 11135
rect 12621 11132 12633 11135
rect 13814 11132 13820 11144
rect 12621 11104 13820 11132
rect 12621 11101 12633 11104
rect 12575 11095 12633 11101
rect 13814 11092 13820 11104
rect 13872 11132 13878 11144
rect 15289 11135 15347 11141
rect 13872 11104 14872 11132
rect 13872 11092 13878 11104
rect 13357 11067 13415 11073
rect 13357 11064 13369 11067
rect 11747 11036 12388 11064
rect 12452 11036 13369 11064
rect 11747 11033 11759 11036
rect 11701 11027 11759 11033
rect 12452 10996 12480 11036
rect 13357 11033 13369 11036
rect 13403 11064 13415 11067
rect 13538 11064 13544 11076
rect 13403 11036 13544 11064
rect 13403 11033 13415 11036
rect 13357 11027 13415 11033
rect 13538 11024 13544 11036
rect 13596 11024 13602 11076
rect 14642 11024 14648 11076
rect 14700 11064 14706 11076
rect 14737 11067 14795 11073
rect 14737 11064 14749 11067
rect 14700 11036 14749 11064
rect 14700 11024 14706 11036
rect 14737 11033 14749 11036
rect 14783 11033 14795 11067
rect 14844 11064 14872 11104
rect 15289 11101 15301 11135
rect 15335 11101 15347 11135
rect 15470 11132 15476 11144
rect 15431 11104 15476 11132
rect 15289 11095 15347 11101
rect 15304 11064 15332 11095
rect 15470 11092 15476 11104
rect 15528 11132 15534 11144
rect 15528 11104 16712 11132
rect 15528 11092 15534 11104
rect 16298 11064 16304 11076
rect 14844 11036 15332 11064
rect 16259 11036 16304 11064
rect 14737 11027 14795 11033
rect 16298 11024 16304 11036
rect 16356 11024 16362 11076
rect 16684 11064 16712 11104
rect 16758 11092 16764 11144
rect 16816 11132 16822 11144
rect 17034 11132 17040 11144
rect 16816 11104 16861 11132
rect 16947 11104 17040 11132
rect 16816 11092 16822 11104
rect 17034 11092 17040 11104
rect 17092 11092 17098 11144
rect 18156 11141 18184 11172
rect 18322 11160 18328 11212
rect 18380 11200 18386 11212
rect 18417 11203 18475 11209
rect 18417 11200 18429 11203
rect 18380 11172 18429 11200
rect 18380 11160 18386 11172
rect 18417 11169 18429 11172
rect 18463 11169 18475 11203
rect 18417 11163 18475 11169
rect 19426 11160 19432 11212
rect 19484 11200 19490 11212
rect 20530 11200 20536 11212
rect 19484 11172 20536 11200
rect 19484 11160 19490 11172
rect 20530 11160 20536 11172
rect 20588 11160 20594 11212
rect 20806 11160 20812 11212
rect 20864 11200 20870 11212
rect 22005 11203 22063 11209
rect 22005 11200 22017 11203
rect 20864 11172 22017 11200
rect 20864 11160 20870 11172
rect 22005 11169 22017 11172
rect 22051 11169 22063 11203
rect 22005 11163 22063 11169
rect 23109 11203 23167 11209
rect 23109 11169 23121 11203
rect 23155 11200 23167 11203
rect 23934 11200 23940 11212
rect 23155 11172 23940 11200
rect 23155 11169 23167 11172
rect 23109 11163 23167 11169
rect 23934 11160 23940 11172
rect 23992 11160 23998 11212
rect 27617 11203 27675 11209
rect 27617 11169 27629 11203
rect 27663 11200 27675 11203
rect 27982 11200 27988 11212
rect 27663 11172 27988 11200
rect 27663 11169 27675 11172
rect 27617 11163 27675 11169
rect 27982 11160 27988 11172
rect 28040 11160 28046 11212
rect 28166 11200 28172 11212
rect 28127 11172 28172 11200
rect 28166 11160 28172 11172
rect 28224 11160 28230 11212
rect 28626 11160 28632 11212
rect 28684 11200 28690 11212
rect 29932 11200 29960 11240
rect 28684 11172 29960 11200
rect 28684 11160 28690 11172
rect 30466 11160 30472 11212
rect 30524 11200 30530 11212
rect 30561 11203 30619 11209
rect 30561 11200 30573 11203
rect 30524 11172 30573 11200
rect 30524 11160 30530 11172
rect 30561 11169 30573 11172
rect 30607 11169 30619 11203
rect 31726 11200 31754 11240
rect 32858 11228 32864 11240
rect 32916 11228 32922 11280
rect 33594 11200 33600 11212
rect 31726 11172 32352 11200
rect 30561 11163 30619 11169
rect 17957 11135 18015 11141
rect 17957 11101 17969 11135
rect 18003 11101 18015 11135
rect 17957 11095 18015 11101
rect 18141 11135 18199 11141
rect 18141 11101 18153 11135
rect 18187 11101 18199 11135
rect 18141 11095 18199 11101
rect 17052 11064 17080 11092
rect 16684 11036 17080 11064
rect 17972 11064 18000 11095
rect 18230 11092 18236 11144
rect 18288 11132 18294 11144
rect 19889 11135 19947 11141
rect 18288 11104 18333 11132
rect 18288 11092 18294 11104
rect 19889 11101 19901 11135
rect 19935 11101 19947 11135
rect 20070 11132 20076 11144
rect 20031 11104 20076 11132
rect 19889 11095 19947 11101
rect 18322 11064 18328 11076
rect 17972 11036 18328 11064
rect 18322 11024 18328 11036
rect 18380 11024 18386 11076
rect 18598 11024 18604 11076
rect 18656 11064 18662 11076
rect 18693 11067 18751 11073
rect 18693 11064 18705 11067
rect 18656 11036 18705 11064
rect 18656 11024 18662 11036
rect 18693 11033 18705 11036
rect 18739 11033 18751 11067
rect 19904 11064 19932 11095
rect 20070 11092 20076 11104
rect 20128 11092 20134 11144
rect 20717 11135 20775 11141
rect 20717 11101 20729 11135
rect 20763 11101 20775 11135
rect 20717 11095 20775 11101
rect 20901 11135 20959 11141
rect 20901 11101 20913 11135
rect 20947 11101 20959 11135
rect 22186 11132 22192 11144
rect 22147 11104 22192 11132
rect 20901 11095 20959 11101
rect 20254 11064 20260 11076
rect 19904 11036 20260 11064
rect 18693 11027 18751 11033
rect 20254 11024 20260 11036
rect 20312 11064 20318 11076
rect 20732 11064 20760 11095
rect 20312 11036 20760 11064
rect 20312 11024 20318 11036
rect 20806 11024 20812 11076
rect 20864 11064 20870 11076
rect 20916 11064 20944 11095
rect 22186 11092 22192 11104
rect 22244 11092 22250 11144
rect 23842 11092 23848 11144
rect 23900 11132 23906 11144
rect 24581 11135 24639 11141
rect 24581 11132 24593 11135
rect 23900 11104 24593 11132
rect 23900 11092 23906 11104
rect 24581 11101 24593 11104
rect 24627 11101 24639 11135
rect 24762 11132 24768 11144
rect 24723 11104 24768 11132
rect 24581 11095 24639 11101
rect 20864 11036 20944 11064
rect 20864 11024 20870 11036
rect 22554 11024 22560 11076
rect 22612 11064 22618 11076
rect 22925 11067 22983 11073
rect 22925 11064 22937 11067
rect 22612 11036 22937 11064
rect 22612 11024 22618 11036
rect 22925 11033 22937 11036
rect 22971 11064 22983 11067
rect 23661 11067 23719 11073
rect 23661 11064 23673 11067
rect 22971 11036 23673 11064
rect 22971 11033 22983 11036
rect 22925 11027 22983 11033
rect 23661 11033 23673 11036
rect 23707 11033 23719 11067
rect 23661 11027 23719 11033
rect 16942 10996 16948 11008
rect 11624 10968 12480 10996
rect 16903 10968 16948 10996
rect 16942 10956 16948 10968
rect 17000 10956 17006 11008
rect 24596 10996 24624 11095
rect 24762 11092 24768 11104
rect 24820 11092 24826 11144
rect 24946 11132 24952 11144
rect 24907 11104 24952 11132
rect 24946 11092 24952 11104
rect 25004 11092 25010 11144
rect 25038 11092 25044 11144
rect 25096 11132 25102 11144
rect 25777 11135 25835 11141
rect 25777 11132 25789 11135
rect 25096 11104 25789 11132
rect 25096 11092 25102 11104
rect 25777 11101 25789 11104
rect 25823 11132 25835 11135
rect 26050 11132 26056 11144
rect 25823 11104 26056 11132
rect 25823 11101 25835 11104
rect 25777 11095 25835 11101
rect 26050 11092 26056 11104
rect 26108 11092 26114 11144
rect 27154 11092 27160 11144
rect 27212 11132 27218 11144
rect 27341 11135 27399 11141
rect 27341 11132 27353 11135
rect 27212 11104 27353 11132
rect 27212 11092 27218 11104
rect 27341 11101 27353 11104
rect 27387 11101 27399 11135
rect 27341 11095 27399 11101
rect 30190 11092 30196 11144
rect 30248 11132 30254 11144
rect 30285 11135 30343 11141
rect 30285 11132 30297 11135
rect 30248 11104 30297 11132
rect 30248 11092 30254 11104
rect 30285 11101 30297 11104
rect 30331 11101 30343 11135
rect 32214 11132 32220 11144
rect 32175 11104 32220 11132
rect 30285 11095 30343 11101
rect 32214 11092 32220 11104
rect 32272 11092 32278 11144
rect 32324 11141 32352 11172
rect 32738 11172 33600 11200
rect 32310 11135 32368 11141
rect 32310 11101 32322 11135
rect 32356 11101 32368 11135
rect 32490 11132 32496 11144
rect 32451 11104 32496 11132
rect 32310 11095 32368 11101
rect 32490 11092 32496 11104
rect 32548 11092 32554 11144
rect 32738 11141 32766 11172
rect 33594 11160 33600 11172
rect 33652 11160 33658 11212
rect 32723 11135 32781 11141
rect 32723 11101 32735 11135
rect 32769 11101 32781 11135
rect 32723 11095 32781 11101
rect 33226 11092 33232 11144
rect 33284 11132 33290 11144
rect 33321 11135 33379 11141
rect 33321 11132 33333 11135
rect 33284 11104 33333 11132
rect 33284 11092 33290 11104
rect 33321 11101 33333 11104
rect 33367 11101 33379 11135
rect 33321 11095 33379 11101
rect 33505 11135 33563 11141
rect 33505 11101 33517 11135
rect 33551 11132 33563 11135
rect 33962 11132 33968 11144
rect 33551 11104 33968 11132
rect 33551 11101 33563 11104
rect 33505 11095 33563 11101
rect 33962 11092 33968 11104
rect 34020 11092 34026 11144
rect 34164 11141 34192 11308
rect 36814 11296 36820 11348
rect 36872 11336 36878 11348
rect 37093 11339 37151 11345
rect 37093 11336 37105 11339
rect 36872 11308 37105 11336
rect 36872 11296 36878 11308
rect 37093 11305 37105 11308
rect 37139 11305 37151 11339
rect 40402 11336 40408 11348
rect 37093 11299 37151 11305
rect 38028 11308 40408 11336
rect 36078 11228 36084 11280
rect 36136 11268 36142 11280
rect 38028 11268 38056 11308
rect 40402 11296 40408 11308
rect 40460 11296 40466 11348
rect 36136 11240 38056 11268
rect 36136 11228 36142 11240
rect 34422 11160 34428 11212
rect 34480 11200 34486 11212
rect 35897 11203 35955 11209
rect 34480 11172 35388 11200
rect 34480 11160 34486 11172
rect 34149 11135 34207 11141
rect 34149 11101 34161 11135
rect 34195 11132 34207 11135
rect 34974 11132 34980 11144
rect 34195 11104 34980 11132
rect 34195 11101 34207 11104
rect 34149 11095 34207 11101
rect 34974 11092 34980 11104
rect 35032 11092 35038 11144
rect 35069 11135 35127 11141
rect 35069 11101 35081 11135
rect 35115 11101 35127 11135
rect 35069 11095 35127 11101
rect 24673 11067 24731 11073
rect 24673 11033 24685 11067
rect 24719 11064 24731 11067
rect 25130 11064 25136 11076
rect 24719 11036 25136 11064
rect 24719 11033 24731 11036
rect 24673 11027 24731 11033
rect 25130 11024 25136 11036
rect 25188 11024 25194 11076
rect 25958 11064 25964 11076
rect 25919 11036 25964 11064
rect 25958 11024 25964 11036
rect 26016 11024 26022 11076
rect 26145 11067 26203 11073
rect 26145 11033 26157 11067
rect 26191 11064 26203 11067
rect 26234 11064 26240 11076
rect 26191 11036 26240 11064
rect 26191 11033 26203 11036
rect 26145 11027 26203 11033
rect 26234 11024 26240 11036
rect 26292 11024 26298 11076
rect 26878 11024 26884 11076
rect 26936 11064 26942 11076
rect 27522 11064 27528 11076
rect 26936 11036 27528 11064
rect 26936 11024 26942 11036
rect 27522 11024 27528 11036
rect 27580 11064 27586 11076
rect 28997 11067 29055 11073
rect 28997 11064 29009 11067
rect 27580 11036 29009 11064
rect 27580 11024 27586 11036
rect 28997 11033 29009 11036
rect 29043 11033 29055 11067
rect 28997 11027 29055 11033
rect 32585 11067 32643 11073
rect 32585 11033 32597 11067
rect 32631 11064 32643 11067
rect 33410 11064 33416 11076
rect 32631 11036 33272 11064
rect 33371 11036 33416 11064
rect 32631 11033 32643 11036
rect 32585 11027 32643 11033
rect 29178 10996 29184 11008
rect 24596 10968 29184 10996
rect 29178 10956 29184 10968
rect 29236 10956 29242 11008
rect 29362 10956 29368 11008
rect 29420 10996 29426 11008
rect 29914 10996 29920 11008
rect 29420 10968 29920 10996
rect 29420 10956 29426 10968
rect 29914 10956 29920 10968
rect 29972 10956 29978 11008
rect 33244 10996 33272 11036
rect 33410 11024 33416 11036
rect 33468 11024 33474 11076
rect 34606 11064 34612 11076
rect 33520 11036 34612 11064
rect 33520 10996 33548 11036
rect 34606 11024 34612 11036
rect 34664 11024 34670 11076
rect 35084 11064 35112 11095
rect 35158 11092 35164 11144
rect 35216 11132 35222 11144
rect 35360 11141 35388 11172
rect 35897 11169 35909 11203
rect 35943 11200 35955 11203
rect 37366 11200 37372 11212
rect 35943 11172 37372 11200
rect 35943 11169 35955 11172
rect 35897 11163 35955 11169
rect 37366 11160 37372 11172
rect 37424 11160 37430 11212
rect 35345 11135 35403 11141
rect 35216 11104 35261 11132
rect 35216 11092 35222 11104
rect 35345 11101 35357 11135
rect 35391 11101 35403 11135
rect 35345 11095 35403 11101
rect 35802 11092 35808 11144
rect 35860 11132 35866 11144
rect 38933 11135 38991 11141
rect 38933 11132 38945 11135
rect 35860 11104 38945 11132
rect 35860 11092 35866 11104
rect 38933 11101 38945 11104
rect 38979 11132 38991 11135
rect 39022 11132 39028 11144
rect 38979 11104 39028 11132
rect 38979 11101 38991 11104
rect 38933 11095 38991 11101
rect 39022 11092 39028 11104
rect 39080 11092 39086 11144
rect 35434 11064 35440 11076
rect 35084 11036 35440 11064
rect 35434 11024 35440 11036
rect 35492 11024 35498 11076
rect 36078 11064 36084 11076
rect 36039 11036 36084 11064
rect 36078 11024 36084 11036
rect 36136 11024 36142 11076
rect 36265 11067 36323 11073
rect 36265 11033 36277 11067
rect 36311 11064 36323 11067
rect 36354 11064 36360 11076
rect 36311 11036 36360 11064
rect 36311 11033 36323 11036
rect 36265 11027 36323 11033
rect 36354 11024 36360 11036
rect 36412 11064 36418 11076
rect 36725 11067 36783 11073
rect 36725 11064 36737 11067
rect 36412 11036 36737 11064
rect 36412 11024 36418 11036
rect 36725 11033 36737 11036
rect 36771 11033 36783 11067
rect 36906 11064 36912 11076
rect 36867 11036 36912 11064
rect 36725 11027 36783 11033
rect 36906 11024 36912 11036
rect 36964 11064 36970 11076
rect 36964 11036 37228 11064
rect 36964 11024 36970 11036
rect 34698 10996 34704 11008
rect 33244 10968 33548 10996
rect 34659 10968 34704 10996
rect 34698 10956 34704 10968
rect 34756 10956 34762 11008
rect 37200 10996 37228 11036
rect 37274 11024 37280 11076
rect 37332 11064 37338 11076
rect 38666 11067 38724 11073
rect 38666 11064 38678 11067
rect 37332 11036 38678 11064
rect 37332 11024 37338 11036
rect 38666 11033 38678 11036
rect 38712 11033 38724 11067
rect 38666 11027 38724 11033
rect 37553 10999 37611 11005
rect 37553 10996 37565 10999
rect 37200 10968 37565 10996
rect 37553 10965 37565 10968
rect 37599 10965 37611 10999
rect 37553 10959 37611 10965
rect 1104 10906 68816 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 50294 10906
rect 50346 10854 50358 10906
rect 50410 10854 50422 10906
rect 50474 10854 50486 10906
rect 50538 10854 50550 10906
rect 50602 10854 68816 10906
rect 1104 10832 68816 10854
rect 1397 10795 1455 10801
rect 1397 10761 1409 10795
rect 1443 10792 1455 10795
rect 1486 10792 1492 10804
rect 1443 10764 1492 10792
rect 1443 10761 1455 10764
rect 1397 10755 1455 10761
rect 1486 10752 1492 10764
rect 1544 10752 1550 10804
rect 5074 10752 5080 10804
rect 5132 10792 5138 10804
rect 5169 10795 5227 10801
rect 5169 10792 5181 10795
rect 5132 10764 5181 10792
rect 5132 10752 5138 10764
rect 5169 10761 5181 10764
rect 5215 10761 5227 10795
rect 6822 10792 6828 10804
rect 5169 10755 5227 10761
rect 5920 10764 6828 10792
rect 5920 10668 5948 10764
rect 6822 10752 6828 10764
rect 6880 10752 6886 10804
rect 8481 10795 8539 10801
rect 8481 10761 8493 10795
rect 8527 10792 8539 10795
rect 9858 10792 9864 10804
rect 8527 10764 9864 10792
rect 8527 10761 8539 10764
rect 8481 10755 8539 10761
rect 9858 10752 9864 10764
rect 9916 10752 9922 10804
rect 10226 10792 10232 10804
rect 10187 10764 10232 10792
rect 10226 10752 10232 10764
rect 10284 10752 10290 10804
rect 14553 10795 14611 10801
rect 14553 10792 14565 10795
rect 12452 10764 14565 10792
rect 11698 10724 11704 10736
rect 9600 10696 11704 10724
rect 1765 10659 1823 10665
rect 1765 10625 1777 10659
rect 1811 10656 1823 10659
rect 2498 10656 2504 10668
rect 1811 10628 2504 10656
rect 1811 10625 1823 10628
rect 1765 10619 1823 10625
rect 2498 10616 2504 10628
rect 2556 10616 2562 10668
rect 4706 10656 4712 10668
rect 4667 10628 4712 10656
rect 4706 10616 4712 10628
rect 4764 10656 4770 10668
rect 5399 10659 5457 10665
rect 5399 10656 5411 10659
rect 4764 10628 5411 10656
rect 4764 10616 4770 10628
rect 5399 10625 5411 10628
rect 5445 10625 5457 10659
rect 5534 10656 5540 10668
rect 5495 10628 5540 10656
rect 5399 10619 5457 10625
rect 5534 10616 5540 10628
rect 5592 10616 5598 10668
rect 5626 10616 5632 10668
rect 5684 10656 5690 10668
rect 5813 10659 5871 10665
rect 5684 10628 5729 10656
rect 5684 10616 5690 10628
rect 5813 10625 5825 10659
rect 5859 10656 5871 10659
rect 5902 10656 5908 10668
rect 5859 10628 5908 10656
rect 5859 10625 5871 10628
rect 5813 10619 5871 10625
rect 5902 10616 5908 10628
rect 5960 10616 5966 10668
rect 6641 10659 6699 10665
rect 6641 10625 6653 10659
rect 6687 10656 6699 10659
rect 6822 10656 6828 10668
rect 6687 10628 6828 10656
rect 6687 10625 6699 10628
rect 6641 10619 6699 10625
rect 6822 10616 6828 10628
rect 6880 10616 6886 10668
rect 7098 10656 7104 10668
rect 7059 10628 7104 10656
rect 7098 10616 7104 10628
rect 7156 10616 7162 10668
rect 7374 10665 7380 10668
rect 7368 10619 7380 10665
rect 7432 10656 7438 10668
rect 7432 10628 7468 10656
rect 7374 10616 7380 10619
rect 7432 10616 7438 10628
rect 8478 10616 8484 10668
rect 8536 10656 8542 10668
rect 8846 10656 8852 10668
rect 8536 10628 8852 10656
rect 8536 10616 8542 10628
rect 8846 10616 8852 10628
rect 8904 10656 8910 10668
rect 8941 10659 8999 10665
rect 8941 10656 8953 10659
rect 8904 10628 8953 10656
rect 8904 10616 8910 10628
rect 8941 10625 8953 10628
rect 8987 10625 8999 10659
rect 8941 10619 8999 10625
rect 9125 10659 9183 10665
rect 9125 10625 9137 10659
rect 9171 10656 9183 10659
rect 9490 10656 9496 10668
rect 9171 10628 9496 10656
rect 9171 10625 9183 10628
rect 9125 10619 9183 10625
rect 9490 10616 9496 10628
rect 9548 10616 9554 10668
rect 9600 10665 9628 10696
rect 11698 10684 11704 10696
rect 11756 10684 11762 10736
rect 11790 10684 11796 10736
rect 11848 10724 11854 10736
rect 12342 10724 12348 10736
rect 11848 10696 12348 10724
rect 11848 10684 11854 10696
rect 9585 10659 9643 10665
rect 9585 10625 9597 10659
rect 9631 10625 9643 10659
rect 9585 10619 9643 10625
rect 9674 10616 9680 10668
rect 9732 10656 9738 10668
rect 9769 10659 9827 10665
rect 9769 10656 9781 10659
rect 9732 10628 9781 10656
rect 9732 10616 9738 10628
rect 9769 10625 9781 10628
rect 9815 10625 9827 10659
rect 9769 10619 9827 10625
rect 9861 10659 9919 10665
rect 9861 10625 9873 10659
rect 9907 10625 9919 10659
rect 9861 10619 9919 10625
rect 1857 10591 1915 10597
rect 1857 10557 1869 10591
rect 1903 10588 1915 10591
rect 1946 10588 1952 10600
rect 1903 10560 1952 10588
rect 1903 10557 1915 10560
rect 1857 10551 1915 10557
rect 1946 10548 1952 10560
rect 2004 10548 2010 10600
rect 9876 10588 9904 10619
rect 9950 10616 9956 10668
rect 10008 10656 10014 10668
rect 10778 10656 10784 10668
rect 10008 10628 10053 10656
rect 10739 10628 10784 10656
rect 10008 10616 10014 10628
rect 10778 10616 10784 10628
rect 10836 10616 10842 10668
rect 11146 10616 11152 10668
rect 11204 10656 11210 10668
rect 11882 10656 11888 10668
rect 11204 10628 11888 10656
rect 11204 10616 11210 10628
rect 11882 10616 11888 10628
rect 11940 10616 11946 10668
rect 12066 10656 12072 10668
rect 12027 10628 12072 10656
rect 12066 10616 12072 10628
rect 12124 10616 12130 10668
rect 12176 10665 12204 10696
rect 12342 10684 12348 10696
rect 12400 10684 12406 10736
rect 12161 10659 12219 10665
rect 12161 10625 12173 10659
rect 12207 10625 12219 10659
rect 12161 10619 12219 10625
rect 12250 10616 12256 10668
rect 12308 10656 12314 10668
rect 12452 10656 12480 10764
rect 14553 10761 14565 10764
rect 14599 10792 14611 10795
rect 16942 10792 16948 10804
rect 14599 10764 16948 10792
rect 14599 10761 14611 10764
rect 14553 10755 14611 10761
rect 16942 10752 16948 10764
rect 17000 10752 17006 10804
rect 17221 10795 17279 10801
rect 17221 10761 17233 10795
rect 17267 10792 17279 10795
rect 17310 10792 17316 10804
rect 17267 10764 17316 10792
rect 17267 10761 17279 10764
rect 17221 10755 17279 10761
rect 17310 10752 17316 10764
rect 17368 10752 17374 10804
rect 22186 10752 22192 10804
rect 22244 10792 22250 10804
rect 22373 10795 22431 10801
rect 22373 10792 22385 10795
rect 22244 10764 22385 10792
rect 22244 10752 22250 10764
rect 22373 10761 22385 10764
rect 22419 10761 22431 10795
rect 22373 10755 22431 10761
rect 25317 10795 25375 10801
rect 25317 10761 25329 10795
rect 25363 10792 25375 10795
rect 25958 10792 25964 10804
rect 25363 10764 25964 10792
rect 25363 10761 25375 10764
rect 25317 10755 25375 10761
rect 25958 10752 25964 10764
rect 26016 10752 26022 10804
rect 26050 10752 26056 10804
rect 26108 10752 26114 10804
rect 27430 10792 27436 10804
rect 27391 10764 27436 10792
rect 27430 10752 27436 10764
rect 27488 10752 27494 10804
rect 28350 10752 28356 10804
rect 28408 10792 28414 10804
rect 28408 10764 32352 10792
rect 28408 10752 28414 10764
rect 12529 10727 12587 10733
rect 12529 10693 12541 10727
rect 12575 10724 12587 10727
rect 13418 10727 13476 10733
rect 13418 10724 13430 10727
rect 12575 10696 13430 10724
rect 12575 10693 12587 10696
rect 12529 10687 12587 10693
rect 13418 10693 13430 10696
rect 13464 10693 13476 10727
rect 13418 10687 13476 10693
rect 24204 10727 24262 10733
rect 24204 10693 24216 10727
rect 24250 10724 24262 10727
rect 25777 10727 25835 10733
rect 25777 10724 25789 10727
rect 24250 10696 25789 10724
rect 24250 10693 24262 10696
rect 24204 10687 24262 10693
rect 25777 10693 25789 10696
rect 25823 10693 25835 10727
rect 26068 10724 26096 10752
rect 27065 10727 27123 10733
rect 27065 10724 27077 10727
rect 26068 10696 27077 10724
rect 25777 10687 25835 10693
rect 27065 10693 27077 10696
rect 27111 10693 27123 10727
rect 27065 10687 27123 10693
rect 27249 10727 27307 10733
rect 27249 10693 27261 10727
rect 27295 10724 27307 10727
rect 27706 10724 27712 10736
rect 27295 10696 27712 10724
rect 27295 10693 27307 10696
rect 27249 10687 27307 10693
rect 27706 10684 27712 10696
rect 27764 10724 27770 10736
rect 28902 10724 28908 10736
rect 27764 10696 28908 10724
rect 27764 10684 27770 10696
rect 28902 10684 28908 10696
rect 28960 10684 28966 10736
rect 13170 10656 13176 10668
rect 12308 10628 12480 10656
rect 13131 10628 13176 10656
rect 12308 10616 12314 10628
rect 13170 10616 13176 10628
rect 13228 10616 13234 10668
rect 18417 10659 18475 10665
rect 18417 10625 18429 10659
rect 18463 10656 18475 10659
rect 18506 10656 18512 10668
rect 18463 10628 18512 10656
rect 18463 10625 18475 10628
rect 18417 10619 18475 10625
rect 18506 10616 18512 10628
rect 18564 10616 18570 10668
rect 22189 10659 22247 10665
rect 22189 10625 22201 10659
rect 22235 10656 22247 10659
rect 22278 10656 22284 10668
rect 22235 10628 22284 10656
rect 22235 10625 22247 10628
rect 22189 10619 22247 10625
rect 22278 10616 22284 10628
rect 22336 10616 22342 10668
rect 25314 10616 25320 10668
rect 25372 10656 25378 10668
rect 25590 10656 25596 10668
rect 25372 10628 25596 10656
rect 25372 10616 25378 10628
rect 25590 10616 25596 10628
rect 25648 10656 25654 10668
rect 26053 10659 26111 10665
rect 26053 10656 26065 10659
rect 25648 10628 26065 10656
rect 25648 10616 25654 10628
rect 26053 10625 26065 10628
rect 26099 10625 26111 10659
rect 26053 10619 26111 10625
rect 26145 10659 26203 10665
rect 26145 10625 26157 10659
rect 26191 10625 26203 10659
rect 26145 10619 26203 10625
rect 9876 10560 9996 10588
rect 9968 10532 9996 10560
rect 11606 10548 11612 10600
rect 11664 10588 11670 10600
rect 13188 10588 13216 10616
rect 11664 10560 13216 10588
rect 18141 10591 18199 10597
rect 11664 10548 11670 10560
rect 18141 10557 18153 10591
rect 18187 10588 18199 10591
rect 18322 10588 18328 10600
rect 18187 10560 18328 10588
rect 18187 10557 18199 10560
rect 18141 10551 18199 10557
rect 18322 10548 18328 10560
rect 18380 10548 18386 10600
rect 20441 10591 20499 10597
rect 20441 10557 20453 10591
rect 20487 10588 20499 10591
rect 20530 10588 20536 10600
rect 20487 10560 20536 10588
rect 20487 10557 20499 10560
rect 20441 10551 20499 10557
rect 20530 10548 20536 10560
rect 20588 10548 20594 10600
rect 20717 10591 20775 10597
rect 20717 10557 20729 10591
rect 20763 10588 20775 10591
rect 23382 10588 23388 10600
rect 20763 10560 23388 10588
rect 20763 10557 20775 10560
rect 20717 10551 20775 10557
rect 23382 10548 23388 10560
rect 23440 10548 23446 10600
rect 23937 10591 23995 10597
rect 23937 10557 23949 10591
rect 23983 10557 23995 10591
rect 26160 10588 26188 10619
rect 26234 10616 26240 10668
rect 26292 10656 26298 10668
rect 26292 10628 26337 10656
rect 26292 10616 26298 10628
rect 26418 10616 26424 10668
rect 26476 10656 26482 10668
rect 27893 10659 27951 10665
rect 26476 10628 26521 10656
rect 26476 10616 26482 10628
rect 27893 10625 27905 10659
rect 27939 10656 27951 10659
rect 27982 10656 27988 10668
rect 27939 10628 27988 10656
rect 27939 10625 27951 10628
rect 27893 10619 27951 10625
rect 27982 10616 27988 10628
rect 28040 10616 28046 10668
rect 29007 10665 29035 10764
rect 29089 10727 29147 10733
rect 29089 10693 29101 10727
rect 29135 10724 29147 10727
rect 30098 10724 30104 10736
rect 29135 10696 30104 10724
rect 29135 10693 29147 10696
rect 29089 10687 29147 10693
rect 30098 10684 30104 10696
rect 30156 10684 30162 10736
rect 28992 10659 29050 10665
rect 28992 10625 29004 10659
rect 29038 10625 29050 10659
rect 28992 10619 29050 10625
rect 29181 10659 29239 10665
rect 29181 10625 29193 10659
rect 29227 10625 29239 10659
rect 29362 10656 29368 10668
rect 29323 10628 29368 10656
rect 29181 10619 29239 10625
rect 26786 10588 26792 10600
rect 26160 10560 26792 10588
rect 23937 10551 23995 10557
rect 9950 10480 9956 10532
rect 10008 10480 10014 10532
rect 2498 10452 2504 10464
rect 2459 10424 2504 10452
rect 2498 10412 2504 10424
rect 2556 10412 2562 10464
rect 5442 10412 5448 10464
rect 5500 10452 5506 10464
rect 6457 10455 6515 10461
rect 6457 10452 6469 10455
rect 5500 10424 6469 10452
rect 5500 10412 5506 10424
rect 6457 10421 6469 10424
rect 6503 10421 6515 10455
rect 6457 10415 6515 10421
rect 7282 10412 7288 10464
rect 7340 10452 7346 10464
rect 9033 10455 9091 10461
rect 9033 10452 9045 10455
rect 7340 10424 9045 10452
rect 7340 10412 7346 10424
rect 9033 10421 9045 10424
rect 9079 10421 9091 10455
rect 9033 10415 9091 10421
rect 9122 10412 9128 10464
rect 9180 10452 9186 10464
rect 10870 10452 10876 10464
rect 9180 10424 10876 10452
rect 9180 10412 9186 10424
rect 10870 10412 10876 10424
rect 10928 10412 10934 10464
rect 15194 10452 15200 10464
rect 15155 10424 15200 10452
rect 15194 10412 15200 10424
rect 15252 10412 15258 10464
rect 17310 10412 17316 10464
rect 17368 10452 17374 10464
rect 22646 10452 22652 10464
rect 17368 10424 22652 10452
rect 17368 10412 17374 10424
rect 22646 10412 22652 10424
rect 22704 10412 22710 10464
rect 23014 10412 23020 10464
rect 23072 10452 23078 10464
rect 23201 10455 23259 10461
rect 23201 10452 23213 10455
rect 23072 10424 23213 10452
rect 23072 10412 23078 10424
rect 23201 10421 23213 10424
rect 23247 10452 23259 10455
rect 23290 10452 23296 10464
rect 23247 10424 23296 10452
rect 23247 10421 23259 10424
rect 23201 10415 23259 10421
rect 23290 10412 23296 10424
rect 23348 10412 23354 10464
rect 23952 10452 23980 10551
rect 26786 10548 26792 10560
rect 26844 10548 26850 10600
rect 29196 10588 29224 10619
rect 29362 10616 29368 10628
rect 29420 10616 29426 10668
rect 29454 10616 29460 10668
rect 29512 10656 29518 10668
rect 30193 10659 30251 10665
rect 29512 10628 29557 10656
rect 29512 10616 29518 10628
rect 30193 10625 30205 10659
rect 30239 10625 30251 10659
rect 30374 10656 30380 10668
rect 30335 10628 30380 10656
rect 30193 10619 30251 10625
rect 30208 10588 30236 10619
rect 30374 10616 30380 10628
rect 30432 10616 30438 10668
rect 30990 10665 31018 10764
rect 31113 10727 31171 10733
rect 31113 10693 31125 10727
rect 31159 10724 31171 10727
rect 31938 10724 31944 10736
rect 31159 10696 31944 10724
rect 31159 10693 31171 10696
rect 31113 10687 31171 10693
rect 31938 10684 31944 10696
rect 31996 10684 32002 10736
rect 30977 10659 31035 10665
rect 30977 10625 30989 10659
rect 31023 10625 31035 10659
rect 30977 10619 31035 10625
rect 31205 10659 31263 10665
rect 31205 10625 31217 10659
rect 31251 10625 31263 10659
rect 31205 10619 31263 10625
rect 31388 10659 31446 10665
rect 31388 10625 31400 10659
rect 31434 10625 31446 10659
rect 31388 10619 31446 10625
rect 31220 10588 31248 10619
rect 29196 10560 31248 10588
rect 31404 10588 31432 10619
rect 31478 10616 31484 10668
rect 31536 10656 31542 10668
rect 32324 10665 32352 10764
rect 33042 10752 33048 10804
rect 33100 10792 33106 10804
rect 34057 10795 34115 10801
rect 33100 10764 33916 10792
rect 33100 10752 33106 10764
rect 32401 10727 32459 10733
rect 32401 10693 32413 10727
rect 32447 10724 32459 10727
rect 33134 10724 33140 10736
rect 32447 10696 33140 10724
rect 32447 10693 32459 10696
rect 32401 10687 32459 10693
rect 33134 10684 33140 10696
rect 33192 10684 33198 10736
rect 33888 10733 33916 10764
rect 34057 10761 34069 10795
rect 34103 10792 34115 10795
rect 35158 10792 35164 10804
rect 34103 10764 35164 10792
rect 34103 10761 34115 10764
rect 34057 10755 34115 10761
rect 35158 10752 35164 10764
rect 35216 10752 35222 10804
rect 40402 10792 40408 10804
rect 40363 10764 40408 10792
rect 40402 10752 40408 10764
rect 40460 10752 40466 10804
rect 41325 10795 41383 10801
rect 41325 10761 41337 10795
rect 41371 10792 41383 10795
rect 42426 10792 42432 10804
rect 41371 10764 42432 10792
rect 41371 10761 41383 10764
rect 41325 10755 41383 10761
rect 42426 10752 42432 10764
rect 42484 10752 42490 10804
rect 33689 10727 33747 10733
rect 33689 10693 33701 10727
rect 33735 10724 33747 10727
rect 33873 10727 33931 10733
rect 33735 10696 33824 10724
rect 33735 10693 33747 10696
rect 33689 10687 33747 10693
rect 32309 10659 32367 10665
rect 31536 10628 31581 10656
rect 31536 10616 31542 10628
rect 32309 10625 32321 10659
rect 32355 10625 32367 10659
rect 32309 10619 32367 10625
rect 32493 10659 32551 10665
rect 32493 10625 32505 10659
rect 32539 10625 32551 10659
rect 32493 10619 32551 10625
rect 32677 10659 32735 10665
rect 32677 10625 32689 10659
rect 32723 10656 32735 10659
rect 33594 10656 33600 10668
rect 32723 10628 33600 10656
rect 32723 10625 32735 10628
rect 32677 10619 32735 10625
rect 31754 10588 31760 10600
rect 31404 10560 31760 10588
rect 27154 10480 27160 10532
rect 27212 10520 27218 10532
rect 29196 10520 29224 10560
rect 30834 10520 30840 10532
rect 27212 10492 29224 10520
rect 30795 10492 30840 10520
rect 27212 10480 27218 10492
rect 30834 10480 30840 10492
rect 30892 10480 30898 10532
rect 31220 10520 31248 10560
rect 31754 10548 31760 10560
rect 31812 10548 31818 10600
rect 32508 10588 32536 10619
rect 33594 10616 33600 10628
rect 33652 10616 33658 10668
rect 33796 10600 33824 10696
rect 33873 10693 33885 10727
rect 33919 10693 33931 10727
rect 33873 10687 33931 10693
rect 33778 10588 33784 10600
rect 31956 10560 32536 10588
rect 33060 10560 33784 10588
rect 31956 10520 31984 10560
rect 32122 10520 32128 10532
rect 31220 10492 31984 10520
rect 32083 10492 32128 10520
rect 32122 10480 32128 10492
rect 32180 10480 32186 10532
rect 24210 10452 24216 10464
rect 23952 10424 24216 10452
rect 24210 10412 24216 10424
rect 24268 10412 24274 10464
rect 28074 10452 28080 10464
rect 28035 10424 28080 10452
rect 28074 10412 28080 10424
rect 28132 10412 28138 10464
rect 28810 10452 28816 10464
rect 28771 10424 28816 10452
rect 28810 10412 28816 10424
rect 28868 10412 28874 10464
rect 30282 10452 30288 10464
rect 30243 10424 30288 10452
rect 30282 10412 30288 10424
rect 30340 10412 30346 10464
rect 31110 10412 31116 10464
rect 31168 10452 31174 10464
rect 33060 10452 33088 10560
rect 33778 10548 33784 10560
rect 33836 10548 33842 10600
rect 33888 10520 33916 10687
rect 34698 10684 34704 10736
rect 34756 10724 34762 10736
rect 35722 10727 35780 10733
rect 35722 10724 35734 10727
rect 34756 10696 35734 10724
rect 34756 10684 34762 10696
rect 35722 10693 35734 10696
rect 35768 10693 35780 10727
rect 40420 10724 40448 10752
rect 35722 10687 35780 10693
rect 35820 10696 36492 10724
rect 40420 10696 41184 10724
rect 34790 10616 34796 10668
rect 34848 10656 34854 10668
rect 35820 10656 35848 10696
rect 34848 10628 35848 10656
rect 34848 10616 34854 10628
rect 35894 10616 35900 10668
rect 35952 10656 35958 10668
rect 36464 10665 36492 10696
rect 35989 10659 36047 10665
rect 35989 10656 36001 10659
rect 35952 10628 36001 10656
rect 35952 10616 35958 10628
rect 35989 10625 36001 10628
rect 36035 10625 36047 10659
rect 35989 10619 36047 10625
rect 36449 10659 36507 10665
rect 36449 10625 36461 10659
rect 36495 10625 36507 10659
rect 36449 10619 36507 10625
rect 36630 10616 36636 10668
rect 36688 10656 36694 10668
rect 37182 10656 37188 10668
rect 36688 10628 37188 10656
rect 36688 10616 36694 10628
rect 37182 10616 37188 10628
rect 37240 10656 37246 10668
rect 37737 10659 37795 10665
rect 37737 10656 37749 10659
rect 37240 10628 37749 10656
rect 37240 10616 37246 10628
rect 37737 10625 37749 10628
rect 37783 10625 37795 10659
rect 37737 10619 37795 10625
rect 37918 10616 37924 10668
rect 37976 10656 37982 10668
rect 38013 10659 38071 10665
rect 38013 10656 38025 10659
rect 37976 10628 38025 10656
rect 37976 10616 37982 10628
rect 38013 10625 38025 10628
rect 38059 10625 38071 10659
rect 39022 10656 39028 10668
rect 38983 10628 39028 10656
rect 38013 10619 38071 10625
rect 39022 10616 39028 10628
rect 39080 10616 39086 10668
rect 39114 10616 39120 10668
rect 39172 10656 39178 10668
rect 39281 10659 39339 10665
rect 39281 10656 39293 10659
rect 39172 10628 39293 10656
rect 39172 10616 39178 10628
rect 39281 10625 39293 10628
rect 39327 10625 39339 10659
rect 39281 10619 39339 10625
rect 39850 10616 39856 10668
rect 39908 10656 39914 10668
rect 41156 10665 41184 10696
rect 40865 10659 40923 10665
rect 40865 10656 40877 10659
rect 39908 10628 40877 10656
rect 39908 10616 39914 10628
rect 40865 10625 40877 10628
rect 40911 10625 40923 10659
rect 40865 10619 40923 10625
rect 41141 10659 41199 10665
rect 41141 10625 41153 10659
rect 41187 10625 41199 10659
rect 41141 10619 41199 10625
rect 40954 10588 40960 10600
rect 40915 10560 40960 10588
rect 40954 10548 40960 10560
rect 41012 10548 41018 10600
rect 34609 10523 34667 10529
rect 34609 10520 34621 10523
rect 33888 10492 34621 10520
rect 34609 10489 34621 10492
rect 34655 10489 34667 10523
rect 34609 10483 34667 10489
rect 31168 10424 33088 10452
rect 33229 10455 33287 10461
rect 31168 10412 31174 10424
rect 33229 10421 33241 10455
rect 33275 10452 33287 10455
rect 34238 10452 34244 10464
rect 33275 10424 34244 10452
rect 33275 10421 33287 10424
rect 33229 10415 33287 10421
rect 34238 10412 34244 10424
rect 34296 10452 34302 10464
rect 35342 10452 35348 10464
rect 34296 10424 35348 10452
rect 34296 10412 34302 10424
rect 35342 10412 35348 10424
rect 35400 10412 35406 10464
rect 36354 10412 36360 10464
rect 36412 10452 36418 10464
rect 36633 10455 36691 10461
rect 36633 10452 36645 10455
rect 36412 10424 36645 10452
rect 36412 10412 36418 10424
rect 36633 10421 36645 10424
rect 36679 10421 36691 10455
rect 40862 10452 40868 10464
rect 40823 10424 40868 10452
rect 36633 10415 36691 10421
rect 40862 10412 40868 10424
rect 40920 10412 40926 10464
rect 1104 10362 68816 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 65654 10362
rect 65706 10310 65718 10362
rect 65770 10310 65782 10362
rect 65834 10310 65846 10362
rect 65898 10310 65910 10362
rect 65962 10310 68816 10362
rect 1104 10288 68816 10310
rect 5169 10251 5227 10257
rect 5169 10217 5181 10251
rect 5215 10248 5227 10251
rect 6638 10248 6644 10260
rect 5215 10220 6644 10248
rect 5215 10217 5227 10220
rect 5169 10211 5227 10217
rect 6638 10208 6644 10220
rect 6696 10208 6702 10260
rect 7374 10208 7380 10260
rect 7432 10248 7438 10260
rect 7469 10251 7527 10257
rect 7469 10248 7481 10251
rect 7432 10220 7481 10248
rect 7432 10208 7438 10220
rect 7469 10217 7481 10220
rect 7515 10217 7527 10251
rect 7469 10211 7527 10217
rect 7558 10208 7564 10260
rect 7616 10248 7622 10260
rect 11885 10251 11943 10257
rect 11885 10248 11897 10251
rect 7616 10220 11897 10248
rect 7616 10208 7622 10220
rect 11885 10217 11897 10220
rect 11931 10217 11943 10251
rect 12250 10248 12256 10260
rect 12211 10220 12256 10248
rect 11885 10211 11943 10217
rect 12250 10208 12256 10220
rect 12308 10208 12314 10260
rect 13262 10248 13268 10260
rect 12406 10220 13268 10248
rect 6914 10140 6920 10192
rect 6972 10180 6978 10192
rect 6972 10152 7880 10180
rect 6972 10140 6978 10152
rect 3786 10112 3792 10124
rect 3747 10084 3792 10112
rect 3786 10072 3792 10084
rect 3844 10072 3850 10124
rect 5534 10072 5540 10124
rect 5592 10112 5598 10124
rect 5592 10084 6040 10112
rect 5592 10072 5598 10084
rect 6012 10053 6040 10084
rect 5905 10047 5963 10053
rect 5905 10044 5917 10047
rect 5828 10016 5917 10044
rect 4056 9979 4114 9985
rect 4056 9945 4068 9979
rect 4102 9976 4114 9979
rect 5629 9979 5687 9985
rect 5629 9976 5641 9979
rect 4102 9948 5641 9976
rect 4102 9945 4114 9948
rect 4056 9939 4114 9945
rect 5629 9945 5641 9948
rect 5675 9945 5687 9979
rect 5629 9939 5687 9945
rect 5828 9908 5856 10016
rect 5905 10013 5917 10016
rect 5951 10013 5963 10047
rect 5905 10007 5963 10013
rect 5997 10047 6055 10053
rect 5997 10013 6009 10047
rect 6043 10013 6055 10047
rect 5997 10007 6055 10013
rect 6012 9976 6040 10007
rect 6086 10004 6092 10056
rect 6144 10044 6150 10056
rect 6144 10016 6189 10044
rect 6144 10004 6150 10016
rect 6270 10004 6276 10056
rect 6328 10044 6334 10056
rect 6822 10044 6828 10056
rect 6328 10016 6373 10044
rect 6735 10016 6828 10044
rect 6328 10004 6334 10016
rect 6822 10004 6828 10016
rect 6880 10044 6886 10056
rect 7722 10053 7728 10056
rect 7699 10047 7728 10053
rect 6880 10016 7604 10044
rect 6880 10004 6886 10016
rect 6914 9976 6920 9988
rect 6012 9948 6920 9976
rect 6914 9936 6920 9948
rect 6972 9936 6978 9988
rect 6086 9908 6092 9920
rect 5828 9880 6092 9908
rect 6086 9868 6092 9880
rect 6144 9868 6150 9920
rect 7009 9911 7067 9917
rect 7009 9877 7021 9911
rect 7055 9908 7067 9911
rect 7098 9908 7104 9920
rect 7055 9880 7104 9908
rect 7055 9877 7067 9880
rect 7009 9871 7067 9877
rect 7098 9868 7104 9880
rect 7156 9868 7162 9920
rect 7576 9908 7604 10016
rect 7699 10013 7711 10047
rect 7699 10007 7728 10013
rect 7722 10004 7728 10007
rect 7780 10004 7786 10056
rect 7852 10053 7880 10152
rect 10318 10112 10324 10124
rect 9968 10084 10324 10112
rect 7834 10047 7892 10053
rect 7834 10013 7846 10047
rect 7880 10013 7892 10047
rect 7834 10007 7892 10013
rect 7929 10047 7987 10053
rect 7929 10013 7941 10047
rect 7975 10013 7987 10047
rect 7929 10007 7987 10013
rect 7944 9976 7972 10007
rect 8110 10004 8116 10056
rect 8168 10044 8174 10056
rect 8938 10044 8944 10056
rect 8168 10016 8213 10044
rect 8899 10016 8944 10044
rect 8168 10004 8174 10016
rect 8938 10004 8944 10016
rect 8996 10004 9002 10056
rect 9125 10047 9183 10053
rect 9125 10013 9137 10047
rect 9171 10044 9183 10047
rect 9858 10044 9864 10056
rect 9171 10016 9864 10044
rect 9171 10013 9183 10016
rect 9125 10007 9183 10013
rect 9858 10004 9864 10016
rect 9916 10004 9922 10056
rect 9968 10053 9996 10084
rect 10318 10072 10324 10084
rect 10376 10112 10382 10124
rect 10686 10112 10692 10124
rect 10376 10084 10692 10112
rect 10376 10072 10382 10084
rect 10686 10072 10692 10084
rect 10744 10072 10750 10124
rect 11422 10112 11428 10124
rect 11383 10084 11428 10112
rect 11422 10072 11428 10084
rect 11480 10072 11486 10124
rect 12406 10112 12434 10220
rect 13262 10208 13268 10220
rect 13320 10248 13326 10260
rect 17129 10251 17187 10257
rect 13320 10220 14504 10248
rect 13320 10208 13326 10220
rect 13630 10140 13636 10192
rect 13688 10180 13694 10192
rect 13688 10152 14412 10180
rect 13688 10140 13694 10152
rect 12084 10084 12434 10112
rect 9953 10047 10011 10053
rect 9953 10013 9965 10047
rect 9999 10013 10011 10047
rect 10134 10044 10140 10056
rect 10095 10016 10140 10044
rect 9953 10007 10011 10013
rect 10134 10004 10140 10016
rect 10192 10004 10198 10056
rect 11146 10044 11152 10056
rect 11107 10016 11152 10044
rect 11146 10004 11152 10016
rect 11204 10004 11210 10056
rect 11882 10004 11888 10056
rect 11940 10044 11946 10056
rect 12084 10053 12112 10084
rect 12069 10047 12127 10053
rect 12069 10044 12081 10047
rect 11940 10016 12081 10044
rect 11940 10004 11946 10016
rect 12069 10013 12081 10016
rect 12115 10013 12127 10047
rect 12069 10007 12127 10013
rect 12250 10004 12256 10056
rect 12308 10044 12314 10056
rect 14090 10044 14096 10056
rect 12308 10016 12434 10044
rect 14051 10016 14096 10044
rect 12308 10004 12314 10016
rect 9309 9979 9367 9985
rect 9309 9976 9321 9979
rect 7944 9948 9321 9976
rect 9309 9945 9321 9948
rect 9355 9945 9367 9979
rect 10318 9976 10324 9988
rect 9309 9939 9367 9945
rect 9646 9948 10324 9976
rect 9646 9908 9674 9948
rect 10318 9936 10324 9948
rect 10376 9936 10382 9988
rect 12406 9976 12434 10016
rect 14090 10004 14096 10016
rect 14148 10004 14154 10056
rect 14182 10004 14188 10056
rect 14240 10044 14246 10056
rect 14384 10053 14412 10152
rect 14476 10112 14504 10220
rect 17129 10217 17141 10251
rect 17175 10248 17187 10251
rect 17310 10248 17316 10260
rect 17175 10220 17316 10248
rect 17175 10217 17187 10220
rect 17129 10211 17187 10217
rect 17144 10112 17172 10211
rect 17310 10208 17316 10220
rect 17368 10208 17374 10260
rect 20070 10208 20076 10260
rect 20128 10208 20134 10260
rect 20346 10208 20352 10260
rect 20404 10248 20410 10260
rect 21269 10251 21327 10257
rect 21269 10248 21281 10251
rect 20404 10220 21281 10248
rect 20404 10208 20410 10220
rect 21269 10217 21281 10220
rect 21315 10217 21327 10251
rect 21269 10211 21327 10217
rect 23477 10251 23535 10257
rect 23477 10217 23489 10251
rect 23523 10248 23535 10251
rect 25590 10248 25596 10260
rect 23523 10220 25596 10248
rect 23523 10217 23535 10220
rect 23477 10211 23535 10217
rect 25590 10208 25596 10220
rect 25648 10208 25654 10260
rect 26050 10208 26056 10260
rect 26108 10248 26114 10260
rect 26329 10251 26387 10257
rect 26329 10248 26341 10251
rect 26108 10220 26341 10248
rect 26108 10208 26114 10220
rect 26329 10217 26341 10220
rect 26375 10217 26387 10251
rect 26329 10211 26387 10217
rect 28997 10251 29055 10257
rect 28997 10217 29009 10251
rect 29043 10248 29055 10251
rect 29454 10248 29460 10260
rect 29043 10220 29460 10248
rect 29043 10217 29055 10220
rect 28997 10211 29055 10217
rect 29454 10208 29460 10220
rect 29512 10208 29518 10260
rect 30101 10251 30159 10257
rect 30101 10217 30113 10251
rect 30147 10248 30159 10251
rect 31478 10248 31484 10260
rect 30147 10220 31484 10248
rect 30147 10217 30159 10220
rect 30101 10211 30159 10217
rect 31478 10208 31484 10220
rect 31536 10208 31542 10260
rect 33689 10251 33747 10257
rect 33689 10217 33701 10251
rect 33735 10248 33747 10251
rect 34790 10248 34796 10260
rect 33735 10220 34796 10248
rect 33735 10217 33747 10220
rect 33689 10211 33747 10217
rect 34790 10208 34796 10220
rect 34848 10208 34854 10260
rect 35621 10251 35679 10257
rect 35621 10217 35633 10251
rect 35667 10248 35679 10251
rect 35802 10248 35808 10260
rect 35667 10220 35808 10248
rect 35667 10217 35679 10220
rect 35621 10211 35679 10217
rect 35802 10208 35808 10220
rect 35860 10208 35866 10260
rect 37737 10251 37795 10257
rect 37737 10217 37749 10251
rect 37783 10248 37795 10251
rect 39114 10248 39120 10260
rect 37783 10220 39120 10248
rect 37783 10217 37795 10220
rect 37737 10211 37795 10217
rect 39114 10208 39120 10220
rect 39172 10208 39178 10260
rect 20088 10180 20116 10208
rect 22741 10183 22799 10189
rect 20088 10152 20392 10180
rect 20364 10124 20392 10152
rect 22741 10149 22753 10183
rect 22787 10180 22799 10183
rect 23842 10180 23848 10192
rect 22787 10152 23848 10180
rect 22787 10149 22799 10152
rect 22741 10143 22799 10149
rect 23842 10140 23848 10152
rect 23900 10140 23906 10192
rect 26418 10140 26424 10192
rect 26476 10180 26482 10192
rect 26476 10152 29868 10180
rect 26476 10140 26482 10152
rect 20070 10112 20076 10124
rect 14476 10084 16344 10112
rect 14369 10047 14427 10053
rect 14240 10016 14285 10044
rect 14240 10004 14246 10016
rect 14369 10013 14381 10047
rect 14415 10013 14427 10047
rect 14369 10007 14427 10013
rect 14461 10047 14519 10053
rect 14461 10013 14473 10047
rect 14507 10044 14519 10047
rect 15470 10044 15476 10056
rect 14507 10016 15476 10044
rect 14507 10013 14519 10016
rect 14461 10007 14519 10013
rect 15470 10004 15476 10016
rect 15528 10004 15534 10056
rect 16316 10053 16344 10084
rect 16500 10084 17172 10112
rect 20031 10084 20076 10112
rect 16500 10053 16528 10084
rect 20070 10072 20076 10084
rect 20128 10072 20134 10124
rect 20346 10072 20352 10124
rect 20404 10072 20410 10124
rect 20714 10112 20720 10124
rect 20675 10084 20720 10112
rect 20714 10072 20720 10084
rect 20772 10072 20778 10124
rect 27341 10115 27399 10121
rect 27341 10081 27353 10115
rect 27387 10112 27399 10115
rect 27430 10112 27436 10124
rect 27387 10084 27436 10112
rect 27387 10081 27399 10084
rect 27341 10075 27399 10081
rect 27430 10072 27436 10084
rect 27488 10072 27494 10124
rect 29840 10112 29868 10152
rect 29914 10140 29920 10192
rect 29972 10180 29978 10192
rect 36541 10183 36599 10189
rect 36541 10180 36553 10183
rect 29972 10152 33180 10180
rect 29972 10140 29978 10152
rect 32030 10112 32036 10124
rect 28644 10084 29776 10112
rect 29840 10084 31892 10112
rect 31943 10084 32036 10112
rect 16209 10047 16267 10053
rect 16209 10013 16221 10047
rect 16255 10013 16267 10047
rect 16209 10007 16267 10013
rect 16301 10047 16359 10053
rect 16301 10013 16313 10047
rect 16347 10013 16359 10047
rect 16301 10007 16359 10013
rect 16485 10047 16543 10053
rect 16485 10013 16497 10047
rect 16531 10013 16543 10047
rect 16485 10007 16543 10013
rect 16577 10047 16635 10053
rect 16577 10013 16589 10047
rect 16623 10044 16635 10047
rect 16666 10044 16672 10056
rect 16623 10016 16672 10044
rect 16623 10013 16635 10016
rect 16577 10007 16635 10013
rect 14550 9976 14556 9988
rect 12406 9948 14556 9976
rect 14550 9936 14556 9948
rect 14608 9936 14614 9988
rect 7576 9880 9674 9908
rect 9769 9911 9827 9917
rect 9769 9877 9781 9911
rect 9815 9908 9827 9911
rect 9858 9908 9864 9920
rect 9815 9880 9864 9908
rect 9815 9877 9827 9880
rect 9769 9871 9827 9877
rect 9858 9868 9864 9880
rect 9916 9868 9922 9920
rect 14645 9911 14703 9917
rect 14645 9877 14657 9911
rect 14691 9908 14703 9911
rect 14826 9908 14832 9920
rect 14691 9880 14832 9908
rect 14691 9877 14703 9880
rect 14645 9871 14703 9877
rect 14826 9868 14832 9880
rect 14884 9868 14890 9920
rect 15194 9908 15200 9920
rect 15155 9880 15200 9908
rect 15194 9868 15200 9880
rect 15252 9868 15258 9920
rect 16022 9908 16028 9920
rect 15983 9880 16028 9908
rect 16022 9868 16028 9880
rect 16080 9868 16086 9920
rect 16224 9908 16252 10007
rect 16666 10004 16672 10016
rect 16724 10004 16730 10056
rect 18141 10047 18199 10053
rect 18141 10044 18153 10047
rect 17052 10016 18153 10044
rect 16850 9908 16856 9920
rect 16224 9880 16856 9908
rect 16850 9868 16856 9880
rect 16908 9908 16914 9920
rect 17052 9908 17080 10016
rect 18141 10013 18153 10016
rect 18187 10013 18199 10047
rect 18414 10044 18420 10056
rect 18375 10016 18420 10044
rect 18141 10007 18199 10013
rect 18414 10004 18420 10016
rect 18472 10004 18478 10056
rect 19981 10047 20039 10053
rect 19981 10013 19993 10047
rect 20027 10044 20039 10047
rect 20162 10044 20168 10056
rect 20027 10016 20168 10044
rect 20027 10013 20039 10016
rect 19981 10007 20039 10013
rect 20162 10004 20168 10016
rect 20220 10004 20226 10056
rect 20257 10047 20315 10053
rect 20257 10013 20269 10047
rect 20303 10044 20315 10047
rect 20530 10044 20536 10056
rect 20303 10016 20536 10044
rect 20303 10013 20315 10016
rect 20257 10007 20315 10013
rect 20530 10004 20536 10016
rect 20588 10004 20594 10056
rect 20625 10047 20683 10053
rect 20625 10013 20637 10047
rect 20671 10044 20683 10047
rect 20806 10044 20812 10056
rect 20671 10016 20812 10044
rect 20671 10013 20683 10016
rect 20625 10007 20683 10013
rect 20806 10004 20812 10016
rect 20864 10004 20870 10056
rect 20898 10004 20904 10056
rect 20956 10044 20962 10056
rect 21453 10047 21511 10053
rect 21453 10044 21465 10047
rect 20956 10016 21465 10044
rect 20956 10004 20962 10016
rect 21453 10013 21465 10016
rect 21499 10013 21511 10047
rect 21453 10007 21511 10013
rect 21545 10047 21603 10053
rect 21545 10013 21557 10047
rect 21591 10013 21603 10047
rect 22373 10047 22431 10053
rect 22373 10044 22385 10047
rect 21545 10007 21603 10013
rect 22066 10016 22385 10044
rect 19334 9936 19340 9988
rect 19392 9976 19398 9988
rect 19392 9948 20208 9976
rect 19392 9936 19398 9948
rect 20180 9920 20208 9948
rect 20346 9936 20352 9988
rect 20404 9976 20410 9988
rect 21560 9976 21588 10007
rect 20404 9948 21588 9976
rect 20404 9936 20410 9948
rect 19978 9908 19984 9920
rect 16908 9880 17080 9908
rect 19939 9880 19984 9908
rect 16908 9868 16914 9880
rect 19978 9868 19984 9880
rect 20036 9868 20042 9920
rect 20162 9868 20168 9920
rect 20220 9908 20226 9920
rect 22066 9908 22094 10016
rect 22373 10013 22385 10016
rect 22419 10013 22431 10047
rect 22373 10007 22431 10013
rect 22557 10047 22615 10053
rect 22557 10013 22569 10047
rect 22603 10013 22615 10047
rect 23290 10044 23296 10056
rect 23251 10016 23296 10044
rect 22557 10007 22615 10013
rect 22278 9936 22284 9988
rect 22336 9976 22342 9988
rect 22572 9976 22600 10007
rect 23290 10004 23296 10016
rect 23348 10004 23354 10056
rect 26513 10047 26571 10053
rect 26513 10013 26525 10047
rect 26559 10044 26571 10047
rect 27154 10044 27160 10056
rect 26559 10016 27016 10044
rect 27115 10016 27160 10044
rect 26559 10013 26571 10016
rect 26513 10007 26571 10013
rect 26988 9985 27016 10016
rect 27154 10004 27160 10016
rect 27212 10004 27218 10056
rect 27801 10047 27859 10053
rect 27801 10013 27813 10047
rect 27847 10013 27859 10047
rect 28442 10044 28448 10056
rect 28403 10016 28448 10044
rect 27801 10007 27859 10013
rect 22336 9948 22600 9976
rect 26973 9979 27031 9985
rect 22336 9936 22342 9948
rect 26973 9945 26985 9979
rect 27019 9976 27031 9979
rect 27816 9976 27844 10007
rect 28442 10004 28448 10016
rect 28500 10004 28506 10056
rect 28534 10004 28540 10056
rect 28592 10044 28598 10056
rect 28644 10053 28672 10084
rect 28629 10047 28687 10053
rect 28629 10044 28641 10047
rect 28592 10016 28641 10044
rect 28592 10004 28598 10016
rect 28629 10013 28641 10016
rect 28675 10013 28687 10047
rect 28629 10007 28687 10013
rect 28813 10047 28871 10053
rect 28813 10013 28825 10047
rect 28859 10044 28871 10047
rect 28859 10016 28948 10044
rect 28859 10013 28871 10016
rect 28813 10007 28871 10013
rect 28718 9976 28724 9988
rect 27019 9948 27844 9976
rect 28679 9948 28724 9976
rect 27019 9945 27031 9948
rect 26973 9939 27031 9945
rect 28718 9936 28724 9948
rect 28776 9936 28782 9988
rect 28920 9976 28948 10016
rect 28994 10004 29000 10056
rect 29052 10044 29058 10056
rect 29748 10053 29776 10084
rect 29549 10047 29607 10053
rect 29549 10044 29561 10047
rect 29052 10016 29561 10044
rect 29052 10004 29058 10016
rect 29549 10013 29561 10016
rect 29595 10013 29607 10047
rect 29549 10007 29607 10013
rect 29733 10047 29791 10053
rect 29733 10013 29745 10047
rect 29779 10013 29791 10047
rect 29914 10044 29920 10056
rect 29875 10016 29920 10044
rect 29733 10007 29791 10013
rect 29914 10004 29920 10016
rect 29972 10004 29978 10056
rect 30653 10047 30711 10053
rect 30653 10013 30665 10047
rect 30699 10044 30711 10047
rect 31202 10044 31208 10056
rect 30699 10016 31208 10044
rect 30699 10013 30711 10016
rect 30653 10007 30711 10013
rect 31202 10004 31208 10016
rect 31260 10004 31266 10056
rect 31297 10047 31355 10053
rect 31297 10013 31309 10047
rect 31343 10044 31355 10047
rect 31754 10044 31760 10056
rect 31343 10016 31760 10044
rect 31343 10013 31355 10016
rect 31297 10007 31355 10013
rect 31754 10004 31760 10016
rect 31812 10004 31818 10056
rect 31864 10044 31892 10084
rect 32030 10072 32036 10084
rect 32088 10112 32094 10124
rect 32582 10112 32588 10124
rect 32088 10084 32588 10112
rect 32088 10072 32094 10084
rect 32582 10072 32588 10084
rect 32640 10072 32646 10124
rect 33152 10044 33180 10152
rect 35866 10152 36553 10180
rect 33318 10112 33324 10124
rect 33279 10084 33324 10112
rect 33318 10072 33324 10084
rect 33376 10072 33382 10124
rect 33686 10072 33692 10124
rect 33744 10112 33750 10124
rect 35866 10112 35894 10152
rect 36541 10149 36553 10152
rect 36587 10180 36599 10183
rect 36587 10152 37688 10180
rect 36587 10149 36599 10152
rect 36541 10143 36599 10149
rect 37550 10112 37556 10124
rect 33744 10084 35894 10112
rect 37108 10084 37556 10112
rect 33744 10072 33750 10084
rect 33502 10044 33508 10056
rect 31864 10016 32076 10044
rect 33152 10016 33508 10044
rect 29178 9976 29184 9988
rect 28920 9948 29184 9976
rect 29178 9936 29184 9948
rect 29236 9936 29242 9988
rect 29822 9936 29828 9988
rect 29880 9976 29886 9988
rect 31110 9976 31116 9988
rect 29880 9948 29925 9976
rect 31023 9948 31116 9976
rect 29880 9936 29886 9948
rect 31110 9936 31116 9948
rect 31168 9936 31174 9988
rect 25130 9908 25136 9920
rect 20220 9880 22094 9908
rect 25043 9880 25136 9908
rect 20220 9868 20226 9880
rect 25130 9868 25136 9880
rect 25188 9908 25194 9920
rect 25314 9908 25320 9920
rect 25188 9880 25320 9908
rect 25188 9868 25194 9880
rect 25314 9868 25320 9880
rect 25372 9868 25378 9920
rect 27985 9911 28043 9917
rect 27985 9877 27997 9911
rect 28031 9908 28043 9911
rect 29914 9908 29920 9920
rect 28031 9880 29920 9908
rect 28031 9877 28043 9880
rect 27985 9871 28043 9877
rect 29914 9868 29920 9880
rect 29972 9908 29978 9920
rect 31128 9908 31156 9936
rect 29972 9880 31156 9908
rect 31481 9911 31539 9917
rect 29972 9868 29978 9880
rect 31481 9877 31493 9911
rect 31527 9908 31539 9911
rect 31938 9908 31944 9920
rect 31527 9880 31944 9908
rect 31527 9877 31539 9880
rect 31481 9871 31539 9877
rect 31938 9868 31944 9880
rect 31996 9868 32002 9920
rect 32048 9908 32076 10016
rect 33502 10004 33508 10016
rect 33560 10004 33566 10056
rect 33778 10004 33784 10056
rect 33836 10044 33842 10056
rect 34698 10044 34704 10056
rect 33836 10016 34704 10044
rect 33836 10004 33842 10016
rect 34698 10004 34704 10016
rect 34756 10004 34762 10056
rect 37108 10053 37136 10084
rect 37550 10072 37556 10084
rect 37608 10072 37614 10124
rect 37093 10047 37151 10053
rect 37093 10013 37105 10047
rect 37139 10013 37151 10047
rect 37274 10044 37280 10056
rect 37235 10016 37280 10044
rect 37093 10007 37151 10013
rect 37274 10004 37280 10016
rect 37332 10004 37338 10056
rect 37369 10047 37427 10053
rect 37369 10013 37381 10047
rect 37415 10013 37427 10047
rect 37369 10007 37427 10013
rect 37461 10047 37519 10053
rect 37461 10013 37473 10047
rect 37507 10044 37519 10047
rect 37660 10044 37688 10152
rect 68094 10044 68100 10056
rect 37507 10016 37688 10044
rect 68055 10016 68100 10044
rect 37507 10013 37519 10016
rect 37461 10007 37519 10013
rect 34790 9936 34796 9988
rect 34848 9976 34854 9988
rect 34885 9979 34943 9985
rect 34885 9976 34897 9979
rect 34848 9948 34897 9976
rect 34848 9936 34854 9948
rect 34885 9945 34897 9948
rect 34931 9945 34943 9979
rect 34885 9939 34943 9945
rect 37182 9936 37188 9988
rect 37240 9976 37246 9988
rect 37384 9976 37412 10007
rect 68094 10004 68100 10016
rect 68152 10004 68158 10056
rect 37240 9948 37412 9976
rect 37240 9936 37246 9948
rect 32263 9911 32321 9917
rect 32263 9908 32275 9911
rect 32048 9880 32275 9908
rect 32263 9877 32275 9880
rect 32309 9908 32321 9911
rect 33870 9908 33876 9920
rect 32309 9880 33876 9908
rect 32309 9877 32321 9880
rect 32263 9871 32321 9877
rect 33870 9868 33876 9880
rect 33928 9868 33934 9920
rect 35066 9908 35072 9920
rect 35027 9880 35072 9908
rect 35066 9868 35072 9880
rect 35124 9868 35130 9920
rect 38194 9908 38200 9920
rect 38155 9880 38200 9908
rect 38194 9868 38200 9880
rect 38252 9868 38258 9920
rect 39298 9868 39304 9920
rect 39356 9908 39362 9920
rect 39850 9908 39856 9920
rect 39356 9880 39856 9908
rect 39356 9868 39362 9880
rect 39850 9868 39856 9880
rect 39908 9908 39914 9920
rect 40681 9911 40739 9917
rect 40681 9908 40693 9911
rect 39908 9880 40693 9908
rect 39908 9868 39914 9880
rect 40681 9877 40693 9880
rect 40727 9877 40739 9911
rect 40681 9871 40739 9877
rect 1104 9818 68816 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 50294 9818
rect 50346 9766 50358 9818
rect 50410 9766 50422 9818
rect 50474 9766 50486 9818
rect 50538 9766 50550 9818
rect 50602 9766 68816 9818
rect 1104 9744 68816 9766
rect 5166 9664 5172 9716
rect 5224 9704 5230 9716
rect 12250 9704 12256 9716
rect 5224 9676 12256 9704
rect 5224 9664 5230 9676
rect 12250 9664 12256 9676
rect 12308 9664 12314 9716
rect 14550 9664 14556 9716
rect 14608 9704 14614 9716
rect 20530 9704 20536 9716
rect 14608 9676 16988 9704
rect 20491 9676 20536 9704
rect 14608 9664 14614 9676
rect 4985 9639 5043 9645
rect 4985 9605 4997 9639
rect 5031 9636 5043 9639
rect 6086 9636 6092 9648
rect 5031 9608 6092 9636
rect 5031 9605 5043 9608
rect 4985 9599 5043 9605
rect 6086 9596 6092 9608
rect 6144 9596 6150 9648
rect 7745 9639 7803 9645
rect 7745 9605 7757 9639
rect 7791 9636 7803 9639
rect 8294 9636 8300 9648
rect 7791 9608 8300 9636
rect 7791 9605 7803 9608
rect 7745 9599 7803 9605
rect 8294 9596 8300 9608
rect 8352 9636 8358 9648
rect 9125 9639 9183 9645
rect 9125 9636 9137 9639
rect 8352 9608 9137 9636
rect 8352 9596 8358 9608
rect 9125 9605 9137 9608
rect 9171 9636 9183 9639
rect 11422 9636 11428 9648
rect 9171 9608 11428 9636
rect 9171 9605 9183 9608
rect 9125 9599 9183 9605
rect 11422 9596 11428 9608
rect 11480 9596 11486 9648
rect 15194 9636 15200 9648
rect 14292 9608 15200 9636
rect 5442 9568 5448 9580
rect 5403 9540 5448 9568
rect 5442 9528 5448 9540
rect 5500 9528 5506 9580
rect 5629 9571 5687 9577
rect 5629 9537 5641 9571
rect 5675 9568 5687 9571
rect 5718 9568 5724 9580
rect 5675 9540 5724 9568
rect 5675 9537 5687 9540
rect 5629 9531 5687 9537
rect 4433 9503 4491 9509
rect 4433 9469 4445 9503
rect 4479 9500 4491 9503
rect 5644 9500 5672 9531
rect 5718 9528 5724 9540
rect 5776 9528 5782 9580
rect 6914 9568 6920 9580
rect 6875 9540 6920 9568
rect 6914 9528 6920 9540
rect 6972 9528 6978 9580
rect 9585 9571 9643 9577
rect 9585 9537 9597 9571
rect 9631 9568 9643 9571
rect 9674 9568 9680 9580
rect 9631 9540 9680 9568
rect 9631 9537 9643 9540
rect 9585 9531 9643 9537
rect 9674 9528 9680 9540
rect 9732 9528 9738 9580
rect 9766 9528 9772 9580
rect 9824 9568 9830 9580
rect 9953 9571 10011 9577
rect 9824 9540 9869 9568
rect 9824 9528 9830 9540
rect 9953 9537 9965 9571
rect 9999 9568 10011 9571
rect 10318 9568 10324 9580
rect 9999 9540 10324 9568
rect 9999 9537 10011 9540
rect 9953 9531 10011 9537
rect 10318 9528 10324 9540
rect 10376 9528 10382 9580
rect 10502 9568 10508 9580
rect 10428 9540 10508 9568
rect 4479 9472 5672 9500
rect 4479 9469 4491 9472
rect 4433 9463 4491 9469
rect 6546 9460 6552 9512
rect 6604 9500 6610 9512
rect 7193 9503 7251 9509
rect 7193 9500 7205 9503
rect 6604 9472 7205 9500
rect 6604 9460 6610 9472
rect 7193 9469 7205 9472
rect 7239 9500 7251 9503
rect 7282 9500 7288 9512
rect 7239 9472 7288 9500
rect 7239 9469 7251 9472
rect 7193 9463 7251 9469
rect 7282 9460 7288 9472
rect 7340 9460 7346 9512
rect 8389 9503 8447 9509
rect 8389 9469 8401 9503
rect 8435 9500 8447 9503
rect 8754 9500 8760 9512
rect 8435 9472 8760 9500
rect 8435 9469 8447 9472
rect 8389 9463 8447 9469
rect 8754 9460 8760 9472
rect 8812 9460 8818 9512
rect 7098 9392 7104 9444
rect 7156 9432 7162 9444
rect 10428 9432 10456 9540
rect 10502 9528 10508 9540
rect 10560 9568 10566 9580
rect 10597 9571 10655 9577
rect 10597 9568 10609 9571
rect 10560 9540 10609 9568
rect 10560 9528 10566 9540
rect 10597 9537 10609 9540
rect 10643 9537 10655 9571
rect 10778 9568 10784 9580
rect 10739 9540 10784 9568
rect 10597 9531 10655 9537
rect 10778 9528 10784 9540
rect 10836 9528 10842 9580
rect 11146 9568 11152 9580
rect 10888 9540 11152 9568
rect 7156 9404 10456 9432
rect 7156 9392 7162 9404
rect 5626 9324 5632 9376
rect 5684 9364 5690 9376
rect 5813 9367 5871 9373
rect 5813 9364 5825 9367
rect 5684 9336 5825 9364
rect 5684 9324 5690 9336
rect 5813 9333 5825 9336
rect 5859 9333 5871 9367
rect 5813 9327 5871 9333
rect 7742 9324 7748 9376
rect 7800 9364 7806 9376
rect 10888 9364 10916 9540
rect 11146 9528 11152 9540
rect 11204 9568 11210 9580
rect 11780 9577 11838 9583
rect 11974 9577 11980 9580
rect 11517 9571 11575 9577
rect 11517 9568 11529 9571
rect 11204 9540 11529 9568
rect 11204 9528 11210 9540
rect 11517 9537 11529 9540
rect 11563 9537 11575 9571
rect 11680 9571 11738 9577
rect 11680 9568 11692 9571
rect 11517 9531 11575 9537
rect 11624 9540 11692 9568
rect 10965 9503 11023 9509
rect 10965 9469 10977 9503
rect 11011 9500 11023 9503
rect 11624 9500 11652 9540
rect 11680 9537 11692 9540
rect 11726 9537 11738 9571
rect 11780 9543 11792 9577
rect 11826 9568 11838 9577
rect 11931 9571 11980 9577
rect 11826 9543 11839 9568
rect 11780 9537 11839 9543
rect 11680 9531 11738 9537
rect 11011 9472 11652 9500
rect 11011 9469 11023 9472
rect 10965 9463 11023 9469
rect 11811 9444 11839 9537
rect 11931 9537 11943 9571
rect 11977 9537 11980 9571
rect 11931 9531 11980 9537
rect 11974 9528 11980 9531
rect 12032 9528 12038 9580
rect 14292 9577 14320 9608
rect 15194 9596 15200 9608
rect 15252 9596 15258 9648
rect 14277 9571 14335 9577
rect 14277 9568 14289 9571
rect 12636 9540 14289 9568
rect 12636 9500 12664 9540
rect 14277 9537 14289 9540
rect 14323 9537 14335 9571
rect 14734 9568 14740 9580
rect 14695 9540 14740 9568
rect 14277 9531 14335 9537
rect 14734 9528 14740 9540
rect 14792 9528 14798 9580
rect 14921 9571 14979 9577
rect 14921 9537 14933 9571
rect 14967 9568 14979 9571
rect 15289 9571 15347 9577
rect 14967 9540 15240 9568
rect 14967 9537 14979 9540
rect 14921 9531 14979 9537
rect 11992 9472 12664 9500
rect 11790 9392 11796 9444
rect 11848 9392 11854 9444
rect 7800 9336 10916 9364
rect 7800 9324 7806 9336
rect 11422 9324 11428 9376
rect 11480 9364 11486 9376
rect 11992 9364 12020 9472
rect 12710 9460 12716 9512
rect 12768 9500 12774 9512
rect 13449 9503 13507 9509
rect 13449 9500 13461 9503
rect 12768 9472 13461 9500
rect 12768 9460 12774 9472
rect 13449 9469 13461 9472
rect 13495 9469 13507 9503
rect 13449 9463 13507 9469
rect 14826 9460 14832 9512
rect 14884 9500 14890 9512
rect 15007 9503 15065 9509
rect 15007 9500 15019 9503
rect 14884 9472 15019 9500
rect 14884 9460 14890 9472
rect 15007 9469 15019 9472
rect 15053 9469 15065 9503
rect 15007 9463 15065 9469
rect 15105 9503 15163 9509
rect 15105 9469 15117 9503
rect 15151 9469 15163 9503
rect 15212 9500 15240 9540
rect 15289 9537 15301 9571
rect 15335 9568 15347 9571
rect 15470 9568 15476 9580
rect 15335 9540 15476 9568
rect 15335 9537 15347 9540
rect 15289 9531 15347 9537
rect 15470 9528 15476 9540
rect 15528 9528 15534 9580
rect 16850 9568 16856 9580
rect 16811 9540 16856 9568
rect 16850 9528 16856 9540
rect 16908 9528 16914 9580
rect 16960 9577 16988 9676
rect 20530 9664 20536 9676
rect 20588 9664 20594 9716
rect 20806 9664 20812 9716
rect 20864 9664 20870 9716
rect 25593 9707 25651 9713
rect 25593 9673 25605 9707
rect 25639 9704 25651 9707
rect 25682 9704 25688 9716
rect 25639 9676 25688 9704
rect 25639 9673 25651 9676
rect 25593 9667 25651 9673
rect 25682 9664 25688 9676
rect 25740 9664 25746 9716
rect 26421 9707 26479 9713
rect 26421 9673 26433 9707
rect 26467 9704 26479 9707
rect 27430 9704 27436 9716
rect 26467 9676 27436 9704
rect 26467 9673 26479 9676
rect 26421 9667 26479 9673
rect 18414 9596 18420 9648
rect 18472 9636 18478 9648
rect 19337 9639 19395 9645
rect 19337 9636 19349 9639
rect 18472 9608 19349 9636
rect 18472 9596 18478 9608
rect 19337 9605 19349 9608
rect 19383 9605 19395 9639
rect 20824 9636 20852 9664
rect 21266 9636 21272 9648
rect 19337 9599 19395 9605
rect 20732 9608 21272 9636
rect 16945 9571 17003 9577
rect 16945 9537 16957 9571
rect 16991 9537 17003 9571
rect 17126 9568 17132 9580
rect 17087 9540 17132 9568
rect 16945 9531 17003 9537
rect 17126 9528 17132 9540
rect 17184 9528 17190 9580
rect 17218 9528 17224 9580
rect 17276 9568 17282 9580
rect 18509 9571 18567 9577
rect 17276 9540 17321 9568
rect 17276 9528 17282 9540
rect 18509 9537 18521 9571
rect 18555 9537 18567 9571
rect 18509 9531 18567 9537
rect 18693 9571 18751 9577
rect 18693 9537 18705 9571
rect 18739 9537 18751 9571
rect 18693 9531 18751 9537
rect 15212 9472 18368 9500
rect 15105 9463 15163 9469
rect 12526 9392 12532 9444
rect 12584 9432 12590 9444
rect 15120 9432 15148 9463
rect 12584 9404 15148 9432
rect 12584 9392 12590 9404
rect 15378 9392 15384 9444
rect 15436 9432 15442 9444
rect 16669 9435 16727 9441
rect 16669 9432 16681 9435
rect 15436 9404 16681 9432
rect 15436 9392 15442 9404
rect 16669 9401 16681 9404
rect 16715 9401 16727 9435
rect 18230 9432 18236 9444
rect 18191 9404 18236 9432
rect 16669 9395 16727 9401
rect 18230 9392 18236 9404
rect 18288 9392 18294 9444
rect 12158 9364 12164 9376
rect 11480 9336 12020 9364
rect 12119 9336 12164 9364
rect 11480 9324 11486 9336
rect 12158 9324 12164 9336
rect 12216 9324 12222 9376
rect 15473 9367 15531 9373
rect 15473 9333 15485 9367
rect 15519 9364 15531 9367
rect 15654 9364 15660 9376
rect 15519 9336 15660 9364
rect 15519 9333 15531 9336
rect 15473 9327 15531 9333
rect 15654 9324 15660 9336
rect 15712 9324 15718 9376
rect 18340 9364 18368 9472
rect 18524 9444 18552 9531
rect 18708 9500 18736 9531
rect 18782 9528 18788 9580
rect 18840 9568 18846 9580
rect 19521 9571 19579 9577
rect 18840 9540 18885 9568
rect 18840 9528 18846 9540
rect 19521 9537 19533 9571
rect 19567 9568 19579 9571
rect 19978 9568 19984 9580
rect 19567 9540 19984 9568
rect 19567 9537 19579 9540
rect 19521 9531 19579 9537
rect 19334 9500 19340 9512
rect 18708 9472 19340 9500
rect 19334 9460 19340 9472
rect 19392 9500 19398 9512
rect 19536 9500 19564 9531
rect 19978 9528 19984 9540
rect 20036 9528 20042 9580
rect 20732 9577 20760 9608
rect 21266 9596 21272 9608
rect 21324 9596 21330 9648
rect 22554 9636 22560 9648
rect 22515 9608 22560 9636
rect 22554 9596 22560 9608
rect 22612 9596 22618 9648
rect 24486 9645 24492 9648
rect 24480 9636 24492 9645
rect 23400 9608 24164 9636
rect 24447 9608 24492 9636
rect 23400 9580 23428 9608
rect 20717 9571 20775 9577
rect 20717 9537 20729 9571
rect 20763 9537 20775 9571
rect 20717 9531 20775 9537
rect 20806 9528 20812 9580
rect 20864 9568 20870 9580
rect 22189 9571 22247 9577
rect 22189 9568 22201 9571
rect 20864 9540 22201 9568
rect 20864 9528 20870 9540
rect 22189 9537 22201 9540
rect 22235 9537 22247 9571
rect 22189 9531 22247 9537
rect 22278 9528 22284 9580
rect 22336 9568 22342 9580
rect 22373 9571 22431 9577
rect 22373 9568 22385 9571
rect 22336 9540 22385 9568
rect 22336 9528 22342 9540
rect 22373 9537 22385 9540
rect 22419 9537 22431 9571
rect 23382 9568 23388 9580
rect 23295 9540 23388 9568
rect 22373 9531 22431 9537
rect 23382 9528 23388 9540
rect 23440 9528 23446 9580
rect 23569 9571 23627 9577
rect 23569 9537 23581 9571
rect 23615 9568 23627 9571
rect 24026 9568 24032 9580
rect 23615 9540 24032 9568
rect 23615 9537 23627 9540
rect 23569 9531 23627 9537
rect 24026 9528 24032 9540
rect 24084 9528 24090 9580
rect 24136 9568 24164 9608
rect 24480 9599 24492 9608
rect 24486 9596 24492 9599
rect 24544 9596 24550 9648
rect 26436 9568 26464 9667
rect 27430 9664 27436 9676
rect 27488 9664 27494 9716
rect 34422 9704 34428 9716
rect 33888 9676 34428 9704
rect 30282 9636 30288 9648
rect 27908 9608 30288 9636
rect 24136 9540 26464 9568
rect 26786 9528 26792 9580
rect 26844 9568 26850 9580
rect 27908 9577 27936 9608
rect 27617 9571 27675 9577
rect 27617 9568 27629 9571
rect 26844 9540 27629 9568
rect 26844 9528 26850 9540
rect 27617 9537 27629 9540
rect 27663 9537 27675 9571
rect 27617 9531 27675 9537
rect 27893 9571 27951 9577
rect 27893 9537 27905 9571
rect 27939 9537 27951 9571
rect 29086 9568 29092 9580
rect 29047 9540 29092 9568
rect 27893 9531 27951 9537
rect 29086 9528 29092 9540
rect 29144 9528 29150 9580
rect 29270 9568 29276 9580
rect 29231 9540 29276 9568
rect 29270 9528 29276 9540
rect 29328 9528 29334 9580
rect 29380 9577 29408 9608
rect 30282 9596 30288 9608
rect 30340 9596 30346 9648
rect 30558 9636 30564 9648
rect 30392 9608 30564 9636
rect 29365 9571 29423 9577
rect 29365 9537 29377 9571
rect 29411 9537 29423 9571
rect 29365 9531 29423 9537
rect 29457 9571 29515 9577
rect 29457 9537 29469 9571
rect 29503 9568 29515 9571
rect 30392 9568 30420 9608
rect 30558 9596 30564 9608
rect 30616 9636 30622 9648
rect 33686 9636 33692 9648
rect 30616 9608 33692 9636
rect 30616 9596 30622 9608
rect 33686 9596 33692 9608
rect 33744 9596 33750 9648
rect 33888 9580 33916 9676
rect 34422 9664 34428 9676
rect 34480 9664 34486 9716
rect 35066 9636 35072 9648
rect 34072 9608 35072 9636
rect 30742 9568 30748 9580
rect 29503 9540 30420 9568
rect 30655 9540 30748 9568
rect 29503 9537 29515 9540
rect 29457 9531 29515 9537
rect 19392 9472 19564 9500
rect 19705 9503 19763 9509
rect 19392 9460 19398 9472
rect 19705 9469 19717 9503
rect 19751 9500 19763 9503
rect 20990 9500 20996 9512
rect 19751 9472 20996 9500
rect 19751 9469 19763 9472
rect 19705 9463 19763 9469
rect 18506 9432 18512 9444
rect 18419 9404 18512 9432
rect 18506 9392 18512 9404
rect 18564 9432 18570 9444
rect 19720 9432 19748 9463
rect 20990 9460 20996 9472
rect 21048 9460 21054 9512
rect 24210 9500 24216 9512
rect 24171 9472 24216 9500
rect 24210 9460 24216 9472
rect 24268 9460 24274 9512
rect 28629 9503 28687 9509
rect 28629 9469 28641 9503
rect 28675 9500 28687 9503
rect 29472 9500 29500 9531
rect 30742 9528 30748 9540
rect 30800 9568 30806 9580
rect 33045 9571 33103 9577
rect 30800 9540 31754 9568
rect 30800 9528 30806 9540
rect 31021 9503 31079 9509
rect 31021 9500 31033 9503
rect 28675 9472 29500 9500
rect 30208 9472 31033 9500
rect 28675 9469 28687 9472
rect 28629 9463 28687 9469
rect 18564 9404 19748 9432
rect 18564 9392 18570 9404
rect 29086 9392 29092 9444
rect 29144 9432 29150 9444
rect 30208 9432 30236 9472
rect 31021 9469 31033 9472
rect 31067 9500 31079 9503
rect 31110 9500 31116 9512
rect 31067 9472 31116 9500
rect 31067 9469 31079 9472
rect 31021 9463 31079 9469
rect 31110 9460 31116 9472
rect 31168 9460 31174 9512
rect 31726 9500 31754 9540
rect 33045 9537 33057 9571
rect 33091 9568 33103 9571
rect 33502 9568 33508 9580
rect 33091 9540 33508 9568
rect 33091 9537 33103 9540
rect 33045 9531 33103 9537
rect 33502 9528 33508 9540
rect 33560 9568 33566 9580
rect 33560 9540 33824 9568
rect 33560 9528 33566 9540
rect 32030 9500 32036 9512
rect 31726 9472 32036 9500
rect 32030 9460 32036 9472
rect 32088 9460 32094 9512
rect 33321 9503 33379 9509
rect 33321 9469 33333 9503
rect 33367 9469 33379 9503
rect 33796 9500 33824 9540
rect 33870 9528 33876 9580
rect 33928 9568 33934 9580
rect 34072 9577 34100 9608
rect 35066 9596 35072 9608
rect 35124 9596 35130 9648
rect 35434 9636 35440 9648
rect 35268 9608 35440 9636
rect 34057 9571 34115 9577
rect 33928 9540 34021 9568
rect 33928 9528 33934 9540
rect 34057 9537 34069 9571
rect 34103 9537 34115 9571
rect 34057 9531 34115 9537
rect 34149 9571 34207 9577
rect 34149 9537 34161 9571
rect 34195 9537 34207 9571
rect 34149 9531 34207 9537
rect 34164 9500 34192 9531
rect 34238 9528 34244 9580
rect 34296 9568 34302 9580
rect 34296 9540 34341 9568
rect 34296 9528 34302 9540
rect 34422 9528 34428 9580
rect 34480 9568 34486 9580
rect 34977 9571 35035 9577
rect 34977 9568 34989 9571
rect 34480 9540 34989 9568
rect 34480 9528 34486 9540
rect 34977 9537 34989 9540
rect 35023 9537 35035 9571
rect 35158 9568 35164 9580
rect 35119 9540 35164 9568
rect 34977 9531 35035 9537
rect 35158 9528 35164 9540
rect 35216 9528 35222 9580
rect 35268 9577 35296 9608
rect 35434 9596 35440 9608
rect 35492 9596 35498 9648
rect 36725 9639 36783 9645
rect 36725 9605 36737 9639
rect 36771 9636 36783 9639
rect 38289 9639 38347 9645
rect 36771 9608 37872 9636
rect 36771 9605 36783 9608
rect 36725 9599 36783 9605
rect 35253 9571 35311 9577
rect 35253 9537 35265 9571
rect 35299 9537 35311 9571
rect 35253 9531 35311 9537
rect 35345 9571 35403 9577
rect 35345 9537 35357 9571
rect 35391 9568 35403 9571
rect 35802 9568 35808 9580
rect 35391 9540 35808 9568
rect 35391 9537 35403 9540
rect 35345 9531 35403 9537
rect 35268 9500 35296 9531
rect 35802 9528 35808 9540
rect 35860 9528 35866 9580
rect 36354 9568 36360 9580
rect 36315 9540 36360 9568
rect 36354 9528 36360 9540
rect 36412 9528 36418 9580
rect 36541 9571 36599 9577
rect 36541 9537 36553 9571
rect 36587 9537 36599 9571
rect 36541 9531 36599 9537
rect 33796 9472 35296 9500
rect 33321 9463 33379 9469
rect 29144 9404 30236 9432
rect 29144 9392 29150 9404
rect 30282 9392 30288 9444
rect 30340 9432 30346 9444
rect 33226 9432 33232 9444
rect 30340 9404 33232 9432
rect 30340 9392 30346 9404
rect 33226 9392 33232 9404
rect 33284 9432 33290 9444
rect 33336 9432 33364 9463
rect 35710 9460 35716 9512
rect 35768 9500 35774 9512
rect 36556 9500 36584 9531
rect 37182 9528 37188 9580
rect 37240 9568 37246 9580
rect 37550 9568 37556 9580
rect 37240 9540 37556 9568
rect 37240 9528 37246 9540
rect 37550 9528 37556 9540
rect 37608 9568 37614 9580
rect 37844 9577 37872 9608
rect 38289 9605 38301 9639
rect 38335 9636 38347 9639
rect 39178 9639 39236 9645
rect 39178 9636 39190 9639
rect 38335 9608 39190 9636
rect 38335 9605 38347 9608
rect 38289 9599 38347 9605
rect 39178 9605 39190 9608
rect 39224 9605 39236 9639
rect 39178 9599 39236 9605
rect 37645 9571 37703 9577
rect 37645 9568 37657 9571
rect 37608 9540 37657 9568
rect 37608 9528 37614 9540
rect 37645 9537 37657 9540
rect 37691 9537 37703 9571
rect 37645 9531 37703 9537
rect 37829 9571 37887 9577
rect 37829 9537 37841 9571
rect 37875 9537 37887 9571
rect 37829 9531 37887 9537
rect 37921 9528 37927 9580
rect 37979 9571 37985 9580
rect 38059 9571 38117 9577
rect 37979 9543 38021 9571
rect 37979 9528 37985 9543
rect 38059 9537 38071 9571
rect 38105 9568 38117 9571
rect 38194 9568 38200 9580
rect 38105 9540 38200 9568
rect 38105 9537 38117 9540
rect 38059 9531 38117 9537
rect 38194 9528 38200 9540
rect 38252 9528 38258 9580
rect 35768 9472 36584 9500
rect 35768 9460 35774 9472
rect 33284 9404 33364 9432
rect 36556 9432 36584 9472
rect 38562 9460 38568 9512
rect 38620 9500 38626 9512
rect 38933 9503 38991 9509
rect 38933 9500 38945 9503
rect 38620 9472 38945 9500
rect 38620 9460 38626 9472
rect 38933 9469 38945 9472
rect 38979 9469 38991 9503
rect 38933 9463 38991 9469
rect 36556 9404 37412 9432
rect 33284 9392 33290 9404
rect 21082 9364 21088 9376
rect 18340 9336 21088 9364
rect 21082 9324 21088 9336
rect 21140 9324 21146 9376
rect 23753 9367 23811 9373
rect 23753 9333 23765 9367
rect 23799 9364 23811 9367
rect 24578 9364 24584 9376
rect 23799 9336 24584 9364
rect 23799 9333 23811 9336
rect 23753 9327 23811 9333
rect 24578 9324 24584 9336
rect 24636 9324 24642 9376
rect 29730 9364 29736 9376
rect 29691 9336 29736 9364
rect 29730 9324 29736 9336
rect 29788 9324 29794 9376
rect 34517 9367 34575 9373
rect 34517 9333 34529 9367
rect 34563 9364 34575 9367
rect 35526 9364 35532 9376
rect 34563 9336 35532 9364
rect 34563 9333 34575 9336
rect 34517 9327 34575 9333
rect 35526 9324 35532 9336
rect 35584 9324 35590 9376
rect 35621 9367 35679 9373
rect 35621 9333 35633 9367
rect 35667 9364 35679 9367
rect 37090 9364 37096 9376
rect 35667 9336 37096 9364
rect 35667 9333 35679 9336
rect 35621 9327 35679 9333
rect 37090 9324 37096 9336
rect 37148 9324 37154 9376
rect 37384 9364 37412 9404
rect 40313 9367 40371 9373
rect 40313 9364 40325 9367
rect 37384 9336 40325 9364
rect 40313 9333 40325 9336
rect 40359 9364 40371 9367
rect 40862 9364 40868 9376
rect 40359 9336 40868 9364
rect 40359 9333 40371 9336
rect 40313 9327 40371 9333
rect 40862 9324 40868 9336
rect 40920 9324 40926 9376
rect 1104 9274 68816 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 65654 9274
rect 65706 9222 65718 9274
rect 65770 9222 65782 9274
rect 65834 9222 65846 9274
rect 65898 9222 65910 9274
rect 65962 9222 68816 9274
rect 1104 9200 68816 9222
rect 1946 9160 1952 9172
rect 1907 9132 1952 9160
rect 1946 9120 1952 9132
rect 2004 9120 2010 9172
rect 5166 9160 5172 9172
rect 5127 9132 5172 9160
rect 5166 9120 5172 9132
rect 5224 9120 5230 9172
rect 10318 9160 10324 9172
rect 10279 9132 10324 9160
rect 10318 9120 10324 9132
rect 10376 9120 10382 9172
rect 13262 9160 13268 9172
rect 13223 9132 13268 9160
rect 13262 9120 13268 9132
rect 13320 9120 13326 9172
rect 14182 9120 14188 9172
rect 14240 9160 14246 9172
rect 14240 9132 15976 9160
rect 14240 9120 14246 9132
rect 11790 9092 11796 9104
rect 10060 9064 11796 9092
rect 6733 9027 6791 9033
rect 6733 8993 6745 9027
rect 6779 9024 6791 9027
rect 9769 9027 9827 9033
rect 9769 9024 9781 9027
rect 6779 8996 9781 9024
rect 6779 8993 6791 8996
rect 6733 8987 6791 8993
rect 9769 8993 9781 8996
rect 9815 9024 9827 9027
rect 9858 9024 9864 9036
rect 9815 8996 9864 9024
rect 9815 8993 9827 8996
rect 9769 8987 9827 8993
rect 9858 8984 9864 8996
rect 9916 8984 9922 9036
rect 2317 8959 2375 8965
rect 2317 8925 2329 8959
rect 2363 8956 2375 8959
rect 2774 8956 2780 8968
rect 2363 8928 2780 8956
rect 2363 8925 2375 8928
rect 2317 8919 2375 8925
rect 2774 8916 2780 8928
rect 2832 8916 2838 8968
rect 3510 8916 3516 8968
rect 3568 8956 3574 8968
rect 3789 8959 3847 8965
rect 3789 8956 3801 8959
rect 3568 8928 3801 8956
rect 3568 8916 3574 8928
rect 3789 8925 3801 8928
rect 3835 8925 3847 8959
rect 3789 8919 3847 8925
rect 5258 8916 5264 8968
rect 5316 8956 5322 8968
rect 6457 8959 6515 8965
rect 6457 8956 6469 8959
rect 5316 8928 6469 8956
rect 5316 8916 5322 8928
rect 6457 8925 6469 8928
rect 6503 8925 6515 8959
rect 6457 8919 6515 8925
rect 6914 8916 6920 8968
rect 6972 8956 6978 8968
rect 7742 8956 7748 8968
rect 6972 8928 7748 8956
rect 6972 8916 6978 8928
rect 7742 8916 7748 8928
rect 7800 8916 7806 8968
rect 7926 8956 7932 8968
rect 7887 8928 7932 8956
rect 7926 8916 7932 8928
rect 7984 8916 7990 8968
rect 8021 8959 8079 8965
rect 8021 8925 8033 8959
rect 8067 8925 8079 8959
rect 8021 8919 8079 8925
rect 2133 8891 2191 8897
rect 2133 8857 2145 8891
rect 2179 8888 2191 8891
rect 2222 8888 2228 8900
rect 2179 8860 2228 8888
rect 2179 8857 2191 8860
rect 2133 8851 2191 8857
rect 2222 8848 2228 8860
rect 2280 8848 2286 8900
rect 2406 8848 2412 8900
rect 2464 8888 2470 8900
rect 4056 8891 4114 8897
rect 2464 8860 4016 8888
rect 2464 8848 2470 8860
rect 2774 8780 2780 8832
rect 2832 8820 2838 8832
rect 2869 8823 2927 8829
rect 2869 8820 2881 8823
rect 2832 8792 2881 8820
rect 2832 8780 2838 8792
rect 2869 8789 2881 8792
rect 2915 8820 2927 8823
rect 3050 8820 3056 8832
rect 2915 8792 3056 8820
rect 2915 8789 2927 8792
rect 2869 8783 2927 8789
rect 3050 8780 3056 8792
rect 3108 8780 3114 8832
rect 3988 8820 4016 8860
rect 4056 8857 4068 8891
rect 4102 8888 4114 8891
rect 5074 8888 5080 8900
rect 4102 8860 5080 8888
rect 4102 8857 4114 8860
rect 4056 8851 4114 8857
rect 5074 8848 5080 8860
rect 5132 8848 5138 8900
rect 8036 8888 8064 8919
rect 8110 8916 8116 8968
rect 8168 8956 8174 8968
rect 9493 8959 9551 8965
rect 8168 8928 8213 8956
rect 8168 8916 8174 8928
rect 9493 8925 9505 8959
rect 9539 8956 9551 8959
rect 10060 8956 10088 9064
rect 11790 9052 11796 9064
rect 11848 9052 11854 9104
rect 15948 9092 15976 9132
rect 17126 9120 17132 9172
rect 17184 9160 17190 9172
rect 17221 9163 17279 9169
rect 17221 9160 17233 9163
rect 17184 9132 17233 9160
rect 17184 9120 17190 9132
rect 17221 9129 17233 9132
rect 17267 9129 17279 9163
rect 17221 9123 17279 9129
rect 17494 9120 17500 9172
rect 17552 9160 17558 9172
rect 18049 9163 18107 9169
rect 17552 9132 18000 9160
rect 17552 9120 17558 9132
rect 17865 9095 17923 9101
rect 17865 9092 17877 9095
rect 15948 9064 17877 9092
rect 17865 9061 17877 9064
rect 17911 9061 17923 9095
rect 17972 9092 18000 9132
rect 18049 9129 18061 9163
rect 18095 9160 18107 9163
rect 18506 9160 18512 9172
rect 18095 9132 18512 9160
rect 18095 9129 18107 9132
rect 18049 9123 18107 9129
rect 18506 9120 18512 9132
rect 18564 9120 18570 9172
rect 20070 9160 20076 9172
rect 20031 9132 20076 9160
rect 20070 9120 20076 9132
rect 20128 9120 20134 9172
rect 23293 9163 23351 9169
rect 23293 9160 23305 9163
rect 22066 9132 23305 9160
rect 22066 9092 22094 9132
rect 23293 9129 23305 9132
rect 23339 9160 23351 9163
rect 23382 9160 23388 9172
rect 23339 9132 23388 9160
rect 23339 9129 23351 9132
rect 23293 9123 23351 9129
rect 23382 9120 23388 9132
rect 23440 9120 23446 9172
rect 27065 9163 27123 9169
rect 25700 9132 26740 9160
rect 17972 9064 22094 9092
rect 22649 9095 22707 9101
rect 17865 9055 17923 9061
rect 22649 9061 22661 9095
rect 22695 9092 22707 9095
rect 25700 9092 25728 9132
rect 22695 9064 25728 9092
rect 22695 9061 22707 9064
rect 22649 9055 22707 9061
rect 11606 8984 11612 9036
rect 11664 9024 11670 9036
rect 11885 9027 11943 9033
rect 11885 9024 11897 9027
rect 11664 8996 11897 9024
rect 11664 8984 11670 8996
rect 11885 8993 11897 8996
rect 11931 8993 11943 9027
rect 11885 8987 11943 8993
rect 15933 9027 15991 9033
rect 15933 8993 15945 9027
rect 15979 9024 15991 9027
rect 16206 9024 16212 9036
rect 15979 8996 16212 9024
rect 15979 8993 15991 8996
rect 15933 8987 15991 8993
rect 16206 8984 16212 8996
rect 16264 8984 16270 9036
rect 20441 9027 20499 9033
rect 19444 8996 20300 9024
rect 9539 8928 10088 8956
rect 9539 8925 9551 8928
rect 9493 8919 9551 8925
rect 9508 8888 9536 8919
rect 10134 8916 10140 8968
rect 10192 8956 10198 8968
rect 10229 8959 10287 8965
rect 10229 8956 10241 8959
rect 10192 8928 10241 8956
rect 10192 8916 10198 8928
rect 10229 8925 10241 8928
rect 10275 8925 10287 8959
rect 10229 8919 10287 8925
rect 10413 8959 10471 8965
rect 10413 8925 10425 8959
rect 10459 8956 10471 8959
rect 10686 8956 10692 8968
rect 10459 8928 10692 8956
rect 10459 8925 10471 8928
rect 10413 8919 10471 8925
rect 8036 8860 9536 8888
rect 10244 8888 10272 8919
rect 10686 8916 10692 8928
rect 10744 8916 10750 8968
rect 12158 8965 12164 8968
rect 12152 8956 12164 8965
rect 12119 8928 12164 8956
rect 12152 8919 12164 8928
rect 12158 8916 12164 8919
rect 12216 8916 12222 8968
rect 15654 8916 15660 8968
rect 15712 8965 15718 8968
rect 15712 8956 15724 8965
rect 19334 8956 19340 8968
rect 15712 8928 15757 8956
rect 18340 8928 19340 8956
rect 15712 8919 15724 8928
rect 15712 8916 15718 8919
rect 18040 8891 18098 8897
rect 10244 8860 18000 8888
rect 7006 8820 7012 8832
rect 3988 8792 7012 8820
rect 7006 8780 7012 8792
rect 7064 8780 7070 8832
rect 7282 8820 7288 8832
rect 7243 8792 7288 8820
rect 7282 8780 7288 8792
rect 7340 8780 7346 8832
rect 8386 8820 8392 8832
rect 8347 8792 8392 8820
rect 8386 8780 8392 8792
rect 8444 8780 8450 8832
rect 10778 8780 10784 8832
rect 10836 8820 10842 8832
rect 11146 8820 11152 8832
rect 10836 8792 11152 8820
rect 10836 8780 10842 8792
rect 11146 8780 11152 8792
rect 11204 8780 11210 8832
rect 13354 8780 13360 8832
rect 13412 8820 13418 8832
rect 14553 8823 14611 8829
rect 14553 8820 14565 8823
rect 13412 8792 14565 8820
rect 13412 8780 13418 8792
rect 14553 8789 14565 8792
rect 14599 8820 14611 8823
rect 15470 8820 15476 8832
rect 14599 8792 15476 8820
rect 14599 8789 14611 8792
rect 14553 8783 14611 8789
rect 15470 8780 15476 8792
rect 15528 8780 15534 8832
rect 17972 8820 18000 8860
rect 18040 8857 18052 8891
rect 18086 8888 18098 8891
rect 18340 8888 18368 8928
rect 19334 8916 19340 8928
rect 19392 8916 19398 8968
rect 19444 8965 19472 8996
rect 19429 8959 19487 8965
rect 19429 8925 19441 8959
rect 19475 8925 19487 8959
rect 19429 8919 19487 8925
rect 19613 8959 19671 8965
rect 19613 8925 19625 8959
rect 19659 8956 19671 8959
rect 20162 8956 20168 8968
rect 19659 8928 20168 8956
rect 19659 8925 19671 8928
rect 19613 8919 19671 8925
rect 20162 8916 20168 8928
rect 20220 8916 20226 8968
rect 20272 8965 20300 8996
rect 20441 8993 20453 9027
rect 20487 9024 20499 9027
rect 20806 9024 20812 9036
rect 20487 8996 20812 9024
rect 20487 8993 20499 8996
rect 20441 8987 20499 8993
rect 20806 8984 20812 8996
rect 20864 8984 20870 9036
rect 20257 8959 20315 8965
rect 20257 8925 20269 8959
rect 20303 8956 20315 8959
rect 20346 8956 20352 8968
rect 20303 8928 20352 8956
rect 20303 8925 20315 8928
rect 20257 8919 20315 8925
rect 20346 8916 20352 8928
rect 20404 8916 20410 8968
rect 20533 8959 20591 8965
rect 20533 8925 20545 8959
rect 20579 8956 20591 8959
rect 20622 8956 20628 8968
rect 20579 8928 20628 8956
rect 20579 8925 20591 8928
rect 20533 8919 20591 8925
rect 20622 8916 20628 8928
rect 20680 8916 20686 8968
rect 22557 8959 22615 8965
rect 22557 8956 22569 8959
rect 21192 8928 22569 8956
rect 21192 8900 21220 8928
rect 22557 8925 22569 8928
rect 22603 8956 22615 8959
rect 23106 8956 23112 8968
rect 22603 8928 23112 8956
rect 22603 8925 22615 8928
rect 22557 8919 22615 8925
rect 23106 8916 23112 8928
rect 23164 8916 23170 8968
rect 18086 8860 18368 8888
rect 18417 8891 18475 8897
rect 18086 8857 18098 8860
rect 18040 8851 18098 8857
rect 18417 8857 18429 8891
rect 18463 8888 18475 8891
rect 18782 8888 18788 8900
rect 18463 8860 18788 8888
rect 18463 8857 18475 8860
rect 18417 8851 18475 8857
rect 18432 8820 18460 8851
rect 18782 8848 18788 8860
rect 18840 8888 18846 8900
rect 19245 8891 19303 8897
rect 19245 8888 19257 8891
rect 18840 8860 19257 8888
rect 18840 8848 18846 8860
rect 19245 8857 19257 8860
rect 19291 8857 19303 8891
rect 21174 8888 21180 8900
rect 21135 8860 21180 8888
rect 19245 8851 19303 8857
rect 21174 8848 21180 8860
rect 21232 8848 21238 8900
rect 21634 8848 21640 8900
rect 21692 8888 21698 8900
rect 21913 8891 21971 8897
rect 21913 8888 21925 8891
rect 21692 8860 21925 8888
rect 21692 8848 21698 8860
rect 21913 8857 21925 8860
rect 21959 8888 21971 8891
rect 23216 8888 23244 9064
rect 24210 8984 24216 9036
rect 24268 9024 24274 9036
rect 26712 9024 26740 9132
rect 27065 9129 27077 9163
rect 27111 9160 27123 9163
rect 27706 9160 27712 9172
rect 27111 9132 27712 9160
rect 27111 9129 27123 9132
rect 27065 9123 27123 9129
rect 27706 9120 27712 9132
rect 27764 9160 27770 9172
rect 28994 9160 29000 9172
rect 27764 9132 29000 9160
rect 27764 9120 27770 9132
rect 28994 9120 29000 9132
rect 29052 9120 29058 9172
rect 29270 9120 29276 9172
rect 29328 9160 29334 9172
rect 29549 9163 29607 9169
rect 29549 9160 29561 9163
rect 29328 9132 29561 9160
rect 29328 9120 29334 9132
rect 29549 9129 29561 9132
rect 29595 9129 29607 9163
rect 29549 9123 29607 9129
rect 36354 9120 36360 9172
rect 36412 9160 36418 9172
rect 36412 9132 38332 9160
rect 36412 9120 36418 9132
rect 29822 9052 29828 9104
rect 29880 9092 29886 9104
rect 35710 9092 35716 9104
rect 29880 9064 35716 9092
rect 29880 9052 29886 9064
rect 35710 9052 35716 9064
rect 35768 9052 35774 9104
rect 35802 9052 35808 9104
rect 35860 9092 35866 9104
rect 36633 9095 36691 9101
rect 36633 9092 36645 9095
rect 35860 9064 36645 9092
rect 35860 9052 35866 9064
rect 36633 9061 36645 9064
rect 36679 9092 36691 9095
rect 36679 9064 37596 9092
rect 36679 9061 36691 9064
rect 36633 9055 36691 9061
rect 30742 9024 30748 9036
rect 24268 8996 25807 9024
rect 26712 8996 27660 9024
rect 24268 8984 24274 8996
rect 25685 8959 25743 8965
rect 25685 8956 25697 8959
rect 21959 8860 23244 8888
rect 23584 8928 25697 8956
rect 21959 8857 21971 8860
rect 21913 8851 21971 8857
rect 17972 8792 18460 8820
rect 19150 8780 19156 8832
rect 19208 8820 19214 8832
rect 20070 8820 20076 8832
rect 19208 8792 20076 8820
rect 19208 8780 19214 8792
rect 20070 8780 20076 8792
rect 20128 8820 20134 8832
rect 21821 8823 21879 8829
rect 21821 8820 21833 8823
rect 20128 8792 21833 8820
rect 20128 8780 20134 8792
rect 21821 8789 21833 8792
rect 21867 8789 21879 8823
rect 21821 8783 21879 8789
rect 22094 8780 22100 8832
rect 22152 8820 22158 8832
rect 23584 8820 23612 8928
rect 25685 8925 25697 8928
rect 25731 8925 25743 8959
rect 25779 8956 25807 8996
rect 27246 8956 27252 8968
rect 25779 8928 27252 8956
rect 25685 8919 25743 8925
rect 27246 8916 27252 8928
rect 27304 8956 27310 8968
rect 27525 8959 27583 8965
rect 27525 8956 27537 8959
rect 27304 8928 27537 8956
rect 27304 8916 27310 8928
rect 27525 8925 27537 8928
rect 27571 8925 27583 8959
rect 27632 8956 27660 8996
rect 28552 8996 30236 9024
rect 30703 8996 30748 9024
rect 28552 8956 28580 8996
rect 30208 8968 30236 8996
rect 30742 8984 30748 8996
rect 30800 8984 30806 9036
rect 30834 8984 30840 9036
rect 30892 9024 30898 9036
rect 31846 9024 31852 9036
rect 30892 8996 31852 9024
rect 30892 8984 30898 8996
rect 31846 8984 31852 8996
rect 31904 8984 31910 9036
rect 33502 9024 33508 9036
rect 32048 8996 33508 9024
rect 27632 8928 28580 8956
rect 27525 8919 27583 8925
rect 29362 8916 29368 8968
rect 29420 8956 29426 8968
rect 29733 8959 29791 8965
rect 29733 8956 29745 8959
rect 29420 8928 29745 8956
rect 29420 8916 29426 8928
rect 29733 8925 29745 8928
rect 29779 8925 29791 8959
rect 29914 8956 29920 8968
rect 29875 8928 29920 8956
rect 29733 8919 29791 8925
rect 24581 8891 24639 8897
rect 24581 8857 24593 8891
rect 24627 8857 24639 8891
rect 24581 8851 24639 8857
rect 23842 8820 23848 8832
rect 22152 8792 23612 8820
rect 23803 8792 23848 8820
rect 22152 8780 22158 8792
rect 23842 8780 23848 8792
rect 23900 8780 23906 8832
rect 24302 8780 24308 8832
rect 24360 8820 24366 8832
rect 24397 8823 24455 8829
rect 24397 8820 24409 8823
rect 24360 8792 24409 8820
rect 24360 8780 24366 8792
rect 24397 8789 24409 8792
rect 24443 8789 24455 8823
rect 24397 8783 24455 8789
rect 24486 8780 24492 8832
rect 24544 8820 24550 8832
rect 24596 8820 24624 8851
rect 24670 8848 24676 8900
rect 24728 8888 24734 8900
rect 24765 8891 24823 8897
rect 24765 8888 24777 8891
rect 24728 8860 24777 8888
rect 24728 8848 24734 8860
rect 24765 8857 24777 8860
rect 24811 8857 24823 8891
rect 24765 8851 24823 8857
rect 25774 8848 25780 8900
rect 25832 8888 25838 8900
rect 27798 8897 27804 8900
rect 25930 8891 25988 8897
rect 25930 8888 25942 8891
rect 25832 8860 25942 8888
rect 25832 8848 25838 8860
rect 25930 8857 25942 8860
rect 25976 8857 25988 8891
rect 25930 8851 25988 8857
rect 27792 8851 27804 8897
rect 27856 8888 27862 8900
rect 29748 8888 29776 8919
rect 29914 8916 29920 8928
rect 29972 8916 29978 8968
rect 30190 8916 30196 8968
rect 30248 8956 30254 8968
rect 30469 8959 30527 8965
rect 30469 8956 30481 8959
rect 30248 8928 30481 8956
rect 30248 8916 30254 8928
rect 30469 8925 30481 8928
rect 30515 8925 30527 8959
rect 30469 8919 30527 8925
rect 31110 8916 31116 8968
rect 31168 8956 31174 8968
rect 31757 8959 31815 8965
rect 31757 8956 31769 8959
rect 31168 8928 31769 8956
rect 31168 8916 31174 8928
rect 31757 8925 31769 8928
rect 31803 8925 31815 8959
rect 31938 8956 31944 8968
rect 31899 8928 31944 8956
rect 31757 8919 31815 8925
rect 31938 8916 31944 8928
rect 31996 8916 32002 8968
rect 32048 8965 32076 8996
rect 32033 8959 32091 8965
rect 32033 8925 32045 8959
rect 32079 8925 32091 8959
rect 32033 8919 32091 8925
rect 32125 8959 32183 8965
rect 32125 8925 32137 8959
rect 32171 8925 32183 8959
rect 33226 8956 33232 8968
rect 33187 8928 33232 8956
rect 32125 8919 32183 8925
rect 31018 8888 31024 8900
rect 27856 8860 27892 8888
rect 29748 8860 31024 8888
rect 27798 8848 27804 8851
rect 27856 8848 27862 8860
rect 31018 8848 31024 8860
rect 31076 8848 31082 8900
rect 31478 8848 31484 8900
rect 31536 8888 31542 8900
rect 32140 8888 32168 8919
rect 33226 8916 33232 8928
rect 33284 8916 33290 8968
rect 33336 8965 33364 8996
rect 33502 8984 33508 8996
rect 33560 8984 33566 9036
rect 33321 8959 33379 8965
rect 33321 8925 33333 8959
rect 33367 8925 33379 8959
rect 33321 8919 33379 8925
rect 33410 8916 33416 8968
rect 33468 8956 33474 8968
rect 33597 8959 33655 8965
rect 33468 8928 33513 8956
rect 33468 8916 33474 8928
rect 33597 8925 33609 8959
rect 33643 8956 33655 8959
rect 33870 8956 33876 8968
rect 33643 8928 33876 8956
rect 33643 8925 33655 8928
rect 33597 8919 33655 8925
rect 33870 8916 33876 8928
rect 33928 8916 33934 8968
rect 33980 8928 37136 8956
rect 33980 8888 34008 8928
rect 34514 8888 34520 8900
rect 31536 8860 32168 8888
rect 32232 8860 34008 8888
rect 34072 8860 34520 8888
rect 31536 8848 31542 8860
rect 28442 8820 28448 8832
rect 24544 8792 28448 8820
rect 24544 8780 24550 8792
rect 28442 8780 28448 8792
rect 28500 8780 28506 8832
rect 28810 8780 28816 8832
rect 28868 8820 28874 8832
rect 28905 8823 28963 8829
rect 28905 8820 28917 8823
rect 28868 8792 28917 8820
rect 28868 8780 28874 8792
rect 28905 8789 28917 8792
rect 28951 8789 28963 8823
rect 28905 8783 28963 8789
rect 31846 8780 31852 8832
rect 31904 8820 31910 8832
rect 32232 8820 32260 8860
rect 34072 8832 34100 8860
rect 34514 8848 34520 8860
rect 34572 8888 34578 8900
rect 35161 8891 35219 8897
rect 35161 8888 35173 8891
rect 34572 8860 35173 8888
rect 34572 8848 34578 8860
rect 35161 8857 35173 8860
rect 35207 8857 35219 8891
rect 35161 8851 35219 8857
rect 35710 8848 35716 8900
rect 35768 8888 35774 8900
rect 35897 8891 35955 8897
rect 35897 8888 35909 8891
rect 35768 8860 35909 8888
rect 35768 8848 35774 8860
rect 35897 8857 35909 8860
rect 35943 8857 35955 8891
rect 37108 8888 37136 8928
rect 37182 8916 37188 8968
rect 37240 8956 37246 8968
rect 37366 8956 37372 8968
rect 37240 8928 37285 8956
rect 37327 8928 37372 8956
rect 37240 8916 37246 8928
rect 37366 8916 37372 8928
rect 37424 8916 37430 8968
rect 37568 8965 37596 9064
rect 37829 9027 37887 9033
rect 37829 8993 37841 9027
rect 37875 9024 37887 9027
rect 38194 9024 38200 9036
rect 37875 8996 38200 9024
rect 37875 8993 37887 8996
rect 37829 8987 37887 8993
rect 38194 8984 38200 8996
rect 38252 8984 38258 9036
rect 38304 8965 38332 9132
rect 37461 8959 37519 8965
rect 37461 8925 37473 8959
rect 37507 8925 37519 8959
rect 37461 8919 37519 8925
rect 37553 8959 37611 8965
rect 37553 8925 37565 8959
rect 37599 8925 37611 8959
rect 37553 8919 37611 8925
rect 38289 8959 38347 8965
rect 38289 8925 38301 8959
rect 38335 8925 38347 8959
rect 38289 8919 38347 8925
rect 37476 8888 37504 8919
rect 37918 8888 37924 8900
rect 37108 8860 37412 8888
rect 37476 8860 37924 8888
rect 35897 8851 35955 8857
rect 32398 8820 32404 8832
rect 31904 8792 32260 8820
rect 32359 8792 32404 8820
rect 31904 8780 31910 8792
rect 32398 8780 32404 8792
rect 32456 8780 32462 8832
rect 32953 8823 33011 8829
rect 32953 8789 32965 8823
rect 32999 8820 33011 8823
rect 33042 8820 33048 8832
rect 32999 8792 33048 8820
rect 32999 8789 33011 8792
rect 32953 8783 33011 8789
rect 33042 8780 33048 8792
rect 33100 8780 33106 8832
rect 34054 8820 34060 8832
rect 34015 8792 34060 8820
rect 34054 8780 34060 8792
rect 34112 8780 34118 8832
rect 37384 8820 37412 8860
rect 37918 8848 37924 8860
rect 37976 8848 37982 8900
rect 38473 8891 38531 8897
rect 38473 8857 38485 8891
rect 38519 8888 38531 8891
rect 39117 8891 39175 8897
rect 39117 8888 39129 8891
rect 38519 8860 39129 8888
rect 38519 8857 38531 8860
rect 38473 8851 38531 8857
rect 39117 8857 39129 8860
rect 39163 8888 39175 8891
rect 39298 8888 39304 8900
rect 39163 8860 39304 8888
rect 39163 8857 39175 8860
rect 39117 8851 39175 8857
rect 38488 8820 38516 8851
rect 39298 8848 39304 8860
rect 39356 8848 39362 8900
rect 38654 8820 38660 8832
rect 37384 8792 38516 8820
rect 38615 8792 38660 8820
rect 38654 8780 38660 8792
rect 38712 8780 38718 8832
rect 1104 8730 68816 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 50294 8730
rect 50346 8678 50358 8730
rect 50410 8678 50422 8730
rect 50474 8678 50486 8730
rect 50538 8678 50550 8730
rect 50602 8678 68816 8730
rect 1104 8656 68816 8678
rect 2038 8576 2044 8628
rect 2096 8616 2102 8628
rect 2096 8588 5028 8616
rect 2096 8576 2102 8588
rect 2053 8548 2081 8576
rect 3510 8548 3516 8560
rect 2053 8520 2084 8548
rect 1854 8440 1860 8492
rect 1912 8483 1918 8492
rect 2056 8489 2084 8520
rect 2792 8520 3516 8548
rect 1949 8483 2007 8489
rect 1912 8455 1961 8483
rect 1912 8440 1918 8455
rect 1949 8449 1961 8455
rect 1995 8449 2007 8483
rect 1949 8443 2007 8449
rect 2041 8483 2099 8489
rect 2041 8449 2053 8483
rect 2087 8449 2099 8483
rect 2041 8443 2099 8449
rect 2154 8483 2212 8489
rect 2154 8449 2166 8483
rect 2200 8480 2212 8483
rect 2317 8483 2375 8489
rect 2200 8449 2222 8480
rect 2154 8443 2222 8449
rect 2317 8449 2329 8483
rect 2363 8480 2375 8483
rect 2406 8480 2412 8492
rect 2363 8452 2412 8480
rect 2363 8449 2375 8452
rect 2317 8443 2375 8449
rect 2194 8356 2222 8443
rect 2406 8440 2412 8452
rect 2464 8440 2470 8492
rect 2792 8489 2820 8520
rect 3510 8508 3516 8520
rect 3568 8508 3574 8560
rect 5000 8548 5028 8588
rect 5074 8576 5080 8628
rect 5132 8616 5138 8628
rect 5169 8619 5227 8625
rect 5169 8616 5181 8619
rect 5132 8588 5181 8616
rect 5132 8576 5138 8588
rect 5169 8585 5181 8588
rect 5215 8585 5227 8619
rect 5169 8579 5227 8585
rect 5626 8576 5632 8628
rect 5684 8576 5690 8628
rect 7926 8576 7932 8628
rect 7984 8616 7990 8628
rect 8113 8619 8171 8625
rect 8113 8616 8125 8619
rect 7984 8588 8125 8616
rect 7984 8576 7990 8588
rect 8113 8585 8125 8588
rect 8159 8585 8171 8619
rect 14366 8616 14372 8628
rect 8113 8579 8171 8585
rect 8220 8588 14372 8616
rect 5258 8548 5264 8560
rect 5000 8520 5264 8548
rect 5258 8508 5264 8520
rect 5316 8548 5322 8560
rect 5316 8520 5580 8548
rect 5316 8508 5322 8520
rect 2777 8483 2835 8489
rect 2777 8449 2789 8483
rect 2823 8449 2835 8483
rect 3033 8483 3091 8489
rect 3033 8480 3045 8483
rect 2777 8443 2835 8449
rect 2884 8452 3045 8480
rect 2884 8412 2912 8452
rect 3033 8449 3045 8452
rect 3079 8449 3091 8483
rect 3033 8443 3091 8449
rect 5166 8440 5172 8492
rect 5224 8480 5230 8492
rect 5552 8489 5580 8520
rect 5649 8489 5677 8576
rect 7006 8508 7012 8560
rect 7064 8548 7070 8560
rect 8220 8548 8248 8588
rect 14366 8576 14372 8588
rect 14424 8576 14430 8628
rect 17034 8616 17040 8628
rect 14568 8588 17040 8616
rect 7064 8520 8248 8548
rect 7064 8508 7070 8520
rect 8386 8508 8392 8560
rect 8444 8548 8450 8560
rect 9002 8551 9060 8557
rect 9002 8548 9014 8551
rect 8444 8520 9014 8548
rect 8444 8508 8450 8520
rect 9002 8517 9014 8520
rect 9048 8517 9060 8551
rect 14568 8548 14596 8588
rect 17034 8576 17040 8588
rect 17092 8576 17098 8628
rect 19242 8616 19248 8628
rect 19076 8588 19248 8616
rect 9002 8511 9060 8517
rect 9140 8520 14596 8548
rect 14645 8551 14703 8557
rect 5399 8483 5457 8489
rect 5399 8480 5411 8483
rect 5224 8452 5411 8480
rect 5224 8440 5230 8452
rect 5399 8449 5411 8452
rect 5445 8449 5457 8483
rect 5399 8443 5457 8449
rect 5537 8483 5595 8489
rect 5537 8449 5549 8483
rect 5583 8449 5595 8483
rect 5537 8443 5595 8449
rect 5629 8483 5687 8489
rect 5629 8449 5641 8483
rect 5675 8449 5687 8483
rect 5629 8443 5687 8449
rect 5813 8483 5871 8489
rect 5813 8449 5825 8483
rect 5859 8480 5871 8483
rect 6914 8480 6920 8492
rect 5859 8452 6920 8480
rect 5859 8449 5871 8452
rect 5813 8443 5871 8449
rect 6914 8440 6920 8452
rect 6972 8440 6978 8492
rect 7098 8440 7104 8492
rect 7156 8480 7162 8492
rect 7745 8483 7803 8489
rect 7745 8480 7757 8483
rect 7156 8452 7757 8480
rect 7156 8440 7162 8452
rect 7745 8449 7757 8452
rect 7791 8449 7803 8483
rect 7926 8480 7932 8492
rect 7887 8452 7932 8480
rect 7745 8443 7803 8449
rect 7926 8440 7932 8452
rect 7984 8440 7990 8492
rect 9140 8480 9168 8520
rect 14645 8517 14657 8551
rect 14691 8548 14703 8551
rect 15010 8548 15016 8560
rect 14691 8520 15016 8548
rect 14691 8517 14703 8520
rect 14645 8511 14703 8517
rect 15010 8508 15016 8520
rect 15068 8508 15074 8560
rect 16500 8520 18552 8548
rect 14458 8480 14464 8492
rect 8036 8452 9168 8480
rect 14419 8452 14464 8480
rect 2130 8304 2136 8356
rect 2188 8316 2222 8356
rect 2792 8384 2912 8412
rect 2188 8304 2194 8316
rect 1673 8279 1731 8285
rect 1673 8245 1685 8279
rect 1719 8276 1731 8279
rect 2792 8276 2820 8384
rect 5902 8372 5908 8424
rect 5960 8412 5966 8424
rect 7006 8412 7012 8424
rect 5960 8384 7012 8412
rect 5960 8372 5966 8384
rect 7006 8372 7012 8384
rect 7064 8372 7070 8424
rect 7285 8415 7343 8421
rect 7285 8381 7297 8415
rect 7331 8412 7343 8415
rect 7466 8412 7472 8424
rect 7331 8384 7472 8412
rect 7331 8381 7343 8384
rect 7285 8375 7343 8381
rect 7466 8372 7472 8384
rect 7524 8372 7530 8424
rect 3786 8304 3792 8356
rect 3844 8344 3850 8356
rect 4157 8347 4215 8353
rect 4157 8344 4169 8347
rect 3844 8316 4169 8344
rect 3844 8304 3850 8316
rect 4157 8313 4169 8316
rect 4203 8344 4215 8347
rect 8036 8344 8064 8452
rect 14458 8440 14464 8452
rect 14516 8440 14522 8492
rect 14737 8483 14795 8489
rect 14737 8449 14749 8483
rect 14783 8480 14795 8483
rect 15102 8480 15108 8492
rect 14783 8452 15108 8480
rect 14783 8449 14795 8452
rect 14737 8443 14795 8449
rect 15102 8440 15108 8452
rect 15160 8440 15166 8492
rect 8754 8412 8760 8424
rect 8715 8384 8760 8412
rect 8754 8372 8760 8384
rect 8812 8372 8818 8424
rect 14366 8372 14372 8424
rect 14424 8412 14430 8424
rect 16500 8412 16528 8520
rect 16758 8440 16764 8492
rect 16816 8480 16822 8492
rect 16925 8483 16983 8489
rect 16925 8480 16937 8483
rect 16816 8452 16937 8480
rect 16816 8440 16822 8452
rect 16925 8449 16937 8452
rect 16971 8449 16983 8483
rect 16925 8443 16983 8449
rect 16666 8412 16672 8424
rect 14424 8384 16528 8412
rect 16627 8384 16672 8412
rect 14424 8372 14430 8384
rect 16666 8372 16672 8384
rect 16724 8372 16730 8424
rect 4203 8316 8064 8344
rect 4203 8313 4215 8316
rect 4157 8307 4215 8313
rect 8110 8304 8116 8356
rect 8168 8344 8174 8356
rect 10137 8347 10195 8353
rect 10137 8344 10149 8347
rect 8168 8316 8800 8344
rect 8168 8304 8174 8316
rect 1719 8248 2820 8276
rect 8772 8276 8800 8316
rect 9692 8316 10149 8344
rect 9692 8276 9720 8316
rect 10137 8313 10149 8316
rect 10183 8344 10195 8347
rect 13630 8344 13636 8356
rect 10183 8316 13636 8344
rect 10183 8313 10195 8316
rect 10137 8307 10195 8313
rect 13630 8304 13636 8316
rect 13688 8304 13694 8356
rect 15286 8304 15292 8356
rect 15344 8344 15350 8356
rect 15381 8347 15439 8353
rect 15381 8344 15393 8347
rect 15344 8316 15393 8344
rect 15344 8304 15350 8316
rect 15381 8313 15393 8316
rect 15427 8313 15439 8347
rect 16117 8347 16175 8353
rect 16117 8344 16129 8347
rect 15381 8307 15439 8313
rect 15488 8316 16129 8344
rect 8772 8248 9720 8276
rect 1719 8245 1731 8248
rect 1673 8239 1731 8245
rect 9766 8236 9772 8288
rect 9824 8276 9830 8288
rect 10686 8276 10692 8288
rect 9824 8248 10692 8276
rect 9824 8236 9830 8248
rect 10686 8236 10692 8248
rect 10744 8236 10750 8288
rect 14277 8279 14335 8285
rect 14277 8245 14289 8279
rect 14323 8276 14335 8279
rect 14734 8276 14740 8288
rect 14323 8248 14740 8276
rect 14323 8245 14335 8248
rect 14277 8239 14335 8245
rect 14734 8236 14740 8248
rect 14792 8236 14798 8288
rect 14826 8236 14832 8288
rect 14884 8276 14890 8288
rect 15488 8276 15516 8316
rect 16117 8313 16129 8316
rect 16163 8313 16175 8347
rect 18049 8347 18107 8353
rect 18049 8344 18061 8347
rect 16117 8307 16175 8313
rect 17604 8316 18061 8344
rect 14884 8248 15516 8276
rect 14884 8236 14890 8248
rect 17402 8236 17408 8288
rect 17460 8276 17466 8288
rect 17604 8276 17632 8316
rect 18049 8313 18061 8316
rect 18095 8313 18107 8347
rect 18524 8344 18552 8520
rect 18690 8440 18696 8492
rect 18748 8480 18754 8492
rect 18785 8483 18843 8489
rect 18785 8480 18797 8483
rect 18748 8452 18797 8480
rect 18748 8440 18754 8452
rect 18785 8449 18797 8452
rect 18831 8449 18843 8483
rect 18966 8480 18972 8492
rect 18927 8452 18972 8480
rect 18785 8443 18843 8449
rect 18800 8412 18828 8443
rect 18966 8440 18972 8452
rect 19024 8440 19030 8492
rect 19076 8489 19104 8588
rect 19242 8576 19248 8588
rect 19300 8576 19306 8628
rect 23385 8619 23443 8625
rect 23385 8585 23397 8619
rect 23431 8616 23443 8619
rect 24486 8616 24492 8628
rect 23431 8588 24492 8616
rect 23431 8585 23443 8588
rect 23385 8579 23443 8585
rect 24486 8576 24492 8588
rect 24544 8576 24550 8628
rect 25314 8576 25320 8628
rect 25372 8616 25378 8628
rect 30834 8616 30840 8628
rect 25372 8588 30840 8616
rect 25372 8576 25378 8588
rect 30834 8576 30840 8588
rect 30892 8576 30898 8628
rect 31478 8616 31484 8628
rect 31439 8588 31484 8616
rect 31478 8576 31484 8588
rect 31536 8576 31542 8628
rect 34054 8616 34060 8628
rect 31726 8588 34060 8616
rect 20070 8548 20076 8560
rect 20031 8520 20076 8548
rect 20070 8508 20076 8520
rect 20128 8548 20134 8560
rect 22272 8551 22330 8557
rect 20128 8520 21036 8548
rect 20128 8508 20134 8520
rect 19061 8483 19119 8489
rect 19061 8449 19073 8483
rect 19107 8449 19119 8483
rect 19061 8443 19119 8449
rect 19150 8440 19156 8492
rect 19208 8480 19214 8492
rect 21008 8489 21036 8520
rect 22272 8517 22284 8551
rect 22318 8548 22330 8551
rect 23845 8551 23903 8557
rect 23845 8548 23857 8551
rect 22318 8520 23857 8548
rect 22318 8517 22330 8520
rect 22272 8511 22330 8517
rect 23845 8517 23857 8520
rect 23891 8517 23903 8551
rect 24394 8548 24400 8560
rect 23845 8511 23903 8517
rect 24228 8520 24400 8548
rect 20993 8483 21051 8489
rect 19208 8452 19253 8480
rect 19208 8440 19214 8452
rect 20993 8449 21005 8483
rect 21039 8449 21051 8483
rect 20993 8443 21051 8449
rect 22005 8483 22063 8489
rect 22005 8449 22017 8483
rect 22051 8480 22063 8483
rect 22094 8480 22100 8492
rect 22051 8452 22100 8480
rect 22051 8449 22063 8452
rect 22005 8443 22063 8449
rect 22094 8440 22100 8452
rect 22152 8440 22158 8492
rect 23566 8440 23572 8492
rect 23624 8480 23630 8492
rect 24228 8489 24256 8520
rect 24394 8508 24400 8520
rect 24452 8508 24458 8560
rect 27522 8508 27528 8560
rect 27580 8548 27586 8560
rect 28537 8551 28595 8557
rect 28537 8548 28549 8551
rect 27580 8520 28549 8548
rect 27580 8508 27586 8520
rect 28537 8517 28549 8520
rect 28583 8548 28595 8551
rect 29917 8551 29975 8557
rect 29917 8548 29929 8551
rect 28583 8520 29929 8548
rect 28583 8517 28595 8520
rect 28537 8511 28595 8517
rect 29917 8517 29929 8520
rect 29963 8548 29975 8551
rect 31726 8548 31754 8588
rect 34054 8576 34060 8588
rect 34112 8576 34118 8628
rect 34606 8576 34612 8628
rect 34664 8616 34670 8628
rect 35069 8619 35127 8625
rect 34664 8588 35020 8616
rect 34664 8576 34670 8588
rect 29963 8520 31754 8548
rect 29963 8517 29975 8520
rect 29917 8511 29975 8517
rect 32398 8508 32404 8560
rect 32456 8548 32462 8560
rect 33238 8551 33296 8557
rect 33238 8548 33250 8551
rect 32456 8520 33250 8548
rect 32456 8508 32462 8520
rect 33238 8517 33250 8520
rect 33284 8517 33296 8551
rect 34698 8548 34704 8560
rect 34659 8520 34704 8548
rect 33238 8511 33296 8517
rect 34698 8508 34704 8520
rect 34756 8508 34762 8560
rect 24121 8483 24179 8489
rect 24121 8480 24133 8483
rect 23624 8452 24133 8480
rect 23624 8440 23630 8452
rect 24121 8449 24133 8452
rect 24167 8449 24179 8483
rect 24121 8443 24179 8449
rect 24213 8483 24271 8489
rect 24213 8449 24225 8483
rect 24259 8449 24271 8483
rect 24213 8443 24271 8449
rect 24302 8440 24308 8492
rect 24360 8480 24366 8492
rect 24489 8483 24547 8489
rect 24360 8452 24405 8480
rect 24360 8440 24366 8452
rect 24489 8449 24501 8483
rect 24535 8449 24547 8483
rect 25130 8480 25136 8492
rect 25091 8452 25136 8480
rect 24489 8443 24547 8449
rect 19889 8415 19947 8421
rect 19889 8412 19901 8415
rect 18800 8384 19901 8412
rect 19889 8381 19901 8384
rect 19935 8381 19947 8415
rect 19889 8375 19947 8381
rect 23842 8372 23848 8424
rect 23900 8412 23906 8424
rect 24504 8412 24532 8443
rect 25130 8440 25136 8452
rect 25188 8440 25194 8492
rect 25317 8483 25375 8489
rect 25317 8449 25329 8483
rect 25363 8480 25375 8483
rect 27706 8480 27712 8492
rect 25363 8452 27712 8480
rect 25363 8449 25375 8452
rect 25317 8443 25375 8449
rect 27706 8440 27712 8452
rect 27764 8440 27770 8492
rect 33594 8440 33600 8492
rect 33652 8480 33658 8492
rect 34146 8480 34152 8492
rect 33652 8452 34152 8480
rect 33652 8440 33658 8452
rect 34146 8440 34152 8452
rect 34204 8440 34210 8492
rect 34885 8483 34943 8489
rect 34885 8480 34897 8483
rect 34624 8452 34897 8480
rect 23900 8384 24532 8412
rect 23900 8372 23906 8384
rect 29178 8372 29184 8424
rect 29236 8412 29242 8424
rect 29273 8415 29331 8421
rect 29273 8412 29285 8415
rect 29236 8384 29285 8412
rect 29236 8372 29242 8384
rect 29273 8381 29285 8384
rect 29319 8381 29331 8415
rect 33502 8412 33508 8424
rect 33463 8384 33508 8412
rect 29273 8375 29331 8381
rect 33502 8372 33508 8384
rect 33560 8372 33566 8424
rect 27798 8344 27804 8356
rect 18524 8316 21220 8344
rect 18049 8307 18107 8313
rect 19426 8276 19432 8288
rect 17460 8248 17632 8276
rect 19387 8248 19432 8276
rect 17460 8236 17466 8248
rect 19426 8236 19432 8248
rect 19484 8236 19490 8288
rect 21192 8285 21220 8316
rect 23124 8316 25636 8344
rect 27759 8316 27804 8344
rect 21177 8279 21235 8285
rect 21177 8245 21189 8279
rect 21223 8276 21235 8279
rect 23124 8276 23152 8316
rect 21223 8248 23152 8276
rect 21223 8245 21235 8248
rect 21177 8239 21235 8245
rect 25222 8236 25228 8288
rect 25280 8276 25286 8288
rect 25501 8279 25559 8285
rect 25501 8276 25513 8279
rect 25280 8248 25513 8276
rect 25280 8236 25286 8248
rect 25501 8245 25513 8248
rect 25547 8245 25559 8279
rect 25608 8276 25636 8316
rect 27798 8304 27804 8316
rect 27856 8344 27862 8356
rect 27982 8344 27988 8356
rect 27856 8316 27988 8344
rect 27856 8304 27862 8316
rect 27982 8304 27988 8316
rect 28040 8304 28046 8356
rect 34624 8344 34652 8452
rect 34885 8449 34897 8452
rect 34931 8449 34943 8483
rect 34992 8480 35020 8588
rect 35069 8585 35081 8619
rect 35115 8616 35127 8619
rect 35342 8616 35348 8628
rect 35115 8588 35348 8616
rect 35115 8585 35127 8588
rect 35069 8579 35127 8585
rect 35342 8576 35348 8588
rect 35400 8576 35406 8628
rect 36725 8619 36783 8625
rect 36725 8585 36737 8619
rect 36771 8616 36783 8619
rect 37366 8616 37372 8628
rect 36771 8588 37372 8616
rect 36771 8585 36783 8588
rect 36725 8579 36783 8585
rect 37366 8576 37372 8588
rect 37424 8576 37430 8628
rect 38654 8616 38660 8628
rect 37568 8588 38660 8616
rect 36354 8548 36360 8560
rect 36315 8520 36360 8548
rect 36354 8508 36360 8520
rect 36412 8508 36418 8560
rect 37568 8495 37596 8588
rect 38654 8576 38660 8588
rect 38712 8576 38718 8628
rect 38194 8508 38200 8560
rect 38252 8548 38258 8560
rect 39086 8551 39144 8557
rect 39086 8548 39098 8551
rect 38252 8520 39098 8548
rect 38252 8508 38258 8520
rect 39086 8517 39098 8520
rect 39132 8517 39144 8551
rect 39086 8511 39144 8517
rect 36538 8480 36544 8492
rect 34992 8452 36544 8480
rect 34885 8443 34943 8449
rect 34900 8412 34928 8443
rect 36538 8440 36544 8452
rect 36596 8440 36602 8492
rect 37182 8440 37188 8492
rect 37240 8480 37246 8492
rect 37548 8489 37606 8495
rect 37369 8483 37427 8489
rect 37369 8480 37381 8483
rect 37240 8452 37381 8480
rect 37240 8440 37246 8452
rect 37369 8449 37381 8452
rect 37415 8449 37427 8483
rect 37548 8455 37560 8489
rect 37594 8455 37606 8489
rect 37548 8449 37606 8455
rect 37645 8483 37703 8489
rect 37645 8449 37657 8483
rect 37691 8449 37703 8483
rect 37369 8443 37427 8449
rect 37645 8443 37703 8449
rect 35802 8412 35808 8424
rect 34900 8384 35808 8412
rect 35802 8372 35808 8384
rect 35860 8372 35866 8424
rect 37660 8412 37688 8443
rect 37754 8440 37760 8492
rect 37812 8489 37818 8492
rect 37812 8483 37841 8489
rect 37829 8449 37841 8483
rect 37812 8443 37841 8449
rect 37812 8440 37818 8443
rect 38010 8440 38016 8492
rect 38068 8480 38074 8492
rect 40954 8480 40960 8492
rect 38068 8452 40960 8480
rect 38068 8440 38074 8452
rect 37660 8384 37872 8412
rect 37844 8356 37872 8384
rect 37918 8372 37924 8424
rect 37976 8412 37982 8424
rect 38562 8412 38568 8424
rect 37976 8384 38568 8412
rect 37976 8372 37982 8384
rect 38562 8372 38568 8384
rect 38620 8412 38626 8424
rect 38841 8415 38899 8421
rect 38841 8412 38853 8415
rect 38620 8384 38853 8412
rect 38620 8372 38626 8384
rect 38841 8381 38853 8384
rect 38887 8381 38899 8415
rect 38841 8375 38899 8381
rect 32048 8316 32352 8344
rect 28718 8276 28724 8288
rect 25608 8248 28724 8276
rect 25501 8239 25559 8245
rect 28718 8236 28724 8248
rect 28776 8236 28782 8288
rect 31570 8236 31576 8288
rect 31628 8276 31634 8288
rect 32048 8276 32076 8316
rect 31628 8248 32076 8276
rect 31628 8236 31634 8248
rect 32122 8236 32128 8288
rect 32180 8276 32186 8288
rect 32324 8276 32352 8316
rect 33980 8316 34652 8344
rect 33980 8276 34008 8316
rect 37826 8304 37832 8356
rect 37884 8304 37890 8356
rect 40236 8353 40264 8452
rect 40954 8440 40960 8452
rect 41012 8440 41018 8492
rect 40221 8347 40279 8353
rect 40221 8313 40233 8347
rect 40267 8313 40279 8347
rect 40221 8307 40279 8313
rect 67542 8304 67548 8356
rect 67600 8344 67606 8356
rect 67637 8347 67695 8353
rect 67637 8344 67649 8347
rect 67600 8316 67649 8344
rect 67600 8304 67606 8316
rect 67637 8313 67649 8316
rect 67683 8313 67695 8347
rect 67637 8307 67695 8313
rect 32180 8248 32225 8276
rect 32324 8248 34008 8276
rect 32180 8236 32186 8248
rect 34054 8236 34060 8288
rect 34112 8276 34118 8288
rect 34112 8248 34157 8276
rect 34112 8236 34118 8248
rect 34238 8236 34244 8288
rect 34296 8276 34302 8288
rect 37734 8276 37740 8288
rect 34296 8248 37740 8276
rect 34296 8236 34302 8248
rect 37734 8236 37740 8248
rect 37792 8236 37798 8288
rect 38010 8276 38016 8288
rect 37971 8248 38016 8276
rect 38010 8236 38016 8248
rect 38068 8236 38074 8288
rect 1104 8186 68816 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 65654 8186
rect 65706 8134 65718 8186
rect 65770 8134 65782 8186
rect 65834 8134 65846 8186
rect 65898 8134 65910 8186
rect 65962 8134 68816 8186
rect 1104 8112 68816 8134
rect 1854 8032 1860 8084
rect 1912 8072 1918 8084
rect 2498 8072 2504 8084
rect 1912 8044 2504 8072
rect 1912 8032 1918 8044
rect 2498 8032 2504 8044
rect 2556 8072 2562 8084
rect 2777 8075 2835 8081
rect 2777 8072 2789 8075
rect 2556 8044 2789 8072
rect 2556 8032 2562 8044
rect 2777 8041 2789 8044
rect 2823 8072 2835 8075
rect 3786 8072 3792 8084
rect 2823 8044 3792 8072
rect 2823 8041 2835 8044
rect 2777 8035 2835 8041
rect 3786 8032 3792 8044
rect 3844 8032 3850 8084
rect 8662 8032 8668 8084
rect 8720 8072 8726 8084
rect 15562 8072 15568 8084
rect 8720 8044 15568 8072
rect 8720 8032 8726 8044
rect 15562 8032 15568 8044
rect 15620 8032 15626 8084
rect 16669 8075 16727 8081
rect 16669 8041 16681 8075
rect 16715 8072 16727 8075
rect 16758 8072 16764 8084
rect 16715 8044 16764 8072
rect 16715 8041 16727 8044
rect 16669 8035 16727 8041
rect 16758 8032 16764 8044
rect 16816 8032 16822 8084
rect 18693 8075 18751 8081
rect 18693 8041 18705 8075
rect 18739 8072 18751 8075
rect 18966 8072 18972 8084
rect 18739 8044 18972 8072
rect 18739 8041 18751 8044
rect 18693 8035 18751 8041
rect 18966 8032 18972 8044
rect 19024 8032 19030 8084
rect 25685 8075 25743 8081
rect 25685 8041 25697 8075
rect 25731 8072 25743 8075
rect 25774 8072 25780 8084
rect 25731 8044 25780 8072
rect 25731 8041 25743 8044
rect 25685 8035 25743 8041
rect 25774 8032 25780 8044
rect 25832 8032 25838 8084
rect 28629 8075 28687 8081
rect 28629 8041 28641 8075
rect 28675 8072 28687 8075
rect 28902 8072 28908 8084
rect 28675 8044 28908 8072
rect 28675 8041 28687 8044
rect 28629 8035 28687 8041
rect 28902 8032 28908 8044
rect 28960 8032 28966 8084
rect 31018 8072 31024 8084
rect 30979 8044 31024 8072
rect 31018 8032 31024 8044
rect 31076 8032 31082 8084
rect 31665 8075 31723 8081
rect 31665 8041 31677 8075
rect 31711 8072 31723 8075
rect 31754 8072 31760 8084
rect 31711 8044 31760 8072
rect 31711 8041 31723 8044
rect 31665 8035 31723 8041
rect 31754 8032 31760 8044
rect 31812 8072 31818 8084
rect 32122 8072 32128 8084
rect 31812 8044 32128 8072
rect 31812 8032 31818 8044
rect 32122 8032 32128 8044
rect 32180 8032 32186 8084
rect 33502 8072 33508 8084
rect 32784 8044 33508 8072
rect 5994 7964 6000 8016
rect 6052 8004 6058 8016
rect 6052 7976 8524 8004
rect 6052 7964 6058 7976
rect 2130 7896 2136 7948
rect 2188 7936 2194 7948
rect 2225 7939 2283 7945
rect 2225 7936 2237 7939
rect 2188 7908 2237 7936
rect 2188 7896 2194 7908
rect 2225 7905 2237 7908
rect 2271 7905 2283 7939
rect 2225 7899 2283 7905
rect 6270 7896 6276 7948
rect 6328 7936 6334 7948
rect 6825 7939 6883 7945
rect 6825 7936 6837 7939
rect 6328 7908 6837 7936
rect 6328 7896 6334 7908
rect 6825 7905 6837 7908
rect 6871 7905 6883 7939
rect 8496 7936 8524 7976
rect 8570 7964 8576 8016
rect 8628 8004 8634 8016
rect 11146 8004 11152 8016
rect 8628 7976 11152 8004
rect 8628 7964 8634 7976
rect 11146 7964 11152 7976
rect 11204 7964 11210 8016
rect 14642 7964 14648 8016
rect 14700 7964 14706 8016
rect 9766 7936 9772 7948
rect 8496 7908 9772 7936
rect 6825 7899 6883 7905
rect 9766 7896 9772 7908
rect 9824 7896 9830 7948
rect 1762 7828 1768 7880
rect 1820 7868 1826 7880
rect 1857 7871 1915 7877
rect 1857 7868 1869 7871
rect 1820 7840 1869 7868
rect 1820 7828 1826 7840
rect 1857 7837 1869 7840
rect 1903 7868 1915 7871
rect 5442 7868 5448 7880
rect 1903 7840 5448 7868
rect 1903 7837 1915 7840
rect 1857 7831 1915 7837
rect 5442 7828 5448 7840
rect 5500 7828 5506 7880
rect 6549 7871 6607 7877
rect 6549 7837 6561 7871
rect 6595 7868 6607 7871
rect 7466 7868 7472 7880
rect 6595 7840 7472 7868
rect 6595 7837 6607 7840
rect 6549 7831 6607 7837
rect 7466 7828 7472 7840
rect 7524 7828 7530 7880
rect 12529 7871 12587 7877
rect 12529 7837 12541 7871
rect 12575 7868 12587 7871
rect 12710 7868 12716 7880
rect 12575 7840 12716 7868
rect 12575 7837 12587 7840
rect 12529 7831 12587 7837
rect 12710 7828 12716 7840
rect 12768 7828 12774 7880
rect 14660 7877 14688 7964
rect 15746 7896 15752 7948
rect 15804 7936 15810 7948
rect 21634 7936 21640 7948
rect 15804 7908 18552 7936
rect 21595 7908 21640 7936
rect 15804 7896 15810 7908
rect 18524 7880 18552 7908
rect 21634 7896 21640 7908
rect 21692 7896 21698 7948
rect 25774 7936 25780 7948
rect 25056 7908 25780 7936
rect 14553 7871 14611 7877
rect 14553 7837 14565 7871
rect 14599 7837 14611 7871
rect 14553 7831 14611 7837
rect 14642 7871 14700 7877
rect 14642 7837 14654 7871
rect 14688 7837 14700 7871
rect 14642 7831 14700 7837
rect 2041 7803 2099 7809
rect 2041 7769 2053 7803
rect 2087 7800 2099 7803
rect 2314 7800 2320 7812
rect 2087 7772 2320 7800
rect 2087 7769 2099 7772
rect 2041 7763 2099 7769
rect 2314 7760 2320 7772
rect 2372 7760 2378 7812
rect 5718 7800 5724 7812
rect 5679 7772 5724 7800
rect 5718 7760 5724 7772
rect 5776 7760 5782 7812
rect 5905 7803 5963 7809
rect 5905 7769 5917 7803
rect 5951 7800 5963 7803
rect 6454 7800 6460 7812
rect 5951 7772 6460 7800
rect 5951 7769 5963 7772
rect 5905 7763 5963 7769
rect 6454 7760 6460 7772
rect 6512 7760 6518 7812
rect 7926 7760 7932 7812
rect 7984 7800 7990 7812
rect 8941 7803 8999 7809
rect 8941 7800 8953 7803
rect 7984 7772 8953 7800
rect 7984 7760 7990 7772
rect 8941 7769 8953 7772
rect 8987 7769 8999 7803
rect 12250 7800 12256 7812
rect 12308 7809 12314 7812
rect 12220 7772 12256 7800
rect 8941 7763 8999 7769
rect 12250 7760 12256 7772
rect 12308 7763 12320 7809
rect 12308 7760 12314 7763
rect 5537 7735 5595 7741
rect 5537 7701 5549 7735
rect 5583 7732 5595 7735
rect 5994 7732 6000 7744
rect 5583 7704 6000 7732
rect 5583 7701 5595 7704
rect 5537 7695 5595 7701
rect 5994 7692 6000 7704
rect 6052 7692 6058 7744
rect 8297 7735 8355 7741
rect 8297 7701 8309 7735
rect 8343 7732 8355 7735
rect 8386 7732 8392 7744
rect 8343 7704 8392 7732
rect 8343 7701 8355 7704
rect 8297 7695 8355 7701
rect 8386 7692 8392 7704
rect 8444 7732 8450 7744
rect 9306 7732 9312 7744
rect 8444 7704 9312 7732
rect 8444 7692 8450 7704
rect 9306 7692 9312 7704
rect 9364 7692 9370 7744
rect 13541 7735 13599 7741
rect 13541 7701 13553 7735
rect 13587 7732 13599 7735
rect 13814 7732 13820 7744
rect 13587 7704 13820 7732
rect 13587 7701 13599 7704
rect 13541 7695 13599 7701
rect 13814 7692 13820 7704
rect 13872 7692 13878 7744
rect 14274 7732 14280 7744
rect 14235 7704 14280 7732
rect 14274 7692 14280 7704
rect 14332 7692 14338 7744
rect 14568 7732 14596 7831
rect 14734 7828 14740 7880
rect 14792 7868 14798 7880
rect 14921 7871 14979 7877
rect 14792 7840 14837 7868
rect 14792 7828 14798 7840
rect 14921 7837 14933 7871
rect 14967 7837 14979 7871
rect 15562 7868 15568 7880
rect 15523 7840 15568 7868
rect 14921 7831 14979 7837
rect 14936 7800 14964 7831
rect 15562 7828 15568 7840
rect 15620 7828 15626 7880
rect 16025 7871 16083 7877
rect 16025 7837 16037 7871
rect 16071 7837 16083 7871
rect 16025 7831 16083 7837
rect 16209 7871 16267 7877
rect 16209 7837 16221 7871
rect 16255 7837 16267 7871
rect 16209 7831 16267 7837
rect 16040 7800 16068 7831
rect 16114 7800 16120 7812
rect 14936 7772 16120 7800
rect 16114 7760 16120 7772
rect 16172 7760 16178 7812
rect 16224 7800 16252 7831
rect 16298 7828 16304 7880
rect 16356 7868 16362 7880
rect 16439 7871 16497 7877
rect 16356 7840 16401 7868
rect 16356 7828 16362 7840
rect 16439 7837 16451 7871
rect 16485 7868 16497 7871
rect 16758 7868 16764 7880
rect 16485 7840 16764 7868
rect 16485 7837 16497 7840
rect 16439 7831 16497 7837
rect 16758 7828 16764 7840
rect 16816 7828 16822 7880
rect 17126 7868 17132 7880
rect 17087 7840 17132 7868
rect 17126 7828 17132 7840
rect 17184 7828 17190 7880
rect 17402 7868 17408 7880
rect 17363 7840 17408 7868
rect 17402 7828 17408 7840
rect 17460 7828 17466 7880
rect 18230 7868 18236 7880
rect 18143 7840 18236 7868
rect 18230 7828 18236 7840
rect 18288 7828 18294 7880
rect 18506 7868 18512 7880
rect 18419 7840 18512 7868
rect 18506 7828 18512 7840
rect 18564 7828 18570 7880
rect 19797 7871 19855 7877
rect 19797 7837 19809 7871
rect 19843 7868 19855 7871
rect 19886 7868 19892 7880
rect 19843 7840 19892 7868
rect 19843 7837 19855 7840
rect 19797 7831 19855 7837
rect 19886 7828 19892 7840
rect 19944 7828 19950 7880
rect 21082 7828 21088 7880
rect 21140 7868 21146 7880
rect 25056 7877 25084 7908
rect 25774 7896 25780 7908
rect 25832 7936 25838 7948
rect 26145 7939 26203 7945
rect 26145 7936 26157 7939
rect 25832 7908 26157 7936
rect 25832 7896 25838 7908
rect 26145 7905 26157 7908
rect 26191 7905 26203 7939
rect 28534 7936 28540 7948
rect 28495 7908 28540 7936
rect 26145 7899 26203 7905
rect 28534 7896 28540 7908
rect 28592 7896 28598 7948
rect 31294 7896 31300 7948
rect 31352 7936 31358 7948
rect 31570 7936 31576 7948
rect 31352 7908 31576 7936
rect 31352 7896 31358 7908
rect 31570 7896 31576 7908
rect 31628 7896 31634 7948
rect 21913 7871 21971 7877
rect 21913 7868 21925 7871
rect 21140 7840 21925 7868
rect 21140 7828 21146 7840
rect 21913 7837 21925 7840
rect 21959 7837 21971 7871
rect 25041 7871 25099 7877
rect 25041 7868 25053 7871
rect 21913 7831 21971 7837
rect 23860 7840 25053 7868
rect 17589 7803 17647 7809
rect 17589 7800 17601 7803
rect 16224 7772 17601 7800
rect 17589 7769 17601 7772
rect 17635 7769 17647 7803
rect 18248 7800 18276 7828
rect 23860 7812 23888 7840
rect 25041 7837 25053 7840
rect 25087 7837 25099 7871
rect 25222 7868 25228 7880
rect 25183 7840 25228 7868
rect 25041 7831 25099 7837
rect 25222 7828 25228 7840
rect 25280 7828 25286 7880
rect 25317 7871 25375 7877
rect 25317 7837 25329 7871
rect 25363 7837 25375 7871
rect 25317 7831 25375 7837
rect 19242 7800 19248 7812
rect 18248 7772 19248 7800
rect 17589 7763 17647 7769
rect 19242 7760 19248 7772
rect 19300 7760 19306 7812
rect 19426 7760 19432 7812
rect 19484 7800 19490 7812
rect 20042 7803 20100 7809
rect 20042 7800 20054 7803
rect 19484 7772 20054 7800
rect 19484 7760 19490 7772
rect 20042 7769 20054 7772
rect 20088 7769 20100 7803
rect 20042 7763 20100 7769
rect 22186 7760 22192 7812
rect 22244 7800 22250 7812
rect 23842 7800 23848 7812
rect 22244 7772 23848 7800
rect 22244 7760 22250 7772
rect 23842 7760 23848 7772
rect 23900 7760 23906 7812
rect 24670 7760 24676 7812
rect 24728 7800 24734 7812
rect 25332 7800 25360 7831
rect 25406 7828 25412 7880
rect 25464 7868 25470 7880
rect 28629 7871 28687 7877
rect 25464 7840 25509 7868
rect 25464 7828 25470 7840
rect 28629 7837 28641 7871
rect 28675 7837 28687 7871
rect 28629 7831 28687 7837
rect 28350 7800 28356 7812
rect 24728 7772 25360 7800
rect 28311 7772 28356 7800
rect 24728 7760 24734 7772
rect 28350 7760 28356 7772
rect 28408 7760 28414 7812
rect 28442 7760 28448 7812
rect 28500 7800 28506 7812
rect 28644 7800 28672 7831
rect 29178 7828 29184 7880
rect 29236 7868 29242 7880
rect 29641 7871 29699 7877
rect 29641 7868 29653 7871
rect 29236 7840 29653 7868
rect 29236 7828 29242 7840
rect 29641 7837 29653 7840
rect 29687 7837 29699 7871
rect 29641 7831 29699 7837
rect 29730 7828 29736 7880
rect 29788 7868 29794 7880
rect 29897 7871 29955 7877
rect 29897 7868 29909 7871
rect 29788 7840 29909 7868
rect 29788 7828 29794 7840
rect 29897 7837 29909 7840
rect 29943 7837 29955 7871
rect 29897 7831 29955 7837
rect 31018 7828 31024 7880
rect 31076 7868 31082 7880
rect 32784 7877 32812 8044
rect 33502 8032 33508 8044
rect 33560 8072 33566 8084
rect 34146 8072 34152 8084
rect 33560 8044 33732 8072
rect 34107 8044 34152 8072
rect 33560 8032 33566 8044
rect 33704 8004 33732 8044
rect 34146 8032 34152 8044
rect 34204 8032 34210 8084
rect 35802 8032 35808 8084
rect 35860 8072 35866 8084
rect 35989 8075 36047 8081
rect 35989 8072 36001 8075
rect 35860 8044 36001 8072
rect 35860 8032 35866 8044
rect 35989 8041 36001 8044
rect 36035 8041 36047 8075
rect 39298 8072 39304 8084
rect 39259 8044 39304 8072
rect 35989 8035 36047 8041
rect 39298 8032 39304 8044
rect 39356 8032 39362 8084
rect 34514 8004 34520 8016
rect 33704 7976 34520 8004
rect 34514 7964 34520 7976
rect 34572 7964 34578 8016
rect 33042 7877 33048 7880
rect 31757 7871 31815 7877
rect 31757 7868 31769 7871
rect 31076 7840 31769 7868
rect 31076 7828 31082 7840
rect 31757 7837 31769 7840
rect 31803 7837 31815 7871
rect 31757 7831 31815 7837
rect 32769 7871 32827 7877
rect 32769 7837 32781 7871
rect 32815 7837 32827 7871
rect 32769 7831 32827 7837
rect 33036 7831 33048 7877
rect 33100 7868 33106 7880
rect 33100 7840 33136 7868
rect 33042 7828 33048 7831
rect 33100 7828 33106 7840
rect 35710 7828 35716 7880
rect 35768 7868 35774 7880
rect 37369 7871 37427 7877
rect 37369 7868 37381 7871
rect 35768 7840 37381 7868
rect 35768 7828 35774 7840
rect 37369 7837 37381 7840
rect 37415 7868 37427 7871
rect 37918 7868 37924 7880
rect 37415 7840 37924 7868
rect 37415 7837 37427 7840
rect 37369 7831 37427 7837
rect 37918 7828 37924 7840
rect 37976 7828 37982 7880
rect 38010 7828 38016 7880
rect 38068 7868 38074 7880
rect 38177 7871 38235 7877
rect 38177 7868 38189 7871
rect 38068 7840 38189 7868
rect 38068 7828 38074 7840
rect 38177 7837 38189 7840
rect 38223 7837 38235 7871
rect 38177 7831 38235 7837
rect 28500 7772 28672 7800
rect 28500 7760 28506 7772
rect 29546 7760 29552 7812
rect 29604 7800 29610 7812
rect 31481 7803 31539 7809
rect 31481 7800 31493 7803
rect 29604 7772 31493 7800
rect 29604 7760 29610 7772
rect 31481 7769 31493 7772
rect 31527 7800 31539 7803
rect 31527 7772 32904 7800
rect 31527 7769 31539 7772
rect 31481 7763 31539 7769
rect 14918 7732 14924 7744
rect 14568 7704 14924 7732
rect 14918 7692 14924 7704
rect 14976 7692 14982 7744
rect 15010 7692 15016 7744
rect 15068 7732 15074 7744
rect 17221 7735 17279 7741
rect 17221 7732 17233 7735
rect 15068 7704 17233 7732
rect 15068 7692 15074 7704
rect 17221 7701 17233 7704
rect 17267 7701 17279 7735
rect 18322 7732 18328 7744
rect 18283 7704 18328 7732
rect 17221 7695 17279 7701
rect 18322 7692 18328 7704
rect 18380 7692 18386 7744
rect 18506 7692 18512 7744
rect 18564 7732 18570 7744
rect 21177 7735 21235 7741
rect 21177 7732 21189 7735
rect 18564 7704 21189 7732
rect 18564 7692 18570 7704
rect 21177 7701 21189 7704
rect 21223 7701 21235 7735
rect 21177 7695 21235 7701
rect 23106 7692 23112 7744
rect 23164 7732 23170 7744
rect 23201 7735 23259 7741
rect 23201 7732 23213 7735
rect 23164 7704 23213 7732
rect 23164 7692 23170 7704
rect 23201 7701 23213 7704
rect 23247 7732 23259 7735
rect 23566 7732 23572 7744
rect 23247 7704 23572 7732
rect 23247 7701 23259 7704
rect 23201 7695 23259 7701
rect 23566 7692 23572 7704
rect 23624 7692 23630 7744
rect 24118 7692 24124 7744
rect 24176 7732 24182 7744
rect 24486 7732 24492 7744
rect 24176 7704 24492 7732
rect 24176 7692 24182 7704
rect 24486 7692 24492 7704
rect 24544 7732 24550 7744
rect 26142 7732 26148 7744
rect 24544 7704 26148 7732
rect 24544 7692 24550 7704
rect 26142 7692 26148 7704
rect 26200 7692 26206 7744
rect 28813 7735 28871 7741
rect 28813 7701 28825 7735
rect 28859 7732 28871 7735
rect 29822 7732 29828 7744
rect 28859 7704 29828 7732
rect 28859 7701 28871 7704
rect 28813 7695 28871 7701
rect 29822 7692 29828 7704
rect 29880 7692 29886 7744
rect 31938 7732 31944 7744
rect 31899 7704 31944 7732
rect 31938 7692 31944 7704
rect 31996 7692 32002 7744
rect 32876 7732 32904 7772
rect 37090 7760 37096 7812
rect 37148 7809 37154 7812
rect 37148 7800 37160 7809
rect 37148 7772 37193 7800
rect 37148 7763 37160 7772
rect 37148 7760 37154 7763
rect 34790 7732 34796 7744
rect 32876 7704 34796 7732
rect 34790 7692 34796 7704
rect 34848 7692 34854 7744
rect 1104 7642 68816 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 50294 7642
rect 50346 7590 50358 7642
rect 50410 7590 50422 7642
rect 50474 7590 50486 7642
rect 50538 7590 50550 7642
rect 50602 7590 68816 7642
rect 1104 7568 68816 7590
rect 2406 7528 2412 7540
rect 2367 7500 2412 7528
rect 2406 7488 2412 7500
rect 2464 7488 2470 7540
rect 5537 7531 5595 7537
rect 5537 7497 5549 7531
rect 5583 7528 5595 7531
rect 5718 7528 5724 7540
rect 5583 7500 5724 7528
rect 5583 7497 5595 7500
rect 5537 7491 5595 7497
rect 5718 7488 5724 7500
rect 5776 7488 5782 7540
rect 8662 7528 8668 7540
rect 6656 7500 8668 7528
rect 4172 7432 6224 7460
rect 3510 7352 3516 7404
rect 3568 7392 3574 7404
rect 4172 7401 4200 7432
rect 4157 7395 4215 7401
rect 4157 7392 4169 7395
rect 3568 7364 4169 7392
rect 3568 7352 3574 7364
rect 4157 7361 4169 7364
rect 4203 7361 4215 7395
rect 4157 7355 4215 7361
rect 4424 7395 4482 7401
rect 4424 7361 4436 7395
rect 4470 7392 4482 7395
rect 5534 7392 5540 7404
rect 4470 7364 5540 7392
rect 4470 7361 4482 7364
rect 4424 7355 4482 7361
rect 5534 7352 5540 7364
rect 5592 7352 5598 7404
rect 6196 7324 6224 7432
rect 6454 7392 6460 7404
rect 6415 7364 6460 7392
rect 6454 7352 6460 7364
rect 6512 7352 6518 7404
rect 6656 7401 6684 7500
rect 8662 7488 8668 7500
rect 8720 7488 8726 7540
rect 9766 7528 9772 7540
rect 9727 7500 9772 7528
rect 9766 7488 9772 7500
rect 9824 7488 9830 7540
rect 12250 7528 12256 7540
rect 12211 7500 12256 7528
rect 12250 7488 12256 7500
rect 12308 7488 12314 7540
rect 13078 7488 13084 7540
rect 13136 7528 13142 7540
rect 18322 7528 18328 7540
rect 13136 7500 18328 7528
rect 13136 7488 13142 7500
rect 8754 7460 8760 7472
rect 7300 7432 8760 7460
rect 7300 7401 7328 7432
rect 8754 7420 8760 7432
rect 8812 7420 8818 7472
rect 11146 7420 11152 7472
rect 11204 7460 11210 7472
rect 12980 7463 13038 7469
rect 11204 7432 12112 7460
rect 11204 7420 11210 7432
rect 7558 7401 7564 7404
rect 6641 7395 6699 7401
rect 6641 7361 6653 7395
rect 6687 7361 6699 7395
rect 6641 7355 6699 7361
rect 7285 7395 7343 7401
rect 7285 7361 7297 7395
rect 7331 7361 7343 7395
rect 7285 7355 7343 7361
rect 7552 7355 7564 7401
rect 7616 7392 7622 7404
rect 11514 7392 11520 7404
rect 7616 7364 7652 7392
rect 11475 7364 11520 7392
rect 7300 7324 7328 7355
rect 7558 7352 7564 7355
rect 7616 7352 7622 7364
rect 11514 7352 11520 7364
rect 11572 7352 11578 7404
rect 11698 7392 11704 7404
rect 11659 7364 11704 7392
rect 11698 7352 11704 7364
rect 11756 7352 11762 7404
rect 12084 7401 12112 7432
rect 12980 7429 12992 7463
rect 13026 7460 13038 7463
rect 14274 7460 14280 7472
rect 13026 7432 14280 7460
rect 13026 7429 13038 7432
rect 12980 7423 13038 7429
rect 14274 7420 14280 7432
rect 14332 7420 14338 7472
rect 12069 7395 12127 7401
rect 12069 7361 12081 7395
rect 12115 7361 12127 7395
rect 12069 7355 12127 7361
rect 12636 7364 14596 7392
rect 6196 7296 7328 7324
rect 11606 7284 11612 7336
rect 11664 7324 11670 7336
rect 11793 7327 11851 7333
rect 11793 7324 11805 7327
rect 11664 7296 11805 7324
rect 11664 7284 11670 7296
rect 11793 7293 11805 7296
rect 11839 7293 11851 7327
rect 11793 7287 11851 7293
rect 11885 7327 11943 7333
rect 11885 7293 11897 7327
rect 11931 7324 11943 7327
rect 12526 7324 12532 7336
rect 11931 7296 12532 7324
rect 11931 7293 11943 7296
rect 11885 7287 11943 7293
rect 12526 7284 12532 7296
rect 12584 7284 12590 7336
rect 6104 7228 7236 7256
rect 2314 7148 2320 7200
rect 2372 7188 2378 7200
rect 3053 7191 3111 7197
rect 3053 7188 3065 7191
rect 2372 7160 3065 7188
rect 2372 7148 2378 7160
rect 3053 7157 3065 7160
rect 3099 7188 3111 7191
rect 6104 7188 6132 7228
rect 3099 7160 6132 7188
rect 6825 7191 6883 7197
rect 3099 7157 3111 7160
rect 3053 7151 3111 7157
rect 6825 7157 6837 7191
rect 6871 7188 6883 7191
rect 7098 7188 7104 7200
rect 6871 7160 7104 7188
rect 6871 7157 6883 7160
rect 6825 7151 6883 7157
rect 7098 7148 7104 7160
rect 7156 7148 7162 7200
rect 7208 7188 7236 7228
rect 9030 7216 9036 7268
rect 9088 7256 9094 7268
rect 9217 7259 9275 7265
rect 9217 7256 9229 7259
rect 9088 7228 9229 7256
rect 9088 7216 9094 7228
rect 9217 7225 9229 7228
rect 9263 7256 9275 7259
rect 12636 7256 12664 7364
rect 12710 7284 12716 7336
rect 12768 7324 12774 7336
rect 12768 7296 12861 7324
rect 12768 7284 12774 7296
rect 9263 7228 12664 7256
rect 9263 7225 9275 7228
rect 9217 7219 9275 7225
rect 7926 7188 7932 7200
rect 7208 7160 7932 7188
rect 7926 7148 7932 7160
rect 7984 7148 7990 7200
rect 10226 7188 10232 7200
rect 10187 7160 10232 7188
rect 10226 7148 10232 7160
rect 10284 7148 10290 7200
rect 10965 7191 11023 7197
rect 10965 7157 10977 7191
rect 11011 7188 11023 7191
rect 11330 7188 11336 7200
rect 11011 7160 11336 7188
rect 11011 7157 11023 7160
rect 10965 7151 11023 7157
rect 11330 7148 11336 7160
rect 11388 7148 11394 7200
rect 12728 7188 12756 7284
rect 14568 7256 14596 7364
rect 14660 7324 14688 7500
rect 18322 7488 18328 7500
rect 18380 7528 18386 7540
rect 19426 7528 19432 7540
rect 18380 7500 19432 7528
rect 18380 7488 18386 7500
rect 19426 7488 19432 7500
rect 19484 7488 19490 7540
rect 19981 7531 20039 7537
rect 19981 7497 19993 7531
rect 20027 7528 20039 7531
rect 20070 7528 20076 7540
rect 20027 7500 20076 7528
rect 20027 7497 20039 7500
rect 19981 7491 20039 7497
rect 20070 7488 20076 7500
rect 20128 7528 20134 7540
rect 20441 7531 20499 7537
rect 20441 7528 20453 7531
rect 20128 7500 20453 7528
rect 20128 7488 20134 7500
rect 20441 7497 20453 7500
rect 20487 7497 20499 7531
rect 20441 7491 20499 7497
rect 25590 7488 25596 7540
rect 25648 7528 25654 7540
rect 29273 7531 29331 7537
rect 25648 7500 28856 7528
rect 25648 7488 25654 7500
rect 21269 7463 21327 7469
rect 21269 7460 21281 7463
rect 14844 7432 21281 7460
rect 14737 7327 14795 7333
rect 14737 7324 14749 7327
rect 14660 7296 14749 7324
rect 14737 7293 14749 7296
rect 14783 7293 14795 7327
rect 14737 7287 14795 7293
rect 14844 7256 14872 7432
rect 21269 7429 21281 7432
rect 21315 7460 21327 7463
rect 22186 7460 22192 7472
rect 21315 7432 22192 7460
rect 21315 7429 21327 7432
rect 21269 7423 21327 7429
rect 22186 7420 22192 7432
rect 22244 7420 22250 7472
rect 22554 7460 22560 7472
rect 22388 7432 22560 7460
rect 19150 7352 19156 7404
rect 19208 7392 19214 7404
rect 19245 7395 19303 7401
rect 19245 7392 19257 7395
rect 19208 7364 19257 7392
rect 19208 7352 19214 7364
rect 19245 7361 19257 7364
rect 19291 7361 19303 7395
rect 21082 7392 21088 7404
rect 21043 7364 21088 7392
rect 19245 7355 19303 7361
rect 21082 7352 21088 7364
rect 21140 7352 21146 7404
rect 22388 7401 22416 7432
rect 22554 7420 22560 7432
rect 22612 7460 22618 7472
rect 24302 7460 24308 7472
rect 22612 7432 24308 7460
rect 22612 7420 22618 7432
rect 24302 7420 24308 7432
rect 24360 7420 24366 7472
rect 26421 7463 26479 7469
rect 24688 7432 26096 7460
rect 22281 7395 22339 7401
rect 22281 7361 22293 7395
rect 22327 7361 22339 7395
rect 22281 7355 22339 7361
rect 22373 7395 22431 7401
rect 22373 7361 22385 7395
rect 22419 7361 22431 7395
rect 22373 7355 22431 7361
rect 15010 7324 15016 7336
rect 14971 7296 15016 7324
rect 15010 7284 15016 7296
rect 15068 7284 15074 7336
rect 16758 7284 16764 7336
rect 16816 7324 16822 7336
rect 18969 7327 19027 7333
rect 18969 7324 18981 7327
rect 16816 7296 18981 7324
rect 16816 7284 16822 7296
rect 18969 7293 18981 7296
rect 19015 7293 19027 7327
rect 22296 7324 22324 7355
rect 22462 7352 22468 7404
rect 22520 7392 22526 7404
rect 22520 7364 22565 7392
rect 22520 7352 22526 7364
rect 22646 7352 22652 7404
rect 22704 7392 22710 7404
rect 24394 7392 24400 7404
rect 22704 7364 22749 7392
rect 24355 7364 24400 7392
rect 22704 7352 22710 7364
rect 24394 7352 24400 7364
rect 24452 7352 24458 7404
rect 24688 7336 24716 7432
rect 25774 7392 25780 7404
rect 25735 7364 25780 7392
rect 25774 7352 25780 7364
rect 25832 7352 25838 7404
rect 26068 7401 26096 7432
rect 26421 7429 26433 7463
rect 26467 7460 26479 7463
rect 26467 7432 26924 7460
rect 26467 7429 26479 7432
rect 26421 7423 26479 7429
rect 25961 7395 26019 7401
rect 25961 7361 25973 7395
rect 26007 7361 26019 7395
rect 25961 7355 26019 7361
rect 26053 7395 26111 7401
rect 26053 7361 26065 7395
rect 26099 7361 26111 7395
rect 26053 7355 26111 7361
rect 23109 7327 23167 7333
rect 23109 7324 23121 7327
rect 22296 7296 23121 7324
rect 18969 7287 19027 7293
rect 14568 7228 14872 7256
rect 13722 7188 13728 7200
rect 12728 7160 13728 7188
rect 13722 7148 13728 7160
rect 13780 7148 13786 7200
rect 14093 7191 14151 7197
rect 14093 7157 14105 7191
rect 14139 7188 14151 7191
rect 14458 7188 14464 7200
rect 14139 7160 14464 7188
rect 14139 7157 14151 7160
rect 14093 7151 14151 7157
rect 14458 7148 14464 7160
rect 14516 7148 14522 7200
rect 14734 7148 14740 7200
rect 14792 7188 14798 7200
rect 15028 7188 15056 7284
rect 22388 7268 22416 7296
rect 23109 7293 23121 7296
rect 23155 7324 23167 7327
rect 23290 7324 23296 7336
rect 23155 7296 23296 7324
rect 23155 7293 23167 7296
rect 23109 7287 23167 7293
rect 23290 7284 23296 7296
rect 23348 7284 23354 7336
rect 24670 7324 24676 7336
rect 24631 7296 24676 7324
rect 24670 7284 24676 7296
rect 24728 7284 24734 7336
rect 16482 7216 16488 7268
rect 16540 7256 16546 7268
rect 17681 7259 17739 7265
rect 17681 7256 17693 7259
rect 16540 7228 17693 7256
rect 16540 7216 16546 7228
rect 17681 7225 17693 7228
rect 17727 7225 17739 7259
rect 17681 7219 17739 7225
rect 22370 7216 22376 7268
rect 22428 7216 22434 7268
rect 25976 7256 26004 7355
rect 26142 7352 26148 7404
rect 26200 7392 26206 7404
rect 26896 7392 26924 7432
rect 28828 7401 28856 7500
rect 29273 7497 29285 7531
rect 29319 7497 29331 7531
rect 29273 7491 29331 7497
rect 32861 7531 32919 7537
rect 32861 7497 32873 7531
rect 32907 7528 32919 7531
rect 33226 7528 33232 7540
rect 32907 7500 33232 7528
rect 32907 7497 32919 7500
rect 32861 7491 32919 7497
rect 27229 7395 27287 7401
rect 27229 7392 27241 7395
rect 26200 7364 26245 7392
rect 26896 7364 27241 7392
rect 26200 7352 26206 7364
rect 27229 7361 27241 7364
rect 27275 7361 27287 7395
rect 27229 7355 27287 7361
rect 28813 7395 28871 7401
rect 28813 7361 28825 7395
rect 28859 7361 28871 7395
rect 28813 7355 28871 7361
rect 29089 7395 29147 7401
rect 29089 7361 29101 7395
rect 29135 7361 29147 7395
rect 29288 7392 29316 7491
rect 33226 7488 33232 7500
rect 33284 7488 33290 7540
rect 34701 7531 34759 7537
rect 34701 7497 34713 7531
rect 34747 7528 34759 7531
rect 34790 7528 34796 7540
rect 34747 7500 34796 7528
rect 34747 7497 34759 7500
rect 34701 7491 34759 7497
rect 34790 7488 34796 7500
rect 34848 7488 34854 7540
rect 37369 7531 37427 7537
rect 37369 7497 37381 7531
rect 37415 7528 37427 7531
rect 37734 7528 37740 7540
rect 37415 7500 37740 7528
rect 37415 7497 37427 7500
rect 37369 7491 37427 7497
rect 37734 7488 37740 7500
rect 37792 7488 37798 7540
rect 34514 7420 34520 7472
rect 34572 7460 34578 7472
rect 35710 7460 35716 7472
rect 34572 7432 35716 7460
rect 34572 7420 34578 7432
rect 35710 7420 35716 7432
rect 35768 7460 35774 7472
rect 35768 7432 36124 7460
rect 35768 7420 35774 7432
rect 29733 7395 29791 7401
rect 29733 7392 29745 7395
rect 29288 7364 29745 7392
rect 29089 7355 29147 7361
rect 29733 7361 29745 7364
rect 29779 7361 29791 7395
rect 29733 7355 29791 7361
rect 26234 7284 26240 7336
rect 26292 7324 26298 7336
rect 26970 7324 26976 7336
rect 26292 7296 26976 7324
rect 26292 7284 26298 7296
rect 26970 7284 26976 7296
rect 27028 7284 27034 7336
rect 28258 7284 28264 7336
rect 28316 7324 28322 7336
rect 28902 7324 28908 7336
rect 28316 7296 28908 7324
rect 28316 7284 28322 7296
rect 28902 7284 28908 7296
rect 28960 7324 28966 7336
rect 28997 7327 29055 7333
rect 28997 7324 29009 7327
rect 28960 7296 29009 7324
rect 28960 7284 28966 7296
rect 28997 7293 29009 7296
rect 29043 7293 29055 7327
rect 29104 7324 29132 7355
rect 29822 7352 29828 7404
rect 29880 7392 29886 7404
rect 29880 7364 29925 7392
rect 29880 7352 29886 7364
rect 35526 7352 35532 7404
rect 35584 7392 35590 7404
rect 36096 7401 36124 7432
rect 35814 7395 35872 7401
rect 35814 7392 35826 7395
rect 35584 7364 35826 7392
rect 35584 7352 35590 7364
rect 35814 7361 35826 7364
rect 35860 7361 35872 7395
rect 35814 7355 35872 7361
rect 36081 7395 36139 7401
rect 36081 7361 36093 7395
rect 36127 7361 36139 7395
rect 36081 7355 36139 7361
rect 30650 7324 30656 7336
rect 29104 7296 30656 7324
rect 28997 7287 29055 7293
rect 30650 7284 30656 7296
rect 30708 7284 30714 7336
rect 26602 7256 26608 7268
rect 25976 7228 26608 7256
rect 26602 7216 26608 7228
rect 26660 7216 26666 7268
rect 28092 7228 29776 7256
rect 14792 7160 15056 7188
rect 14792 7148 14798 7160
rect 15838 7148 15844 7200
rect 15896 7188 15902 7200
rect 16025 7191 16083 7197
rect 16025 7188 16037 7191
rect 15896 7160 16037 7188
rect 15896 7148 15902 7160
rect 16025 7157 16037 7160
rect 16071 7157 16083 7191
rect 16025 7151 16083 7157
rect 16942 7148 16948 7200
rect 17000 7188 17006 7200
rect 17037 7191 17095 7197
rect 17037 7188 17049 7191
rect 17000 7160 17049 7188
rect 17000 7148 17006 7160
rect 17037 7157 17049 7160
rect 17083 7157 17095 7191
rect 17037 7151 17095 7157
rect 22005 7191 22063 7197
rect 22005 7157 22017 7191
rect 22051 7188 22063 7191
rect 22186 7188 22192 7200
rect 22051 7160 22192 7188
rect 22051 7157 22063 7160
rect 22005 7151 22063 7157
rect 22186 7148 22192 7160
rect 22244 7148 22250 7200
rect 23750 7148 23756 7200
rect 23808 7188 23814 7200
rect 23845 7191 23903 7197
rect 23845 7188 23857 7191
rect 23808 7160 23857 7188
rect 23808 7148 23814 7160
rect 23845 7157 23857 7160
rect 23891 7188 23903 7191
rect 24854 7188 24860 7200
rect 23891 7160 24860 7188
rect 23891 7157 23903 7160
rect 23845 7151 23903 7157
rect 24854 7148 24860 7160
rect 24912 7188 24918 7200
rect 25406 7188 25412 7200
rect 24912 7160 25412 7188
rect 24912 7148 24918 7160
rect 25406 7148 25412 7160
rect 25464 7148 25470 7200
rect 27338 7148 27344 7200
rect 27396 7188 27402 7200
rect 28092 7188 28120 7228
rect 27396 7160 28120 7188
rect 28353 7191 28411 7197
rect 27396 7148 27402 7160
rect 28353 7157 28365 7191
rect 28399 7188 28411 7191
rect 28534 7188 28540 7200
rect 28399 7160 28540 7188
rect 28399 7157 28411 7160
rect 28353 7151 28411 7157
rect 28534 7148 28540 7160
rect 28592 7148 28598 7200
rect 29089 7191 29147 7197
rect 29089 7157 29101 7191
rect 29135 7188 29147 7191
rect 29638 7188 29644 7200
rect 29135 7160 29644 7188
rect 29135 7157 29147 7160
rect 29089 7151 29147 7157
rect 29638 7148 29644 7160
rect 29696 7148 29702 7200
rect 29748 7197 29776 7228
rect 29733 7191 29791 7197
rect 29733 7157 29745 7191
rect 29779 7157 29791 7191
rect 29733 7151 29791 7157
rect 30101 7191 30159 7197
rect 30101 7157 30113 7191
rect 30147 7188 30159 7191
rect 30926 7188 30932 7200
rect 30147 7160 30932 7188
rect 30147 7157 30159 7160
rect 30101 7151 30159 7157
rect 30926 7148 30932 7160
rect 30984 7148 30990 7200
rect 1104 7098 68816 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 65654 7098
rect 65706 7046 65718 7098
rect 65770 7046 65782 7098
rect 65834 7046 65846 7098
rect 65898 7046 65910 7098
rect 65962 7046 68816 7098
rect 1104 7024 68816 7046
rect 7558 6984 7564 6996
rect 7519 6956 7564 6984
rect 7558 6944 7564 6956
rect 7616 6944 7622 6996
rect 11330 6984 11336 6996
rect 7668 6956 11336 6984
rect 4062 6876 4068 6928
rect 4120 6916 4126 6928
rect 6178 6916 6184 6928
rect 4120 6888 6184 6916
rect 4120 6876 4126 6888
rect 6178 6876 6184 6888
rect 6236 6916 6242 6928
rect 7668 6916 7696 6956
rect 11330 6944 11336 6956
rect 11388 6944 11394 6996
rect 11606 6984 11612 6996
rect 11567 6956 11612 6984
rect 11606 6944 11612 6956
rect 11664 6944 11670 6996
rect 12342 6944 12348 6996
rect 12400 6984 12406 6996
rect 12526 6984 12532 6996
rect 12400 6956 12532 6984
rect 12400 6944 12406 6956
rect 12526 6944 12532 6956
rect 12584 6944 12590 6996
rect 18690 6984 18696 6996
rect 16592 6956 18696 6984
rect 6236 6888 7696 6916
rect 6236 6876 6242 6888
rect 11514 6876 11520 6928
rect 11572 6916 11578 6928
rect 12250 6916 12256 6928
rect 11572 6888 12256 6916
rect 11572 6876 11578 6888
rect 12250 6876 12256 6888
rect 12308 6916 12314 6928
rect 16592 6916 16620 6956
rect 18690 6944 18696 6956
rect 18748 6944 18754 6996
rect 26970 6944 26976 6996
rect 27028 6984 27034 6996
rect 29178 6984 29184 6996
rect 27028 6956 29184 6984
rect 27028 6944 27034 6956
rect 29178 6944 29184 6956
rect 29236 6944 29242 6996
rect 29638 6944 29644 6996
rect 29696 6984 29702 6996
rect 30193 6987 30251 6993
rect 30193 6984 30205 6987
rect 29696 6956 30205 6984
rect 29696 6944 29702 6956
rect 30193 6953 30205 6956
rect 30239 6953 30251 6987
rect 31846 6984 31852 6996
rect 31807 6956 31852 6984
rect 30193 6947 30251 6953
rect 31846 6944 31852 6956
rect 31904 6944 31910 6996
rect 16758 6916 16764 6928
rect 12308 6888 16620 6916
rect 16684 6888 16764 6916
rect 12308 6876 12314 6888
rect 5534 6848 5540 6860
rect 5495 6820 5540 6848
rect 5534 6808 5540 6820
rect 5592 6808 5598 6860
rect 8662 6848 8668 6860
rect 6932 6820 8668 6848
rect 1765 6783 1823 6789
rect 1765 6749 1777 6783
rect 1811 6749 1823 6783
rect 1946 6780 1952 6792
rect 1907 6752 1952 6780
rect 1765 6743 1823 6749
rect 1780 6644 1808 6743
rect 1946 6740 1952 6752
rect 2004 6740 2010 6792
rect 2038 6740 2044 6792
rect 2096 6780 2102 6792
rect 2179 6783 2237 6789
rect 2096 6752 2141 6780
rect 2096 6740 2102 6752
rect 2179 6749 2191 6783
rect 2225 6780 2237 6783
rect 2869 6783 2927 6789
rect 2869 6780 2881 6783
rect 2225 6752 2881 6780
rect 2225 6749 2237 6752
rect 2179 6743 2237 6749
rect 2869 6749 2881 6752
rect 2915 6780 2927 6783
rect 3050 6780 3056 6792
rect 2915 6752 3056 6780
rect 2915 6749 2927 6752
rect 2869 6743 2927 6749
rect 3050 6740 3056 6752
rect 3108 6780 3114 6792
rect 4062 6780 4068 6792
rect 3108 6752 4068 6780
rect 3108 6740 3114 6752
rect 4062 6740 4068 6752
rect 4120 6740 4126 6792
rect 5718 6740 5724 6792
rect 5776 6780 5782 6792
rect 5813 6783 5871 6789
rect 5813 6780 5825 6783
rect 5776 6752 5825 6780
rect 5776 6740 5782 6752
rect 5813 6749 5825 6752
rect 5859 6749 5871 6783
rect 5813 6743 5871 6749
rect 5905 6783 5963 6789
rect 5905 6749 5917 6783
rect 5951 6749 5963 6783
rect 5905 6743 5963 6749
rect 2409 6715 2467 6721
rect 2409 6681 2421 6715
rect 2455 6712 2467 6715
rect 2958 6712 2964 6724
rect 2455 6684 2964 6712
rect 2455 6681 2467 6684
rect 2409 6675 2467 6681
rect 2958 6672 2964 6684
rect 3016 6672 3022 6724
rect 5920 6712 5948 6743
rect 5994 6740 6000 6792
rect 6052 6780 6058 6792
rect 6181 6783 6239 6789
rect 6052 6752 6097 6780
rect 6052 6740 6058 6752
rect 6181 6749 6193 6783
rect 6227 6780 6239 6783
rect 6270 6780 6276 6792
rect 6227 6752 6276 6780
rect 6227 6749 6239 6752
rect 6181 6743 6239 6749
rect 6270 6740 6276 6752
rect 6328 6740 6334 6792
rect 6932 6789 6960 6820
rect 8662 6808 8668 6820
rect 8720 6808 8726 6860
rect 8754 6808 8760 6860
rect 8812 6848 8818 6860
rect 9125 6851 9183 6857
rect 9125 6848 9137 6851
rect 8812 6820 9137 6848
rect 8812 6808 8818 6820
rect 9125 6817 9137 6820
rect 9171 6817 9183 6851
rect 9125 6811 9183 6817
rect 13541 6851 13599 6857
rect 13541 6817 13553 6851
rect 13587 6848 13599 6851
rect 15010 6848 15016 6860
rect 13587 6820 15016 6848
rect 13587 6817 13599 6820
rect 13541 6811 13599 6817
rect 15010 6808 15016 6820
rect 15068 6808 15074 6860
rect 16574 6848 16580 6860
rect 16408 6820 16580 6848
rect 6917 6783 6975 6789
rect 6917 6749 6929 6783
rect 6963 6749 6975 6783
rect 7098 6780 7104 6792
rect 7059 6752 7104 6780
rect 6917 6743 6975 6749
rect 7098 6740 7104 6752
rect 7156 6740 7162 6792
rect 7193 6783 7251 6789
rect 7193 6749 7205 6783
rect 7239 6749 7251 6783
rect 7193 6743 7251 6749
rect 6730 6712 6736 6724
rect 5920 6684 6736 6712
rect 6730 6672 6736 6684
rect 6788 6712 6794 6724
rect 7208 6712 7236 6743
rect 7282 6740 7288 6792
rect 7340 6780 7346 6792
rect 7340 6752 7385 6780
rect 7340 6740 7346 6752
rect 7466 6740 7472 6792
rect 7524 6780 7530 6792
rect 11054 6780 11060 6792
rect 7524 6752 10640 6780
rect 11015 6752 11060 6780
rect 7524 6740 7530 6752
rect 6788 6684 7236 6712
rect 6788 6672 6794 6684
rect 9214 6672 9220 6724
rect 9272 6712 9278 6724
rect 9370 6715 9428 6721
rect 9370 6712 9382 6715
rect 9272 6684 9382 6712
rect 9272 6672 9278 6684
rect 9370 6681 9382 6684
rect 9416 6681 9428 6715
rect 9370 6675 9428 6681
rect 2498 6644 2504 6656
rect 1780 6616 2504 6644
rect 2498 6604 2504 6616
rect 2556 6644 2562 6656
rect 3510 6644 3516 6656
rect 2556 6616 3516 6644
rect 2556 6604 2562 6616
rect 3510 6604 3516 6616
rect 3568 6644 3574 6656
rect 3789 6647 3847 6653
rect 3789 6644 3801 6647
rect 3568 6616 3801 6644
rect 3568 6604 3574 6616
rect 3789 6613 3801 6616
rect 3835 6613 3847 6647
rect 8294 6644 8300 6656
rect 8255 6616 8300 6644
rect 3789 6607 3847 6613
rect 8294 6604 8300 6616
rect 8352 6604 8358 6656
rect 10410 6604 10416 6656
rect 10468 6644 10474 6656
rect 10505 6647 10563 6653
rect 10505 6644 10517 6647
rect 10468 6616 10517 6644
rect 10468 6604 10474 6616
rect 10505 6613 10517 6616
rect 10551 6613 10563 6647
rect 10612 6644 10640 6752
rect 11054 6740 11060 6752
rect 11112 6740 11118 6792
rect 11149 6783 11207 6789
rect 11149 6749 11161 6783
rect 11195 6749 11207 6783
rect 11330 6780 11336 6792
rect 11291 6752 11336 6780
rect 11149 6743 11207 6749
rect 11164 6712 11192 6743
rect 11330 6740 11336 6752
rect 11388 6740 11394 6792
rect 11422 6740 11428 6792
rect 11480 6780 11486 6792
rect 12253 6783 12311 6789
rect 11480 6752 11525 6780
rect 11480 6740 11486 6752
rect 12253 6749 12265 6783
rect 12299 6780 12311 6783
rect 12897 6783 12955 6789
rect 12897 6780 12909 6783
rect 12299 6752 12909 6780
rect 12299 6749 12311 6752
rect 12253 6743 12311 6749
rect 12897 6749 12909 6752
rect 12943 6780 12955 6783
rect 13998 6780 14004 6792
rect 12943 6752 14004 6780
rect 12943 6749 12955 6752
rect 12897 6743 12955 6749
rect 13998 6740 14004 6752
rect 14056 6740 14062 6792
rect 14274 6740 14280 6792
rect 14332 6780 14338 6792
rect 14369 6783 14427 6789
rect 14369 6780 14381 6783
rect 14332 6752 14381 6780
rect 14332 6740 14338 6752
rect 14369 6749 14381 6752
rect 14415 6749 14427 6783
rect 14369 6743 14427 6749
rect 14645 6783 14703 6789
rect 14645 6749 14657 6783
rect 14691 6780 14703 6783
rect 15654 6780 15660 6792
rect 14691 6752 15660 6780
rect 14691 6749 14703 6752
rect 14645 6743 14703 6749
rect 12434 6712 12440 6724
rect 11164 6684 12440 6712
rect 12434 6672 12440 6684
rect 12492 6672 12498 6724
rect 12342 6644 12348 6656
rect 10612 6616 12348 6644
rect 10505 6607 10563 6613
rect 12342 6604 12348 6616
rect 12400 6604 12406 6656
rect 12713 6647 12771 6653
rect 12713 6613 12725 6647
rect 12759 6644 12771 6647
rect 12802 6644 12808 6656
rect 12759 6616 12808 6644
rect 12759 6613 12771 6616
rect 12713 6607 12771 6613
rect 12802 6604 12808 6616
rect 12860 6604 12866 6656
rect 14384 6644 14412 6743
rect 15654 6740 15660 6752
rect 15712 6780 15718 6792
rect 16114 6780 16120 6792
rect 15712 6752 16120 6780
rect 15712 6740 15718 6752
rect 16114 6740 16120 6752
rect 16172 6740 16178 6792
rect 16298 6780 16304 6792
rect 16259 6752 16304 6780
rect 16298 6740 16304 6752
rect 16356 6740 16362 6792
rect 16408 6789 16436 6820
rect 16574 6808 16580 6820
rect 16632 6808 16638 6860
rect 16393 6783 16451 6789
rect 16393 6749 16405 6783
rect 16439 6749 16451 6783
rect 16393 6743 16451 6749
rect 16485 6783 16543 6789
rect 16485 6749 16497 6783
rect 16531 6780 16543 6783
rect 16684 6780 16712 6888
rect 16758 6876 16764 6888
rect 16816 6876 16822 6928
rect 28902 6876 28908 6928
rect 28960 6916 28966 6928
rect 28960 6888 30420 6916
rect 28960 6876 28966 6888
rect 19150 6808 19156 6860
rect 19208 6848 19214 6860
rect 19337 6851 19395 6857
rect 19337 6848 19349 6851
rect 19208 6820 19349 6848
rect 19208 6808 19214 6820
rect 19337 6817 19349 6820
rect 19383 6817 19395 6851
rect 19978 6848 19984 6860
rect 19939 6820 19984 6848
rect 19337 6811 19395 6817
rect 19978 6808 19984 6820
rect 20036 6808 20042 6860
rect 22094 6808 22100 6860
rect 22152 6848 22158 6860
rect 22152 6820 22197 6848
rect 22152 6808 22158 6820
rect 24394 6808 24400 6860
rect 24452 6848 24458 6860
rect 24489 6851 24547 6857
rect 24489 6848 24501 6851
rect 24452 6820 24501 6848
rect 24452 6808 24458 6820
rect 24489 6817 24501 6820
rect 24535 6817 24547 6851
rect 26602 6848 26608 6860
rect 26563 6820 26608 6848
rect 24489 6811 24547 6817
rect 26602 6808 26608 6820
rect 26660 6808 26666 6860
rect 30392 6857 30420 6888
rect 30377 6851 30435 6857
rect 30377 6817 30389 6851
rect 30423 6848 30435 6851
rect 30558 6848 30564 6860
rect 30423 6820 30564 6848
rect 30423 6817 30435 6820
rect 30377 6811 30435 6817
rect 30558 6808 30564 6820
rect 30616 6808 30622 6860
rect 30926 6808 30932 6860
rect 30984 6848 30990 6860
rect 30984 6820 35388 6848
rect 30984 6808 30990 6820
rect 16531 6752 16712 6780
rect 16531 6749 16543 6752
rect 16485 6743 16543 6749
rect 14918 6672 14924 6724
rect 14976 6712 14982 6724
rect 16500 6712 16528 6743
rect 17218 6740 17224 6792
rect 17276 6780 17282 6792
rect 17313 6783 17371 6789
rect 17313 6780 17325 6783
rect 17276 6752 17325 6780
rect 17276 6740 17282 6752
rect 17313 6749 17325 6752
rect 17359 6749 17371 6783
rect 17954 6780 17960 6792
rect 17915 6752 17960 6780
rect 17313 6743 17371 6749
rect 17954 6740 17960 6752
rect 18012 6740 18018 6792
rect 19242 6780 19248 6792
rect 19203 6752 19248 6780
rect 19242 6740 19248 6752
rect 19300 6740 19306 6792
rect 19426 6780 19432 6792
rect 19387 6752 19432 6780
rect 19426 6740 19432 6752
rect 19484 6740 19490 6792
rect 21082 6780 21088 6792
rect 19996 6752 21088 6780
rect 19996 6712 20024 6752
rect 21082 6740 21088 6752
rect 21140 6740 21146 6792
rect 22186 6740 22192 6792
rect 22244 6780 22250 6792
rect 22353 6783 22411 6789
rect 22353 6780 22365 6783
rect 22244 6752 22365 6780
rect 22244 6740 22250 6752
rect 22353 6749 22365 6752
rect 22399 6749 22411 6783
rect 22353 6743 22411 6749
rect 24302 6740 24308 6792
rect 24360 6780 24366 6792
rect 24765 6783 24823 6789
rect 24765 6780 24777 6783
rect 24360 6752 24777 6780
rect 24360 6740 24366 6752
rect 24765 6749 24777 6752
rect 24811 6749 24823 6783
rect 24765 6743 24823 6749
rect 14976 6684 16528 6712
rect 16684 6684 20024 6712
rect 14976 6672 14982 6684
rect 16684 6644 16712 6684
rect 20070 6672 20076 6724
rect 20128 6712 20134 6724
rect 20226 6715 20284 6721
rect 20226 6712 20238 6715
rect 20128 6684 20238 6712
rect 20128 6672 20134 6684
rect 20226 6681 20238 6684
rect 20272 6681 20284 6715
rect 20226 6675 20284 6681
rect 14384 6616 16712 6644
rect 16761 6647 16819 6653
rect 16761 6613 16773 6647
rect 16807 6644 16819 6647
rect 16850 6644 16856 6656
rect 16807 6616 16856 6644
rect 16807 6613 16819 6616
rect 16761 6607 16819 6613
rect 16850 6604 16856 6616
rect 16908 6604 16914 6656
rect 18506 6604 18512 6656
rect 18564 6644 18570 6656
rect 18601 6647 18659 6653
rect 18601 6644 18613 6647
rect 18564 6616 18613 6644
rect 18564 6604 18570 6616
rect 18601 6613 18613 6616
rect 18647 6613 18659 6647
rect 18601 6607 18659 6613
rect 20346 6604 20352 6656
rect 20404 6644 20410 6656
rect 21361 6647 21419 6653
rect 21361 6644 21373 6647
rect 20404 6616 21373 6644
rect 20404 6604 20410 6616
rect 21361 6613 21373 6616
rect 21407 6613 21419 6647
rect 21361 6607 21419 6613
rect 23477 6647 23535 6653
rect 23477 6613 23489 6647
rect 23523 6644 23535 6647
rect 23658 6644 23664 6656
rect 23523 6616 23664 6644
rect 23523 6613 23535 6616
rect 23477 6607 23535 6613
rect 23658 6604 23664 6616
rect 23716 6604 23722 6656
rect 24780 6644 24808 6743
rect 25130 6740 25136 6792
rect 25188 6780 25194 6792
rect 26237 6783 26295 6789
rect 26237 6780 26249 6783
rect 25188 6752 26249 6780
rect 25188 6740 25194 6752
rect 26237 6749 26249 6752
rect 26283 6749 26295 6783
rect 26237 6743 26295 6749
rect 29822 6740 29828 6792
rect 29880 6780 29886 6792
rect 30193 6783 30251 6789
rect 30193 6780 30205 6783
rect 29880 6752 30205 6780
rect 29880 6740 29886 6752
rect 30193 6749 30205 6752
rect 30239 6749 30251 6783
rect 30193 6743 30251 6749
rect 30469 6783 30527 6789
rect 30469 6749 30481 6783
rect 30515 6780 30527 6783
rect 30650 6780 30656 6792
rect 30515 6752 30656 6780
rect 30515 6749 30527 6752
rect 30469 6743 30527 6749
rect 30650 6740 30656 6752
rect 30708 6740 30714 6792
rect 32030 6780 32036 6792
rect 31991 6752 32036 6780
rect 32030 6740 32036 6752
rect 32088 6740 32094 6792
rect 32125 6783 32183 6789
rect 32125 6749 32137 6783
rect 32171 6780 32183 6783
rect 32214 6780 32220 6792
rect 32171 6752 32220 6780
rect 32171 6749 32183 6752
rect 32125 6743 32183 6749
rect 32214 6740 32220 6752
rect 32272 6740 32278 6792
rect 34790 6740 34796 6792
rect 34848 6780 34854 6792
rect 35360 6789 35388 6820
rect 34885 6783 34943 6789
rect 34885 6780 34897 6783
rect 34848 6752 34897 6780
rect 34848 6740 34854 6752
rect 34885 6749 34897 6752
rect 34931 6749 34943 6783
rect 34885 6743 34943 6749
rect 35161 6783 35219 6789
rect 35161 6749 35173 6783
rect 35207 6749 35219 6783
rect 35161 6743 35219 6749
rect 35345 6783 35403 6789
rect 35345 6749 35357 6783
rect 35391 6749 35403 6783
rect 68094 6780 68100 6792
rect 68055 6752 68100 6780
rect 35345 6743 35403 6749
rect 26421 6715 26479 6721
rect 26421 6681 26433 6715
rect 26467 6712 26479 6715
rect 28534 6712 28540 6724
rect 26467 6684 28540 6712
rect 26467 6681 26479 6684
rect 26421 6675 26479 6681
rect 28534 6672 28540 6684
rect 28592 6672 28598 6724
rect 31849 6715 31907 6721
rect 31849 6681 31861 6715
rect 31895 6712 31907 6715
rect 31938 6712 31944 6724
rect 31895 6684 31944 6712
rect 31895 6681 31907 6684
rect 31849 6675 31907 6681
rect 31938 6672 31944 6684
rect 31996 6672 32002 6724
rect 35176 6712 35204 6743
rect 68094 6740 68100 6752
rect 68152 6740 68158 6792
rect 32324 6684 35204 6712
rect 28258 6644 28264 6656
rect 24780 6616 28264 6644
rect 28258 6604 28264 6616
rect 28316 6604 28322 6656
rect 30653 6647 30711 6653
rect 30653 6613 30665 6647
rect 30699 6644 30711 6647
rect 31662 6644 31668 6656
rect 30699 6616 31668 6644
rect 30699 6613 30711 6616
rect 30653 6607 30711 6613
rect 31662 6604 31668 6616
rect 31720 6604 31726 6656
rect 32324 6653 32352 6684
rect 32309 6647 32367 6653
rect 32309 6613 32321 6647
rect 32355 6613 32367 6647
rect 32309 6607 32367 6613
rect 33778 6604 33784 6656
rect 33836 6644 33842 6656
rect 34701 6647 34759 6653
rect 34701 6644 34713 6647
rect 33836 6616 34713 6644
rect 33836 6604 33842 6616
rect 34701 6613 34713 6616
rect 34747 6613 34759 6647
rect 34701 6607 34759 6613
rect 1104 6554 68816 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 50294 6554
rect 50346 6502 50358 6554
rect 50410 6502 50422 6554
rect 50474 6502 50486 6554
rect 50538 6502 50550 6554
rect 50602 6502 68816 6554
rect 1104 6480 68816 6502
rect 1946 6400 1952 6452
rect 2004 6440 2010 6452
rect 2133 6443 2191 6449
rect 2133 6440 2145 6443
rect 2004 6412 2145 6440
rect 2004 6400 2010 6412
rect 2133 6409 2145 6412
rect 2179 6409 2191 6443
rect 4062 6440 4068 6452
rect 4023 6412 4068 6440
rect 2133 6403 2191 6409
rect 4062 6400 4068 6412
rect 4120 6400 4126 6452
rect 6454 6440 6460 6452
rect 6415 6412 6460 6440
rect 6454 6400 6460 6412
rect 6512 6440 6518 6452
rect 9214 6440 9220 6452
rect 6512 6412 7788 6440
rect 6512 6400 6518 6412
rect 1762 6372 1768 6384
rect 1723 6344 1768 6372
rect 1762 6332 1768 6344
rect 1820 6332 1826 6384
rect 2774 6372 2780 6384
rect 2700 6344 2780 6372
rect 2700 6313 2728 6344
rect 2774 6332 2780 6344
rect 2832 6372 2838 6384
rect 3418 6372 3424 6384
rect 2832 6344 3424 6372
rect 2832 6332 2838 6344
rect 3418 6332 3424 6344
rect 3476 6332 3482 6384
rect 7760 6381 7788 6412
rect 7944 6412 8892 6440
rect 9175 6412 9220 6440
rect 7944 6381 7972 6412
rect 7745 6375 7803 6381
rect 7745 6341 7757 6375
rect 7791 6341 7803 6375
rect 7745 6335 7803 6341
rect 7929 6375 7987 6381
rect 7929 6341 7941 6375
rect 7975 6341 7987 6375
rect 7929 6335 7987 6341
rect 8113 6375 8171 6381
rect 8113 6341 8125 6375
rect 8159 6372 8171 6375
rect 8864 6372 8892 6412
rect 9214 6400 9220 6412
rect 9272 6400 9278 6452
rect 9766 6400 9772 6452
rect 9824 6440 9830 6452
rect 9824 6412 10548 6440
rect 9824 6400 9830 6412
rect 10410 6372 10416 6384
rect 8159 6344 8800 6372
rect 8864 6344 10416 6372
rect 8159 6341 8171 6344
rect 8113 6335 8171 6341
rect 2958 6313 2964 6316
rect 1949 6307 2007 6313
rect 1949 6273 1961 6307
rect 1995 6273 2007 6307
rect 1949 6267 2007 6273
rect 2685 6307 2743 6313
rect 2685 6273 2697 6307
rect 2731 6273 2743 6307
rect 2685 6267 2743 6273
rect 2952 6267 2964 6313
rect 3016 6304 3022 6316
rect 3016 6276 3052 6304
rect 1964 6168 1992 6267
rect 2958 6264 2964 6267
rect 3016 6264 3022 6276
rect 5810 6264 5816 6316
rect 5868 6304 5874 6316
rect 6638 6304 6644 6316
rect 5868 6276 6644 6304
rect 5868 6264 5874 6276
rect 6638 6264 6644 6276
rect 6696 6264 6702 6316
rect 8573 6307 8631 6313
rect 8573 6273 8585 6307
rect 8619 6304 8631 6307
rect 8662 6304 8668 6316
rect 8619 6276 8668 6304
rect 8619 6273 8631 6276
rect 8573 6267 8631 6273
rect 8662 6264 8668 6276
rect 8720 6264 8726 6316
rect 8772 6313 8800 6344
rect 10410 6332 10416 6344
rect 10468 6332 10474 6384
rect 10520 6372 10548 6412
rect 10594 6400 10600 6452
rect 10652 6440 10658 6452
rect 14918 6440 14924 6452
rect 10652 6412 12940 6440
rect 10652 6400 10658 6412
rect 10870 6372 10876 6384
rect 10520 6344 10876 6372
rect 10870 6332 10876 6344
rect 10928 6332 10934 6384
rect 12434 6372 12440 6384
rect 11650 6344 12440 6372
rect 8757 6307 8815 6313
rect 8757 6273 8769 6307
rect 8803 6273 8815 6307
rect 8757 6267 8815 6273
rect 8849 6307 8907 6313
rect 8849 6273 8861 6307
rect 8895 6273 8907 6307
rect 8849 6267 8907 6273
rect 8941 6307 8999 6313
rect 8941 6273 8953 6307
rect 8987 6273 8999 6307
rect 8941 6267 8999 6273
rect 6730 6196 6736 6248
rect 6788 6236 6794 6248
rect 8864 6236 8892 6267
rect 6788 6208 8892 6236
rect 8956 6236 8984 6267
rect 9122 6264 9128 6316
rect 9180 6304 9186 6316
rect 11054 6304 11060 6316
rect 9180 6276 11060 6304
rect 9180 6264 9186 6276
rect 11054 6264 11060 6276
rect 11112 6304 11118 6316
rect 11650 6313 11678 6344
rect 12434 6332 12440 6344
rect 12492 6332 12498 6384
rect 11609 6307 11678 6313
rect 11112 6294 11468 6304
rect 11507 6297 11565 6303
rect 11507 6294 11519 6297
rect 11112 6276 11519 6294
rect 11112 6264 11118 6276
rect 11440 6266 11519 6276
rect 11507 6263 11519 6266
rect 11553 6263 11565 6297
rect 11609 6273 11621 6307
rect 11655 6273 11678 6307
rect 11720 6307 11778 6313
rect 11720 6304 11732 6307
rect 11609 6267 11678 6273
rect 11624 6266 11678 6267
rect 11716 6273 11732 6304
rect 11766 6273 11778 6307
rect 11716 6267 11778 6273
rect 11882 6307 11940 6313
rect 11882 6273 11894 6307
rect 11928 6304 11940 6307
rect 11974 6304 11980 6316
rect 11928 6276 11980 6304
rect 11928 6273 11940 6276
rect 11882 6267 11940 6273
rect 11507 6257 11565 6263
rect 9214 6236 9220 6248
rect 8956 6208 9220 6236
rect 6788 6196 6794 6208
rect 1964 6140 2360 6168
rect 2332 6100 2360 6140
rect 8294 6128 8300 6180
rect 8352 6168 8358 6180
rect 8662 6168 8668 6180
rect 8352 6140 8668 6168
rect 8352 6128 8358 6140
rect 8662 6128 8668 6140
rect 8720 6168 8726 6180
rect 8956 6168 8984 6208
rect 9214 6196 9220 6208
rect 9272 6196 9278 6248
rect 9861 6239 9919 6245
rect 9861 6205 9873 6239
rect 9907 6236 9919 6239
rect 11238 6236 11244 6248
rect 9907 6208 11244 6236
rect 9907 6205 9919 6208
rect 9861 6199 9919 6205
rect 11238 6196 11244 6208
rect 11296 6196 11302 6248
rect 8720 6140 8984 6168
rect 8720 6128 8726 6140
rect 11422 6128 11428 6180
rect 11480 6168 11486 6180
rect 11716 6168 11744 6267
rect 11974 6264 11980 6276
rect 12032 6264 12038 6316
rect 12158 6264 12164 6316
rect 12216 6304 12222 6316
rect 12805 6307 12863 6313
rect 12805 6304 12817 6307
rect 12216 6276 12817 6304
rect 12216 6264 12222 6276
rect 12805 6273 12817 6276
rect 12851 6273 12863 6307
rect 12805 6267 12863 6273
rect 12529 6239 12587 6245
rect 12529 6205 12541 6239
rect 12575 6236 12587 6239
rect 12912 6236 12940 6412
rect 14200 6412 14924 6440
rect 14200 6313 14228 6412
rect 14918 6400 14924 6412
rect 14976 6400 14982 6452
rect 16114 6400 16120 6452
rect 16172 6440 16178 6452
rect 19337 6443 19395 6449
rect 16172 6412 19288 6440
rect 16172 6400 16178 6412
rect 16022 6372 16028 6384
rect 14292 6344 16028 6372
rect 14292 6313 14320 6344
rect 16022 6332 16028 6344
rect 16080 6332 16086 6384
rect 16666 6332 16672 6384
rect 16724 6372 16730 6384
rect 16724 6344 17816 6372
rect 16724 6332 16730 6344
rect 14185 6307 14243 6313
rect 14185 6273 14197 6307
rect 14231 6273 14243 6307
rect 14185 6267 14243 6273
rect 14277 6307 14335 6313
rect 14277 6273 14289 6307
rect 14323 6273 14335 6307
rect 14277 6267 14335 6273
rect 14366 6264 14372 6316
rect 14424 6304 14430 6316
rect 14553 6307 14611 6313
rect 14424 6276 14469 6304
rect 14424 6264 14430 6276
rect 14553 6273 14565 6307
rect 14599 6273 14611 6307
rect 14553 6267 14611 6273
rect 14090 6236 14096 6248
rect 12575 6208 14096 6236
rect 12575 6205 12587 6208
rect 12529 6199 12587 6205
rect 14090 6196 14096 6208
rect 14148 6196 14154 6248
rect 14568 6236 14596 6267
rect 14918 6264 14924 6316
rect 14976 6304 14982 6316
rect 15243 6307 15301 6313
rect 15243 6304 15255 6307
rect 14976 6276 15255 6304
rect 14976 6264 14982 6276
rect 15243 6273 15255 6276
rect 15289 6273 15301 6307
rect 15378 6304 15384 6316
rect 15339 6276 15384 6304
rect 15243 6267 15301 6273
rect 15378 6264 15384 6276
rect 15436 6264 15442 6316
rect 15470 6264 15476 6316
rect 15528 6304 15534 6316
rect 15528 6276 15573 6304
rect 15528 6264 15534 6276
rect 15654 6264 15660 6316
rect 15712 6304 15718 6316
rect 16776 6313 16804 6344
rect 16761 6307 16819 6313
rect 15712 6276 15757 6304
rect 15712 6264 15718 6276
rect 16761 6273 16773 6307
rect 16807 6273 16819 6307
rect 16761 6267 16819 6273
rect 16850 6264 16856 6316
rect 16908 6304 16914 6316
rect 17017 6307 17075 6313
rect 17017 6304 17029 6307
rect 16908 6276 17029 6304
rect 16908 6264 16914 6276
rect 17017 6273 17029 6276
rect 17063 6273 17075 6307
rect 17017 6267 17075 6273
rect 15672 6236 15700 6264
rect 14568 6208 15700 6236
rect 17788 6236 17816 6344
rect 18598 6332 18604 6384
rect 18656 6372 18662 6384
rect 18656 6344 19012 6372
rect 18656 6332 18662 6344
rect 18690 6304 18696 6316
rect 18651 6276 18696 6304
rect 18690 6264 18696 6276
rect 18748 6264 18754 6316
rect 18874 6304 18880 6316
rect 18835 6276 18880 6304
rect 18874 6264 18880 6276
rect 18932 6264 18938 6316
rect 18984 6313 19012 6344
rect 18969 6307 19027 6313
rect 18969 6273 18981 6307
rect 19015 6273 19027 6307
rect 18969 6267 19027 6273
rect 19061 6307 19119 6313
rect 19061 6273 19073 6307
rect 19107 6304 19119 6307
rect 19150 6304 19156 6316
rect 19107 6276 19156 6304
rect 19107 6273 19119 6276
rect 19061 6267 19119 6273
rect 19150 6264 19156 6276
rect 19208 6264 19214 6316
rect 19260 6304 19288 6412
rect 19337 6409 19349 6443
rect 19383 6440 19395 6443
rect 20070 6440 20076 6452
rect 19383 6412 20076 6440
rect 19383 6409 19395 6412
rect 19337 6403 19395 6409
rect 20070 6400 20076 6412
rect 20128 6400 20134 6452
rect 22462 6400 22468 6452
rect 22520 6440 22526 6452
rect 23109 6443 23167 6449
rect 23109 6440 23121 6443
rect 22520 6412 23121 6440
rect 22520 6400 22526 6412
rect 23109 6409 23121 6412
rect 23155 6409 23167 6443
rect 23109 6403 23167 6409
rect 23474 6400 23480 6452
rect 23532 6440 23538 6452
rect 25593 6443 25651 6449
rect 25593 6440 25605 6443
rect 23532 6412 25605 6440
rect 23532 6400 23538 6412
rect 25593 6409 25605 6412
rect 25639 6409 25651 6443
rect 25593 6403 25651 6409
rect 27617 6443 27675 6449
rect 27617 6409 27629 6443
rect 27663 6440 27675 6443
rect 27706 6440 27712 6452
rect 27663 6412 27712 6440
rect 27663 6409 27675 6412
rect 27617 6403 27675 6409
rect 23293 6375 23351 6381
rect 23293 6341 23305 6375
rect 23339 6372 23351 6375
rect 23658 6372 23664 6384
rect 23339 6344 23664 6372
rect 23339 6341 23351 6344
rect 23293 6335 23351 6341
rect 23658 6332 23664 6344
rect 23716 6332 23722 6384
rect 24210 6332 24216 6384
rect 24268 6372 24274 6384
rect 24489 6375 24547 6381
rect 24489 6372 24501 6375
rect 24268 6344 24501 6372
rect 24268 6332 24274 6344
rect 24489 6341 24501 6344
rect 24535 6341 24547 6375
rect 24489 6335 24547 6341
rect 24578 6332 24584 6384
rect 24636 6372 24642 6384
rect 24636 6344 25452 6372
rect 24636 6332 24642 6344
rect 19797 6307 19855 6313
rect 19797 6304 19809 6307
rect 19260 6276 19809 6304
rect 19797 6273 19809 6276
rect 19843 6273 19855 6307
rect 19797 6267 19855 6273
rect 21082 6264 21088 6316
rect 21140 6304 21146 6316
rect 21821 6307 21879 6313
rect 21821 6304 21833 6307
rect 21140 6276 21833 6304
rect 21140 6264 21146 6276
rect 21821 6273 21833 6276
rect 21867 6273 21879 6307
rect 21821 6267 21879 6273
rect 22097 6307 22155 6313
rect 22097 6273 22109 6307
rect 22143 6304 22155 6307
rect 22186 6304 22192 6316
rect 22143 6276 22192 6304
rect 22143 6273 22155 6276
rect 22097 6267 22155 6273
rect 22186 6264 22192 6276
rect 22244 6304 22250 6316
rect 22646 6304 22652 6316
rect 22244 6276 22652 6304
rect 22244 6264 22250 6276
rect 22646 6264 22652 6276
rect 22704 6264 22710 6316
rect 23474 6304 23480 6316
rect 23435 6276 23480 6304
rect 23474 6264 23480 6276
rect 23532 6264 23538 6316
rect 19978 6236 19984 6248
rect 17788 6208 19984 6236
rect 19978 6196 19984 6208
rect 20036 6196 20042 6248
rect 23676 6236 23704 6332
rect 24762 6304 24768 6316
rect 24675 6276 24768 6304
rect 24762 6264 24768 6276
rect 24820 6304 24826 6316
rect 24946 6304 24952 6316
rect 24820 6276 24952 6304
rect 24820 6264 24826 6276
rect 24946 6264 24952 6276
rect 25004 6264 25010 6316
rect 25424 6313 25452 6344
rect 25409 6307 25467 6313
rect 25409 6273 25421 6307
rect 25455 6273 25467 6307
rect 25608 6304 25636 6403
rect 27706 6400 27712 6412
rect 27764 6440 27770 6452
rect 27890 6440 27896 6452
rect 27764 6412 27896 6440
rect 27764 6400 27770 6412
rect 27890 6400 27896 6412
rect 27948 6400 27954 6452
rect 30561 6443 30619 6449
rect 30561 6409 30573 6443
rect 30607 6440 30619 6443
rect 30650 6440 30656 6452
rect 30607 6412 30656 6440
rect 30607 6409 30619 6412
rect 30561 6403 30619 6409
rect 30650 6400 30656 6412
rect 30708 6400 30714 6452
rect 31573 6443 31631 6449
rect 31573 6409 31585 6443
rect 31619 6440 31631 6443
rect 31846 6440 31852 6452
rect 31619 6412 31852 6440
rect 31619 6409 31631 6412
rect 31573 6403 31631 6409
rect 31846 6400 31852 6412
rect 31904 6400 31910 6452
rect 32030 6400 32036 6452
rect 32088 6440 32094 6452
rect 32401 6443 32459 6449
rect 32401 6440 32413 6443
rect 32088 6412 32413 6440
rect 32088 6400 32094 6412
rect 32401 6409 32413 6412
rect 32447 6409 32459 6443
rect 32401 6403 32459 6409
rect 34517 6443 34575 6449
rect 34517 6409 34529 6443
rect 34563 6440 34575 6443
rect 34563 6412 35296 6440
rect 34563 6409 34575 6412
rect 34517 6403 34575 6409
rect 27908 6304 27936 6400
rect 28077 6375 28135 6381
rect 28077 6341 28089 6375
rect 28123 6372 28135 6375
rect 29426 6375 29484 6381
rect 29426 6372 29438 6375
rect 28123 6344 29438 6372
rect 28123 6341 28135 6344
rect 28077 6335 28135 6341
rect 29426 6341 29438 6344
rect 29472 6341 29484 6375
rect 33686 6372 33692 6384
rect 29426 6335 29484 6341
rect 32600 6344 33692 6372
rect 28353 6307 28411 6313
rect 28353 6304 28365 6307
rect 25608 6276 27844 6304
rect 27908 6276 28365 6304
rect 25409 6267 25467 6273
rect 24581 6239 24639 6245
rect 24581 6236 24593 6239
rect 23676 6208 24593 6236
rect 24581 6205 24593 6208
rect 24627 6205 24639 6239
rect 27816 6236 27844 6276
rect 28353 6273 28365 6276
rect 28399 6273 28411 6307
rect 28353 6267 28411 6273
rect 28442 6307 28500 6313
rect 28442 6273 28454 6307
rect 28488 6273 28500 6307
rect 28442 6267 28500 6273
rect 28074 6236 28080 6248
rect 27816 6208 28080 6236
rect 24581 6199 24639 6205
rect 28074 6196 28080 6208
rect 28132 6196 28138 6248
rect 28258 6196 28264 6248
rect 28316 6236 28322 6248
rect 28457 6236 28485 6267
rect 28534 6264 28540 6316
rect 28592 6313 28598 6316
rect 28592 6304 28600 6313
rect 28721 6307 28779 6313
rect 28592 6276 28637 6304
rect 28592 6267 28600 6276
rect 28721 6273 28733 6307
rect 28767 6304 28779 6307
rect 28994 6304 29000 6316
rect 28767 6276 29000 6304
rect 28767 6273 28779 6276
rect 28721 6267 28779 6273
rect 28592 6264 28598 6267
rect 28994 6264 29000 6276
rect 29052 6264 29058 6316
rect 29178 6304 29184 6316
rect 29139 6276 29184 6304
rect 29178 6264 29184 6276
rect 29236 6264 29242 6316
rect 32600 6313 32628 6344
rect 33686 6332 33692 6344
rect 33744 6332 33750 6384
rect 35268 6381 35296 6412
rect 35253 6375 35311 6381
rect 35253 6341 35265 6375
rect 35299 6341 35311 6375
rect 36722 6372 36728 6384
rect 36478 6344 36728 6372
rect 35253 6335 35311 6341
rect 36722 6332 36728 6344
rect 36780 6332 36786 6384
rect 31205 6307 31263 6313
rect 31205 6304 31217 6307
rect 29288 6276 31217 6304
rect 28316 6208 28485 6236
rect 28316 6196 28322 6208
rect 28810 6196 28816 6248
rect 28868 6236 28874 6248
rect 29288 6236 29316 6276
rect 31205 6273 31217 6276
rect 31251 6273 31263 6307
rect 31205 6267 31263 6273
rect 32585 6307 32643 6313
rect 32585 6273 32597 6307
rect 32631 6273 32643 6307
rect 32585 6267 32643 6273
rect 32674 6264 32680 6316
rect 32732 6304 32738 6316
rect 32950 6304 32956 6316
rect 32732 6276 32956 6304
rect 32732 6264 32738 6276
rect 32950 6264 32956 6276
rect 33008 6264 33014 6316
rect 33778 6304 33784 6316
rect 33739 6276 33784 6304
rect 33778 6264 33784 6276
rect 33836 6264 33842 6316
rect 37734 6264 37740 6316
rect 37792 6304 37798 6316
rect 38381 6307 38439 6313
rect 38381 6304 38393 6307
rect 37792 6276 38393 6304
rect 37792 6264 37798 6276
rect 38381 6273 38393 6276
rect 38427 6273 38439 6307
rect 38381 6267 38439 6273
rect 39209 6307 39267 6313
rect 39209 6273 39221 6307
rect 39255 6304 39267 6307
rect 39390 6304 39396 6316
rect 39255 6276 39396 6304
rect 39255 6273 39267 6276
rect 39209 6267 39267 6273
rect 39390 6264 39396 6276
rect 39448 6264 39454 6316
rect 31110 6236 31116 6248
rect 28868 6208 29316 6236
rect 31071 6208 31116 6236
rect 28868 6196 28874 6208
rect 31110 6196 31116 6208
rect 31168 6196 31174 6248
rect 11480 6140 11744 6168
rect 11480 6128 11486 6140
rect 12342 6128 12348 6180
rect 12400 6168 12406 6180
rect 14274 6168 14280 6180
rect 12400 6140 14280 6168
rect 12400 6128 12406 6140
rect 14274 6128 14280 6140
rect 14332 6128 14338 6180
rect 26050 6168 26056 6180
rect 24780 6140 26056 6168
rect 3050 6100 3056 6112
rect 2332 6072 3056 6100
rect 3050 6060 3056 6072
rect 3108 6060 3114 6112
rect 5810 6100 5816 6112
rect 5771 6072 5816 6100
rect 5810 6060 5816 6072
rect 5868 6060 5874 6112
rect 7282 6100 7288 6112
rect 7195 6072 7288 6100
rect 7282 6060 7288 6072
rect 7340 6100 7346 6112
rect 9950 6100 9956 6112
rect 7340 6072 9956 6100
rect 7340 6060 7346 6072
rect 9950 6060 9956 6072
rect 10008 6060 10014 6112
rect 10413 6103 10471 6109
rect 10413 6069 10425 6103
rect 10459 6100 10471 6103
rect 11606 6100 11612 6112
rect 10459 6072 11612 6100
rect 10459 6069 10471 6072
rect 10413 6063 10471 6069
rect 11606 6060 11612 6072
rect 11664 6060 11670 6112
rect 12066 6100 12072 6112
rect 12027 6072 12072 6100
rect 12066 6060 12072 6072
rect 12124 6060 12130 6112
rect 13906 6100 13912 6112
rect 13867 6072 13912 6100
rect 13906 6060 13912 6072
rect 13964 6060 13970 6112
rect 13998 6060 14004 6112
rect 14056 6100 14062 6112
rect 14642 6100 14648 6112
rect 14056 6072 14648 6100
rect 14056 6060 14062 6072
rect 14642 6060 14648 6072
rect 14700 6060 14706 6112
rect 15013 6103 15071 6109
rect 15013 6069 15025 6103
rect 15059 6100 15071 6103
rect 15194 6100 15200 6112
rect 15059 6072 15200 6100
rect 15059 6069 15071 6072
rect 15013 6063 15071 6069
rect 15194 6060 15200 6072
rect 15252 6060 15258 6112
rect 16390 6060 16396 6112
rect 16448 6100 16454 6112
rect 18141 6103 18199 6109
rect 18141 6100 18153 6103
rect 16448 6072 18153 6100
rect 16448 6060 16454 6072
rect 18141 6069 18153 6072
rect 18187 6069 18199 6103
rect 20438 6100 20444 6112
rect 20399 6072 20444 6100
rect 18141 6063 18199 6069
rect 20438 6060 20444 6072
rect 20496 6060 20502 6112
rect 20898 6060 20904 6112
rect 20956 6100 20962 6112
rect 24780 6109 24808 6140
rect 26050 6128 26056 6140
rect 26108 6128 26114 6180
rect 32692 6168 32720 6264
rect 33042 6236 33048 6248
rect 33003 6208 33048 6236
rect 33042 6196 33048 6208
rect 33100 6196 33106 6248
rect 33505 6239 33563 6245
rect 33505 6205 33517 6239
rect 33551 6205 33563 6239
rect 33505 6199 33563 6205
rect 30116 6140 32720 6168
rect 20993 6103 21051 6109
rect 20993 6100 21005 6103
rect 20956 6072 21005 6100
rect 20956 6060 20962 6072
rect 20993 6069 21005 6072
rect 21039 6069 21051 6103
rect 20993 6063 21051 6069
rect 24765 6103 24823 6109
rect 24765 6069 24777 6103
rect 24811 6069 24823 6103
rect 24946 6100 24952 6112
rect 24907 6072 24952 6100
rect 24765 6063 24823 6069
rect 24946 6060 24952 6072
rect 25004 6060 25010 6112
rect 27614 6060 27620 6112
rect 27672 6100 27678 6112
rect 28350 6100 28356 6112
rect 27672 6072 28356 6100
rect 27672 6060 27678 6072
rect 28350 6060 28356 6072
rect 28408 6100 28414 6112
rect 30116 6100 30144 6140
rect 28408 6072 30144 6100
rect 28408 6060 28414 6072
rect 33226 6060 33232 6112
rect 33284 6100 33290 6112
rect 33520 6100 33548 6199
rect 34514 6196 34520 6248
rect 34572 6236 34578 6248
rect 34977 6239 35035 6245
rect 34977 6236 34989 6239
rect 34572 6208 34989 6236
rect 34572 6196 34578 6208
rect 34977 6205 34989 6208
rect 35023 6205 35035 6239
rect 34977 6199 35035 6205
rect 36262 6196 36268 6248
rect 36320 6236 36326 6248
rect 38105 6239 38163 6245
rect 38105 6236 38117 6239
rect 36320 6208 38117 6236
rect 36320 6196 36326 6208
rect 38105 6205 38117 6208
rect 38151 6205 38163 6239
rect 38105 6199 38163 6205
rect 36262 6100 36268 6112
rect 33284 6072 36268 6100
rect 33284 6060 33290 6072
rect 36262 6060 36268 6072
rect 36320 6060 36326 6112
rect 36722 6100 36728 6112
rect 36683 6072 36728 6100
rect 36722 6060 36728 6072
rect 36780 6060 36786 6112
rect 1104 6010 68816 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 65654 6010
rect 65706 5958 65718 6010
rect 65770 5958 65782 6010
rect 65834 5958 65846 6010
rect 65898 5958 65910 6010
rect 65962 5958 68816 6010
rect 1104 5936 68816 5958
rect 2774 5896 2780 5908
rect 1872 5868 2780 5896
rect 1872 5769 1900 5868
rect 2774 5856 2780 5868
rect 2832 5856 2838 5908
rect 3234 5896 3240 5908
rect 3147 5868 3240 5896
rect 3234 5856 3240 5868
rect 3292 5896 3298 5908
rect 9030 5896 9036 5908
rect 3292 5868 8892 5896
rect 8991 5868 9036 5896
rect 3292 5856 3298 5868
rect 5810 5788 5816 5840
rect 5868 5828 5874 5840
rect 8110 5828 8116 5840
rect 5868 5800 8116 5828
rect 5868 5788 5874 5800
rect 8110 5788 8116 5800
rect 8168 5788 8174 5840
rect 8864 5828 8892 5868
rect 9030 5856 9036 5868
rect 9088 5856 9094 5908
rect 9677 5899 9735 5905
rect 9677 5865 9689 5899
rect 9723 5896 9735 5899
rect 12618 5896 12624 5908
rect 9723 5868 12624 5896
rect 9723 5865 9735 5868
rect 9677 5859 9735 5865
rect 12618 5856 12624 5868
rect 12676 5856 12682 5908
rect 16117 5899 16175 5905
rect 16117 5865 16129 5899
rect 16163 5896 16175 5899
rect 16298 5896 16304 5908
rect 16163 5868 16304 5896
rect 16163 5865 16175 5868
rect 16117 5859 16175 5865
rect 16298 5856 16304 5868
rect 16356 5856 16362 5908
rect 18874 5856 18880 5908
rect 18932 5896 18938 5908
rect 19705 5899 19763 5905
rect 19705 5896 19717 5899
rect 18932 5868 19717 5896
rect 18932 5856 18938 5868
rect 19705 5865 19717 5868
rect 19751 5865 19763 5899
rect 19705 5859 19763 5865
rect 24946 5856 24952 5908
rect 25004 5896 25010 5908
rect 28445 5899 28503 5905
rect 25004 5868 28396 5896
rect 25004 5856 25010 5868
rect 24673 5831 24731 5837
rect 8864 5800 11928 5828
rect 1857 5763 1915 5769
rect 1857 5729 1869 5763
rect 1903 5729 1915 5763
rect 6730 5760 6736 5772
rect 1857 5723 1915 5729
rect 5736 5732 6736 5760
rect 4893 5695 4951 5701
rect 4893 5661 4905 5695
rect 4939 5692 4951 5695
rect 5626 5692 5632 5704
rect 4939 5664 5632 5692
rect 4939 5661 4951 5664
rect 4893 5655 4951 5661
rect 5626 5652 5632 5664
rect 5684 5652 5690 5704
rect 5736 5701 5764 5732
rect 6730 5720 6736 5732
rect 6788 5760 6794 5772
rect 6788 5732 8156 5760
rect 6788 5720 6794 5732
rect 5721 5695 5779 5701
rect 5721 5661 5733 5695
rect 5767 5661 5779 5695
rect 5721 5655 5779 5661
rect 5810 5652 5816 5704
rect 5868 5692 5874 5704
rect 5997 5695 6055 5701
rect 5868 5664 5913 5692
rect 5868 5652 5874 5664
rect 5997 5661 6009 5695
rect 6043 5692 6055 5695
rect 6270 5692 6276 5704
rect 6043 5664 6276 5692
rect 6043 5661 6055 5664
rect 5997 5655 6055 5661
rect 6270 5652 6276 5664
rect 6328 5652 6334 5704
rect 6457 5695 6515 5701
rect 6457 5661 6469 5695
rect 6503 5692 6515 5695
rect 6546 5692 6552 5704
rect 6503 5664 6552 5692
rect 6503 5661 6515 5664
rect 6457 5655 6515 5661
rect 6546 5652 6552 5664
rect 6604 5692 6610 5704
rect 6822 5692 6828 5704
rect 6604 5664 6828 5692
rect 6604 5652 6610 5664
rect 6822 5652 6828 5664
rect 6880 5652 6886 5704
rect 7926 5652 7932 5704
rect 7984 5692 7990 5704
rect 8128 5701 8156 5732
rect 8021 5695 8079 5701
rect 8021 5692 8033 5695
rect 7984 5664 8033 5692
rect 7984 5652 7990 5664
rect 8021 5661 8033 5664
rect 8067 5661 8079 5695
rect 8021 5655 8079 5661
rect 8113 5695 8171 5701
rect 8113 5661 8125 5695
rect 8159 5661 8171 5695
rect 8113 5655 8171 5661
rect 8202 5652 8208 5704
rect 8260 5692 8266 5704
rect 8389 5695 8447 5701
rect 8260 5664 8305 5692
rect 8260 5652 8266 5664
rect 8389 5661 8401 5695
rect 8435 5661 8447 5695
rect 10410 5692 10416 5704
rect 10371 5664 10416 5692
rect 8389 5655 8447 5661
rect 1854 5584 1860 5636
rect 1912 5624 1918 5636
rect 2102 5627 2160 5633
rect 2102 5624 2114 5627
rect 1912 5596 2114 5624
rect 1912 5584 1918 5596
rect 2102 5593 2114 5596
rect 2148 5593 2160 5627
rect 6288 5624 6316 5652
rect 8404 5624 8432 5655
rect 10410 5652 10416 5664
rect 10468 5652 10474 5704
rect 11149 5695 11207 5701
rect 11149 5661 11161 5695
rect 11195 5661 11207 5695
rect 11790 5692 11796 5704
rect 11751 5664 11796 5692
rect 11149 5655 11207 5661
rect 6288 5596 8432 5624
rect 11164 5624 11192 5655
rect 11790 5652 11796 5664
rect 11848 5652 11854 5704
rect 11900 5701 11928 5800
rect 24673 5797 24685 5831
rect 24719 5828 24731 5831
rect 25130 5828 25136 5840
rect 24719 5800 25136 5828
rect 24719 5797 24731 5800
rect 24673 5791 24731 5797
rect 25130 5788 25136 5800
rect 25188 5788 25194 5840
rect 27614 5828 27620 5840
rect 27575 5800 27620 5828
rect 27614 5788 27620 5800
rect 27672 5788 27678 5840
rect 12434 5760 12440 5772
rect 12084 5732 12440 5760
rect 12084 5701 12112 5732
rect 12434 5720 12440 5732
rect 12492 5760 12498 5772
rect 14829 5763 14887 5769
rect 12492 5732 13124 5760
rect 12492 5720 12498 5732
rect 11885 5695 11943 5701
rect 11885 5661 11897 5695
rect 11931 5661 11943 5695
rect 11885 5655 11943 5661
rect 12069 5695 12127 5701
rect 12069 5661 12081 5695
rect 12115 5661 12127 5695
rect 12069 5655 12127 5661
rect 12158 5652 12164 5704
rect 12216 5692 12222 5704
rect 13096 5701 13124 5732
rect 14829 5729 14841 5763
rect 14875 5760 14887 5763
rect 15102 5760 15108 5772
rect 14875 5732 15108 5760
rect 14875 5729 14887 5732
rect 14829 5723 14887 5729
rect 15102 5720 15108 5732
rect 15160 5760 15166 5772
rect 20346 5760 20352 5772
rect 15160 5732 16620 5760
rect 15160 5720 15166 5732
rect 12805 5695 12863 5701
rect 12805 5692 12817 5695
rect 12216 5664 12817 5692
rect 12216 5652 12222 5664
rect 12805 5661 12817 5664
rect 12851 5661 12863 5695
rect 12805 5655 12863 5661
rect 13081 5695 13139 5701
rect 13081 5661 13093 5695
rect 13127 5692 13139 5695
rect 14182 5692 14188 5704
rect 13127 5664 14188 5692
rect 13127 5661 13139 5664
rect 13081 5655 13139 5661
rect 14182 5652 14188 5664
rect 14240 5652 14246 5704
rect 14274 5652 14280 5704
rect 14332 5692 14338 5704
rect 14553 5695 14611 5701
rect 14553 5692 14565 5695
rect 14332 5664 14565 5692
rect 14332 5652 14338 5664
rect 14553 5661 14565 5664
rect 14599 5661 14611 5695
rect 14553 5655 14611 5661
rect 16301 5695 16359 5701
rect 16301 5661 16313 5695
rect 16347 5692 16359 5695
rect 16390 5692 16396 5704
rect 16347 5664 16396 5692
rect 16347 5661 16359 5664
rect 16301 5655 16359 5661
rect 12342 5624 12348 5636
rect 11164 5596 12348 5624
rect 2102 5587 2160 5593
rect 12342 5584 12348 5596
rect 12400 5584 12406 5636
rect 5350 5556 5356 5568
rect 5311 5528 5356 5556
rect 5350 5516 5356 5528
rect 5408 5516 5414 5568
rect 7742 5556 7748 5568
rect 7703 5528 7748 5556
rect 7742 5516 7748 5528
rect 7800 5516 7806 5568
rect 10229 5559 10287 5565
rect 10229 5525 10241 5559
rect 10275 5556 10287 5559
rect 10778 5556 10784 5568
rect 10275 5528 10784 5556
rect 10275 5525 10287 5528
rect 10229 5519 10287 5525
rect 10778 5516 10784 5528
rect 10836 5516 10842 5568
rect 10965 5559 11023 5565
rect 10965 5525 10977 5559
rect 11011 5556 11023 5559
rect 11514 5556 11520 5568
rect 11011 5528 11520 5556
rect 11011 5525 11023 5528
rect 10965 5519 11023 5525
rect 11514 5516 11520 5528
rect 11572 5516 11578 5568
rect 11609 5559 11667 5565
rect 11609 5525 11621 5559
rect 11655 5556 11667 5559
rect 11974 5556 11980 5568
rect 11655 5528 11980 5556
rect 11655 5525 11667 5528
rect 11609 5519 11667 5525
rect 11974 5516 11980 5528
rect 12032 5516 12038 5568
rect 12526 5516 12532 5568
rect 12584 5556 12590 5568
rect 12897 5559 12955 5565
rect 12897 5556 12909 5559
rect 12584 5528 12909 5556
rect 12584 5516 12590 5528
rect 12897 5525 12909 5528
rect 12943 5525 12955 5559
rect 14568 5556 14596 5655
rect 16390 5652 16396 5664
rect 16448 5652 16454 5704
rect 16592 5701 16620 5732
rect 19536 5732 20352 5760
rect 16577 5695 16635 5701
rect 16577 5661 16589 5695
rect 16623 5692 16635 5695
rect 17126 5692 17132 5704
rect 16623 5664 17132 5692
rect 16623 5661 16635 5664
rect 16577 5655 16635 5661
rect 17126 5652 17132 5664
rect 17184 5652 17190 5704
rect 17313 5695 17371 5701
rect 17313 5661 17325 5695
rect 17359 5692 17371 5695
rect 17494 5692 17500 5704
rect 17359 5664 17500 5692
rect 17359 5661 17371 5664
rect 17313 5655 17371 5661
rect 17494 5652 17500 5664
rect 17552 5652 17558 5704
rect 17770 5692 17776 5704
rect 17731 5664 17776 5692
rect 17770 5652 17776 5664
rect 17828 5652 17834 5704
rect 18322 5652 18328 5704
rect 18380 5692 18386 5704
rect 18417 5695 18475 5701
rect 18417 5692 18429 5695
rect 18380 5664 18429 5692
rect 18380 5652 18386 5664
rect 18417 5661 18429 5664
rect 18463 5661 18475 5695
rect 19242 5692 19248 5704
rect 19155 5664 19248 5692
rect 18417 5655 18475 5661
rect 19242 5652 19248 5664
rect 19300 5652 19306 5704
rect 19337 5695 19395 5701
rect 19337 5661 19349 5695
rect 19383 5692 19395 5695
rect 19426 5692 19432 5704
rect 19383 5664 19432 5692
rect 19383 5661 19395 5664
rect 19337 5655 19395 5661
rect 19426 5652 19432 5664
rect 19484 5652 19490 5704
rect 19536 5701 19564 5732
rect 20346 5720 20352 5732
rect 20404 5720 20410 5772
rect 20714 5720 20720 5772
rect 20772 5760 20778 5772
rect 20809 5763 20867 5769
rect 20809 5760 20821 5763
rect 20772 5732 20821 5760
rect 20772 5720 20778 5732
rect 20809 5729 20821 5732
rect 20855 5729 20867 5763
rect 20809 5723 20867 5729
rect 22646 5720 22652 5772
rect 22704 5760 22710 5772
rect 26234 5760 26240 5772
rect 22704 5732 26240 5760
rect 22704 5720 22710 5732
rect 26234 5720 26240 5732
rect 26292 5720 26298 5772
rect 19521 5695 19579 5701
rect 19521 5661 19533 5695
rect 19567 5661 19579 5695
rect 19521 5655 19579 5661
rect 19978 5652 19984 5704
rect 20036 5692 20042 5704
rect 20165 5695 20223 5701
rect 20165 5692 20177 5695
rect 20036 5664 20177 5692
rect 20036 5652 20042 5664
rect 20165 5661 20177 5664
rect 20211 5661 20223 5695
rect 20438 5692 20444 5704
rect 20399 5664 20444 5692
rect 20165 5655 20223 5661
rect 20438 5652 20444 5664
rect 20496 5652 20502 5704
rect 20625 5695 20683 5701
rect 20625 5661 20637 5695
rect 20671 5692 20683 5695
rect 24489 5695 24547 5701
rect 20671 5664 20760 5692
rect 20671 5661 20683 5664
rect 20625 5655 20683 5661
rect 14734 5584 14740 5636
rect 14792 5624 14798 5636
rect 16485 5627 16543 5633
rect 16485 5624 16497 5627
rect 14792 5596 16497 5624
rect 14792 5584 14798 5596
rect 16485 5593 16497 5596
rect 16531 5593 16543 5627
rect 16485 5587 16543 5593
rect 19260 5556 19288 5652
rect 20732 5636 20760 5664
rect 24489 5661 24501 5695
rect 24535 5692 24547 5695
rect 24578 5692 24584 5704
rect 24535 5664 24584 5692
rect 24535 5661 24547 5664
rect 24489 5655 24547 5661
rect 24578 5652 24584 5664
rect 24636 5652 24642 5704
rect 25130 5652 25136 5704
rect 25188 5692 25194 5704
rect 25409 5695 25467 5701
rect 25409 5692 25421 5695
rect 25188 5664 25421 5692
rect 25188 5652 25194 5664
rect 25409 5661 25421 5664
rect 25455 5661 25467 5695
rect 25409 5655 25467 5661
rect 25593 5695 25651 5701
rect 25593 5661 25605 5695
rect 25639 5692 25651 5695
rect 27632 5692 27660 5788
rect 28368 5760 28396 5868
rect 28445 5865 28457 5899
rect 28491 5896 28503 5899
rect 28534 5896 28540 5908
rect 28491 5868 28540 5896
rect 28491 5865 28503 5868
rect 28445 5859 28503 5865
rect 28534 5856 28540 5868
rect 28592 5856 28598 5908
rect 31941 5899 31999 5905
rect 31941 5865 31953 5899
rect 31987 5865 31999 5899
rect 31941 5859 31999 5865
rect 32585 5899 32643 5905
rect 32585 5865 32597 5899
rect 32631 5896 32643 5899
rect 33042 5896 33048 5908
rect 32631 5868 33048 5896
rect 32631 5865 32643 5868
rect 32585 5859 32643 5865
rect 31956 5828 31984 5859
rect 33042 5856 33048 5868
rect 33100 5856 33106 5908
rect 36262 5896 36268 5908
rect 36223 5868 36268 5896
rect 36262 5856 36268 5868
rect 36320 5856 36326 5908
rect 37734 5896 37740 5908
rect 37695 5868 37740 5896
rect 37734 5856 37740 5868
rect 37792 5856 37798 5908
rect 31956 5800 32720 5828
rect 31849 5763 31907 5769
rect 31849 5760 31861 5763
rect 28368 5732 31861 5760
rect 31849 5729 31861 5732
rect 31895 5760 31907 5763
rect 32214 5760 32220 5772
rect 31895 5732 32220 5760
rect 31895 5729 31907 5732
rect 31849 5723 31907 5729
rect 32214 5720 32220 5732
rect 32272 5720 32278 5772
rect 32692 5760 32720 5800
rect 32766 5788 32772 5840
rect 32824 5828 32830 5840
rect 32824 5800 33916 5828
rect 32824 5788 32830 5800
rect 33045 5763 33103 5769
rect 32692 5732 32904 5760
rect 32876 5704 32904 5732
rect 33045 5729 33057 5763
rect 33091 5760 33103 5763
rect 33686 5760 33692 5772
rect 33091 5732 33692 5760
rect 33091 5729 33103 5732
rect 33045 5723 33103 5729
rect 33686 5720 33692 5732
rect 33744 5720 33750 5772
rect 33888 5760 33916 5800
rect 33888 5732 34008 5760
rect 28074 5692 28080 5704
rect 25639 5664 27660 5692
rect 28035 5664 28080 5692
rect 25639 5661 25651 5664
rect 25593 5655 25651 5661
rect 28074 5652 28080 5664
rect 28132 5652 28138 5704
rect 28261 5695 28319 5701
rect 28261 5661 28273 5695
rect 28307 5692 28319 5695
rect 30650 5692 30656 5704
rect 28307 5664 30656 5692
rect 28307 5661 28319 5664
rect 28261 5655 28319 5661
rect 30650 5652 30656 5664
rect 30708 5652 30714 5704
rect 31662 5692 31668 5704
rect 31623 5664 31668 5692
rect 31662 5652 31668 5664
rect 31720 5652 31726 5704
rect 31941 5695 31999 5701
rect 31941 5661 31953 5695
rect 31987 5692 31999 5695
rect 32582 5692 32588 5704
rect 31987 5664 32588 5692
rect 31987 5661 31999 5664
rect 31941 5655 31999 5661
rect 32582 5652 32588 5664
rect 32640 5692 32646 5704
rect 32769 5695 32827 5701
rect 32769 5692 32781 5695
rect 32640 5664 32781 5692
rect 32640 5652 32646 5664
rect 32769 5661 32781 5664
rect 32815 5661 32827 5695
rect 32769 5655 32827 5661
rect 32858 5652 32864 5704
rect 32916 5692 32922 5704
rect 33134 5692 33140 5704
rect 32916 5664 33009 5692
rect 33095 5664 33140 5692
rect 32916 5652 32922 5664
rect 33134 5652 33140 5664
rect 33192 5652 33198 5704
rect 33980 5701 34008 5732
rect 33873 5695 33931 5701
rect 33873 5661 33885 5695
rect 33919 5661 33931 5695
rect 33873 5655 33931 5661
rect 33965 5695 34023 5701
rect 33965 5661 33977 5695
rect 34011 5661 34023 5695
rect 33965 5655 34023 5661
rect 20714 5584 20720 5636
rect 20772 5584 20778 5636
rect 26510 5633 26516 5636
rect 26504 5587 26516 5633
rect 26568 5624 26574 5636
rect 33888 5624 33916 5655
rect 34054 5652 34060 5704
rect 34112 5692 34118 5704
rect 36262 5692 36268 5704
rect 34112 5664 36268 5692
rect 34112 5652 34118 5664
rect 36262 5652 36268 5664
rect 36320 5652 36326 5704
rect 36446 5692 36452 5704
rect 36407 5664 36452 5692
rect 36446 5652 36452 5664
rect 36504 5652 36510 5704
rect 37553 5695 37611 5701
rect 37553 5661 37565 5695
rect 37599 5661 37611 5695
rect 68094 5692 68100 5704
rect 68055 5664 68100 5692
rect 37553 5655 37611 5661
rect 36170 5624 36176 5636
rect 26568 5596 26604 5624
rect 33888 5596 36176 5624
rect 26510 5584 26516 5587
rect 26568 5584 26574 5596
rect 36170 5584 36176 5596
rect 36228 5624 36234 5636
rect 37568 5624 37596 5655
rect 68094 5652 68100 5664
rect 68152 5652 68158 5704
rect 36228 5596 37596 5624
rect 36228 5584 36234 5596
rect 14568 5528 19288 5556
rect 12897 5519 12955 5525
rect 20438 5516 20444 5568
rect 20496 5556 20502 5568
rect 21269 5559 21327 5565
rect 21269 5556 21281 5559
rect 20496 5528 21281 5556
rect 20496 5516 20502 5528
rect 21269 5525 21281 5528
rect 21315 5525 21327 5559
rect 21269 5519 21327 5525
rect 25777 5559 25835 5565
rect 25777 5525 25789 5559
rect 25823 5556 25835 5559
rect 25958 5556 25964 5568
rect 25823 5528 25964 5556
rect 25823 5525 25835 5528
rect 25777 5519 25835 5525
rect 25958 5516 25964 5528
rect 26016 5516 26022 5568
rect 32125 5559 32183 5565
rect 32125 5525 32137 5559
rect 32171 5556 32183 5559
rect 32766 5556 32772 5568
rect 32171 5528 32772 5556
rect 32171 5525 32183 5528
rect 32125 5519 32183 5525
rect 32766 5516 32772 5528
rect 32824 5516 32830 5568
rect 32858 5516 32864 5568
rect 32916 5556 32922 5568
rect 34054 5556 34060 5568
rect 32916 5528 34060 5556
rect 32916 5516 32922 5528
rect 34054 5516 34060 5528
rect 34112 5516 34118 5568
rect 34149 5559 34207 5565
rect 34149 5525 34161 5559
rect 34195 5556 34207 5559
rect 34698 5556 34704 5568
rect 34195 5528 34704 5556
rect 34195 5525 34207 5528
rect 34149 5519 34207 5525
rect 34698 5516 34704 5528
rect 34756 5516 34762 5568
rect 1104 5466 68816 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 50294 5466
rect 50346 5414 50358 5466
rect 50410 5414 50422 5466
rect 50474 5414 50486 5466
rect 50538 5414 50550 5466
rect 50602 5414 68816 5466
rect 1104 5392 68816 5414
rect 1854 5352 1860 5364
rect 1815 5324 1860 5352
rect 1854 5312 1860 5324
rect 1912 5312 1918 5364
rect 3510 5352 3516 5364
rect 3471 5324 3516 5352
rect 3510 5312 3516 5324
rect 3568 5312 3574 5364
rect 5810 5312 5816 5364
rect 5868 5352 5874 5364
rect 6365 5355 6423 5361
rect 6365 5352 6377 5355
rect 5868 5324 6377 5352
rect 5868 5312 5874 5324
rect 6365 5321 6377 5324
rect 6411 5321 6423 5355
rect 6365 5315 6423 5321
rect 7653 5355 7711 5361
rect 7653 5321 7665 5355
rect 7699 5352 7711 5355
rect 8202 5352 8208 5364
rect 7699 5324 8208 5352
rect 7699 5321 7711 5324
rect 7653 5315 7711 5321
rect 8202 5312 8208 5324
rect 8260 5312 8266 5364
rect 9674 5352 9680 5364
rect 8312 5324 9680 5352
rect 3234 5284 3240 5296
rect 2148 5256 3240 5284
rect 2148 5225 2176 5256
rect 3234 5244 3240 5256
rect 3292 5244 3298 5296
rect 2133 5219 2191 5225
rect 2133 5185 2145 5219
rect 2179 5185 2191 5219
rect 2133 5179 2191 5185
rect 2225 5219 2283 5225
rect 2225 5185 2237 5219
rect 2271 5185 2283 5219
rect 2225 5179 2283 5185
rect 2038 5108 2044 5160
rect 2096 5148 2102 5160
rect 2240 5148 2268 5179
rect 2314 5176 2320 5228
rect 2372 5216 2378 5228
rect 2372 5188 2417 5216
rect 2372 5176 2378 5188
rect 2498 5176 2504 5228
rect 2556 5216 2562 5228
rect 3528 5216 3556 5312
rect 4332 5287 4390 5293
rect 4332 5253 4344 5287
rect 4378 5284 4390 5287
rect 5350 5284 5356 5296
rect 4378 5256 5356 5284
rect 4378 5253 4390 5256
rect 4332 5247 4390 5253
rect 5350 5244 5356 5256
rect 5408 5244 5414 5296
rect 6454 5244 6460 5296
rect 6512 5284 6518 5296
rect 6733 5287 6791 5293
rect 6733 5284 6745 5287
rect 6512 5256 6745 5284
rect 6512 5244 6518 5256
rect 6733 5253 6745 5256
rect 6779 5284 6791 5287
rect 7285 5287 7343 5293
rect 7285 5284 7297 5287
rect 6779 5256 7297 5284
rect 6779 5253 6791 5256
rect 6733 5247 6791 5253
rect 7285 5253 7297 5256
rect 7331 5253 7343 5287
rect 8312 5284 8340 5324
rect 9674 5312 9680 5324
rect 9732 5312 9738 5364
rect 9766 5312 9772 5364
rect 9824 5352 9830 5364
rect 10962 5352 10968 5364
rect 9824 5324 10968 5352
rect 9824 5312 9830 5324
rect 10962 5312 10968 5324
rect 11020 5312 11026 5364
rect 11606 5312 11612 5364
rect 11664 5352 11670 5364
rect 13262 5352 13268 5364
rect 11664 5324 13268 5352
rect 11664 5312 11670 5324
rect 13262 5312 13268 5324
rect 13320 5312 13326 5364
rect 14185 5355 14243 5361
rect 14185 5321 14197 5355
rect 14231 5352 14243 5355
rect 14366 5352 14372 5364
rect 14231 5324 14372 5352
rect 14231 5321 14243 5324
rect 14185 5315 14243 5321
rect 14366 5312 14372 5324
rect 14424 5312 14430 5364
rect 14553 5355 14611 5361
rect 14553 5321 14565 5355
rect 14599 5352 14611 5355
rect 14734 5352 14740 5364
rect 14599 5324 14740 5352
rect 14599 5321 14611 5324
rect 14553 5315 14611 5321
rect 14734 5312 14740 5324
rect 14792 5352 14798 5364
rect 15197 5355 15255 5361
rect 15197 5352 15209 5355
rect 14792 5324 15209 5352
rect 14792 5312 14798 5324
rect 15197 5321 15209 5324
rect 15243 5321 15255 5355
rect 15197 5315 15255 5321
rect 15470 5312 15476 5364
rect 15528 5352 15534 5364
rect 15565 5355 15623 5361
rect 15565 5352 15577 5355
rect 15528 5324 15577 5352
rect 15528 5312 15534 5324
rect 15565 5321 15577 5324
rect 15611 5321 15623 5355
rect 15565 5315 15623 5321
rect 17497 5355 17555 5361
rect 17497 5321 17509 5355
rect 17543 5352 17555 5355
rect 19334 5352 19340 5364
rect 17543 5324 19340 5352
rect 17543 5321 17555 5324
rect 17497 5315 17555 5321
rect 19334 5312 19340 5324
rect 19392 5312 19398 5364
rect 19797 5355 19855 5361
rect 19797 5321 19809 5355
rect 19843 5352 19855 5355
rect 20254 5352 20260 5364
rect 19843 5324 20260 5352
rect 19843 5321 19855 5324
rect 19797 5315 19855 5321
rect 20254 5312 20260 5324
rect 20312 5312 20318 5364
rect 20806 5352 20812 5364
rect 20767 5324 20812 5352
rect 20806 5312 20812 5324
rect 20864 5312 20870 5364
rect 22189 5355 22247 5361
rect 22189 5321 22201 5355
rect 22235 5352 22247 5355
rect 22830 5352 22836 5364
rect 22235 5324 22836 5352
rect 22235 5321 22247 5324
rect 22189 5315 22247 5321
rect 22830 5312 22836 5324
rect 22888 5312 22894 5364
rect 24029 5355 24087 5361
rect 24029 5321 24041 5355
rect 24075 5352 24087 5355
rect 24210 5352 24216 5364
rect 24075 5324 24216 5352
rect 24075 5321 24087 5324
rect 24029 5315 24087 5321
rect 24210 5312 24216 5324
rect 24268 5312 24274 5364
rect 26421 5355 26479 5361
rect 26421 5321 26433 5355
rect 26467 5352 26479 5355
rect 26510 5352 26516 5364
rect 26467 5324 26516 5352
rect 26467 5321 26479 5324
rect 26421 5315 26479 5321
rect 26510 5312 26516 5324
rect 26568 5312 26574 5364
rect 31021 5355 31079 5361
rect 31021 5321 31033 5355
rect 31067 5352 31079 5355
rect 31110 5352 31116 5364
rect 31067 5324 31116 5352
rect 31067 5321 31079 5324
rect 31021 5315 31079 5321
rect 31110 5312 31116 5324
rect 31168 5312 31174 5364
rect 34790 5312 34796 5364
rect 34848 5352 34854 5364
rect 34885 5355 34943 5361
rect 34885 5352 34897 5355
rect 34848 5324 34897 5352
rect 34848 5312 34854 5324
rect 34885 5321 34897 5324
rect 34931 5321 34943 5355
rect 36170 5352 36176 5364
rect 36131 5324 36176 5352
rect 34885 5315 34943 5321
rect 36170 5312 36176 5324
rect 36228 5312 36234 5364
rect 7285 5247 7343 5253
rect 7392 5256 8340 5284
rect 8389 5287 8447 5293
rect 2556 5188 3556 5216
rect 4065 5219 4123 5225
rect 2556 5176 2562 5188
rect 4065 5185 4077 5219
rect 4111 5185 4123 5219
rect 4065 5179 4123 5185
rect 6549 5219 6607 5225
rect 6549 5185 6561 5219
rect 6595 5216 6607 5219
rect 7392 5216 7420 5256
rect 8389 5253 8401 5287
rect 8435 5284 8447 5287
rect 14274 5284 14280 5296
rect 8435 5256 12434 5284
rect 8435 5253 8447 5256
rect 8389 5247 8447 5253
rect 6595 5188 7420 5216
rect 7469 5219 7527 5225
rect 6595 5185 6607 5188
rect 6549 5179 6607 5185
rect 7469 5185 7481 5219
rect 7515 5185 7527 5219
rect 7469 5179 7527 5185
rect 2406 5148 2412 5160
rect 2096 5120 2412 5148
rect 2096 5108 2102 5120
rect 2406 5108 2412 5120
rect 2464 5108 2470 5160
rect 3418 5108 3424 5160
rect 3476 5148 3482 5160
rect 4080 5148 4108 5179
rect 3476 5120 4108 5148
rect 3476 5108 3482 5120
rect 5445 5083 5503 5089
rect 5445 5049 5457 5083
rect 5491 5080 5503 5083
rect 6564 5080 6592 5179
rect 7484 5148 7512 5179
rect 7834 5176 7840 5228
rect 7892 5216 7898 5228
rect 8297 5219 8355 5225
rect 8297 5216 8309 5219
rect 7892 5188 8309 5216
rect 7892 5176 7898 5188
rect 8297 5185 8309 5188
rect 8343 5185 8355 5219
rect 8478 5216 8484 5228
rect 8439 5188 8484 5216
rect 8297 5179 8355 5185
rect 8478 5176 8484 5188
rect 8536 5176 8542 5228
rect 8941 5219 8999 5225
rect 8941 5185 8953 5219
rect 8987 5185 8999 5219
rect 9122 5216 9128 5228
rect 9083 5188 9128 5216
rect 8941 5179 8999 5185
rect 8386 5148 8392 5160
rect 7484 5120 8392 5148
rect 8386 5108 8392 5120
rect 8444 5108 8450 5160
rect 8956 5148 8984 5179
rect 9122 5176 9128 5188
rect 9180 5176 9186 5228
rect 9852 5219 9910 5225
rect 9852 5185 9864 5219
rect 9898 5216 9910 5219
rect 11517 5219 11575 5225
rect 11517 5216 11529 5219
rect 9898 5188 11529 5216
rect 9898 5185 9910 5188
rect 9852 5179 9910 5185
rect 11517 5185 11529 5188
rect 11563 5185 11575 5219
rect 11698 5216 11704 5228
rect 11659 5188 11704 5216
rect 11517 5179 11575 5185
rect 11698 5176 11704 5188
rect 11756 5176 11762 5228
rect 11974 5216 11980 5228
rect 11935 5188 11980 5216
rect 11974 5176 11980 5188
rect 12032 5176 12038 5228
rect 12069 5219 12127 5225
rect 12069 5185 12081 5219
rect 12115 5216 12127 5219
rect 12158 5216 12164 5228
rect 12115 5188 12164 5216
rect 12115 5185 12127 5188
rect 12069 5179 12127 5185
rect 12158 5176 12164 5188
rect 12216 5176 12222 5228
rect 12250 5176 12256 5228
rect 12308 5216 12314 5228
rect 12406 5216 12434 5256
rect 13280 5256 14280 5284
rect 13280 5225 13308 5256
rect 14274 5244 14280 5256
rect 14332 5244 14338 5296
rect 16758 5284 16764 5296
rect 16719 5256 16764 5284
rect 16758 5244 16764 5256
rect 16816 5244 16822 5296
rect 18506 5284 18512 5296
rect 18064 5256 18512 5284
rect 13173 5219 13231 5225
rect 13173 5216 13185 5219
rect 12308 5188 12353 5216
rect 12406 5188 13185 5216
rect 12308 5176 12314 5188
rect 13173 5185 13185 5188
rect 13219 5185 13231 5219
rect 13173 5179 13231 5185
rect 13265 5219 13323 5225
rect 13265 5185 13277 5219
rect 13311 5185 13323 5219
rect 13446 5216 13452 5228
rect 13407 5188 13452 5216
rect 13265 5179 13323 5185
rect 13446 5176 13452 5188
rect 13504 5176 13510 5228
rect 14366 5216 14372 5228
rect 14327 5188 14372 5216
rect 14366 5176 14372 5188
rect 14424 5176 14430 5228
rect 14645 5219 14703 5225
rect 14645 5185 14657 5219
rect 14691 5216 14703 5219
rect 15102 5216 15108 5228
rect 14691 5188 15108 5216
rect 14691 5185 14703 5188
rect 14645 5179 14703 5185
rect 15102 5176 15108 5188
rect 15160 5176 15166 5228
rect 15381 5219 15439 5225
rect 15381 5185 15393 5219
rect 15427 5185 15439 5219
rect 15381 5179 15439 5185
rect 17221 5219 17279 5225
rect 17221 5185 17233 5219
rect 17267 5216 17279 5219
rect 17586 5216 17592 5228
rect 17267 5188 17592 5216
rect 17267 5185 17279 5188
rect 17221 5179 17279 5185
rect 9582 5148 9588 5160
rect 8956 5120 9260 5148
rect 9543 5120 9588 5148
rect 5491 5052 6592 5080
rect 5491 5049 5503 5052
rect 5445 5043 5503 5049
rect 3050 5012 3056 5024
rect 2963 4984 3056 5012
rect 3050 4972 3056 4984
rect 3108 5012 3114 5024
rect 6454 5012 6460 5024
rect 3108 4984 6460 5012
rect 3108 4972 3114 4984
rect 6454 4972 6460 4984
rect 6512 4972 6518 5024
rect 9122 5012 9128 5024
rect 9083 4984 9128 5012
rect 9122 4972 9128 4984
rect 9180 4972 9186 5024
rect 9232 5012 9260 5120
rect 9582 5108 9588 5120
rect 9640 5108 9646 5160
rect 11885 5151 11943 5157
rect 11885 5117 11897 5151
rect 11931 5117 11943 5151
rect 12526 5148 12532 5160
rect 11885 5111 11943 5117
rect 12176 5120 12532 5148
rect 10965 5083 11023 5089
rect 10965 5049 10977 5083
rect 11011 5080 11023 5083
rect 11698 5080 11704 5092
rect 11011 5052 11704 5080
rect 11011 5049 11023 5052
rect 10965 5043 11023 5049
rect 11698 5040 11704 5052
rect 11756 5040 11762 5092
rect 11900 5080 11928 5111
rect 12176 5080 12204 5120
rect 12526 5108 12532 5120
rect 12584 5108 12590 5160
rect 12710 5108 12716 5160
rect 12768 5148 12774 5160
rect 13078 5148 13084 5160
rect 12768 5120 13084 5148
rect 12768 5108 12774 5120
rect 13078 5108 13084 5120
rect 13136 5148 13142 5160
rect 13357 5151 13415 5157
rect 13357 5148 13369 5151
rect 13136 5120 13369 5148
rect 13136 5108 13142 5120
rect 13357 5117 13369 5120
rect 13403 5117 13415 5151
rect 13357 5111 13415 5117
rect 14090 5108 14096 5160
rect 14148 5148 14154 5160
rect 15396 5148 15424 5179
rect 17586 5176 17592 5188
rect 17644 5176 17650 5228
rect 14148 5120 15424 5148
rect 17313 5151 17371 5157
rect 14148 5108 14154 5120
rect 17313 5117 17325 5151
rect 17359 5148 17371 5151
rect 17402 5148 17408 5160
rect 17359 5120 17408 5148
rect 17359 5117 17371 5120
rect 17313 5111 17371 5117
rect 17402 5108 17408 5120
rect 17460 5108 17466 5160
rect 12989 5083 13047 5089
rect 12989 5080 13001 5083
rect 11900 5052 12204 5080
rect 12406 5052 13001 5080
rect 9858 5012 9864 5024
rect 9232 4984 9864 5012
rect 9858 4972 9864 4984
rect 9916 4972 9922 5024
rect 10502 4972 10508 5024
rect 10560 5012 10566 5024
rect 12406 5012 12434 5052
rect 12989 5049 13001 5052
rect 13035 5049 13047 5083
rect 12989 5043 13047 5049
rect 16574 5040 16580 5092
rect 16632 5080 16638 5092
rect 16761 5083 16819 5089
rect 16761 5080 16773 5083
rect 16632 5052 16773 5080
rect 16632 5040 16638 5052
rect 16761 5049 16773 5052
rect 16807 5049 16819 5083
rect 16761 5043 16819 5049
rect 10560 4984 12434 5012
rect 10560 4972 10566 4984
rect 14274 4972 14280 5024
rect 14332 5012 14338 5024
rect 16025 5015 16083 5021
rect 16025 5012 16037 5015
rect 14332 4984 16037 5012
rect 14332 4972 14338 4984
rect 16025 4981 16037 4984
rect 16071 5012 16083 5015
rect 18064 5012 18092 5256
rect 18506 5244 18512 5256
rect 18564 5284 18570 5296
rect 19061 5287 19119 5293
rect 19061 5284 19073 5287
rect 18564 5256 19073 5284
rect 18564 5244 18570 5256
rect 19061 5253 19073 5256
rect 19107 5284 19119 5287
rect 19702 5284 19708 5296
rect 19107 5256 19708 5284
rect 19107 5253 19119 5256
rect 19061 5247 19119 5253
rect 19702 5244 19708 5256
rect 19760 5284 19766 5296
rect 20438 5284 20444 5296
rect 19760 5256 20444 5284
rect 19760 5244 19766 5256
rect 20438 5244 20444 5256
rect 20496 5284 20502 5296
rect 24762 5284 24768 5296
rect 20496 5256 20576 5284
rect 24723 5256 24768 5284
rect 20496 5244 20502 5256
rect 19978 5176 19984 5228
rect 20036 5216 20042 5228
rect 20548 5225 20576 5256
rect 24762 5244 24768 5256
rect 24820 5244 24826 5296
rect 28074 5244 28080 5296
rect 28132 5284 28138 5296
rect 28534 5284 28540 5296
rect 28132 5256 28540 5284
rect 28132 5244 28138 5256
rect 28534 5244 28540 5256
rect 28592 5244 28598 5296
rect 28721 5287 28779 5293
rect 28721 5253 28733 5287
rect 28767 5284 28779 5287
rect 29638 5284 29644 5296
rect 28767 5256 29644 5284
rect 28767 5253 28779 5256
rect 28721 5247 28779 5253
rect 29638 5244 29644 5256
rect 29696 5284 29702 5296
rect 30282 5284 30288 5296
rect 29696 5256 30288 5284
rect 29696 5244 29702 5256
rect 30282 5244 30288 5256
rect 30340 5284 30346 5296
rect 34808 5284 34836 5312
rect 36722 5284 36728 5296
rect 30340 5256 30696 5284
rect 30340 5244 30346 5256
rect 20257 5219 20315 5225
rect 20257 5216 20269 5219
rect 20036 5188 20269 5216
rect 20036 5176 20042 5188
rect 20257 5185 20269 5188
rect 20303 5185 20315 5219
rect 20257 5179 20315 5185
rect 20533 5219 20591 5225
rect 20533 5185 20545 5219
rect 20579 5185 20591 5219
rect 20533 5179 20591 5185
rect 20809 5219 20867 5225
rect 20809 5185 20821 5219
rect 20855 5185 20867 5219
rect 20809 5179 20867 5185
rect 19426 5108 19432 5160
rect 19484 5148 19490 5160
rect 19521 5151 19579 5157
rect 19521 5148 19533 5151
rect 19484 5120 19533 5148
rect 19484 5108 19490 5120
rect 19521 5117 19533 5120
rect 19567 5117 19579 5151
rect 19521 5111 19579 5117
rect 19613 5151 19671 5157
rect 19613 5117 19625 5151
rect 19659 5148 19671 5151
rect 20824 5148 20852 5179
rect 22094 5176 22100 5228
rect 22152 5216 22158 5228
rect 22646 5216 22652 5228
rect 22152 5188 22652 5216
rect 22152 5176 22158 5188
rect 22646 5176 22652 5188
rect 22704 5176 22710 5228
rect 22922 5225 22928 5228
rect 22916 5179 22928 5225
rect 22980 5216 22986 5228
rect 24581 5219 24639 5225
rect 22980 5188 23016 5216
rect 22922 5176 22928 5179
rect 22980 5176 22986 5188
rect 24581 5185 24593 5219
rect 24627 5216 24639 5219
rect 25130 5216 25136 5228
rect 24627 5188 25136 5216
rect 24627 5185 24639 5188
rect 24581 5179 24639 5185
rect 25130 5176 25136 5188
rect 25188 5176 25194 5228
rect 25682 5176 25688 5228
rect 25740 5216 25746 5228
rect 25777 5219 25835 5225
rect 25777 5216 25789 5219
rect 25740 5188 25789 5216
rect 25740 5176 25746 5188
rect 25777 5185 25789 5188
rect 25823 5185 25835 5219
rect 25958 5216 25964 5228
rect 25919 5188 25964 5216
rect 25777 5179 25835 5185
rect 25958 5176 25964 5188
rect 26016 5176 26022 5228
rect 26053 5219 26111 5225
rect 26053 5185 26065 5219
rect 26099 5185 26111 5219
rect 26053 5179 26111 5185
rect 21082 5148 21088 5160
rect 19659 5120 21088 5148
rect 19659 5117 19671 5120
rect 19613 5111 19671 5117
rect 18138 5040 18144 5092
rect 18196 5080 18202 5092
rect 19061 5083 19119 5089
rect 19061 5080 19073 5083
rect 18196 5052 19073 5080
rect 18196 5040 18202 5052
rect 19061 5049 19073 5052
rect 19107 5049 19119 5083
rect 19061 5043 19119 5049
rect 16071 4984 18092 5012
rect 18509 5015 18567 5021
rect 16071 4981 16083 4984
rect 16025 4975 16083 4981
rect 18509 4981 18521 5015
rect 18555 5012 18567 5015
rect 18874 5012 18880 5024
rect 18555 4984 18880 5012
rect 18555 4981 18567 4984
rect 18509 4975 18567 4981
rect 18874 4972 18880 4984
rect 18932 4972 18938 5024
rect 19076 5012 19104 5043
rect 19334 5040 19340 5092
rect 19392 5080 19398 5092
rect 19628 5080 19656 5111
rect 21082 5108 21088 5120
rect 21140 5108 21146 5160
rect 26068 5148 26096 5179
rect 26142 5176 26148 5228
rect 26200 5216 26206 5228
rect 26973 5219 27031 5225
rect 26973 5216 26985 5219
rect 26200 5188 26985 5216
rect 26200 5176 26206 5188
rect 26973 5185 26985 5188
rect 27019 5216 27031 5219
rect 27798 5216 27804 5228
rect 27019 5188 27804 5216
rect 27019 5185 27031 5188
rect 26973 5179 27031 5185
rect 27798 5176 27804 5188
rect 27856 5176 27862 5228
rect 30668 5225 30696 5256
rect 33520 5256 34836 5284
rect 36188 5256 36728 5284
rect 30653 5219 30711 5225
rect 30653 5185 30665 5219
rect 30699 5185 30711 5219
rect 33226 5216 33232 5228
rect 33187 5188 33232 5216
rect 30653 5179 30711 5185
rect 33226 5176 33232 5188
rect 33284 5176 33290 5228
rect 33520 5225 33548 5256
rect 36188 5228 36216 5256
rect 36722 5244 36728 5256
rect 36780 5244 36786 5296
rect 33505 5219 33563 5225
rect 33505 5185 33517 5219
rect 33551 5185 33563 5219
rect 34698 5216 34704 5228
rect 34659 5188 34704 5216
rect 33505 5179 33563 5185
rect 34698 5176 34704 5188
rect 34756 5176 34762 5228
rect 36170 5225 36176 5228
rect 36165 5216 36176 5225
rect 36131 5188 36176 5216
rect 36165 5179 36176 5188
rect 36170 5176 36176 5179
rect 36228 5176 36234 5228
rect 36262 5176 36268 5228
rect 36320 5216 36326 5228
rect 36357 5219 36415 5225
rect 36357 5216 36369 5219
rect 36320 5188 36369 5216
rect 36320 5176 36326 5188
rect 36357 5185 36369 5188
rect 36403 5185 36415 5219
rect 36357 5179 36415 5185
rect 25792 5120 26096 5148
rect 25792 5092 25820 5120
rect 26326 5108 26332 5160
rect 26384 5148 26390 5160
rect 29365 5151 29423 5157
rect 29365 5148 29377 5151
rect 26384 5120 29377 5148
rect 26384 5108 26390 5120
rect 29365 5117 29377 5120
rect 29411 5148 29423 5151
rect 29914 5148 29920 5160
rect 29411 5120 29920 5148
rect 29411 5117 29423 5120
rect 29365 5111 29423 5117
rect 29914 5108 29920 5120
rect 29972 5108 29978 5160
rect 30558 5148 30564 5160
rect 30519 5120 30564 5148
rect 30558 5108 30564 5120
rect 30616 5108 30622 5160
rect 58802 5108 58808 5160
rect 58860 5148 58866 5160
rect 59449 5151 59507 5157
rect 59449 5148 59461 5151
rect 58860 5120 59461 5148
rect 58860 5108 58866 5120
rect 59449 5117 59461 5120
rect 59495 5117 59507 5151
rect 59449 5111 59507 5117
rect 19392 5052 19656 5080
rect 19392 5040 19398 5052
rect 20806 5040 20812 5092
rect 20864 5080 20870 5092
rect 21269 5083 21327 5089
rect 21269 5080 21281 5083
rect 20864 5052 21281 5080
rect 20864 5040 20870 5052
rect 21269 5049 21281 5052
rect 21315 5049 21327 5083
rect 21269 5043 21327 5049
rect 25774 5040 25780 5092
rect 25832 5040 25838 5092
rect 59262 5040 59268 5092
rect 59320 5080 59326 5092
rect 60093 5083 60151 5089
rect 60093 5080 60105 5083
rect 59320 5052 60105 5080
rect 59320 5040 59326 5052
rect 60093 5049 60105 5052
rect 60139 5049 60151 5083
rect 60093 5043 60151 5049
rect 19978 5012 19984 5024
rect 19076 4984 19984 5012
rect 19978 4972 19984 4984
rect 20036 4972 20042 5024
rect 24854 4972 24860 5024
rect 24912 5012 24918 5024
rect 24949 5015 25007 5021
rect 24949 5012 24961 5015
rect 24912 4984 24961 5012
rect 24912 4972 24918 4984
rect 24949 4981 24961 4984
rect 24995 4981 25007 5015
rect 24949 4975 25007 4981
rect 28810 4972 28816 5024
rect 28868 5012 28874 5024
rect 28905 5015 28963 5021
rect 28905 5012 28917 5015
rect 28868 4984 28917 5012
rect 28868 4972 28874 4984
rect 28905 4981 28917 4984
rect 28951 4981 28963 5015
rect 28905 4975 28963 4981
rect 34241 5015 34299 5021
rect 34241 4981 34253 5015
rect 34287 5012 34299 5015
rect 34606 5012 34612 5024
rect 34287 4984 34612 5012
rect 34287 4981 34299 4984
rect 34241 4975 34299 4981
rect 34606 4972 34612 4984
rect 34664 4972 34670 5024
rect 58710 4972 58716 5024
rect 58768 5012 58774 5024
rect 58805 5015 58863 5021
rect 58805 5012 58817 5015
rect 58768 4984 58817 5012
rect 58768 4972 58774 4984
rect 58805 4981 58817 4984
rect 58851 4981 58863 5015
rect 58805 4975 58863 4981
rect 1104 4922 68816 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 65654 4922
rect 65706 4870 65718 4922
rect 65770 4870 65782 4922
rect 65834 4870 65846 4922
rect 65898 4870 65910 4922
rect 65962 4870 68816 4922
rect 1104 4848 68816 4870
rect 2133 4811 2191 4817
rect 2133 4777 2145 4811
rect 2179 4808 2191 4811
rect 2314 4808 2320 4820
rect 2179 4780 2320 4808
rect 2179 4777 2191 4780
rect 2133 4771 2191 4777
rect 2314 4768 2320 4780
rect 2372 4768 2378 4820
rect 3881 4811 3939 4817
rect 3881 4777 3893 4811
rect 3927 4808 3939 4811
rect 3970 4808 3976 4820
rect 3927 4780 3976 4808
rect 3927 4777 3939 4780
rect 3881 4771 3939 4777
rect 3970 4768 3976 4780
rect 4028 4768 4034 4820
rect 5626 4768 5632 4820
rect 5684 4808 5690 4820
rect 8386 4808 8392 4820
rect 5684 4780 7972 4808
rect 8347 4780 8392 4808
rect 5684 4768 5690 4780
rect 7944 4740 7972 4780
rect 8386 4768 8392 4780
rect 8444 4768 8450 4820
rect 9766 4808 9772 4820
rect 8496 4780 9772 4808
rect 8496 4740 8524 4780
rect 9766 4768 9772 4780
rect 9824 4768 9830 4820
rect 10505 4811 10563 4817
rect 10505 4777 10517 4811
rect 10551 4808 10563 4811
rect 10594 4808 10600 4820
rect 10551 4780 10600 4808
rect 10551 4777 10563 4780
rect 10505 4771 10563 4777
rect 10594 4768 10600 4780
rect 10652 4768 10658 4820
rect 11238 4768 11244 4820
rect 11296 4808 11302 4820
rect 12158 4808 12164 4820
rect 11296 4780 12164 4808
rect 11296 4768 11302 4780
rect 12158 4768 12164 4780
rect 12216 4768 12222 4820
rect 14090 4808 14096 4820
rect 14051 4780 14096 4808
rect 14090 4768 14096 4780
rect 14148 4768 14154 4820
rect 21266 4808 21272 4820
rect 18248 4780 21272 4808
rect 7944 4712 8524 4740
rect 9125 4743 9183 4749
rect 9125 4709 9137 4743
rect 9171 4740 9183 4743
rect 11606 4740 11612 4752
rect 9171 4712 11612 4740
rect 9171 4709 9183 4712
rect 9125 4703 9183 4709
rect 11606 4700 11612 4712
rect 11664 4700 11670 4752
rect 12250 4740 12256 4752
rect 11808 4712 12256 4740
rect 2222 4672 2228 4684
rect 1964 4644 2228 4672
rect 1762 4604 1768 4616
rect 1723 4576 1768 4604
rect 1762 4564 1768 4576
rect 1820 4564 1826 4616
rect 1964 4613 1992 4644
rect 2222 4632 2228 4644
rect 2280 4672 2286 4684
rect 5718 4672 5724 4684
rect 2280 4644 5724 4672
rect 2280 4632 2286 4644
rect 5718 4632 5724 4644
rect 5776 4632 5782 4684
rect 11146 4672 11152 4684
rect 8956 4644 11152 4672
rect 1949 4607 2007 4613
rect 1949 4573 1961 4607
rect 1995 4573 2007 4607
rect 2961 4607 3019 4613
rect 2961 4604 2973 4607
rect 1949 4567 2007 4573
rect 2148 4576 2973 4604
rect 1780 4536 1808 4564
rect 2148 4536 2176 4576
rect 2961 4573 2973 4576
rect 3007 4573 3019 4607
rect 2961 4567 3019 4573
rect 5997 4607 6055 4613
rect 5997 4573 6009 4607
rect 6043 4604 6055 4607
rect 6043 4576 6868 4604
rect 6043 4573 6055 4576
rect 5997 4567 6055 4573
rect 1780 4508 2176 4536
rect 2777 4539 2835 4545
rect 2777 4505 2789 4539
rect 2823 4536 2835 4539
rect 3142 4536 3148 4548
rect 2823 4508 3148 4536
rect 2823 4505 2835 4508
rect 2777 4499 2835 4505
rect 3142 4496 3148 4508
rect 3200 4536 3206 4548
rect 3970 4536 3976 4548
rect 3200 4508 3976 4536
rect 3200 4496 3206 4508
rect 3970 4496 3976 4508
rect 4028 4496 4034 4548
rect 4893 4539 4951 4545
rect 4893 4505 4905 4539
rect 4939 4536 4951 4539
rect 6638 4536 6644 4548
rect 4939 4508 6644 4536
rect 4939 4505 4951 4508
rect 4893 4499 4951 4505
rect 6638 4496 6644 4508
rect 6696 4496 6702 4548
rect 6840 4536 6868 4576
rect 6914 4564 6920 4616
rect 6972 4604 6978 4616
rect 7009 4607 7067 4613
rect 7009 4604 7021 4607
rect 6972 4576 7021 4604
rect 6972 4564 6978 4576
rect 7009 4573 7021 4576
rect 7055 4573 7067 4607
rect 7009 4567 7067 4573
rect 7276 4607 7334 4613
rect 7276 4573 7288 4607
rect 7322 4604 7334 4607
rect 7742 4604 7748 4616
rect 7322 4576 7748 4604
rect 7322 4573 7334 4576
rect 7276 4567 7334 4573
rect 7742 4564 7748 4576
rect 7800 4564 7806 4616
rect 8956 4613 8984 4644
rect 11146 4632 11152 4644
rect 11204 4632 11210 4684
rect 8941 4607 8999 4613
rect 8941 4573 8953 4607
rect 8987 4573 8999 4607
rect 8941 4567 8999 4573
rect 9585 4607 9643 4613
rect 9585 4573 9597 4607
rect 9631 4604 9643 4607
rect 10318 4604 10324 4616
rect 9631 4576 9904 4604
rect 10279 4576 10324 4604
rect 9631 4573 9643 4576
rect 9585 4567 9643 4573
rect 8956 4536 8984 4567
rect 6840 4508 8984 4536
rect 2314 4428 2320 4480
rect 2372 4468 2378 4480
rect 2593 4471 2651 4477
rect 2593 4468 2605 4471
rect 2372 4440 2605 4468
rect 2372 4428 2378 4440
rect 2593 4437 2605 4440
rect 2639 4437 2651 4471
rect 2593 4431 2651 4437
rect 5445 4471 5503 4477
rect 5445 4437 5457 4471
rect 5491 4468 5503 4471
rect 5534 4468 5540 4480
rect 5491 4440 5540 4468
rect 5491 4437 5503 4440
rect 5445 4431 5503 4437
rect 5534 4428 5540 4440
rect 5592 4428 5598 4480
rect 6549 4471 6607 4477
rect 6549 4437 6561 4471
rect 6595 4468 6607 4471
rect 9600 4468 9628 4567
rect 9766 4468 9772 4480
rect 6595 4440 9628 4468
rect 9727 4440 9772 4468
rect 6595 4437 6607 4440
rect 6549 4431 6607 4437
rect 9766 4428 9772 4440
rect 9824 4428 9830 4480
rect 9876 4468 9904 4576
rect 10318 4564 10324 4576
rect 10376 4564 10382 4616
rect 11057 4607 11115 4613
rect 11057 4573 11069 4607
rect 11103 4604 11115 4607
rect 11238 4604 11244 4616
rect 11103 4576 11244 4604
rect 11103 4573 11115 4576
rect 11057 4567 11115 4573
rect 11238 4564 11244 4576
rect 11296 4564 11302 4616
rect 11808 4613 11836 4712
rect 12250 4700 12256 4712
rect 12308 4700 12314 4752
rect 12066 4672 12072 4684
rect 12027 4644 12072 4672
rect 12066 4632 12072 4644
rect 12124 4632 12130 4684
rect 12161 4675 12219 4681
rect 12161 4641 12173 4675
rect 12207 4672 12219 4675
rect 12526 4672 12532 4684
rect 12207 4644 12532 4672
rect 12207 4641 12219 4644
rect 12161 4635 12219 4641
rect 12526 4632 12532 4644
rect 12584 4632 12590 4684
rect 14108 4672 14136 4768
rect 16577 4743 16635 4749
rect 16577 4709 16589 4743
rect 16623 4740 16635 4743
rect 18046 4740 18052 4752
rect 16623 4712 18052 4740
rect 16623 4709 16635 4712
rect 16577 4703 16635 4709
rect 18046 4700 18052 4712
rect 18104 4700 18110 4752
rect 18248 4749 18276 4780
rect 21266 4768 21272 4780
rect 21324 4768 21330 4820
rect 22186 4768 22192 4820
rect 22244 4808 22250 4820
rect 22922 4808 22928 4820
rect 22244 4780 22784 4808
rect 22883 4780 22928 4808
rect 22244 4768 22250 4780
rect 18233 4743 18291 4749
rect 18233 4709 18245 4743
rect 18279 4709 18291 4743
rect 18233 4703 18291 4709
rect 18598 4700 18604 4752
rect 18656 4740 18662 4752
rect 21177 4743 21235 4749
rect 21177 4740 21189 4743
rect 18656 4712 21189 4740
rect 18656 4700 18662 4712
rect 21177 4709 21189 4712
rect 21223 4709 21235 4743
rect 21177 4703 21235 4709
rect 22554 4700 22560 4752
rect 22612 4700 22618 4752
rect 13280 4644 14136 4672
rect 15473 4675 15531 4681
rect 11793 4607 11851 4613
rect 11793 4573 11805 4607
rect 11839 4573 11851 4607
rect 11974 4604 11980 4616
rect 11935 4576 11980 4604
rect 11793 4567 11851 4573
rect 11974 4564 11980 4576
rect 12032 4564 12038 4616
rect 12342 4604 12348 4616
rect 12303 4576 12348 4604
rect 12342 4564 12348 4576
rect 12400 4564 12406 4616
rect 10134 4496 10140 4548
rect 10192 4536 10198 4548
rect 10413 4539 10471 4545
rect 10413 4536 10425 4539
rect 10192 4508 10425 4536
rect 10192 4496 10198 4508
rect 10413 4505 10425 4508
rect 10459 4505 10471 4539
rect 10413 4499 10471 4505
rect 10597 4539 10655 4545
rect 10597 4505 10609 4539
rect 10643 4536 10655 4539
rect 10870 4536 10876 4548
rect 10643 4508 10876 4536
rect 10643 4505 10655 4508
rect 10597 4499 10655 4505
rect 10870 4496 10876 4508
rect 10928 4496 10934 4548
rect 11882 4536 11888 4548
rect 10980 4508 11888 4536
rect 10980 4468 11008 4508
rect 11882 4496 11888 4508
rect 11940 4496 11946 4548
rect 13280 4536 13308 4644
rect 15473 4641 15485 4675
rect 15519 4672 15531 4675
rect 16666 4672 16672 4684
rect 15519 4644 16672 4672
rect 15519 4641 15531 4644
rect 15473 4635 15531 4641
rect 13722 4564 13728 4616
rect 13780 4604 13786 4616
rect 15488 4604 15516 4635
rect 16666 4632 16672 4644
rect 16724 4632 16730 4684
rect 17402 4632 17408 4684
rect 17460 4672 17466 4684
rect 17460 4644 18644 4672
rect 17460 4632 17466 4644
rect 13780 4576 15516 4604
rect 17313 4607 17371 4613
rect 13780 4564 13786 4576
rect 17313 4573 17325 4607
rect 17359 4573 17371 4607
rect 17313 4567 17371 4573
rect 17681 4607 17739 4613
rect 17681 4573 17693 4607
rect 17727 4573 17739 4607
rect 17862 4604 17868 4616
rect 17823 4576 17868 4604
rect 17681 4567 17739 4573
rect 11992 4508 13308 4536
rect 13357 4539 13415 4545
rect 11992 4480 12020 4508
rect 13357 4505 13369 4539
rect 13403 4505 13415 4539
rect 13357 4499 13415 4505
rect 9876 4440 11008 4468
rect 11241 4471 11299 4477
rect 11241 4437 11253 4471
rect 11287 4468 11299 4471
rect 11330 4468 11336 4480
rect 11287 4440 11336 4468
rect 11287 4437 11299 4440
rect 11241 4431 11299 4437
rect 11330 4428 11336 4440
rect 11388 4428 11394 4480
rect 11974 4428 11980 4480
rect 12032 4428 12038 4480
rect 12526 4468 12532 4480
rect 12487 4440 12532 4468
rect 12526 4428 12532 4440
rect 12584 4428 12590 4480
rect 13262 4428 13268 4480
rect 13320 4468 13326 4480
rect 13372 4468 13400 4499
rect 15194 4496 15200 4548
rect 15252 4545 15258 4548
rect 15252 4536 15264 4545
rect 15252 4508 15297 4536
rect 15252 4499 15264 4508
rect 15252 4496 15258 4499
rect 16574 4496 16580 4548
rect 16632 4536 16638 4548
rect 17328 4536 17356 4567
rect 17586 4536 17592 4548
rect 16632 4508 17264 4536
rect 17328 4508 17592 4536
rect 16632 4496 16638 4508
rect 13320 4440 13400 4468
rect 13449 4471 13507 4477
rect 13320 4428 13326 4440
rect 13449 4437 13461 4471
rect 13495 4468 13507 4471
rect 16758 4468 16764 4480
rect 13495 4440 16764 4468
rect 13495 4437 13507 4440
rect 13449 4431 13507 4437
rect 16758 4428 16764 4440
rect 16816 4468 16822 4480
rect 17034 4468 17040 4480
rect 16816 4440 17040 4468
rect 16816 4428 16822 4440
rect 17034 4428 17040 4440
rect 17092 4428 17098 4480
rect 17236 4468 17264 4508
rect 17586 4496 17592 4508
rect 17644 4496 17650 4548
rect 17696 4468 17724 4567
rect 17862 4564 17868 4576
rect 17920 4564 17926 4616
rect 18616 4613 18644 4644
rect 19150 4632 19156 4684
rect 19208 4672 19214 4684
rect 20533 4675 20591 4681
rect 20533 4672 20545 4675
rect 19208 4644 20545 4672
rect 19208 4632 19214 4644
rect 20533 4641 20545 4644
rect 20579 4641 20591 4675
rect 20533 4635 20591 4641
rect 18601 4607 18659 4613
rect 18601 4573 18613 4607
rect 18647 4573 18659 4607
rect 18601 4567 18659 4573
rect 19058 4564 19064 4616
rect 19116 4604 19122 4616
rect 19334 4604 19340 4616
rect 19116 4576 19340 4604
rect 19116 4564 19122 4576
rect 19334 4564 19340 4576
rect 19392 4564 19398 4616
rect 19426 4564 19432 4616
rect 19484 4604 19490 4616
rect 19521 4607 19579 4613
rect 19521 4604 19533 4607
rect 19484 4576 19533 4604
rect 19484 4564 19490 4576
rect 19521 4573 19533 4576
rect 19567 4573 19579 4607
rect 19521 4567 19579 4573
rect 19702 4564 19708 4616
rect 19760 4604 19766 4616
rect 19797 4607 19855 4613
rect 19797 4604 19809 4607
rect 19760 4576 19809 4604
rect 19760 4564 19766 4576
rect 19797 4573 19809 4576
rect 19843 4573 19855 4607
rect 19978 4604 19984 4616
rect 19939 4576 19984 4604
rect 19797 4567 19855 4573
rect 19812 4536 19840 4567
rect 19978 4564 19984 4576
rect 20036 4564 20042 4616
rect 22186 4564 22192 4616
rect 22244 4604 22250 4616
rect 22572 4613 22600 4700
rect 22756 4672 22784 4780
rect 22922 4768 22928 4780
rect 22980 4768 22986 4820
rect 23842 4808 23848 4820
rect 23755 4780 23848 4808
rect 23842 4768 23848 4780
rect 23900 4808 23906 4820
rect 24578 4808 24584 4820
rect 23900 4780 24584 4808
rect 23900 4768 23906 4780
rect 24578 4768 24584 4780
rect 24636 4808 24642 4820
rect 25038 4808 25044 4820
rect 24636 4780 25044 4808
rect 24636 4768 24642 4780
rect 25038 4768 25044 4780
rect 25096 4768 25102 4820
rect 28718 4768 28724 4820
rect 28776 4808 28782 4820
rect 28776 4780 28994 4808
rect 28776 4768 28782 4780
rect 28166 4740 28172 4752
rect 26804 4712 28172 4740
rect 22756 4644 25084 4672
rect 22281 4607 22339 4613
rect 22281 4604 22293 4607
rect 22244 4576 22293 4604
rect 22244 4564 22250 4576
rect 22281 4573 22293 4576
rect 22327 4573 22339 4607
rect 22444 4607 22502 4613
rect 22444 4604 22456 4607
rect 22281 4567 22339 4573
rect 22368 4576 22456 4604
rect 20530 4536 20536 4548
rect 19812 4508 20536 4536
rect 20530 4496 20536 4508
rect 20588 4496 20594 4548
rect 17236 4440 17724 4468
rect 19981 4471 20039 4477
rect 19981 4437 19993 4471
rect 20027 4468 20039 4471
rect 20162 4468 20168 4480
rect 20027 4440 20168 4468
rect 20027 4437 20039 4440
rect 19981 4431 20039 4437
rect 20162 4428 20168 4440
rect 20220 4428 20226 4480
rect 22186 4428 22192 4480
rect 22244 4468 22250 4480
rect 22368 4468 22396 4576
rect 22444 4573 22456 4576
rect 22490 4573 22502 4607
rect 22444 4567 22502 4573
rect 22544 4607 22602 4613
rect 22544 4573 22556 4607
rect 22590 4573 22602 4607
rect 22544 4567 22602 4573
rect 22695 4607 22753 4613
rect 22695 4573 22707 4607
rect 22741 4604 22753 4607
rect 22830 4604 22836 4616
rect 22741 4576 22836 4604
rect 22741 4573 22753 4576
rect 22695 4567 22753 4573
rect 22830 4564 22836 4576
rect 22888 4564 22894 4616
rect 24578 4564 24584 4616
rect 24636 4604 24642 4616
rect 24673 4607 24731 4613
rect 24673 4604 24685 4607
rect 24636 4576 24685 4604
rect 24636 4564 24642 4576
rect 24673 4573 24685 4576
rect 24719 4573 24731 4607
rect 24673 4567 24731 4573
rect 24765 4607 24823 4613
rect 24765 4573 24777 4607
rect 24811 4573 24823 4607
rect 24765 4567 24823 4573
rect 24780 4536 24808 4567
rect 24854 4564 24860 4616
rect 24912 4604 24918 4616
rect 25056 4613 25084 4644
rect 25590 4632 25596 4684
rect 25648 4672 25654 4684
rect 26804 4681 26832 4712
rect 28166 4700 28172 4712
rect 28224 4700 28230 4752
rect 28258 4700 28264 4752
rect 28316 4740 28322 4752
rect 28626 4740 28632 4752
rect 28316 4712 28632 4740
rect 28316 4700 28322 4712
rect 28626 4700 28632 4712
rect 28684 4740 28690 4752
rect 28966 4740 28994 4780
rect 30282 4768 30288 4820
rect 30340 4808 30346 4820
rect 31757 4811 31815 4817
rect 31757 4808 31769 4811
rect 30340 4780 31769 4808
rect 30340 4768 30346 4780
rect 31757 4777 31769 4780
rect 31803 4777 31815 4811
rect 31757 4771 31815 4777
rect 36357 4811 36415 4817
rect 36357 4777 36369 4811
rect 36403 4808 36415 4811
rect 36446 4808 36452 4820
rect 36403 4780 36452 4808
rect 36403 4777 36415 4780
rect 36357 4771 36415 4777
rect 36446 4768 36452 4780
rect 36504 4768 36510 4820
rect 32122 4740 32128 4752
rect 28684 4712 28764 4740
rect 28966 4712 32128 4740
rect 28684 4700 28690 4712
rect 26789 4675 26847 4681
rect 26789 4672 26801 4675
rect 25648 4644 26801 4672
rect 25648 4632 25654 4644
rect 25041 4607 25099 4613
rect 24912 4576 24957 4604
rect 24912 4564 24918 4576
rect 25041 4573 25053 4607
rect 25087 4604 25099 4607
rect 25682 4604 25688 4616
rect 25087 4576 25688 4604
rect 25087 4573 25099 4576
rect 25041 4567 25099 4573
rect 25682 4564 25688 4576
rect 25740 4564 25746 4616
rect 25866 4604 25872 4616
rect 25827 4576 25872 4604
rect 25866 4564 25872 4576
rect 25924 4564 25930 4616
rect 26068 4613 26096 4644
rect 26789 4641 26801 4644
rect 26835 4641 26847 4675
rect 26789 4635 26847 4641
rect 25961 4607 26019 4613
rect 25961 4573 25973 4607
rect 26007 4573 26019 4607
rect 25961 4567 26019 4573
rect 26053 4607 26111 4613
rect 26053 4573 26065 4607
rect 26099 4573 26111 4607
rect 27798 4604 27804 4616
rect 27759 4576 27804 4604
rect 26053 4567 26111 4573
rect 25774 4536 25780 4548
rect 24780 4508 25780 4536
rect 24394 4468 24400 4480
rect 22244 4440 22396 4468
rect 24355 4440 24400 4468
rect 22244 4428 22250 4440
rect 24394 4428 24400 4440
rect 24452 4428 24458 4480
rect 24670 4428 24676 4480
rect 24728 4468 24734 4480
rect 24780 4468 24808 4508
rect 25774 4496 25780 4508
rect 25832 4536 25838 4548
rect 25976 4536 26004 4567
rect 27798 4564 27804 4576
rect 27856 4604 27862 4616
rect 28736 4613 28764 4712
rect 32122 4700 32128 4712
rect 32180 4700 32186 4752
rect 36262 4700 36268 4752
rect 36320 4740 36326 4752
rect 37001 4743 37059 4749
rect 37001 4740 37013 4743
rect 36320 4712 37013 4740
rect 36320 4700 36326 4712
rect 37001 4709 37013 4712
rect 37047 4709 37059 4743
rect 37001 4703 37059 4709
rect 57238 4700 57244 4752
rect 57296 4740 57302 4752
rect 57885 4743 57943 4749
rect 57885 4740 57897 4743
rect 57296 4712 57897 4740
rect 57296 4700 57302 4712
rect 57885 4709 57897 4712
rect 57931 4709 57943 4743
rect 57885 4703 57943 4709
rect 58250 4700 58256 4752
rect 58308 4740 58314 4752
rect 59173 4743 59231 4749
rect 59173 4740 59185 4743
rect 58308 4712 59185 4740
rect 58308 4700 58314 4712
rect 59173 4709 59185 4712
rect 59219 4709 59231 4743
rect 59173 4703 59231 4709
rect 28902 4632 28908 4684
rect 28960 4672 28966 4684
rect 36170 4672 36176 4684
rect 28960 4644 29868 4672
rect 28960 4632 28966 4644
rect 28629 4607 28687 4613
rect 27856 4601 28580 4604
rect 28629 4601 28641 4607
rect 27856 4576 28641 4601
rect 27856 4564 27862 4576
rect 28552 4573 28641 4576
rect 28675 4573 28687 4607
rect 28629 4567 28687 4573
rect 28718 4607 28776 4613
rect 28718 4573 28730 4607
rect 28764 4573 28776 4607
rect 28718 4567 28776 4573
rect 28810 4564 28816 4616
rect 28868 4604 28874 4616
rect 28868 4576 28913 4604
rect 28868 4564 28874 4576
rect 28994 4564 29000 4616
rect 29052 4604 29058 4616
rect 29549 4607 29607 4613
rect 29549 4604 29561 4607
rect 29052 4576 29561 4604
rect 29052 4564 29058 4576
rect 29549 4573 29561 4576
rect 29595 4573 29607 4607
rect 29730 4604 29736 4616
rect 29691 4576 29736 4604
rect 29549 4567 29607 4573
rect 29730 4564 29736 4576
rect 29788 4564 29794 4616
rect 29840 4613 29868 4644
rect 33060 4644 36176 4672
rect 29825 4607 29883 4613
rect 29825 4573 29837 4607
rect 29871 4573 29883 4607
rect 29825 4567 29883 4573
rect 29914 4564 29920 4616
rect 29972 4604 29978 4616
rect 29972 4576 30017 4604
rect 29972 4564 29978 4576
rect 32582 4564 32588 4616
rect 32640 4604 32646 4616
rect 33060 4604 33088 4644
rect 36170 4632 36176 4644
rect 36228 4672 36234 4684
rect 36228 4644 36308 4672
rect 36228 4632 36234 4644
rect 32640 4576 33088 4604
rect 33137 4607 33195 4613
rect 32640 4564 32646 4576
rect 33137 4573 33149 4607
rect 33183 4604 33195 4607
rect 34514 4604 34520 4616
rect 33183 4576 34520 4604
rect 33183 4573 33195 4576
rect 33137 4567 33195 4573
rect 34514 4564 34520 4576
rect 34572 4564 34578 4616
rect 36280 4613 36308 4644
rect 58894 4632 58900 4684
rect 58952 4672 58958 4684
rect 60461 4675 60519 4681
rect 60461 4672 60473 4675
rect 58952 4644 60473 4672
rect 58952 4632 58958 4644
rect 60461 4641 60473 4644
rect 60507 4641 60519 4675
rect 60461 4635 60519 4641
rect 36265 4607 36323 4613
rect 36265 4573 36277 4607
rect 36311 4573 36323 4607
rect 36906 4604 36912 4616
rect 36867 4576 36912 4604
rect 36265 4567 36323 4573
rect 36906 4564 36912 4576
rect 36964 4564 36970 4616
rect 57146 4564 57152 4616
rect 57204 4604 57210 4616
rect 57241 4607 57299 4613
rect 57241 4604 57253 4607
rect 57204 4576 57253 4604
rect 57204 4564 57210 4576
rect 57241 4573 57253 4576
rect 57287 4573 57299 4607
rect 57241 4567 57299 4573
rect 57606 4564 57612 4616
rect 57664 4604 57670 4616
rect 58529 4607 58587 4613
rect 58529 4604 58541 4607
rect 57664 4576 58541 4604
rect 57664 4564 57670 4576
rect 58529 4573 58541 4576
rect 58575 4573 58587 4607
rect 58529 4567 58587 4573
rect 25832 4508 26004 4536
rect 26329 4539 26387 4545
rect 25832 4496 25838 4508
rect 26329 4505 26341 4539
rect 26375 4536 26387 4539
rect 27246 4536 27252 4548
rect 26375 4508 27252 4536
rect 26375 4505 26387 4508
rect 26329 4499 26387 4505
rect 27246 4496 27252 4508
rect 27304 4496 27310 4548
rect 28353 4539 28411 4545
rect 28353 4505 28365 4539
rect 28399 4536 28411 4539
rect 32870 4539 32928 4545
rect 32870 4536 32882 4539
rect 28399 4508 32882 4536
rect 28399 4505 28411 4508
rect 28353 4499 28411 4505
rect 32870 4505 32882 4508
rect 32916 4505 32928 4539
rect 32870 4499 32928 4505
rect 24728 4440 24808 4468
rect 30193 4471 30251 4477
rect 24728 4428 24734 4440
rect 30193 4437 30205 4471
rect 30239 4468 30251 4471
rect 30282 4468 30288 4480
rect 30239 4440 30288 4468
rect 30239 4437 30251 4440
rect 30193 4431 30251 4437
rect 30282 4428 30288 4440
rect 30340 4428 30346 4480
rect 1104 4378 68816 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 50294 4378
rect 50346 4326 50358 4378
rect 50410 4326 50422 4378
rect 50474 4326 50486 4378
rect 50538 4326 50550 4378
rect 50602 4326 68816 4378
rect 1104 4304 68816 4326
rect 6822 4264 6828 4276
rect 6748 4236 6828 4264
rect 2406 4196 2412 4208
rect 2240 4168 2412 4196
rect 2130 4128 2136 4140
rect 2091 4100 2136 4128
rect 2130 4088 2136 4100
rect 2188 4088 2194 4140
rect 2240 4137 2268 4168
rect 2406 4156 2412 4168
rect 2464 4156 2470 4208
rect 3418 4196 3424 4208
rect 2976 4168 3424 4196
rect 2225 4131 2283 4137
rect 2225 4097 2237 4131
rect 2271 4097 2283 4131
rect 2225 4091 2283 4097
rect 2314 4088 2320 4140
rect 2372 4128 2378 4140
rect 2372 4100 2417 4128
rect 2372 4088 2378 4100
rect 2498 4088 2504 4140
rect 2556 4128 2562 4140
rect 2976 4137 3004 4168
rect 3418 4156 3424 4168
rect 3476 4156 3482 4208
rect 5626 4196 5632 4208
rect 5587 4168 5632 4196
rect 5626 4156 5632 4168
rect 5684 4156 5690 4208
rect 5813 4199 5871 4205
rect 5813 4165 5825 4199
rect 5859 4196 5871 4199
rect 6546 4196 6552 4208
rect 5859 4168 6552 4196
rect 5859 4165 5871 4168
rect 5813 4159 5871 4165
rect 6546 4156 6552 4168
rect 6604 4156 6610 4208
rect 2961 4131 3019 4137
rect 2556 4100 2601 4128
rect 2556 4088 2562 4100
rect 2961 4097 2973 4131
rect 3007 4097 3019 4131
rect 3217 4131 3275 4137
rect 3217 4128 3229 4131
rect 2961 4091 3019 4097
rect 3068 4100 3229 4128
rect 1857 4063 1915 4069
rect 1857 4029 1869 4063
rect 1903 4060 1915 4063
rect 3068 4060 3096 4100
rect 3217 4097 3229 4100
rect 3263 4097 3275 4131
rect 4982 4128 4988 4140
rect 4943 4100 4988 4128
rect 3217 4091 3275 4097
rect 4982 4088 4988 4100
rect 5040 4088 5046 4140
rect 6638 4128 6644 4140
rect 6599 4100 6644 4128
rect 6638 4088 6644 4100
rect 6696 4088 6702 4140
rect 6748 4137 6776 4236
rect 6822 4224 6828 4236
rect 6880 4224 6886 4276
rect 9674 4224 9680 4276
rect 9732 4264 9738 4276
rect 10226 4264 10232 4276
rect 9732 4236 10232 4264
rect 9732 4224 9738 4236
rect 10226 4224 10232 4236
rect 10284 4264 10290 4276
rect 11790 4264 11796 4276
rect 10284 4236 11796 4264
rect 10284 4224 10290 4236
rect 11790 4224 11796 4236
rect 11848 4224 11854 4276
rect 12069 4267 12127 4273
rect 12069 4233 12081 4267
rect 12115 4264 12127 4267
rect 12342 4264 12348 4276
rect 12115 4236 12348 4264
rect 12115 4233 12127 4236
rect 12069 4227 12127 4233
rect 12342 4224 12348 4236
rect 12400 4224 12406 4276
rect 17221 4267 17279 4273
rect 17221 4233 17233 4267
rect 17267 4264 17279 4267
rect 17267 4236 22094 4264
rect 17267 4233 17279 4236
rect 17221 4227 17279 4233
rect 8938 4196 8944 4208
rect 8899 4168 8944 4196
rect 8938 4156 8944 4168
rect 8996 4156 9002 4208
rect 9508 4168 9812 4196
rect 6733 4131 6791 4137
rect 6733 4097 6745 4131
rect 6779 4097 6791 4131
rect 6733 4091 6791 4097
rect 6825 4131 6883 4137
rect 6825 4097 6837 4131
rect 6871 4097 6883 4131
rect 7006 4128 7012 4140
rect 6967 4100 7012 4128
rect 6825 4091 6883 4097
rect 1903 4032 3096 4060
rect 5445 4063 5503 4069
rect 1903 4029 1915 4032
rect 1857 4023 1915 4029
rect 5445 4029 5457 4063
rect 5491 4060 5503 4063
rect 6840 4060 6868 4091
rect 7006 4088 7012 4100
rect 7064 4088 7070 4140
rect 7469 4131 7527 4137
rect 7469 4097 7481 4131
rect 7515 4097 7527 4131
rect 7469 4091 7527 4097
rect 8389 4131 8447 4137
rect 8389 4097 8401 4131
rect 8435 4128 8447 4131
rect 8570 4128 8576 4140
rect 8435 4100 8576 4128
rect 8435 4097 8447 4100
rect 8389 4091 8447 4097
rect 5491 4032 6868 4060
rect 7484 4060 7512 4091
rect 8570 4088 8576 4100
rect 8628 4088 8634 4140
rect 9508 4128 9536 4168
rect 9674 4128 9680 4140
rect 8680 4100 9536 4128
rect 9635 4100 9680 4128
rect 8680 4060 8708 4100
rect 9674 4088 9680 4100
rect 9732 4088 9738 4140
rect 9784 4128 9812 4168
rect 9858 4156 9864 4208
rect 9916 4196 9922 4208
rect 12434 4196 12440 4208
rect 9916 4168 10364 4196
rect 9916 4156 9922 4168
rect 10226 4128 10232 4140
rect 9784 4100 10232 4128
rect 10226 4088 10232 4100
rect 10284 4088 10290 4140
rect 10336 4137 10364 4168
rect 10888 4168 12440 4196
rect 10321 4131 10379 4137
rect 10321 4097 10333 4131
rect 10367 4097 10379 4131
rect 10502 4128 10508 4140
rect 10463 4100 10508 4128
rect 10321 4091 10379 4097
rect 10502 4088 10508 4100
rect 10560 4088 10566 4140
rect 10781 4131 10839 4137
rect 10781 4097 10793 4131
rect 10827 4128 10839 4131
rect 10888 4128 10916 4168
rect 12434 4156 12440 4168
rect 12492 4156 12498 4208
rect 12526 4156 12532 4208
rect 12584 4196 12590 4208
rect 13182 4199 13240 4205
rect 13182 4196 13194 4199
rect 12584 4168 13194 4196
rect 12584 4156 12590 4168
rect 13182 4165 13194 4168
rect 13228 4165 13240 4199
rect 17402 4196 17408 4208
rect 13182 4159 13240 4165
rect 16868 4168 17408 4196
rect 16868 4140 16896 4168
rect 17402 4156 17408 4168
rect 17460 4156 17466 4208
rect 22066 4196 22094 4236
rect 22186 4224 22192 4276
rect 22244 4264 22250 4276
rect 24210 4264 24216 4276
rect 22244 4236 22289 4264
rect 22480 4236 24216 4264
rect 22244 4224 22250 4236
rect 22278 4196 22284 4208
rect 22066 4168 22284 4196
rect 22278 4156 22284 4168
rect 22336 4156 22342 4208
rect 22373 4199 22431 4205
rect 22373 4165 22385 4199
rect 22419 4196 22431 4199
rect 22480 4196 22508 4236
rect 24210 4224 24216 4236
rect 24268 4224 24274 4276
rect 24762 4264 24768 4276
rect 24723 4236 24768 4264
rect 24762 4224 24768 4236
rect 24820 4224 24826 4276
rect 25777 4267 25835 4273
rect 25777 4233 25789 4267
rect 25823 4264 25835 4267
rect 25866 4264 25872 4276
rect 25823 4236 25872 4264
rect 25823 4233 25835 4236
rect 25777 4227 25835 4233
rect 25866 4224 25872 4236
rect 25924 4224 25930 4276
rect 29181 4267 29239 4273
rect 29181 4233 29193 4267
rect 29227 4264 29239 4267
rect 29730 4264 29736 4276
rect 29227 4236 29736 4264
rect 29227 4233 29239 4236
rect 29181 4227 29239 4233
rect 29730 4224 29736 4236
rect 29788 4224 29794 4276
rect 31389 4267 31447 4273
rect 31389 4233 31401 4267
rect 31435 4233 31447 4267
rect 31389 4227 31447 4233
rect 22419 4168 22508 4196
rect 22557 4199 22615 4205
rect 22419 4165 22431 4168
rect 22373 4159 22431 4165
rect 22557 4165 22569 4199
rect 22603 4196 22615 4199
rect 23474 4196 23480 4208
rect 22603 4168 23480 4196
rect 22603 4165 22615 4168
rect 22557 4159 22615 4165
rect 23474 4156 23480 4168
rect 23532 4156 23538 4208
rect 23652 4199 23710 4205
rect 23652 4165 23664 4199
rect 23698 4196 23710 4199
rect 24394 4196 24400 4208
rect 23698 4168 24400 4196
rect 23698 4165 23710 4168
rect 23652 4159 23710 4165
rect 24394 4156 24400 4168
rect 24452 4156 24458 4208
rect 25130 4156 25136 4208
rect 25188 4196 25194 4208
rect 26145 4199 26203 4205
rect 26145 4196 26157 4199
rect 25188 4168 26157 4196
rect 25188 4156 25194 4168
rect 26145 4165 26157 4168
rect 26191 4165 26203 4199
rect 26145 4159 26203 4165
rect 27080 4168 27384 4196
rect 10827 4100 10916 4128
rect 10965 4131 11023 4137
rect 10827 4097 10839 4100
rect 10781 4091 10839 4097
rect 10965 4097 10977 4131
rect 11011 4128 11023 4131
rect 11054 4128 11060 4140
rect 11011 4100 11060 4128
rect 11011 4097 11023 4100
rect 10965 4091 11023 4097
rect 11054 4088 11060 4100
rect 11112 4088 11118 4140
rect 11609 4131 11667 4137
rect 11609 4097 11621 4131
rect 11655 4128 11667 4131
rect 12894 4128 12900 4140
rect 11655 4100 12900 4128
rect 11655 4097 11667 4100
rect 11609 4091 11667 4097
rect 12894 4088 12900 4100
rect 12952 4128 12958 4140
rect 13449 4131 13507 4137
rect 12952 4100 13400 4128
rect 12952 4088 12958 4100
rect 7484 4032 8708 4060
rect 9125 4063 9183 4069
rect 5491 4029 5503 4032
rect 5445 4023 5503 4029
rect 5534 3952 5540 4004
rect 5592 3992 5598 4004
rect 7484 3992 7512 4032
rect 9125 4029 9137 4063
rect 9171 4060 9183 4063
rect 12434 4060 12440 4072
rect 9171 4032 12440 4060
rect 9171 4029 9183 4032
rect 9125 4023 9183 4029
rect 12434 4020 12440 4032
rect 12492 4020 12498 4072
rect 13372 4060 13400 4100
rect 13449 4097 13461 4131
rect 13495 4128 13507 4131
rect 13538 4128 13544 4140
rect 13495 4100 13544 4128
rect 13495 4097 13507 4100
rect 13449 4091 13507 4097
rect 13538 4088 13544 4100
rect 13596 4128 13602 4140
rect 13722 4128 13728 4140
rect 13596 4100 13728 4128
rect 13596 4088 13602 4100
rect 13722 4088 13728 4100
rect 13780 4088 13786 4140
rect 13814 4088 13820 4140
rect 13872 4128 13878 4140
rect 13909 4131 13967 4137
rect 13909 4128 13921 4131
rect 13872 4100 13921 4128
rect 13872 4088 13878 4100
rect 13909 4097 13921 4100
rect 13955 4097 13967 4131
rect 14918 4128 14924 4140
rect 14879 4100 14924 4128
rect 13909 4091 13967 4097
rect 14918 4088 14924 4100
rect 14976 4088 14982 4140
rect 15381 4131 15439 4137
rect 15381 4097 15393 4131
rect 15427 4097 15439 4131
rect 16850 4128 16856 4140
rect 16763 4100 16856 4128
rect 15381 4091 15439 4097
rect 15396 4060 15424 4091
rect 16850 4088 16856 4100
rect 16908 4088 16914 4140
rect 16945 4131 17003 4137
rect 16945 4097 16957 4131
rect 16991 4097 17003 4131
rect 16945 4091 17003 4097
rect 13372 4032 15424 4060
rect 16574 4020 16580 4072
rect 16632 4060 16638 4072
rect 16960 4060 16988 4091
rect 17034 4088 17040 4140
rect 17092 4128 17098 4140
rect 17221 4131 17279 4137
rect 17221 4128 17233 4131
rect 17092 4100 17233 4128
rect 17092 4088 17098 4100
rect 17221 4097 17233 4100
rect 17267 4128 17279 4131
rect 17862 4128 17868 4140
rect 17267 4100 17868 4128
rect 17267 4097 17279 4100
rect 17221 4091 17279 4097
rect 17862 4088 17868 4100
rect 17920 4088 17926 4140
rect 18230 4088 18236 4140
rect 18288 4128 18294 4140
rect 18325 4131 18383 4137
rect 18325 4128 18337 4131
rect 18288 4100 18337 4128
rect 18288 4088 18294 4100
rect 18325 4097 18337 4100
rect 18371 4097 18383 4131
rect 18325 4091 18383 4097
rect 18969 4131 19027 4137
rect 18969 4097 18981 4131
rect 19015 4128 19027 4131
rect 19015 4100 19288 4128
rect 19015 4097 19027 4100
rect 18969 4091 19027 4097
rect 18690 4060 18696 4072
rect 16632 4032 16988 4060
rect 17052 4032 18696 4060
rect 16632 4020 16638 4032
rect 7650 3992 7656 4004
rect 5592 3964 7512 3992
rect 7611 3964 7656 3992
rect 5592 3952 5598 3964
rect 7650 3952 7656 3964
rect 7708 3952 7714 4004
rect 7742 3952 7748 4004
rect 7800 3992 7806 4004
rect 9861 3995 9919 4001
rect 7800 3964 8340 3992
rect 7800 3952 7806 3964
rect 2130 3884 2136 3936
rect 2188 3924 2194 3936
rect 4341 3927 4399 3933
rect 4341 3924 4353 3927
rect 2188 3896 4353 3924
rect 2188 3884 2194 3896
rect 4341 3893 4353 3896
rect 4387 3924 4399 3927
rect 4614 3924 4620 3936
rect 4387 3896 4620 3924
rect 4387 3893 4399 3896
rect 4341 3887 4399 3893
rect 4614 3884 4620 3896
rect 4672 3884 4678 3936
rect 6362 3924 6368 3936
rect 6323 3896 6368 3924
rect 6362 3884 6368 3896
rect 6420 3884 6426 3936
rect 6546 3884 6552 3936
rect 6604 3924 6610 3936
rect 7558 3924 7564 3936
rect 6604 3896 7564 3924
rect 6604 3884 6610 3896
rect 7558 3884 7564 3896
rect 7616 3884 7622 3936
rect 8202 3924 8208 3936
rect 8163 3896 8208 3924
rect 8202 3884 8208 3896
rect 8260 3884 8266 3936
rect 8312 3924 8340 3964
rect 9861 3961 9873 3995
rect 9907 3992 9919 3995
rect 10962 3992 10968 4004
rect 9907 3964 10968 3992
rect 9907 3961 9919 3964
rect 9861 3955 9919 3961
rect 10962 3952 10968 3964
rect 11020 3952 11026 4004
rect 14737 3995 14795 4001
rect 14737 3992 14749 3995
rect 13464 3964 14749 3992
rect 11238 3924 11244 3936
rect 8312 3896 11244 3924
rect 11238 3884 11244 3896
rect 11296 3884 11302 3936
rect 13078 3884 13084 3936
rect 13136 3924 13142 3936
rect 13464 3924 13492 3964
rect 14737 3961 14749 3964
rect 14783 3961 14795 3995
rect 14737 3955 14795 3961
rect 15378 3952 15384 4004
rect 15436 3992 15442 4004
rect 15565 3995 15623 4001
rect 15565 3992 15577 3995
rect 15436 3964 15577 3992
rect 15436 3952 15442 3964
rect 15565 3961 15577 3964
rect 15611 3992 15623 3995
rect 17052 3992 17080 4032
rect 18690 4020 18696 4032
rect 18748 4020 18754 4072
rect 15611 3964 17080 3992
rect 15611 3961 15623 3964
rect 15565 3955 15623 3961
rect 17586 3952 17592 4004
rect 17644 3992 17650 4004
rect 17681 3995 17739 4001
rect 17681 3992 17693 3995
rect 17644 3964 17693 3992
rect 17644 3952 17650 3964
rect 17681 3961 17693 3964
rect 17727 3961 17739 3995
rect 19260 3992 19288 4100
rect 19334 4088 19340 4140
rect 19392 4128 19398 4140
rect 19613 4131 19671 4137
rect 19613 4128 19625 4131
rect 19392 4100 19625 4128
rect 19392 4088 19398 4100
rect 19613 4097 19625 4100
rect 19659 4097 19671 4131
rect 19613 4091 19671 4097
rect 19978 4088 19984 4140
rect 20036 4128 20042 4140
rect 20257 4131 20315 4137
rect 20257 4128 20269 4131
rect 20036 4100 20269 4128
rect 20036 4088 20042 4100
rect 20257 4097 20269 4100
rect 20303 4097 20315 4131
rect 20530 4128 20536 4140
rect 20491 4100 20536 4128
rect 20257 4091 20315 4097
rect 20530 4088 20536 4100
rect 20588 4088 20594 4140
rect 20806 4088 20812 4140
rect 20864 4128 20870 4140
rect 20901 4131 20959 4137
rect 20901 4128 20913 4131
rect 20864 4100 20913 4128
rect 20864 4088 20870 4100
rect 20901 4097 20913 4100
rect 20947 4097 20959 4131
rect 20901 4091 20959 4097
rect 21082 4088 21088 4140
rect 21140 4128 21146 4140
rect 21269 4131 21327 4137
rect 21269 4128 21281 4131
rect 21140 4100 21281 4128
rect 21140 4088 21146 4100
rect 21269 4097 21281 4100
rect 21315 4097 21327 4131
rect 21269 4091 21327 4097
rect 22646 4088 22652 4140
rect 22704 4128 22710 4140
rect 23385 4131 23443 4137
rect 23385 4128 23397 4131
rect 22704 4100 23397 4128
rect 22704 4088 22710 4100
rect 23385 4097 23397 4100
rect 23431 4097 23443 4131
rect 23385 4091 23443 4097
rect 25961 4131 26019 4137
rect 25961 4097 25973 4131
rect 26007 4128 26019 4131
rect 26050 4128 26056 4140
rect 26007 4100 26056 4128
rect 26007 4097 26019 4100
rect 25961 4091 26019 4097
rect 20622 4020 20628 4072
rect 20680 4060 20686 4072
rect 20993 4063 21051 4069
rect 20993 4060 21005 4063
rect 20680 4032 21005 4060
rect 20680 4020 20686 4032
rect 20993 4029 21005 4032
rect 21039 4029 21051 4063
rect 20993 4023 21051 4029
rect 20898 3992 20904 4004
rect 19260 3964 20904 3992
rect 17681 3955 17739 3961
rect 20640 3936 20668 3964
rect 20898 3952 20904 3964
rect 20956 3952 20962 4004
rect 13136 3896 13492 3924
rect 13136 3884 13142 3896
rect 13630 3884 13636 3936
rect 13688 3924 13694 3936
rect 14090 3924 14096 3936
rect 13688 3896 14096 3924
rect 13688 3884 13694 3896
rect 14090 3884 14096 3896
rect 14148 3884 14154 3936
rect 16666 3884 16672 3936
rect 16724 3924 16730 3936
rect 17954 3924 17960 3936
rect 16724 3896 17960 3924
rect 16724 3884 16730 3896
rect 17954 3884 17960 3896
rect 18012 3884 18018 3936
rect 18506 3924 18512 3936
rect 18467 3896 18512 3924
rect 18506 3884 18512 3896
rect 18564 3884 18570 3936
rect 19153 3927 19211 3933
rect 19153 3893 19165 3927
rect 19199 3924 19211 3927
rect 19426 3924 19432 3936
rect 19199 3896 19432 3924
rect 19199 3893 19211 3896
rect 19153 3887 19211 3893
rect 19426 3884 19432 3896
rect 19484 3884 19490 3936
rect 19797 3927 19855 3933
rect 19797 3893 19809 3927
rect 19843 3924 19855 3927
rect 19978 3924 19984 3936
rect 19843 3896 19984 3924
rect 19843 3893 19855 3896
rect 19797 3887 19855 3893
rect 19978 3884 19984 3896
rect 20036 3884 20042 3936
rect 20622 3884 20628 3936
rect 20680 3884 20686 3936
rect 25976 3924 26004 4091
rect 26050 4088 26056 4100
rect 26108 4088 26114 4140
rect 26234 4088 26240 4140
rect 26292 4128 26298 4140
rect 26973 4131 27031 4137
rect 26973 4128 26985 4131
rect 26292 4100 26985 4128
rect 26292 4088 26298 4100
rect 26973 4097 26985 4100
rect 27019 4128 27031 4131
rect 27080 4128 27108 4168
rect 27246 4137 27252 4140
rect 27240 4128 27252 4137
rect 27019 4100 27108 4128
rect 27207 4100 27252 4128
rect 27019 4097 27031 4100
rect 26973 4091 27031 4097
rect 27240 4091 27252 4100
rect 27246 4088 27252 4091
rect 27304 4088 27310 4140
rect 27356 4128 27384 4168
rect 28534 4156 28540 4208
rect 28592 4196 28598 4208
rect 28813 4199 28871 4205
rect 28813 4196 28825 4199
rect 28592 4168 28825 4196
rect 28592 4156 28598 4168
rect 28813 4165 28825 4168
rect 28859 4165 28871 4199
rect 28813 4159 28871 4165
rect 28997 4199 29055 4205
rect 28997 4165 29009 4199
rect 29043 4196 29055 4199
rect 30558 4196 30564 4208
rect 29043 4168 30564 4196
rect 29043 4165 29055 4168
rect 28997 4159 29055 4165
rect 30558 4156 30564 4168
rect 30616 4196 30622 4208
rect 31404 4196 31432 4227
rect 32122 4224 32128 4276
rect 32180 4264 32186 4276
rect 33689 4267 33747 4273
rect 33689 4264 33701 4267
rect 32180 4236 33701 4264
rect 32180 4224 32186 4236
rect 33689 4233 33701 4236
rect 33735 4264 33747 4267
rect 35989 4267 36047 4273
rect 33735 4236 34652 4264
rect 33735 4233 33747 4236
rect 33689 4227 33747 4233
rect 34514 4196 34520 4208
rect 30616 4168 31432 4196
rect 34256 4168 34520 4196
rect 30616 4156 30622 4168
rect 30282 4137 30288 4140
rect 30276 4128 30288 4137
rect 27356 4100 30052 4128
rect 30243 4100 30288 4128
rect 30024 4069 30052 4100
rect 30276 4091 30288 4100
rect 30282 4088 30288 4091
rect 30340 4088 30346 4140
rect 34256 4137 34284 4168
rect 34514 4156 34520 4168
rect 34572 4156 34578 4208
rect 34624 4196 34652 4236
rect 35989 4233 36001 4267
rect 36035 4264 36047 4267
rect 36906 4264 36912 4276
rect 36035 4236 36912 4264
rect 36035 4233 36047 4236
rect 35989 4227 36047 4233
rect 36906 4224 36912 4236
rect 36964 4224 36970 4276
rect 34624 4168 35006 4196
rect 34241 4131 34299 4137
rect 34241 4097 34253 4131
rect 34287 4097 34299 4131
rect 34241 4091 34299 4097
rect 57974 4088 57980 4140
rect 58032 4128 58038 4140
rect 59817 4131 59875 4137
rect 59817 4128 59829 4131
rect 58032 4100 59829 4128
rect 58032 4088 58038 4100
rect 59817 4097 59829 4100
rect 59863 4097 59875 4131
rect 59817 4091 59875 4097
rect 30009 4063 30067 4069
rect 30009 4029 30021 4063
rect 30055 4029 30067 4063
rect 30009 4023 30067 4029
rect 34517 4063 34575 4069
rect 34517 4029 34529 4063
rect 34563 4060 34575 4063
rect 34606 4060 34612 4072
rect 34563 4032 34612 4060
rect 34563 4029 34575 4032
rect 34517 4023 34575 4029
rect 34606 4020 34612 4032
rect 34664 4020 34670 4072
rect 59170 4020 59176 4072
rect 59228 4060 59234 4072
rect 61105 4063 61163 4069
rect 61105 4060 61117 4063
rect 59228 4032 61117 4060
rect 59228 4020 59234 4032
rect 61105 4029 61117 4032
rect 61151 4029 61163 4063
rect 61105 4023 61163 4029
rect 57514 3952 57520 4004
rect 57572 3992 57578 4004
rect 58529 3995 58587 4001
rect 58529 3992 58541 3995
rect 57572 3964 58541 3992
rect 57572 3952 57578 3964
rect 58529 3961 58541 3964
rect 58575 3961 58587 3995
rect 58529 3955 58587 3961
rect 58618 3952 58624 4004
rect 58676 3992 58682 4004
rect 60461 3995 60519 4001
rect 60461 3992 60473 3995
rect 58676 3964 60473 3992
rect 58676 3952 58682 3964
rect 60461 3961 60473 3964
rect 60507 3961 60519 3995
rect 60461 3955 60519 3961
rect 28353 3927 28411 3933
rect 28353 3924 28365 3927
rect 25976 3896 28365 3924
rect 28353 3893 28365 3896
rect 28399 3924 28411 3927
rect 30006 3924 30012 3936
rect 28399 3896 30012 3924
rect 28399 3893 28411 3896
rect 28353 3887 28411 3893
rect 30006 3884 30012 3896
rect 30064 3884 30070 3936
rect 56134 3884 56140 3936
rect 56192 3924 56198 3936
rect 56229 3927 56287 3933
rect 56229 3924 56241 3927
rect 56192 3896 56241 3924
rect 56192 3884 56198 3896
rect 56229 3893 56241 3896
rect 56275 3893 56287 3927
rect 56229 3887 56287 3893
rect 56318 3884 56324 3936
rect 56376 3924 56382 3936
rect 56873 3927 56931 3933
rect 56873 3924 56885 3927
rect 56376 3896 56885 3924
rect 56376 3884 56382 3896
rect 56873 3893 56885 3896
rect 56919 3893 56931 3927
rect 56873 3887 56931 3893
rect 56962 3884 56968 3936
rect 57020 3924 57026 3936
rect 57885 3927 57943 3933
rect 57885 3924 57897 3927
rect 57020 3896 57897 3924
rect 57020 3884 57026 3896
rect 57885 3893 57897 3896
rect 57931 3893 57943 3927
rect 57885 3887 57943 3893
rect 58066 3884 58072 3936
rect 58124 3924 58130 3936
rect 59173 3927 59231 3933
rect 59173 3924 59185 3927
rect 58124 3896 59185 3924
rect 58124 3884 58130 3896
rect 59173 3893 59185 3896
rect 59219 3893 59231 3927
rect 67634 3924 67640 3936
rect 67595 3896 67640 3924
rect 59173 3887 59231 3893
rect 67634 3884 67640 3896
rect 67692 3884 67698 3936
rect 1104 3834 68816 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 65654 3834
rect 65706 3782 65718 3834
rect 65770 3782 65782 3834
rect 65834 3782 65846 3834
rect 65898 3782 65910 3834
rect 65962 3782 68816 3834
rect 1104 3760 68816 3782
rect 2222 3720 2228 3732
rect 2183 3692 2228 3720
rect 2222 3680 2228 3692
rect 2280 3680 2286 3732
rect 2498 3680 2504 3732
rect 2556 3720 2562 3732
rect 2777 3723 2835 3729
rect 2777 3720 2789 3723
rect 2556 3692 2789 3720
rect 2556 3680 2562 3692
rect 2777 3689 2789 3692
rect 2823 3689 2835 3723
rect 2777 3683 2835 3689
rect 4709 3723 4767 3729
rect 4709 3689 4721 3723
rect 4755 3720 4767 3723
rect 4755 3692 6960 3720
rect 4755 3689 4767 3692
rect 4709 3683 4767 3689
rect 6932 3584 6960 3692
rect 8202 3680 8208 3732
rect 8260 3720 8266 3732
rect 11330 3720 11336 3732
rect 8260 3692 11336 3720
rect 8260 3680 8266 3692
rect 11330 3680 11336 3692
rect 11388 3680 11394 3732
rect 11606 3720 11612 3732
rect 11567 3692 11612 3720
rect 11606 3680 11612 3692
rect 11664 3680 11670 3732
rect 12434 3680 12440 3732
rect 12492 3720 12498 3732
rect 15841 3723 15899 3729
rect 12492 3692 15792 3720
rect 12492 3680 12498 3692
rect 7193 3655 7251 3661
rect 7193 3621 7205 3655
rect 7239 3652 7251 3655
rect 10965 3655 11023 3661
rect 7239 3624 9352 3652
rect 7239 3621 7251 3624
rect 7193 3615 7251 3621
rect 6932 3556 7052 3584
rect 6282 3519 6340 3525
rect 6282 3485 6294 3519
rect 6328 3485 6340 3519
rect 6282 3479 6340 3485
rect 6549 3519 6607 3525
rect 6549 3485 6561 3519
rect 6595 3516 6607 3519
rect 6914 3516 6920 3528
rect 6595 3488 6920 3516
rect 6595 3485 6607 3488
rect 6549 3479 6607 3485
rect 3418 3408 3424 3460
rect 3476 3448 3482 3460
rect 6288 3448 6316 3479
rect 6362 3448 6368 3460
rect 3476 3420 6224 3448
rect 6288 3420 6368 3448
rect 3476 3408 3482 3420
rect 4154 3380 4160 3392
rect 4115 3352 4160 3380
rect 4154 3340 4160 3352
rect 4212 3340 4218 3392
rect 5169 3383 5227 3389
rect 5169 3349 5181 3383
rect 5215 3380 5227 3383
rect 5626 3380 5632 3392
rect 5215 3352 5632 3380
rect 5215 3349 5227 3352
rect 5169 3343 5227 3349
rect 5626 3340 5632 3352
rect 5684 3340 5690 3392
rect 6196 3380 6224 3420
rect 6362 3408 6368 3420
rect 6420 3408 6426 3460
rect 6564 3380 6592 3479
rect 6914 3476 6920 3488
rect 6972 3476 6978 3528
rect 7024 3525 7052 3556
rect 7558 3544 7564 3596
rect 7616 3584 7622 3596
rect 7616 3556 8064 3584
rect 7616 3544 7622 3556
rect 7009 3519 7067 3525
rect 7009 3485 7021 3519
rect 7055 3516 7067 3519
rect 7742 3516 7748 3528
rect 7055 3488 7748 3516
rect 7055 3485 7067 3488
rect 7009 3479 7067 3485
rect 7742 3476 7748 3488
rect 7800 3476 7806 3528
rect 7834 3476 7840 3528
rect 7892 3516 7898 3528
rect 8036 3525 8064 3556
rect 8021 3519 8079 3525
rect 7892 3488 7937 3516
rect 7892 3476 7898 3488
rect 8021 3485 8033 3519
rect 8067 3485 8079 3519
rect 8021 3479 8079 3485
rect 9030 3476 9036 3528
rect 9088 3516 9094 3528
rect 9125 3519 9183 3525
rect 9125 3516 9137 3519
rect 9088 3488 9137 3516
rect 9088 3476 9094 3488
rect 9125 3485 9137 3488
rect 9171 3485 9183 3519
rect 9125 3479 9183 3485
rect 6730 3408 6736 3460
rect 6788 3448 6794 3460
rect 8570 3448 8576 3460
rect 6788 3420 8576 3448
rect 6788 3408 6794 3420
rect 8570 3408 8576 3420
rect 8628 3408 8634 3460
rect 9324 3448 9352 3624
rect 10965 3621 10977 3655
rect 11011 3621 11023 3655
rect 10965 3615 11023 3621
rect 11793 3655 11851 3661
rect 11793 3621 11805 3655
rect 11839 3652 11851 3655
rect 13446 3652 13452 3664
rect 11839 3624 13452 3652
rect 11839 3621 11851 3624
rect 11793 3615 11851 3621
rect 10980 3584 11008 3615
rect 13446 3612 13452 3624
rect 13504 3612 13510 3664
rect 15102 3652 15108 3664
rect 15063 3624 15108 3652
rect 15102 3612 15108 3624
rect 15160 3612 15166 3664
rect 15764 3652 15792 3692
rect 15841 3689 15853 3723
rect 15887 3720 15899 3723
rect 18230 3720 18236 3732
rect 15887 3692 18236 3720
rect 15887 3689 15899 3692
rect 15841 3683 15899 3689
rect 18230 3680 18236 3692
rect 18288 3720 18294 3732
rect 18414 3720 18420 3732
rect 18288 3692 18420 3720
rect 18288 3680 18294 3692
rect 18414 3680 18420 3692
rect 18472 3680 18478 3732
rect 18690 3680 18696 3732
rect 18748 3720 18754 3732
rect 22370 3720 22376 3732
rect 18748 3692 22376 3720
rect 18748 3680 18754 3692
rect 22370 3680 22376 3692
rect 22428 3680 22434 3732
rect 57790 3680 57796 3732
rect 57848 3720 57854 3732
rect 58066 3720 58072 3732
rect 57848 3692 58072 3720
rect 57848 3680 57854 3692
rect 58066 3680 58072 3692
rect 58124 3680 58130 3732
rect 18138 3652 18144 3664
rect 15764 3624 18144 3652
rect 18138 3612 18144 3624
rect 18196 3612 18202 3664
rect 18506 3612 18512 3664
rect 18564 3652 18570 3664
rect 19981 3655 20039 3661
rect 18564 3624 19564 3652
rect 18564 3612 18570 3624
rect 11054 3584 11060 3596
rect 10967 3556 11060 3584
rect 11054 3544 11060 3556
rect 11112 3584 11118 3596
rect 12805 3587 12863 3593
rect 11112 3556 12434 3584
rect 11112 3544 11118 3556
rect 9582 3516 9588 3528
rect 9543 3488 9588 3516
rect 9582 3476 9588 3488
rect 9640 3476 9646 3528
rect 9858 3525 9864 3528
rect 9852 3516 9864 3525
rect 9819 3488 9864 3516
rect 9852 3479 9864 3488
rect 9858 3476 9864 3479
rect 9916 3476 9922 3528
rect 10686 3476 10692 3528
rect 10744 3516 10750 3528
rect 10870 3516 10876 3528
rect 10744 3488 10876 3516
rect 10744 3476 10750 3488
rect 10870 3476 10876 3488
rect 10928 3476 10934 3528
rect 11606 3476 11612 3528
rect 11664 3516 11670 3528
rect 11882 3516 11888 3528
rect 11664 3488 11888 3516
rect 11664 3476 11670 3488
rect 11882 3476 11888 3488
rect 11940 3476 11946 3528
rect 12406 3516 12434 3556
rect 12805 3553 12817 3587
rect 12851 3584 12863 3587
rect 16574 3584 16580 3596
rect 12851 3556 16580 3584
rect 12851 3553 12863 3556
rect 12805 3547 12863 3553
rect 16574 3544 16580 3556
rect 16632 3584 16638 3596
rect 19426 3584 19432 3596
rect 16632 3556 16712 3584
rect 19387 3556 19432 3584
rect 16632 3544 16638 3556
rect 12986 3516 12992 3528
rect 12406 3488 12992 3516
rect 12986 3476 12992 3488
rect 13044 3476 13050 3528
rect 13354 3476 13360 3528
rect 13412 3516 13418 3528
rect 13541 3519 13599 3525
rect 13541 3516 13553 3519
rect 13412 3488 13553 3516
rect 13412 3476 13418 3488
rect 13541 3485 13553 3488
rect 13587 3485 13599 3519
rect 13541 3479 13599 3485
rect 14553 3519 14611 3525
rect 14553 3485 14565 3519
rect 14599 3485 14611 3519
rect 14553 3479 14611 3485
rect 15289 3519 15347 3525
rect 15289 3485 15301 3519
rect 15335 3516 15347 3519
rect 15378 3516 15384 3528
rect 15335 3488 15384 3516
rect 15335 3485 15347 3488
rect 15289 3479 15347 3485
rect 11425 3451 11483 3457
rect 11425 3448 11437 3451
rect 9324 3420 11437 3448
rect 11425 3417 11437 3420
rect 11471 3417 11483 3451
rect 12618 3448 12624 3460
rect 12579 3420 12624 3448
rect 11425 3411 11483 3417
rect 12618 3408 12624 3420
rect 12676 3448 12682 3460
rect 13446 3448 13452 3460
rect 12676 3420 13452 3448
rect 12676 3408 12682 3420
rect 13446 3408 13452 3420
rect 13504 3408 13510 3460
rect 14561 3448 14589 3479
rect 15378 3476 15384 3488
rect 15436 3516 15442 3528
rect 15838 3516 15844 3528
rect 15436 3488 15844 3516
rect 15436 3476 15442 3488
rect 15838 3476 15844 3488
rect 15896 3476 15902 3528
rect 16298 3516 16304 3528
rect 16259 3488 16304 3516
rect 16298 3476 16304 3488
rect 16356 3476 16362 3528
rect 16684 3525 16712 3556
rect 19426 3544 19432 3556
rect 19484 3544 19490 3596
rect 19536 3593 19564 3624
rect 19981 3621 19993 3655
rect 20027 3652 20039 3655
rect 20070 3652 20076 3664
rect 20027 3624 20076 3652
rect 20027 3621 20039 3624
rect 19981 3615 20039 3621
rect 20070 3612 20076 3624
rect 20128 3612 20134 3664
rect 41138 3612 41144 3664
rect 41196 3652 41202 3664
rect 41785 3655 41843 3661
rect 41785 3652 41797 3655
rect 41196 3624 41797 3652
rect 41196 3612 41202 3624
rect 41785 3621 41797 3624
rect 41831 3621 41843 3655
rect 41785 3615 41843 3621
rect 56502 3612 56508 3664
rect 56560 3652 56566 3664
rect 57885 3655 57943 3661
rect 57885 3652 57897 3655
rect 56560 3624 57897 3652
rect 56560 3612 56566 3624
rect 57885 3621 57897 3624
rect 57931 3621 57943 3655
rect 57885 3615 57943 3621
rect 58342 3612 58348 3664
rect 58400 3652 58406 3664
rect 61105 3655 61163 3661
rect 61105 3652 61117 3655
rect 58400 3624 61117 3652
rect 58400 3612 58406 3624
rect 61105 3621 61117 3624
rect 61151 3621 61163 3655
rect 61105 3615 61163 3621
rect 19521 3587 19579 3593
rect 19521 3553 19533 3587
rect 19567 3553 19579 3587
rect 19521 3547 19579 3553
rect 55766 3544 55772 3596
rect 55824 3584 55830 3596
rect 56597 3587 56655 3593
rect 56597 3584 56609 3587
rect 55824 3556 56609 3584
rect 55824 3544 55830 3556
rect 56597 3553 56609 3556
rect 56643 3553 56655 3587
rect 56597 3547 56655 3553
rect 56778 3544 56784 3596
rect 56836 3584 56842 3596
rect 58529 3587 58587 3593
rect 58529 3584 58541 3587
rect 56836 3556 58541 3584
rect 56836 3544 56842 3556
rect 58529 3553 58541 3556
rect 58575 3553 58587 3587
rect 58529 3547 58587 3553
rect 58986 3544 58992 3596
rect 59044 3584 59050 3596
rect 61749 3587 61807 3593
rect 61749 3584 61761 3587
rect 59044 3556 61761 3584
rect 59044 3544 59050 3556
rect 61749 3553 61761 3556
rect 61795 3553 61807 3587
rect 61749 3547 61807 3553
rect 16485 3519 16543 3525
rect 16485 3485 16497 3519
rect 16531 3485 16543 3519
rect 16485 3479 16543 3485
rect 16669 3519 16727 3525
rect 16669 3485 16681 3519
rect 16715 3485 16727 3519
rect 16850 3516 16856 3528
rect 16811 3488 16856 3516
rect 16669 3479 16727 3485
rect 15746 3448 15752 3460
rect 14561 3420 15752 3448
rect 15746 3408 15752 3420
rect 15804 3408 15810 3460
rect 16500 3448 16528 3479
rect 16850 3476 16856 3488
rect 16908 3516 16914 3528
rect 17034 3516 17040 3528
rect 16908 3488 17040 3516
rect 16908 3476 16914 3488
rect 17034 3476 17040 3488
rect 17092 3476 17098 3528
rect 17129 3519 17187 3525
rect 17129 3485 17141 3519
rect 17175 3516 17187 3519
rect 17586 3516 17592 3528
rect 17175 3488 17592 3516
rect 17175 3485 17187 3488
rect 17129 3479 17187 3485
rect 17586 3476 17592 3488
rect 17644 3476 17650 3528
rect 18049 3519 18107 3525
rect 18049 3485 18061 3519
rect 18095 3485 18107 3519
rect 18049 3479 18107 3485
rect 18693 3519 18751 3525
rect 18693 3485 18705 3519
rect 18739 3516 18751 3519
rect 20162 3516 20168 3528
rect 18739 3488 20168 3516
rect 18739 3485 18751 3488
rect 18693 3479 18751 3485
rect 16758 3448 16764 3460
rect 16500 3420 16764 3448
rect 16758 3408 16764 3420
rect 16816 3408 16822 3460
rect 18064 3448 18092 3479
rect 20162 3476 20168 3488
rect 20220 3476 20226 3528
rect 20438 3476 20444 3528
rect 20496 3516 20502 3528
rect 20533 3519 20591 3525
rect 20533 3516 20545 3519
rect 20496 3488 20545 3516
rect 20496 3476 20502 3488
rect 20533 3485 20545 3488
rect 20579 3485 20591 3519
rect 20533 3479 20591 3485
rect 21542 3476 21548 3528
rect 21600 3516 21606 3528
rect 21637 3519 21695 3525
rect 21637 3516 21649 3519
rect 21600 3488 21649 3516
rect 21600 3476 21606 3488
rect 21637 3485 21649 3488
rect 21683 3485 21695 3519
rect 21637 3479 21695 3485
rect 22370 3476 22376 3528
rect 22428 3516 22434 3528
rect 22465 3519 22523 3525
rect 22465 3516 22477 3519
rect 22428 3488 22477 3516
rect 22428 3476 22434 3488
rect 22465 3485 22477 3488
rect 22511 3485 22523 3519
rect 22465 3479 22523 3485
rect 23474 3476 23480 3528
rect 23532 3516 23538 3528
rect 23569 3519 23627 3525
rect 23569 3516 23581 3519
rect 23532 3488 23581 3516
rect 23532 3476 23538 3488
rect 23569 3485 23581 3488
rect 23615 3485 23627 3519
rect 23569 3479 23627 3485
rect 24302 3476 24308 3528
rect 24360 3516 24366 3528
rect 24397 3519 24455 3525
rect 24397 3516 24409 3519
rect 24360 3488 24409 3516
rect 24360 3476 24366 3488
rect 24397 3485 24409 3488
rect 24443 3485 24455 3519
rect 24397 3479 24455 3485
rect 25130 3476 25136 3528
rect 25188 3516 25194 3528
rect 25225 3519 25283 3525
rect 25225 3516 25237 3519
rect 25188 3488 25237 3516
rect 25188 3476 25194 3488
rect 25225 3485 25237 3488
rect 25271 3485 25283 3519
rect 25225 3479 25283 3485
rect 25958 3476 25964 3528
rect 26016 3516 26022 3528
rect 26053 3519 26111 3525
rect 26053 3516 26065 3519
rect 26016 3488 26065 3516
rect 26016 3476 26022 3488
rect 26053 3485 26065 3488
rect 26099 3485 26111 3519
rect 26053 3479 26111 3485
rect 26786 3476 26792 3528
rect 26844 3516 26850 3528
rect 26881 3519 26939 3525
rect 26881 3516 26893 3519
rect 26844 3488 26893 3516
rect 26844 3476 26850 3488
rect 26881 3485 26893 3488
rect 26927 3485 26939 3519
rect 26881 3479 26939 3485
rect 27614 3476 27620 3528
rect 27672 3516 27678 3528
rect 27709 3519 27767 3525
rect 27709 3516 27721 3519
rect 27672 3488 27721 3516
rect 27672 3476 27678 3488
rect 27709 3485 27721 3488
rect 27755 3485 27767 3519
rect 27709 3479 27767 3485
rect 28718 3476 28724 3528
rect 28776 3516 28782 3528
rect 28813 3519 28871 3525
rect 28813 3516 28825 3519
rect 28776 3488 28825 3516
rect 28776 3476 28782 3488
rect 28813 3485 28825 3488
rect 28859 3485 28871 3519
rect 28813 3479 28871 3485
rect 29822 3476 29828 3528
rect 29880 3516 29886 3528
rect 29917 3519 29975 3525
rect 29917 3516 29929 3519
rect 29880 3488 29929 3516
rect 29880 3476 29886 3488
rect 29917 3485 29929 3488
rect 29963 3485 29975 3519
rect 29917 3479 29975 3485
rect 30650 3476 30656 3528
rect 30708 3516 30714 3528
rect 30745 3519 30803 3525
rect 30745 3516 30757 3519
rect 30708 3488 30757 3516
rect 30708 3476 30714 3488
rect 30745 3485 30757 3488
rect 30791 3485 30803 3519
rect 30745 3479 30803 3485
rect 31478 3476 31484 3528
rect 31536 3516 31542 3528
rect 31573 3519 31631 3525
rect 31573 3516 31585 3519
rect 31536 3488 31585 3516
rect 31536 3476 31542 3488
rect 31573 3485 31585 3488
rect 31619 3485 31631 3519
rect 31573 3479 31631 3485
rect 32306 3476 32312 3528
rect 32364 3516 32370 3528
rect 32401 3519 32459 3525
rect 32401 3516 32413 3519
rect 32364 3488 32413 3516
rect 32364 3476 32370 3488
rect 32401 3485 32413 3488
rect 32447 3485 32459 3519
rect 32401 3479 32459 3485
rect 33134 3476 33140 3528
rect 33192 3516 33198 3528
rect 33229 3519 33287 3525
rect 33229 3516 33241 3519
rect 33192 3488 33241 3516
rect 33192 3476 33198 3488
rect 33229 3485 33241 3488
rect 33275 3485 33287 3519
rect 33229 3479 33287 3485
rect 39206 3476 39212 3528
rect 39264 3516 39270 3528
rect 39853 3519 39911 3525
rect 39853 3516 39865 3519
rect 39264 3488 39865 3516
rect 39264 3476 39270 3488
rect 39853 3485 39865 3488
rect 39899 3485 39911 3519
rect 39853 3479 39911 3485
rect 40034 3476 40040 3528
rect 40092 3516 40098 3528
rect 40497 3519 40555 3525
rect 40497 3516 40509 3519
rect 40092 3488 40509 3516
rect 40092 3476 40098 3488
rect 40497 3485 40509 3488
rect 40543 3485 40555 3519
rect 40497 3479 40555 3485
rect 40862 3476 40868 3528
rect 40920 3516 40926 3528
rect 41141 3519 41199 3525
rect 41141 3516 41153 3519
rect 40920 3488 41153 3516
rect 40920 3476 40926 3488
rect 41141 3485 41153 3488
rect 41187 3485 41199 3519
rect 41141 3479 41199 3485
rect 42518 3476 42524 3528
rect 42576 3516 42582 3528
rect 42613 3519 42671 3525
rect 42613 3516 42625 3519
rect 42576 3488 42625 3516
rect 42576 3476 42582 3488
rect 42613 3485 42625 3488
rect 42659 3485 42671 3519
rect 42613 3479 42671 3485
rect 43070 3476 43076 3528
rect 43128 3516 43134 3528
rect 43257 3519 43315 3525
rect 43257 3516 43269 3519
rect 43128 3488 43269 3516
rect 43128 3476 43134 3488
rect 43257 3485 43269 3488
rect 43303 3485 43315 3519
rect 43257 3479 43315 3485
rect 45002 3476 45008 3528
rect 45060 3516 45066 3528
rect 45097 3519 45155 3525
rect 45097 3516 45109 3519
rect 45060 3488 45109 3516
rect 45060 3476 45066 3488
rect 45097 3485 45109 3488
rect 45143 3485 45155 3519
rect 45097 3479 45155 3485
rect 45278 3476 45284 3528
rect 45336 3516 45342 3528
rect 45741 3519 45799 3525
rect 45741 3516 45753 3519
rect 45336 3488 45753 3516
rect 45336 3476 45342 3488
rect 45741 3485 45753 3488
rect 45787 3485 45799 3519
rect 45741 3479 45799 3485
rect 46106 3476 46112 3528
rect 46164 3516 46170 3528
rect 46385 3519 46443 3525
rect 46385 3516 46397 3519
rect 46164 3488 46397 3516
rect 46164 3476 46170 3488
rect 46385 3485 46397 3488
rect 46431 3485 46443 3519
rect 46385 3479 46443 3485
rect 46934 3476 46940 3528
rect 46992 3516 46998 3528
rect 47029 3519 47087 3525
rect 47029 3516 47041 3519
rect 46992 3488 47041 3516
rect 46992 3476 46998 3488
rect 47029 3485 47041 3488
rect 47075 3485 47087 3519
rect 47029 3479 47087 3485
rect 47762 3476 47768 3528
rect 47820 3516 47826 3528
rect 47857 3519 47915 3525
rect 47857 3516 47869 3519
rect 47820 3488 47869 3516
rect 47820 3476 47826 3488
rect 47857 3485 47869 3488
rect 47903 3485 47915 3519
rect 47857 3479 47915 3485
rect 48866 3476 48872 3528
rect 48924 3516 48930 3528
rect 48961 3519 49019 3525
rect 48961 3516 48973 3519
rect 48924 3488 48973 3516
rect 48924 3476 48930 3488
rect 48961 3485 48973 3488
rect 49007 3485 49019 3519
rect 48961 3479 49019 3485
rect 50154 3476 50160 3528
rect 50212 3516 50218 3528
rect 50341 3519 50399 3525
rect 50341 3516 50353 3519
rect 50212 3488 50353 3516
rect 50212 3476 50218 3488
rect 50341 3485 50353 3488
rect 50387 3485 50399 3519
rect 50341 3479 50399 3485
rect 50798 3476 50804 3528
rect 50856 3516 50862 3528
rect 50985 3519 51043 3525
rect 50985 3516 50997 3519
rect 50856 3488 50997 3516
rect 50856 3476 50862 3488
rect 50985 3485 50997 3488
rect 51031 3485 51043 3519
rect 50985 3479 51043 3485
rect 51350 3476 51356 3528
rect 51408 3516 51414 3528
rect 51629 3519 51687 3525
rect 51629 3516 51641 3519
rect 51408 3488 51641 3516
rect 51408 3476 51414 3488
rect 51629 3485 51641 3488
rect 51675 3485 51687 3519
rect 51629 3479 51687 3485
rect 52730 3476 52736 3528
rect 52788 3516 52794 3528
rect 52825 3519 52883 3525
rect 52825 3516 52837 3519
rect 52788 3488 52837 3516
rect 52788 3476 52794 3488
rect 52825 3485 52837 3488
rect 52871 3485 52883 3519
rect 52825 3479 52883 3485
rect 53006 3476 53012 3528
rect 53064 3516 53070 3528
rect 53469 3519 53527 3525
rect 53469 3516 53481 3519
rect 53064 3488 53481 3516
rect 53064 3476 53070 3488
rect 53469 3485 53481 3488
rect 53515 3485 53527 3519
rect 53469 3479 53527 3485
rect 54662 3476 54668 3528
rect 54720 3516 54726 3528
rect 55309 3519 55367 3525
rect 55309 3516 55321 3519
rect 54720 3488 55321 3516
rect 54720 3476 54726 3488
rect 55309 3485 55321 3488
rect 55355 3485 55367 3519
rect 55309 3479 55367 3485
rect 55490 3476 55496 3528
rect 55548 3516 55554 3528
rect 55953 3519 56011 3525
rect 55953 3516 55965 3519
rect 55548 3488 55965 3516
rect 55548 3476 55554 3488
rect 55953 3485 55965 3488
rect 55999 3485 56011 3519
rect 55953 3479 56011 3485
rect 56226 3476 56232 3528
rect 56284 3516 56290 3528
rect 57241 3519 57299 3525
rect 57241 3516 57253 3519
rect 56284 3488 57253 3516
rect 56284 3476 56290 3488
rect 57241 3485 57253 3488
rect 57287 3485 57299 3519
rect 57241 3479 57299 3485
rect 57330 3476 57336 3528
rect 57388 3516 57394 3528
rect 59173 3519 59231 3525
rect 59173 3516 59185 3519
rect 57388 3488 59185 3516
rect 57388 3476 57394 3488
rect 59173 3485 59185 3488
rect 59219 3485 59231 3519
rect 60458 3516 60464 3528
rect 60419 3488 60464 3516
rect 59173 3479 59231 3485
rect 60458 3476 60464 3488
rect 60516 3476 60522 3528
rect 19426 3448 19432 3460
rect 18064 3420 19432 3448
rect 19426 3408 19432 3420
rect 19484 3408 19490 3460
rect 19978 3448 19984 3460
rect 19939 3420 19984 3448
rect 19978 3408 19984 3420
rect 20036 3408 20042 3460
rect 6196 3352 6592 3380
rect 7374 3340 7380 3392
rect 7432 3380 7438 3392
rect 7653 3383 7711 3389
rect 7653 3380 7665 3383
rect 7432 3352 7665 3380
rect 7432 3340 7438 3352
rect 7653 3349 7665 3352
rect 7699 3349 7711 3383
rect 7653 3343 7711 3349
rect 7742 3340 7748 3392
rect 7800 3380 7806 3392
rect 10686 3380 10692 3392
rect 7800 3352 10692 3380
rect 7800 3340 7806 3352
rect 10686 3340 10692 3352
rect 10744 3340 10750 3392
rect 11054 3340 11060 3392
rect 11112 3380 11118 3392
rect 11238 3380 11244 3392
rect 11112 3352 11244 3380
rect 11112 3340 11118 3352
rect 11238 3340 11244 3352
rect 11296 3340 11302 3392
rect 11635 3383 11693 3389
rect 11635 3349 11647 3383
rect 11681 3380 11693 3383
rect 12250 3380 12256 3392
rect 11681 3352 12256 3380
rect 11681 3349 11693 3352
rect 11635 3343 11693 3349
rect 12250 3340 12256 3352
rect 12308 3340 12314 3392
rect 13357 3383 13415 3389
rect 13357 3349 13369 3383
rect 13403 3380 13415 3383
rect 13630 3380 13636 3392
rect 13403 3352 13636 3380
rect 13403 3349 13415 3352
rect 13357 3343 13415 3349
rect 13630 3340 13636 3352
rect 13688 3340 13694 3392
rect 14182 3340 14188 3392
rect 14240 3380 14246 3392
rect 14369 3383 14427 3389
rect 14369 3380 14381 3383
rect 14240 3352 14381 3380
rect 14240 3340 14246 3352
rect 14369 3349 14381 3352
rect 14415 3349 14427 3383
rect 19242 3380 19248 3392
rect 19203 3352 19248 3380
rect 14369 3343 14427 3349
rect 19242 3340 19248 3352
rect 19300 3340 19306 3392
rect 1104 3290 68816 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 50294 3290
rect 50346 3238 50358 3290
rect 50410 3238 50422 3290
rect 50474 3238 50486 3290
rect 50538 3238 50550 3290
rect 50602 3238 68816 3290
rect 1104 3216 68816 3238
rect 7742 3176 7748 3188
rect 6564 3148 7748 3176
rect 4154 3000 4160 3052
rect 4212 3040 4218 3052
rect 5537 3043 5595 3049
rect 5537 3040 5549 3043
rect 4212 3012 5549 3040
rect 4212 3000 4218 3012
rect 5537 3009 5549 3012
rect 5583 3040 5595 3043
rect 6564 3040 6592 3148
rect 7742 3136 7748 3148
rect 7800 3136 7806 3188
rect 7834 3136 7840 3188
rect 7892 3176 7898 3188
rect 8481 3179 8539 3185
rect 8481 3176 8493 3179
rect 7892 3148 8493 3176
rect 7892 3136 7898 3148
rect 8481 3145 8493 3148
rect 8527 3145 8539 3179
rect 8481 3139 8539 3145
rect 8570 3136 8576 3188
rect 8628 3176 8634 3188
rect 10410 3176 10416 3188
rect 8628 3148 9720 3176
rect 10371 3148 10416 3176
rect 8628 3136 8634 3148
rect 9582 3108 9588 3120
rect 7116 3080 9588 3108
rect 5583 3012 6592 3040
rect 6641 3043 6699 3049
rect 5583 3009 5595 3012
rect 5537 3003 5595 3009
rect 6641 3009 6653 3043
rect 6687 3040 6699 3043
rect 6730 3040 6736 3052
rect 6687 3012 6736 3040
rect 6687 3009 6699 3012
rect 6641 3003 6699 3009
rect 6730 3000 6736 3012
rect 6788 3000 6794 3052
rect 6914 3000 6920 3052
rect 6972 3040 6978 3052
rect 7116 3049 7144 3080
rect 7101 3043 7159 3049
rect 7101 3040 7113 3043
rect 6972 3012 7113 3040
rect 6972 3000 6978 3012
rect 7101 3009 7113 3012
rect 7147 3009 7159 3043
rect 7101 3003 7159 3009
rect 7368 3043 7426 3049
rect 7368 3009 7380 3043
rect 7414 3040 7426 3043
rect 7834 3040 7840 3052
rect 7414 3012 7840 3040
rect 7414 3009 7426 3012
rect 7368 3003 7426 3009
rect 7834 3000 7840 3012
rect 7892 3000 7898 3052
rect 9048 3049 9076 3080
rect 9582 3068 9588 3080
rect 9640 3068 9646 3120
rect 9692 3108 9720 3148
rect 10410 3136 10416 3148
rect 10468 3136 10474 3188
rect 12434 3136 12440 3188
rect 12492 3176 12498 3188
rect 14918 3176 14924 3188
rect 12492 3148 14044 3176
rect 14879 3148 14924 3176
rect 12492 3136 12498 3148
rect 11238 3108 11244 3120
rect 9692 3080 11244 3108
rect 11238 3068 11244 3080
rect 11296 3068 11302 3120
rect 13262 3108 13268 3120
rect 11808 3080 13268 3108
rect 9033 3043 9091 3049
rect 9033 3009 9045 3043
rect 9079 3009 9091 3043
rect 9033 3003 9091 3009
rect 9122 3000 9128 3052
rect 9180 3040 9186 3052
rect 11808 3049 11836 3080
rect 13262 3068 13268 3080
rect 13320 3068 13326 3120
rect 13808 3111 13866 3117
rect 13372 3080 13768 3108
rect 9289 3043 9347 3049
rect 9289 3040 9301 3043
rect 9180 3012 9301 3040
rect 9180 3000 9186 3012
rect 9289 3009 9301 3012
rect 9335 3009 9347 3043
rect 11793 3043 11851 3049
rect 11793 3040 11805 3043
rect 9289 3003 9347 3009
rect 10060 3012 11805 3040
rect 3421 2975 3479 2981
rect 3421 2941 3433 2975
rect 3467 2972 3479 2975
rect 4890 2972 4896 2984
rect 3467 2944 4896 2972
rect 3467 2941 3479 2944
rect 3421 2935 3479 2941
rect 4890 2932 4896 2944
rect 4948 2932 4954 2984
rect 5077 2975 5135 2981
rect 5077 2941 5089 2975
rect 5123 2972 5135 2975
rect 5123 2944 7144 2972
rect 5123 2941 5135 2944
rect 5077 2935 5135 2941
rect 4525 2907 4583 2913
rect 4525 2873 4537 2907
rect 4571 2904 4583 2907
rect 5626 2904 5632 2916
rect 4571 2876 5632 2904
rect 4571 2873 4583 2876
rect 4525 2867 4583 2873
rect 5626 2864 5632 2876
rect 5684 2864 5690 2916
rect 5721 2907 5779 2913
rect 5721 2873 5733 2907
rect 5767 2904 5779 2907
rect 5902 2904 5908 2916
rect 5767 2876 5908 2904
rect 5767 2873 5779 2876
rect 5721 2867 5779 2873
rect 5902 2864 5908 2876
rect 5960 2864 5966 2916
rect 6454 2904 6460 2916
rect 6415 2876 6460 2904
rect 6454 2864 6460 2876
rect 6512 2864 6518 2916
rect 6730 2864 6736 2916
rect 6788 2864 6794 2916
rect 3973 2839 4031 2845
rect 3973 2805 3985 2839
rect 4019 2836 4031 2839
rect 6748 2836 6776 2864
rect 4019 2808 6776 2836
rect 7116 2836 7144 2944
rect 10060 2836 10088 3012
rect 11793 3009 11805 3012
rect 11839 3009 11851 3043
rect 12250 3040 12256 3052
rect 12211 3012 12256 3040
rect 11793 3003 11851 3009
rect 12250 3000 12256 3012
rect 12308 3000 12314 3052
rect 13372 3040 13400 3080
rect 13538 3040 13544 3052
rect 12406 3012 13400 3040
rect 13499 3012 13544 3040
rect 10410 2932 10416 2984
rect 10468 2972 10474 2984
rect 12406 2972 12434 3012
rect 13538 3000 13544 3012
rect 13596 3000 13602 3052
rect 13740 3040 13768 3080
rect 13808 3077 13820 3111
rect 13854 3108 13866 3111
rect 13906 3108 13912 3120
rect 13854 3080 13912 3108
rect 13854 3077 13866 3080
rect 13808 3071 13866 3077
rect 13906 3068 13912 3080
rect 13964 3068 13970 3120
rect 14016 3108 14044 3148
rect 14918 3136 14924 3148
rect 14976 3136 14982 3188
rect 15565 3179 15623 3185
rect 15565 3145 15577 3179
rect 15611 3176 15623 3179
rect 15654 3176 15660 3188
rect 15611 3148 15660 3176
rect 15611 3145 15623 3148
rect 15565 3139 15623 3145
rect 15654 3136 15660 3148
rect 15712 3136 15718 3188
rect 16853 3179 16911 3185
rect 16853 3176 16865 3179
rect 15764 3148 16865 3176
rect 15764 3108 15792 3148
rect 16853 3145 16865 3148
rect 16899 3145 16911 3179
rect 16853 3139 16911 3145
rect 19337 3179 19395 3185
rect 19337 3145 19349 3179
rect 19383 3176 19395 3179
rect 20070 3176 20076 3188
rect 19383 3148 20076 3176
rect 19383 3145 19395 3148
rect 19337 3139 19395 3145
rect 20070 3136 20076 3148
rect 20128 3136 20134 3188
rect 20530 3136 20536 3188
rect 20588 3176 20594 3188
rect 21821 3179 21879 3185
rect 21821 3176 21833 3179
rect 20588 3148 21833 3176
rect 20588 3136 20594 3148
rect 21821 3145 21833 3148
rect 21867 3145 21879 3179
rect 21821 3139 21879 3145
rect 55950 3136 55956 3188
rect 56008 3176 56014 3188
rect 58066 3176 58072 3188
rect 56008 3148 58072 3176
rect 56008 3136 56014 3148
rect 58066 3136 58072 3148
rect 58124 3136 58130 3188
rect 14016 3080 15792 3108
rect 16390 3068 16396 3120
rect 16448 3108 16454 3120
rect 16448 3080 17724 3108
rect 16448 3068 16454 3080
rect 14366 3040 14372 3052
rect 13740 3012 14372 3040
rect 14366 3000 14372 3012
rect 14424 3040 14430 3052
rect 14918 3040 14924 3052
rect 14424 3012 14924 3040
rect 14424 3000 14430 3012
rect 14918 3000 14924 3012
rect 14976 3000 14982 3052
rect 15194 3000 15200 3052
rect 15252 3040 15258 3052
rect 15381 3043 15439 3049
rect 15381 3040 15393 3043
rect 15252 3012 15393 3040
rect 15252 3000 15258 3012
rect 15381 3009 15393 3012
rect 15427 3009 15439 3043
rect 15381 3003 15439 3009
rect 16669 3043 16727 3049
rect 16669 3009 16681 3043
rect 16715 3040 16727 3043
rect 17310 3040 17316 3052
rect 16715 3012 17316 3040
rect 16715 3009 16727 3012
rect 16669 3003 16727 3009
rect 17310 3000 17316 3012
rect 17368 3000 17374 3052
rect 17696 3049 17724 3080
rect 57698 3068 57704 3120
rect 57756 3108 57762 3120
rect 60458 3108 60464 3120
rect 57756 3080 60464 3108
rect 57756 3068 57762 3080
rect 60458 3068 60464 3080
rect 60516 3068 60522 3120
rect 17681 3043 17739 3049
rect 17681 3009 17693 3043
rect 17727 3009 17739 3043
rect 17681 3003 17739 3009
rect 19153 3043 19211 3049
rect 19153 3009 19165 3043
rect 19199 3040 19211 3043
rect 21726 3040 21732 3052
rect 19199 3012 21732 3040
rect 19199 3009 19211 3012
rect 19153 3003 19211 3009
rect 20180 2984 20208 3012
rect 21726 3000 21732 3012
rect 21784 3000 21790 3052
rect 58158 3000 58164 3052
rect 58216 3040 58222 3052
rect 61105 3043 61163 3049
rect 61105 3040 61117 3043
rect 58216 3012 61117 3040
rect 58216 3000 58222 3012
rect 61105 3009 61117 3012
rect 61151 3009 61163 3043
rect 61105 3003 61163 3009
rect 10468 2944 12434 2972
rect 12529 2975 12587 2981
rect 10468 2932 10474 2944
rect 12529 2941 12541 2975
rect 12575 2972 12587 2975
rect 12710 2972 12716 2984
rect 12575 2944 12716 2972
rect 12575 2941 12587 2944
rect 12529 2935 12587 2941
rect 12710 2932 12716 2944
rect 12768 2932 12774 2984
rect 18693 2975 18751 2981
rect 18693 2941 18705 2975
rect 18739 2972 18751 2975
rect 19978 2972 19984 2984
rect 18739 2944 19984 2972
rect 18739 2941 18751 2944
rect 18693 2935 18751 2941
rect 19978 2932 19984 2944
rect 20036 2932 20042 2984
rect 20162 2932 20168 2984
rect 20220 2932 20226 2984
rect 21269 2975 21327 2981
rect 21269 2941 21281 2975
rect 21315 2972 21327 2975
rect 21818 2972 21824 2984
rect 21315 2944 21824 2972
rect 21315 2941 21327 2944
rect 21269 2935 21327 2941
rect 21818 2932 21824 2944
rect 21876 2932 21882 2984
rect 37274 2932 37280 2984
rect 37332 2972 37338 2984
rect 37921 2975 37979 2981
rect 37921 2972 37933 2975
rect 37332 2944 37933 2972
rect 37332 2932 37338 2944
rect 37921 2941 37933 2944
rect 37967 2941 37979 2975
rect 37921 2935 37979 2941
rect 44726 2932 44732 2984
rect 44784 2972 44790 2984
rect 45649 2975 45707 2981
rect 45649 2972 45661 2975
rect 44784 2944 45661 2972
rect 44784 2932 44790 2944
rect 45649 2941 45661 2944
rect 45695 2941 45707 2975
rect 45649 2935 45707 2941
rect 48590 2932 48596 2984
rect 48648 2972 48654 2984
rect 49513 2975 49571 2981
rect 49513 2972 49525 2975
rect 48648 2944 49525 2972
rect 48648 2932 48654 2944
rect 49513 2941 49525 2944
rect 49559 2941 49571 2975
rect 49513 2935 49571 2941
rect 52454 2932 52460 2984
rect 52512 2972 52518 2984
rect 53377 2975 53435 2981
rect 53377 2972 53389 2975
rect 52512 2944 53389 2972
rect 52512 2932 52518 2944
rect 53377 2941 53389 2944
rect 53423 2941 53435 2975
rect 53377 2935 53435 2941
rect 53558 2932 53564 2984
rect 53616 2972 53622 2984
rect 55214 2972 55220 2984
rect 53616 2944 55220 2972
rect 53616 2932 53622 2944
rect 55214 2932 55220 2944
rect 55272 2932 55278 2984
rect 56686 2932 56692 2984
rect 56744 2972 56750 2984
rect 56744 2944 58204 2972
rect 56744 2932 56750 2944
rect 10965 2907 11023 2913
rect 10965 2873 10977 2907
rect 11011 2904 11023 2907
rect 16758 2904 16764 2916
rect 11011 2876 12434 2904
rect 11011 2873 11023 2876
rect 10965 2867 11023 2873
rect 7116 2808 10088 2836
rect 11609 2839 11667 2845
rect 4019 2805 4031 2808
rect 3973 2799 4031 2805
rect 11609 2805 11621 2839
rect 11655 2836 11667 2839
rect 12066 2836 12072 2848
rect 11655 2808 12072 2836
rect 11655 2805 11667 2808
rect 11609 2799 11667 2805
rect 12066 2796 12072 2808
rect 12124 2796 12130 2848
rect 12406 2836 12434 2876
rect 14476 2876 16764 2904
rect 12526 2836 12532 2848
rect 12406 2808 12532 2836
rect 12526 2796 12532 2808
rect 12584 2796 12590 2848
rect 13906 2796 13912 2848
rect 13964 2836 13970 2848
rect 14476 2836 14504 2876
rect 16758 2864 16764 2876
rect 16816 2864 16822 2916
rect 38378 2864 38384 2916
rect 38436 2904 38442 2916
rect 39209 2907 39267 2913
rect 39209 2904 39221 2907
rect 38436 2876 39221 2904
rect 38436 2864 38442 2876
rect 39209 2873 39221 2876
rect 39255 2873 39267 2907
rect 39209 2867 39267 2873
rect 39758 2864 39764 2916
rect 39816 2904 39822 2916
rect 40497 2907 40555 2913
rect 40497 2904 40509 2907
rect 39816 2876 40509 2904
rect 39816 2864 39822 2876
rect 40497 2873 40509 2876
rect 40543 2873 40555 2907
rect 40497 2867 40555 2873
rect 42242 2864 42248 2916
rect 42300 2904 42306 2916
rect 43073 2907 43131 2913
rect 43073 2904 43085 2907
rect 42300 2876 43085 2904
rect 42300 2864 42306 2876
rect 43073 2873 43085 2876
rect 43119 2873 43131 2907
rect 43073 2867 43131 2873
rect 43622 2864 43628 2916
rect 43680 2904 43686 2916
rect 44361 2907 44419 2913
rect 44361 2904 44373 2907
rect 43680 2876 44373 2904
rect 43680 2864 43686 2876
rect 44361 2873 44373 2876
rect 44407 2873 44419 2907
rect 44361 2867 44419 2873
rect 47486 2864 47492 2916
rect 47544 2904 47550 2916
rect 48225 2907 48283 2913
rect 48225 2904 48237 2907
rect 47544 2876 48237 2904
rect 47544 2864 47550 2876
rect 48225 2873 48237 2876
rect 48271 2873 48283 2907
rect 48225 2867 48283 2873
rect 49418 2864 49424 2916
rect 49476 2904 49482 2916
rect 50157 2907 50215 2913
rect 50157 2904 50169 2907
rect 49476 2876 50169 2904
rect 49476 2864 49482 2876
rect 50157 2873 50169 2876
rect 50203 2873 50215 2907
rect 50157 2867 50215 2873
rect 50614 2864 50620 2916
rect 50672 2904 50678 2916
rect 51445 2907 51503 2913
rect 51445 2904 51457 2907
rect 50672 2876 51457 2904
rect 50672 2864 50678 2876
rect 51445 2873 51457 2876
rect 51491 2873 51503 2907
rect 51445 2867 51503 2873
rect 53282 2864 53288 2916
rect 53340 2904 53346 2916
rect 54021 2907 54079 2913
rect 54021 2904 54033 2907
rect 53340 2876 54033 2904
rect 53340 2864 53346 2876
rect 54021 2873 54033 2876
rect 54067 2873 54079 2907
rect 54021 2867 54079 2873
rect 54386 2864 54392 2916
rect 54444 2904 54450 2916
rect 55309 2907 55367 2913
rect 55309 2904 55321 2907
rect 54444 2876 55321 2904
rect 54444 2864 54450 2876
rect 55309 2873 55321 2876
rect 55355 2873 55367 2907
rect 55309 2867 55367 2873
rect 55674 2864 55680 2916
rect 55732 2904 55738 2916
rect 56597 2907 56655 2913
rect 56597 2904 56609 2907
rect 55732 2876 56609 2904
rect 55732 2864 55738 2876
rect 56597 2873 56609 2876
rect 56643 2873 56655 2907
rect 56597 2867 56655 2873
rect 57054 2864 57060 2916
rect 57112 2904 57118 2916
rect 58176 2904 58204 2944
rect 58434 2932 58440 2984
rect 58492 2972 58498 2984
rect 61749 2975 61807 2981
rect 61749 2972 61761 2975
rect 58492 2944 61761 2972
rect 58492 2932 58498 2944
rect 61749 2941 61761 2944
rect 61795 2941 61807 2975
rect 61749 2935 61807 2941
rect 58529 2907 58587 2913
rect 58529 2904 58541 2907
rect 57112 2876 58020 2904
rect 58176 2876 58541 2904
rect 57112 2864 57118 2876
rect 13964 2808 14504 2836
rect 13964 2796 13970 2808
rect 17034 2796 17040 2848
rect 17092 2836 17098 2848
rect 17497 2839 17555 2845
rect 17497 2836 17509 2839
rect 17092 2808 17509 2836
rect 17092 2796 17098 2808
rect 17497 2805 17509 2808
rect 17543 2805 17555 2839
rect 17497 2799 17555 2805
rect 19981 2839 20039 2845
rect 19981 2805 19993 2839
rect 20027 2836 20039 2839
rect 20254 2836 20260 2848
rect 20027 2808 20260 2836
rect 20027 2805 20039 2808
rect 19981 2799 20039 2805
rect 20254 2796 20260 2808
rect 20312 2796 20318 2848
rect 20625 2839 20683 2845
rect 20625 2805 20637 2839
rect 20671 2836 20683 2839
rect 20990 2836 20996 2848
rect 20671 2808 20996 2836
rect 20671 2805 20683 2808
rect 20625 2799 20683 2805
rect 20990 2796 20996 2808
rect 21048 2796 21054 2848
rect 22557 2839 22615 2845
rect 22557 2805 22569 2839
rect 22603 2836 22615 2839
rect 22646 2836 22652 2848
rect 22603 2808 22652 2836
rect 22603 2805 22615 2808
rect 22557 2799 22615 2805
rect 22646 2796 22652 2808
rect 22704 2796 22710 2848
rect 22922 2796 22928 2848
rect 22980 2836 22986 2848
rect 23017 2839 23075 2845
rect 23017 2836 23029 2839
rect 22980 2808 23029 2836
rect 22980 2796 22986 2808
rect 23017 2805 23029 2808
rect 23063 2805 23075 2839
rect 23017 2799 23075 2805
rect 23845 2839 23903 2845
rect 23845 2805 23857 2839
rect 23891 2836 23903 2839
rect 24026 2836 24032 2848
rect 23891 2808 24032 2836
rect 23891 2805 23903 2808
rect 23845 2799 23903 2805
rect 24026 2796 24032 2808
rect 24084 2796 24090 2848
rect 24489 2839 24547 2845
rect 24489 2805 24501 2839
rect 24535 2836 24547 2839
rect 24854 2836 24860 2848
rect 24535 2808 24860 2836
rect 24535 2805 24547 2808
rect 24489 2799 24547 2805
rect 24854 2796 24860 2808
rect 24912 2796 24918 2848
rect 25133 2839 25191 2845
rect 25133 2805 25145 2839
rect 25179 2836 25191 2839
rect 25406 2836 25412 2848
rect 25179 2808 25412 2836
rect 25179 2805 25191 2808
rect 25133 2799 25191 2805
rect 25406 2796 25412 2808
rect 25464 2796 25470 2848
rect 25777 2839 25835 2845
rect 25777 2805 25789 2839
rect 25823 2836 25835 2839
rect 26234 2836 26240 2848
rect 25823 2808 26240 2836
rect 25823 2805 25835 2808
rect 25777 2799 25835 2805
rect 26234 2796 26240 2808
rect 26292 2796 26298 2848
rect 26421 2839 26479 2845
rect 26421 2805 26433 2839
rect 26467 2836 26479 2839
rect 27062 2836 27068 2848
rect 26467 2808 27068 2836
rect 26467 2805 26479 2808
rect 26421 2799 26479 2805
rect 27062 2796 27068 2808
rect 27120 2796 27126 2848
rect 27709 2839 27767 2845
rect 27709 2805 27721 2839
rect 27755 2836 27767 2839
rect 27890 2836 27896 2848
rect 27755 2808 27896 2836
rect 27755 2805 27767 2808
rect 27709 2799 27767 2805
rect 27890 2796 27896 2808
rect 27948 2796 27954 2848
rect 28353 2839 28411 2845
rect 28353 2805 28365 2839
rect 28399 2836 28411 2839
rect 28442 2836 28448 2848
rect 28399 2808 28448 2836
rect 28399 2805 28411 2808
rect 28353 2799 28411 2805
rect 28442 2796 28448 2808
rect 28500 2796 28506 2848
rect 28997 2839 29055 2845
rect 28997 2805 29009 2839
rect 29043 2836 29055 2839
rect 29270 2836 29276 2848
rect 29043 2808 29276 2836
rect 29043 2805 29055 2808
rect 28997 2799 29055 2805
rect 29270 2796 29276 2808
rect 29328 2796 29334 2848
rect 29641 2839 29699 2845
rect 29641 2805 29653 2839
rect 29687 2836 29699 2839
rect 30098 2836 30104 2848
rect 29687 2808 30104 2836
rect 29687 2805 29699 2808
rect 29641 2799 29699 2805
rect 30098 2796 30104 2808
rect 30156 2796 30162 2848
rect 30285 2839 30343 2845
rect 30285 2805 30297 2839
rect 30331 2836 30343 2839
rect 30374 2836 30380 2848
rect 30331 2808 30380 2836
rect 30331 2805 30343 2808
rect 30285 2799 30343 2805
rect 30374 2796 30380 2808
rect 30432 2796 30438 2848
rect 30929 2839 30987 2845
rect 30929 2805 30941 2839
rect 30975 2836 30987 2839
rect 31202 2836 31208 2848
rect 30975 2808 31208 2836
rect 30975 2805 30987 2808
rect 30929 2799 30987 2805
rect 31202 2796 31208 2808
rect 31260 2796 31266 2848
rect 31573 2839 31631 2845
rect 31573 2805 31585 2839
rect 31619 2836 31631 2839
rect 32030 2836 32036 2848
rect 31619 2808 32036 2836
rect 31619 2805 31631 2808
rect 31573 2799 31631 2805
rect 32030 2796 32036 2808
rect 32088 2796 32094 2848
rect 32858 2836 32864 2848
rect 32819 2808 32864 2836
rect 32858 2796 32864 2808
rect 32916 2796 32922 2848
rect 33505 2839 33563 2845
rect 33505 2805 33517 2839
rect 33551 2836 33563 2839
rect 33686 2836 33692 2848
rect 33551 2808 33692 2836
rect 33551 2805 33563 2808
rect 33505 2799 33563 2805
rect 33686 2796 33692 2808
rect 33744 2796 33750 2848
rect 34149 2839 34207 2845
rect 34149 2805 34161 2839
rect 34195 2836 34207 2839
rect 34238 2836 34244 2848
rect 34195 2808 34244 2836
rect 34195 2805 34207 2808
rect 34149 2799 34207 2805
rect 34238 2796 34244 2808
rect 34296 2796 34302 2848
rect 34514 2796 34520 2848
rect 34572 2836 34578 2848
rect 34609 2839 34667 2845
rect 34609 2836 34621 2839
rect 34572 2808 34621 2836
rect 34572 2796 34578 2808
rect 34609 2805 34621 2808
rect 34655 2805 34667 2839
rect 34609 2799 34667 2805
rect 35342 2796 35348 2848
rect 35400 2836 35406 2848
rect 35437 2839 35495 2845
rect 35437 2836 35449 2839
rect 35400 2808 35449 2836
rect 35400 2796 35406 2808
rect 35437 2805 35449 2808
rect 35483 2805 35495 2839
rect 35437 2799 35495 2805
rect 36170 2796 36176 2848
rect 36228 2836 36234 2848
rect 36265 2839 36323 2845
rect 36265 2836 36277 2839
rect 36228 2808 36277 2836
rect 36228 2796 36234 2808
rect 36265 2805 36277 2808
rect 36311 2805 36323 2839
rect 36265 2799 36323 2805
rect 36722 2796 36728 2848
rect 36780 2836 36786 2848
rect 37277 2839 37335 2845
rect 37277 2836 37289 2839
rect 36780 2808 37289 2836
rect 36780 2796 36786 2808
rect 37277 2805 37289 2808
rect 37323 2805 37335 2839
rect 37277 2799 37335 2805
rect 37826 2796 37832 2848
rect 37884 2836 37890 2848
rect 38565 2839 38623 2845
rect 38565 2836 38577 2839
rect 37884 2808 38577 2836
rect 37884 2796 37890 2808
rect 38565 2805 38577 2808
rect 38611 2805 38623 2839
rect 38565 2799 38623 2805
rect 38930 2796 38936 2848
rect 38988 2836 38994 2848
rect 39853 2839 39911 2845
rect 39853 2836 39865 2839
rect 38988 2808 39865 2836
rect 38988 2796 38994 2808
rect 39853 2805 39865 2808
rect 39899 2805 39911 2839
rect 39853 2799 39911 2805
rect 40310 2796 40316 2848
rect 40368 2836 40374 2848
rect 41141 2839 41199 2845
rect 41141 2836 41153 2839
rect 40368 2808 41153 2836
rect 40368 2796 40374 2808
rect 41141 2805 41153 2808
rect 41187 2805 41199 2839
rect 41141 2799 41199 2805
rect 41690 2796 41696 2848
rect 41748 2836 41754 2848
rect 42429 2839 42487 2845
rect 42429 2836 42441 2839
rect 41748 2808 42441 2836
rect 41748 2796 41754 2808
rect 42429 2805 42441 2808
rect 42475 2805 42487 2839
rect 42429 2799 42487 2805
rect 42794 2796 42800 2848
rect 42852 2836 42858 2848
rect 43717 2839 43775 2845
rect 43717 2836 43729 2839
rect 42852 2808 43729 2836
rect 42852 2796 42858 2808
rect 43717 2805 43729 2808
rect 43763 2805 43775 2839
rect 43717 2799 43775 2805
rect 44174 2796 44180 2848
rect 44232 2836 44238 2848
rect 45005 2839 45063 2845
rect 45005 2836 45017 2839
rect 44232 2808 45017 2836
rect 44232 2796 44238 2808
rect 45005 2805 45017 2808
rect 45051 2805 45063 2839
rect 45005 2799 45063 2805
rect 45554 2796 45560 2848
rect 45612 2836 45618 2848
rect 46293 2839 46351 2845
rect 46293 2836 46305 2839
rect 45612 2808 46305 2836
rect 45612 2796 45618 2808
rect 46293 2805 46305 2808
rect 46339 2805 46351 2839
rect 46293 2799 46351 2805
rect 46658 2796 46664 2848
rect 46716 2836 46722 2848
rect 47581 2839 47639 2845
rect 47581 2836 47593 2839
rect 46716 2808 47593 2836
rect 46716 2796 46722 2808
rect 47581 2805 47593 2808
rect 47627 2805 47639 2839
rect 47581 2799 47639 2805
rect 48038 2796 48044 2848
rect 48096 2836 48102 2848
rect 48869 2839 48927 2845
rect 48869 2836 48881 2839
rect 48096 2808 48881 2836
rect 48096 2796 48102 2808
rect 48869 2805 48881 2808
rect 48915 2805 48927 2839
rect 48869 2799 48927 2805
rect 49970 2796 49976 2848
rect 50028 2836 50034 2848
rect 50801 2839 50859 2845
rect 50801 2836 50813 2839
rect 50028 2808 50813 2836
rect 50028 2796 50034 2808
rect 50801 2805 50813 2808
rect 50847 2805 50859 2839
rect 50801 2799 50859 2805
rect 51902 2796 51908 2848
rect 51960 2836 51966 2848
rect 52733 2839 52791 2845
rect 52733 2836 52745 2839
rect 51960 2808 52745 2836
rect 51960 2796 51966 2808
rect 52733 2805 52745 2808
rect 52779 2805 52791 2839
rect 52733 2799 52791 2805
rect 53834 2796 53840 2848
rect 53892 2836 53898 2848
rect 54665 2839 54723 2845
rect 54665 2836 54677 2839
rect 53892 2808 54677 2836
rect 53892 2796 53898 2808
rect 54665 2805 54677 2808
rect 54711 2805 54723 2839
rect 54665 2799 54723 2805
rect 55398 2796 55404 2848
rect 55456 2836 55462 2848
rect 55953 2839 56011 2845
rect 55953 2836 55965 2839
rect 55456 2808 55965 2836
rect 55456 2796 55462 2808
rect 55953 2805 55965 2808
rect 55999 2805 56011 2839
rect 55953 2799 56011 2805
rect 56042 2796 56048 2848
rect 56100 2836 56106 2848
rect 57885 2839 57943 2845
rect 57885 2836 57897 2839
rect 56100 2808 57897 2836
rect 56100 2796 56106 2808
rect 57885 2805 57897 2808
rect 57931 2805 57943 2839
rect 57992 2836 58020 2876
rect 58529 2873 58541 2876
rect 58575 2873 58587 2907
rect 58529 2867 58587 2873
rect 59354 2864 59360 2916
rect 59412 2904 59418 2916
rect 63037 2907 63095 2913
rect 63037 2904 63049 2907
rect 59412 2876 63049 2904
rect 59412 2864 59418 2876
rect 63037 2873 63049 2876
rect 63083 2873 63095 2907
rect 63037 2867 63095 2873
rect 59173 2839 59231 2845
rect 59173 2836 59185 2839
rect 57992 2808 59185 2836
rect 57885 2799 57943 2805
rect 59173 2805 59185 2808
rect 59219 2805 59231 2839
rect 59173 2799 59231 2805
rect 59446 2796 59452 2848
rect 59504 2836 59510 2848
rect 59817 2839 59875 2845
rect 59817 2836 59829 2839
rect 59504 2808 59829 2836
rect 59504 2796 59510 2808
rect 59817 2805 59829 2808
rect 59863 2805 59875 2839
rect 60458 2836 60464 2848
rect 60419 2808 60464 2836
rect 59817 2799 59875 2805
rect 60458 2796 60464 2808
rect 60516 2796 60522 2848
rect 1104 2746 68816 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 65654 2746
rect 65706 2694 65718 2746
rect 65770 2694 65782 2746
rect 65834 2694 65846 2746
rect 65898 2694 65910 2746
rect 65962 2694 68816 2746
rect 1104 2672 68816 2694
rect 7834 2632 7840 2644
rect 7795 2604 7840 2632
rect 7834 2592 7840 2604
rect 7892 2592 7898 2644
rect 9490 2592 9496 2644
rect 9548 2632 9554 2644
rect 11974 2632 11980 2644
rect 9548 2604 11980 2632
rect 9548 2592 9554 2604
rect 11974 2592 11980 2604
rect 12032 2592 12038 2644
rect 12066 2592 12072 2644
rect 12124 2632 12130 2644
rect 12250 2632 12256 2644
rect 12124 2604 12169 2632
rect 12211 2604 12256 2632
rect 12124 2592 12130 2604
rect 12250 2592 12256 2604
rect 12308 2592 12314 2644
rect 16850 2632 16856 2644
rect 12912 2604 16712 2632
rect 16811 2604 16856 2632
rect 9309 2567 9367 2573
rect 9309 2533 9321 2567
rect 9355 2564 9367 2567
rect 12710 2564 12716 2576
rect 9355 2536 12716 2564
rect 9355 2533 9367 2536
rect 9309 2527 9367 2533
rect 12710 2524 12716 2536
rect 12768 2524 12774 2576
rect 3881 2499 3939 2505
rect 3881 2465 3893 2499
rect 3927 2496 3939 2499
rect 3927 2468 6592 2496
rect 3927 2465 3939 2468
rect 3881 2459 3939 2465
rect 4890 2428 4896 2440
rect 4851 2400 4896 2428
rect 4890 2388 4896 2400
rect 4948 2388 4954 2440
rect 6564 2437 6592 2468
rect 6730 2456 6736 2508
rect 6788 2496 6794 2508
rect 8389 2499 8447 2505
rect 6788 2468 7512 2496
rect 6788 2456 6794 2468
rect 6549 2431 6607 2437
rect 6549 2397 6561 2431
rect 6595 2428 6607 2431
rect 6595 2400 6868 2428
rect 6595 2397 6607 2400
rect 6549 2391 6607 2397
rect 3237 2363 3295 2369
rect 3237 2329 3249 2363
rect 3283 2360 3295 2363
rect 5629 2363 5687 2369
rect 5629 2360 5641 2363
rect 3283 2332 5641 2360
rect 3283 2329 3295 2332
rect 3237 2323 3295 2329
rect 5629 2329 5641 2332
rect 5675 2360 5687 2363
rect 6730 2360 6736 2372
rect 5675 2332 6500 2360
rect 6691 2332 6736 2360
rect 5675 2329 5687 2332
rect 5629 2323 5687 2329
rect 4430 2292 4436 2304
rect 4391 2264 4436 2292
rect 4430 2252 4436 2264
rect 4488 2252 4494 2304
rect 5074 2292 5080 2304
rect 5035 2264 5080 2292
rect 5074 2252 5080 2264
rect 5132 2252 5138 2304
rect 5718 2292 5724 2304
rect 5679 2264 5724 2292
rect 5718 2252 5724 2264
rect 5776 2252 5782 2304
rect 6472 2292 6500 2332
rect 6730 2320 6736 2332
rect 6788 2320 6794 2372
rect 6840 2360 6868 2400
rect 7006 2388 7012 2440
rect 7064 2428 7070 2440
rect 7193 2431 7251 2437
rect 7193 2428 7205 2431
rect 7064 2400 7205 2428
rect 7064 2388 7070 2400
rect 7193 2397 7205 2400
rect 7239 2397 7251 2431
rect 7374 2428 7380 2440
rect 7335 2400 7380 2428
rect 7193 2391 7251 2397
rect 7374 2388 7380 2400
rect 7432 2388 7438 2440
rect 7484 2437 7512 2468
rect 8389 2465 8401 2499
rect 8435 2496 8447 2499
rect 11514 2496 11520 2508
rect 8435 2468 11520 2496
rect 8435 2465 8447 2468
rect 8389 2459 8447 2465
rect 11514 2456 11520 2468
rect 11572 2456 11578 2508
rect 7469 2431 7527 2437
rect 7469 2397 7481 2431
rect 7515 2397 7527 2431
rect 7469 2391 7527 2397
rect 7558 2388 7564 2440
rect 7616 2428 7622 2440
rect 9490 2428 9496 2440
rect 7616 2400 7661 2428
rect 9451 2400 9496 2428
rect 7616 2388 7622 2400
rect 9490 2388 9496 2400
rect 9548 2388 9554 2440
rect 9582 2388 9588 2440
rect 9640 2388 9646 2440
rect 10226 2428 10232 2440
rect 10187 2400 10232 2428
rect 10226 2388 10232 2400
rect 10284 2388 10290 2440
rect 10410 2388 10416 2440
rect 10468 2428 10474 2440
rect 10965 2431 11023 2437
rect 10965 2428 10977 2431
rect 10468 2400 10977 2428
rect 10468 2388 10474 2400
rect 10965 2397 10977 2400
rect 11011 2397 11023 2431
rect 10965 2391 11023 2397
rect 12115 2397 12173 2403
rect 9600 2360 9628 2388
rect 6840 2332 9628 2360
rect 10502 2320 10508 2372
rect 10560 2360 10566 2372
rect 11885 2363 11943 2369
rect 11885 2360 11897 2363
rect 10560 2332 11897 2360
rect 10560 2320 10566 2332
rect 11885 2329 11897 2332
rect 11931 2329 11943 2363
rect 12115 2363 12127 2397
rect 12161 2394 12173 2397
rect 12161 2372 12204 2394
rect 12618 2388 12624 2440
rect 12676 2428 12682 2440
rect 12713 2431 12771 2437
rect 12713 2428 12725 2431
rect 12676 2400 12725 2428
rect 12676 2388 12682 2400
rect 12713 2397 12725 2400
rect 12759 2397 12771 2431
rect 12912 2428 12940 2604
rect 12986 2524 12992 2576
rect 13044 2564 13050 2576
rect 13044 2536 13492 2564
rect 13044 2524 13050 2536
rect 12989 2431 13047 2437
rect 12989 2428 13001 2431
rect 12912 2400 13001 2428
rect 12713 2391 12771 2397
rect 12989 2397 13001 2400
rect 13035 2397 13047 2431
rect 12989 2391 13047 2397
rect 12161 2363 12164 2372
rect 12115 2357 12164 2363
rect 11885 2323 11943 2329
rect 12158 2320 12164 2357
rect 12216 2320 12222 2372
rect 13464 2360 13492 2536
rect 14366 2524 14372 2576
rect 14424 2564 14430 2576
rect 14734 2564 14740 2576
rect 14424 2536 14740 2564
rect 14424 2524 14430 2536
rect 14734 2524 14740 2536
rect 14792 2524 14798 2576
rect 16684 2564 16712 2604
rect 16850 2592 16856 2604
rect 16908 2592 16914 2644
rect 17586 2632 17592 2644
rect 17547 2604 17592 2632
rect 17586 2592 17592 2604
rect 17644 2592 17650 2644
rect 18230 2632 18236 2644
rect 18191 2604 18236 2632
rect 18230 2592 18236 2604
rect 18288 2592 18294 2644
rect 19306 2604 21404 2632
rect 17126 2564 17132 2576
rect 16684 2536 17132 2564
rect 17126 2524 17132 2536
rect 17184 2524 17190 2576
rect 19306 2564 19334 2604
rect 17604 2536 19334 2564
rect 20625 2567 20683 2573
rect 14458 2456 14464 2508
rect 14516 2496 14522 2508
rect 14516 2468 16712 2496
rect 14516 2456 14522 2468
rect 14369 2431 14427 2437
rect 14369 2397 14381 2431
rect 14415 2428 14427 2431
rect 14550 2428 14556 2440
rect 14415 2400 14556 2428
rect 14415 2397 14427 2400
rect 14369 2391 14427 2397
rect 14550 2388 14556 2400
rect 14608 2388 14614 2440
rect 14829 2431 14887 2437
rect 14829 2397 14841 2431
rect 14875 2397 14887 2431
rect 14829 2391 14887 2397
rect 14844 2360 14872 2391
rect 14918 2388 14924 2440
rect 14976 2428 14982 2440
rect 16684 2437 16712 2468
rect 15841 2431 15899 2437
rect 15841 2428 15853 2431
rect 14976 2400 15853 2428
rect 14976 2388 14982 2400
rect 15841 2397 15853 2400
rect 15887 2397 15899 2431
rect 15841 2391 15899 2397
rect 16669 2431 16727 2437
rect 16669 2397 16681 2431
rect 16715 2397 16727 2431
rect 16669 2391 16727 2397
rect 13464 2332 14872 2360
rect 15194 2320 15200 2372
rect 15252 2360 15258 2372
rect 17497 2363 17555 2369
rect 17497 2360 17509 2363
rect 15252 2332 17509 2360
rect 15252 2320 15258 2332
rect 17497 2329 17509 2332
rect 17543 2329 17555 2363
rect 17497 2323 17555 2329
rect 9582 2292 9588 2304
rect 6472 2264 9588 2292
rect 9582 2252 9588 2264
rect 9640 2252 9646 2304
rect 10042 2292 10048 2304
rect 10003 2264 10048 2292
rect 10042 2252 10048 2264
rect 10100 2252 10106 2304
rect 10781 2295 10839 2301
rect 10781 2261 10793 2295
rect 10827 2292 10839 2295
rect 12250 2292 12256 2304
rect 10827 2264 12256 2292
rect 10827 2261 10839 2264
rect 10781 2255 10839 2261
rect 12250 2252 12256 2264
rect 12308 2252 12314 2304
rect 14185 2295 14243 2301
rect 14185 2261 14197 2295
rect 14231 2292 14243 2295
rect 14458 2292 14464 2304
rect 14231 2264 14464 2292
rect 14231 2261 14243 2264
rect 14185 2255 14243 2261
rect 14458 2252 14464 2264
rect 14516 2252 14522 2304
rect 14734 2252 14740 2304
rect 14792 2292 14798 2304
rect 15013 2295 15071 2301
rect 15013 2292 15025 2295
rect 14792 2264 15025 2292
rect 14792 2252 14798 2264
rect 15013 2261 15025 2264
rect 15059 2261 15071 2295
rect 15654 2292 15660 2304
rect 15567 2264 15660 2292
rect 15013 2255 15071 2261
rect 15654 2252 15660 2264
rect 15712 2292 15718 2304
rect 17604 2292 17632 2536
rect 20625 2533 20637 2567
rect 20671 2564 20683 2567
rect 21266 2564 21272 2576
rect 20671 2536 21272 2564
rect 20671 2533 20683 2536
rect 20625 2527 20683 2533
rect 21266 2524 21272 2536
rect 21324 2524 21330 2576
rect 21376 2564 21404 2604
rect 21726 2592 21732 2644
rect 21784 2632 21790 2644
rect 21821 2635 21879 2641
rect 21821 2632 21833 2635
rect 21784 2604 21833 2632
rect 21784 2592 21790 2604
rect 21821 2601 21833 2604
rect 21867 2601 21879 2635
rect 23106 2632 23112 2644
rect 21821 2595 21879 2601
rect 22066 2604 23112 2632
rect 22066 2564 22094 2604
rect 23106 2592 23112 2604
rect 23164 2592 23170 2644
rect 55214 2592 55220 2644
rect 55272 2632 55278 2644
rect 55309 2635 55367 2641
rect 55309 2632 55321 2635
rect 55272 2604 55321 2632
rect 55272 2592 55278 2604
rect 55309 2601 55321 2604
rect 55355 2601 55367 2635
rect 55309 2595 55367 2601
rect 57422 2592 57428 2644
rect 57480 2632 57486 2644
rect 61105 2635 61163 2641
rect 61105 2632 61117 2635
rect 57480 2604 61117 2632
rect 57480 2592 57486 2604
rect 61105 2601 61117 2604
rect 61151 2601 61163 2635
rect 61105 2595 61163 2601
rect 21376 2536 22094 2564
rect 22557 2567 22615 2573
rect 22557 2533 22569 2567
rect 22603 2564 22615 2567
rect 23198 2564 23204 2576
rect 22603 2536 23204 2564
rect 22603 2533 22615 2536
rect 22557 2527 22615 2533
rect 23198 2524 23204 2536
rect 23256 2524 23262 2576
rect 28353 2567 28411 2573
rect 28353 2533 28365 2567
rect 28399 2564 28411 2567
rect 28994 2564 29000 2576
rect 28399 2536 29000 2564
rect 28399 2533 28411 2536
rect 28353 2527 28411 2533
rect 28994 2524 29000 2536
rect 29052 2524 29058 2576
rect 30285 2567 30343 2573
rect 30285 2533 30297 2567
rect 30331 2564 30343 2567
rect 30926 2564 30932 2576
rect 30331 2536 30932 2564
rect 30331 2533 30343 2536
rect 30285 2527 30343 2533
rect 30926 2524 30932 2536
rect 30984 2524 30990 2576
rect 40586 2524 40592 2576
rect 40644 2564 40650 2576
rect 42429 2567 42487 2573
rect 42429 2564 42441 2567
rect 40644 2536 42441 2564
rect 40644 2524 40650 2536
rect 42429 2533 42441 2536
rect 42475 2533 42487 2567
rect 42429 2527 42487 2533
rect 44450 2524 44456 2576
rect 44508 2564 44514 2576
rect 46293 2567 46351 2573
rect 46293 2564 46305 2567
rect 44508 2536 46305 2564
rect 44508 2524 44514 2536
rect 46293 2533 46305 2536
rect 46339 2533 46351 2567
rect 46293 2527 46351 2533
rect 48314 2524 48320 2576
rect 48372 2564 48378 2576
rect 50157 2567 50215 2573
rect 50157 2564 50169 2567
rect 48372 2536 50169 2564
rect 48372 2524 48378 2536
rect 50157 2533 50169 2536
rect 50203 2533 50215 2567
rect 50157 2527 50215 2533
rect 52178 2524 52184 2576
rect 52236 2564 52242 2576
rect 54021 2567 54079 2573
rect 54021 2564 54033 2567
rect 52236 2536 54033 2564
rect 52236 2524 52242 2536
rect 54021 2533 54033 2536
rect 54067 2533 54079 2567
rect 54021 2527 54079 2533
rect 55858 2524 55864 2576
rect 55916 2564 55922 2576
rect 57885 2567 57943 2573
rect 57885 2564 57897 2567
rect 55916 2536 57897 2564
rect 55916 2524 55922 2536
rect 57885 2533 57897 2536
rect 57931 2533 57943 2567
rect 57885 2527 57943 2533
rect 58066 2524 58072 2576
rect 58124 2564 58130 2576
rect 58529 2567 58587 2573
rect 58529 2564 58541 2567
rect 58124 2536 58541 2564
rect 58124 2524 58130 2536
rect 58529 2533 58541 2536
rect 58575 2533 58587 2567
rect 58529 2527 58587 2533
rect 60461 2567 60519 2573
rect 60461 2533 60473 2567
rect 60507 2533 60519 2567
rect 60461 2527 60519 2533
rect 18230 2456 18236 2508
rect 18288 2496 18294 2508
rect 25777 2499 25835 2505
rect 18288 2468 24808 2496
rect 18288 2456 18294 2468
rect 18414 2428 18420 2440
rect 18375 2400 18420 2428
rect 18414 2388 18420 2400
rect 18472 2388 18478 2440
rect 19981 2431 20039 2437
rect 19981 2397 19993 2431
rect 20027 2428 20039 2431
rect 20714 2428 20720 2440
rect 20027 2400 20720 2428
rect 20027 2397 20039 2400
rect 19981 2391 20039 2397
rect 20714 2388 20720 2400
rect 20772 2388 20778 2440
rect 21269 2431 21327 2437
rect 21269 2397 21281 2431
rect 21315 2428 21327 2431
rect 22094 2428 22100 2440
rect 21315 2400 22100 2428
rect 21315 2397 21327 2400
rect 21269 2391 21327 2397
rect 22094 2388 22100 2400
rect 22152 2388 22158 2440
rect 23201 2431 23259 2437
rect 23201 2397 23213 2431
rect 23247 2428 23259 2431
rect 23750 2428 23756 2440
rect 23247 2400 23756 2428
rect 23247 2397 23259 2400
rect 23201 2391 23259 2397
rect 23750 2388 23756 2400
rect 23808 2388 23814 2440
rect 23845 2431 23903 2437
rect 23845 2397 23857 2431
rect 23891 2428 23903 2431
rect 24578 2428 24584 2440
rect 23891 2400 24584 2428
rect 23891 2397 23903 2400
rect 23845 2391 23903 2397
rect 24578 2388 24584 2400
rect 24636 2388 24642 2440
rect 18432 2360 18460 2388
rect 24397 2363 24455 2369
rect 24397 2360 24409 2363
rect 18432 2332 24409 2360
rect 24397 2329 24409 2332
rect 24443 2329 24455 2363
rect 24780 2360 24808 2468
rect 25777 2465 25789 2499
rect 25823 2496 25835 2499
rect 26510 2496 26516 2508
rect 25823 2468 26516 2496
rect 25823 2465 25835 2468
rect 25777 2459 25835 2465
rect 26510 2456 26516 2468
rect 26568 2456 26574 2508
rect 36998 2456 37004 2508
rect 37056 2496 37062 2508
rect 37921 2499 37979 2505
rect 37921 2496 37933 2499
rect 37056 2468 37933 2496
rect 37056 2456 37062 2468
rect 37921 2465 37933 2468
rect 37967 2465 37979 2499
rect 37921 2459 37979 2465
rect 38102 2456 38108 2508
rect 38160 2496 38166 2508
rect 39853 2499 39911 2505
rect 39853 2496 39865 2499
rect 38160 2468 39865 2496
rect 38160 2456 38166 2468
rect 39853 2465 39865 2468
rect 39899 2465 39911 2499
rect 39853 2459 39911 2465
rect 41414 2456 41420 2508
rect 41472 2496 41478 2508
rect 43073 2499 43131 2505
rect 43073 2496 43085 2499
rect 41472 2468 43085 2496
rect 41472 2456 41478 2468
rect 43073 2465 43085 2468
rect 43119 2465 43131 2499
rect 43073 2459 43131 2465
rect 43346 2456 43352 2508
rect 43404 2496 43410 2508
rect 45005 2499 45063 2505
rect 45005 2496 45017 2499
rect 43404 2468 45017 2496
rect 43404 2456 43410 2468
rect 45005 2465 45017 2468
rect 45051 2465 45063 2499
rect 45005 2459 45063 2465
rect 46382 2456 46388 2508
rect 46440 2496 46446 2508
rect 48225 2499 48283 2505
rect 48225 2496 48237 2499
rect 46440 2468 48237 2496
rect 46440 2456 46446 2468
rect 48225 2465 48237 2468
rect 48271 2465 48283 2499
rect 48225 2459 48283 2465
rect 49142 2456 49148 2508
rect 49200 2496 49206 2508
rect 50801 2499 50859 2505
rect 50801 2496 50813 2499
rect 49200 2468 50813 2496
rect 49200 2456 49206 2468
rect 50801 2465 50813 2468
rect 50847 2465 50859 2499
rect 50801 2459 50859 2465
rect 51074 2456 51080 2508
rect 51132 2496 51138 2508
rect 52733 2499 52791 2505
rect 52733 2496 52745 2499
rect 51132 2468 52745 2496
rect 51132 2456 51138 2468
rect 52733 2465 52745 2468
rect 52779 2465 52791 2499
rect 52733 2459 52791 2465
rect 54938 2456 54944 2508
rect 54996 2496 55002 2508
rect 56597 2499 56655 2505
rect 56597 2496 56609 2499
rect 54996 2468 56609 2496
rect 54996 2456 55002 2468
rect 56597 2465 56609 2468
rect 56643 2465 56655 2499
rect 60476 2496 60504 2527
rect 63678 2496 63684 2508
rect 60476 2468 60596 2496
rect 63639 2468 63684 2496
rect 56597 2459 56655 2465
rect 25133 2431 25191 2437
rect 25133 2397 25145 2431
rect 25179 2428 25191 2431
rect 25682 2428 25688 2440
rect 25179 2400 25688 2428
rect 25179 2397 25191 2400
rect 25133 2391 25191 2397
rect 25682 2388 25688 2400
rect 25740 2388 25746 2440
rect 26421 2431 26479 2437
rect 26421 2397 26433 2431
rect 26467 2428 26479 2431
rect 27338 2428 27344 2440
rect 26467 2400 27344 2428
rect 26467 2397 26479 2400
rect 26421 2391 26479 2397
rect 27338 2388 27344 2400
rect 27396 2388 27402 2440
rect 27709 2431 27767 2437
rect 27709 2397 27721 2431
rect 27755 2428 27767 2431
rect 28166 2428 28172 2440
rect 27755 2400 28172 2428
rect 27755 2397 27767 2400
rect 27709 2391 27767 2397
rect 28166 2388 28172 2400
rect 28224 2388 28230 2440
rect 28997 2431 29055 2437
rect 28997 2397 29009 2431
rect 29043 2428 29055 2431
rect 29546 2428 29552 2440
rect 29043 2400 29552 2428
rect 29043 2397 29055 2400
rect 28997 2391 29055 2397
rect 29546 2388 29552 2400
rect 29604 2388 29610 2440
rect 30929 2431 30987 2437
rect 30929 2397 30941 2431
rect 30975 2397 30987 2431
rect 30929 2391 30987 2397
rect 31573 2431 31631 2437
rect 31573 2397 31585 2431
rect 31619 2428 31631 2431
rect 32582 2428 32588 2440
rect 31619 2400 32588 2428
rect 31619 2397 31631 2400
rect 31573 2391 31631 2397
rect 30944 2360 30972 2391
rect 32582 2388 32588 2400
rect 32640 2388 32646 2440
rect 32861 2431 32919 2437
rect 32861 2397 32873 2431
rect 32907 2428 32919 2431
rect 33410 2428 33416 2440
rect 32907 2400 33416 2428
rect 32907 2397 32919 2400
rect 32861 2391 32919 2397
rect 33410 2388 33416 2400
rect 33468 2388 33474 2440
rect 33505 2431 33563 2437
rect 33505 2397 33517 2431
rect 33551 2428 33563 2431
rect 33962 2428 33968 2440
rect 33551 2400 33968 2428
rect 33551 2397 33563 2400
rect 33505 2391 33563 2397
rect 33962 2388 33968 2400
rect 34020 2388 34026 2440
rect 34149 2431 34207 2437
rect 34149 2397 34161 2431
rect 34195 2428 34207 2431
rect 34790 2428 34796 2440
rect 34195 2400 34796 2428
rect 34195 2397 34207 2400
rect 34149 2391 34207 2397
rect 34790 2388 34796 2400
rect 34848 2388 34854 2440
rect 34885 2431 34943 2437
rect 34885 2397 34897 2431
rect 34931 2428 34943 2431
rect 35066 2428 35072 2440
rect 34931 2400 35072 2428
rect 34931 2397 34943 2400
rect 34885 2391 34943 2397
rect 35066 2388 35072 2400
rect 35124 2388 35130 2440
rect 35529 2431 35587 2437
rect 35529 2397 35541 2431
rect 35575 2428 35587 2431
rect 35618 2428 35624 2440
rect 35575 2400 35624 2428
rect 35575 2397 35587 2400
rect 35529 2391 35587 2397
rect 35618 2388 35624 2400
rect 35676 2388 35682 2440
rect 35894 2388 35900 2440
rect 35952 2428 35958 2440
rect 35989 2431 36047 2437
rect 35989 2428 36001 2431
rect 35952 2400 36001 2428
rect 35952 2388 35958 2400
rect 35989 2397 36001 2400
rect 36035 2397 36047 2431
rect 35989 2391 36047 2397
rect 36446 2388 36452 2440
rect 36504 2428 36510 2440
rect 37277 2431 37335 2437
rect 37277 2428 37289 2431
rect 36504 2400 37289 2428
rect 36504 2388 36510 2400
rect 37277 2397 37289 2400
rect 37323 2397 37335 2431
rect 37277 2391 37335 2397
rect 37550 2388 37556 2440
rect 37608 2428 37614 2440
rect 38565 2431 38623 2437
rect 38565 2428 38577 2431
rect 37608 2400 38577 2428
rect 37608 2388 37614 2400
rect 38565 2397 38577 2400
rect 38611 2397 38623 2431
rect 38565 2391 38623 2397
rect 38654 2388 38660 2440
rect 38712 2428 38718 2440
rect 40497 2431 40555 2437
rect 40497 2428 40509 2431
rect 38712 2400 40509 2428
rect 38712 2388 38718 2400
rect 40497 2397 40509 2400
rect 40543 2397 40555 2431
rect 40497 2391 40555 2397
rect 41141 2431 41199 2437
rect 41141 2397 41153 2431
rect 41187 2397 41199 2431
rect 41141 2391 41199 2397
rect 31754 2360 31760 2372
rect 24780 2332 26234 2360
rect 30944 2332 31760 2360
rect 24397 2323 24455 2329
rect 19334 2292 19340 2304
rect 15712 2264 17632 2292
rect 19295 2264 19340 2292
rect 15712 2252 15718 2264
rect 19334 2252 19340 2264
rect 19392 2252 19398 2304
rect 26206 2292 26234 2332
rect 31754 2320 31760 2332
rect 31812 2320 31818 2372
rect 39482 2320 39488 2372
rect 39540 2360 39546 2372
rect 41156 2360 41184 2391
rect 41966 2388 41972 2440
rect 42024 2428 42030 2440
rect 43717 2431 43775 2437
rect 43717 2428 43729 2431
rect 42024 2400 43729 2428
rect 42024 2388 42030 2400
rect 43717 2397 43729 2400
rect 43763 2397 43775 2431
rect 45649 2431 45707 2437
rect 45649 2428 45661 2431
rect 43717 2391 43775 2397
rect 45526 2400 45661 2428
rect 39540 2332 41184 2360
rect 39540 2320 39546 2332
rect 43898 2320 43904 2372
rect 43956 2360 43962 2372
rect 45526 2360 45554 2400
rect 45649 2397 45661 2400
rect 45695 2397 45707 2431
rect 45649 2391 45707 2397
rect 45830 2388 45836 2440
rect 45888 2428 45894 2440
rect 47581 2431 47639 2437
rect 47581 2428 47593 2431
rect 45888 2400 47593 2428
rect 45888 2388 45894 2400
rect 47581 2397 47593 2400
rect 47627 2397 47639 2431
rect 47581 2391 47639 2397
rect 48869 2431 48927 2437
rect 48869 2397 48881 2431
rect 48915 2397 48927 2431
rect 48869 2391 48927 2397
rect 43956 2332 45554 2360
rect 43956 2320 43962 2332
rect 47210 2320 47216 2372
rect 47268 2360 47274 2372
rect 48884 2360 48912 2391
rect 49694 2388 49700 2440
rect 49752 2428 49758 2440
rect 51445 2431 51503 2437
rect 51445 2428 51457 2431
rect 49752 2400 51457 2428
rect 49752 2388 49758 2400
rect 51445 2397 51457 2400
rect 51491 2397 51503 2431
rect 51445 2391 51503 2397
rect 51626 2388 51632 2440
rect 51684 2428 51690 2440
rect 53377 2431 53435 2437
rect 53377 2428 53389 2431
rect 51684 2400 53389 2428
rect 51684 2388 51690 2400
rect 53377 2397 53389 2400
rect 53423 2397 53435 2431
rect 53377 2391 53435 2397
rect 55953 2431 56011 2437
rect 55953 2397 55965 2431
rect 55999 2397 56011 2431
rect 55953 2391 56011 2397
rect 47268 2332 48912 2360
rect 47268 2320 47274 2332
rect 54110 2320 54116 2372
rect 54168 2360 54174 2372
rect 55968 2360 55996 2391
rect 56410 2388 56416 2440
rect 56468 2428 56474 2440
rect 59173 2431 59231 2437
rect 59173 2428 59185 2431
rect 56468 2400 59185 2428
rect 56468 2388 56474 2400
rect 59173 2397 59185 2400
rect 59219 2397 59231 2431
rect 59173 2391 59231 2397
rect 54168 2332 55996 2360
rect 54168 2320 54174 2332
rect 27706 2292 27712 2304
rect 26206 2264 27712 2292
rect 27706 2252 27712 2264
rect 27764 2252 27770 2304
rect 56870 2252 56876 2304
rect 56928 2292 56934 2304
rect 60568 2292 60596 2468
rect 63678 2456 63684 2468
rect 63736 2456 63742 2508
rect 61746 2428 61752 2440
rect 61707 2400 61752 2428
rect 61746 2388 61752 2400
rect 61804 2388 61810 2440
rect 63034 2428 63040 2440
rect 62995 2400 63040 2428
rect 63034 2388 63040 2400
rect 63092 2388 63098 2440
rect 67634 2428 67640 2440
rect 67595 2400 67640 2428
rect 67634 2388 67640 2400
rect 67692 2388 67698 2440
rect 56928 2264 60596 2292
rect 56928 2252 56934 2264
rect 1104 2202 68816 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 50294 2202
rect 50346 2150 50358 2202
rect 50410 2150 50422 2202
rect 50474 2150 50486 2202
rect 50538 2150 50550 2202
rect 50602 2150 68816 2202
rect 1104 2128 68816 2150
rect 4430 2048 4436 2100
rect 4488 2088 4494 2100
rect 12618 2088 12624 2100
rect 4488 2060 12624 2088
rect 4488 2048 4494 2060
rect 12618 2048 12624 2060
rect 12676 2048 12682 2100
rect 14550 2048 14556 2100
rect 14608 2088 14614 2100
rect 20346 2088 20352 2100
rect 14608 2060 20352 2088
rect 14608 2048 14614 2060
rect 20346 2048 20352 2060
rect 20404 2048 20410 2100
rect 58066 2048 58072 2100
rect 58124 2088 58130 2100
rect 61746 2088 61752 2100
rect 58124 2060 61752 2088
rect 58124 2048 58130 2060
rect 61746 2048 61752 2060
rect 61804 2048 61810 2100
rect 5074 1980 5080 2032
rect 5132 2020 5138 2032
rect 10134 2020 10140 2032
rect 5132 1992 10140 2020
rect 5132 1980 5138 1992
rect 10134 1980 10140 1992
rect 10192 2020 10198 2032
rect 12066 2020 12072 2032
rect 10192 1992 12072 2020
rect 10192 1980 10198 1992
rect 12066 1980 12072 1992
rect 12124 1980 12130 2032
rect 12986 2020 12992 2032
rect 12406 1992 12992 2020
rect 5626 1912 5632 1964
rect 5684 1952 5690 1964
rect 10226 1952 10232 1964
rect 5684 1924 10232 1952
rect 5684 1912 5690 1924
rect 10226 1912 10232 1924
rect 10284 1952 10290 1964
rect 12406 1952 12434 1992
rect 12986 1980 12992 1992
rect 13044 1980 13050 2032
rect 59078 1980 59084 2032
rect 59136 2020 59142 2032
rect 63678 2020 63684 2032
rect 59136 1992 63684 2020
rect 59136 1980 59142 1992
rect 63678 1980 63684 1992
rect 63736 1980 63742 2032
rect 10284 1924 12434 1952
rect 10284 1912 10290 1924
rect 12526 1912 12532 1964
rect 12584 1952 12590 1964
rect 15194 1952 15200 1964
rect 12584 1924 15200 1952
rect 12584 1912 12590 1924
rect 15194 1912 15200 1924
rect 15252 1912 15258 1964
rect 58526 1912 58532 1964
rect 58584 1952 58590 1964
rect 63034 1952 63040 1964
rect 58584 1924 63040 1952
rect 58584 1912 58590 1924
rect 63034 1912 63040 1924
rect 63092 1912 63098 1964
rect 12158 1844 12164 1896
rect 12216 1884 12222 1896
rect 19242 1884 19248 1896
rect 12216 1856 19248 1884
rect 12216 1844 12222 1856
rect 19242 1844 19248 1856
rect 19300 1844 19306 1896
rect 13538 1776 13544 1828
rect 13596 1816 13602 1828
rect 15378 1816 15384 1828
rect 13596 1788 15384 1816
rect 13596 1776 13602 1788
rect 15378 1776 15384 1788
rect 15436 1776 15442 1828
rect 4890 1708 4896 1760
rect 4948 1748 4954 1760
rect 10870 1748 10876 1760
rect 4948 1720 10876 1748
rect 4948 1708 4954 1720
rect 10870 1708 10876 1720
rect 10928 1708 10934 1760
rect 11974 1708 11980 1760
rect 12032 1748 12038 1760
rect 18414 1748 18420 1760
rect 12032 1720 18420 1748
rect 12032 1708 12038 1720
rect 18414 1708 18420 1720
rect 18472 1708 18478 1760
rect 19334 1708 19340 1760
rect 19392 1748 19398 1760
rect 19794 1748 19800 1760
rect 19392 1720 19800 1748
rect 19392 1708 19398 1720
rect 19794 1708 19800 1720
rect 19852 1708 19858 1760
rect 7558 1640 7564 1692
rect 7616 1680 7622 1692
rect 12802 1680 12808 1692
rect 7616 1652 12808 1680
rect 7616 1640 7622 1652
rect 12802 1640 12808 1652
rect 12860 1640 12866 1692
rect 5718 1572 5724 1624
rect 5776 1612 5782 1624
rect 14274 1612 14280 1624
rect 5776 1584 14280 1612
rect 5776 1572 5782 1584
rect 14274 1572 14280 1584
rect 14332 1572 14338 1624
rect 12250 1504 12256 1556
rect 12308 1544 12314 1556
rect 13354 1544 13360 1556
rect 12308 1516 13360 1544
rect 12308 1504 12314 1516
rect 13354 1504 13360 1516
rect 13412 1504 13418 1556
rect 19702 1504 19708 1556
rect 19760 1544 19766 1556
rect 20070 1544 20076 1556
rect 19760 1516 20076 1544
rect 19760 1504 19766 1516
rect 20070 1504 20076 1516
rect 20128 1504 20134 1556
rect 12066 1436 12072 1488
rect 12124 1476 12130 1488
rect 17034 1476 17040 1488
rect 12124 1448 17040 1476
rect 12124 1436 12130 1448
rect 17034 1436 17040 1448
rect 17092 1436 17098 1488
rect 10318 1368 10324 1420
rect 10376 1408 10382 1420
rect 10962 1408 10968 1420
rect 10376 1380 10968 1408
rect 10376 1368 10382 1380
rect 10962 1368 10968 1380
rect 11020 1368 11026 1420
rect 11790 1368 11796 1420
rect 11848 1408 11854 1420
rect 12250 1408 12256 1420
rect 11848 1380 12256 1408
rect 11848 1368 11854 1380
rect 12250 1368 12256 1380
rect 12308 1368 12314 1420
rect 12526 1368 12532 1420
rect 12584 1408 12590 1420
rect 12584 1380 12940 1408
rect 12584 1368 12590 1380
rect 11146 1300 11152 1352
rect 11204 1340 11210 1352
rect 11422 1340 11428 1352
rect 11204 1312 11428 1340
rect 11204 1300 11210 1312
rect 11422 1300 11428 1312
rect 11480 1300 11486 1352
rect 12912 1216 12940 1380
rect 18506 1368 18512 1420
rect 18564 1408 18570 1420
rect 19242 1408 19248 1420
rect 18564 1380 19248 1408
rect 18564 1368 18570 1380
rect 19242 1368 19248 1380
rect 19300 1368 19306 1420
rect 19518 1368 19524 1420
rect 19576 1408 19582 1420
rect 20622 1408 20628 1420
rect 19576 1380 20628 1408
rect 19576 1368 19582 1380
rect 20622 1368 20628 1380
rect 20680 1368 20686 1420
rect 9582 1164 9588 1216
rect 9640 1204 9646 1216
rect 11146 1204 11152 1216
rect 9640 1176 11152 1204
rect 9640 1164 9646 1176
rect 11146 1164 11152 1176
rect 11204 1164 11210 1216
rect 12894 1164 12900 1216
rect 12952 1164 12958 1216
rect 56778 1164 56784 1216
rect 56836 1204 56842 1216
rect 57054 1204 57060 1216
rect 56836 1176 57060 1204
rect 56836 1164 56842 1176
rect 57054 1164 57060 1176
rect 57112 1164 57118 1216
rect 57054 1028 57060 1080
rect 57112 1068 57118 1080
rect 59446 1068 59452 1080
rect 57112 1040 59452 1068
rect 57112 1028 57118 1040
rect 59446 1028 59452 1040
rect 59504 1028 59510 1080
<< via1 >>
rect 19574 57638 19626 57690
rect 19638 57638 19690 57690
rect 19702 57638 19754 57690
rect 19766 57638 19818 57690
rect 19830 57638 19882 57690
rect 50294 57638 50346 57690
rect 50358 57638 50410 57690
rect 50422 57638 50474 57690
rect 50486 57638 50538 57690
rect 50550 57638 50602 57690
rect 22100 57579 22152 57588
rect 22100 57545 22109 57579
rect 22109 57545 22143 57579
rect 22143 57545 22152 57579
rect 22100 57536 22152 57545
rect 30564 57536 30616 57588
rect 39304 57536 39356 57588
rect 48320 57579 48372 57588
rect 48320 57545 48329 57579
rect 48329 57545 48363 57579
rect 48363 57545 48372 57579
rect 48320 57536 48372 57545
rect 56784 57536 56836 57588
rect 65524 57536 65576 57588
rect 36820 57468 36872 57520
rect 4344 57400 4396 57452
rect 13084 57400 13136 57452
rect 21640 57400 21692 57452
rect 30104 57400 30156 57452
rect 56324 57400 56376 57452
rect 39304 57332 39356 57384
rect 67640 57443 67692 57452
rect 67640 57409 67649 57443
rect 67649 57409 67683 57443
rect 67683 57409 67692 57443
rect 67640 57400 67692 57409
rect 30104 57239 30156 57248
rect 30104 57205 30113 57239
rect 30113 57205 30147 57239
rect 30147 57205 30156 57239
rect 30104 57196 30156 57205
rect 39212 57239 39264 57248
rect 39212 57205 39221 57239
rect 39221 57205 39255 57239
rect 39255 57205 39264 57239
rect 39212 57196 39264 57205
rect 56324 57239 56376 57248
rect 56324 57205 56333 57239
rect 56333 57205 56367 57239
rect 56367 57205 56376 57239
rect 56324 57196 56376 57205
rect 4214 57094 4266 57146
rect 4278 57094 4330 57146
rect 4342 57094 4394 57146
rect 4406 57094 4458 57146
rect 4470 57094 4522 57146
rect 34934 57094 34986 57146
rect 34998 57094 35050 57146
rect 35062 57094 35114 57146
rect 35126 57094 35178 57146
rect 35190 57094 35242 57146
rect 65654 57094 65706 57146
rect 65718 57094 65770 57146
rect 65782 57094 65834 57146
rect 65846 57094 65898 57146
rect 65910 57094 65962 57146
rect 27160 56992 27212 57044
rect 39212 56992 39264 57044
rect 21640 56652 21692 56704
rect 19574 56550 19626 56602
rect 19638 56550 19690 56602
rect 19702 56550 19754 56602
rect 19766 56550 19818 56602
rect 19830 56550 19882 56602
rect 50294 56550 50346 56602
rect 50358 56550 50410 56602
rect 50422 56550 50474 56602
rect 50486 56550 50538 56602
rect 50550 56550 50602 56602
rect 67640 56151 67692 56160
rect 67640 56117 67649 56151
rect 67649 56117 67683 56151
rect 67683 56117 67692 56151
rect 67640 56108 67692 56117
rect 4214 56006 4266 56058
rect 4278 56006 4330 56058
rect 4342 56006 4394 56058
rect 4406 56006 4458 56058
rect 4470 56006 4522 56058
rect 34934 56006 34986 56058
rect 34998 56006 35050 56058
rect 35062 56006 35114 56058
rect 35126 56006 35178 56058
rect 35190 56006 35242 56058
rect 65654 56006 65706 56058
rect 65718 56006 65770 56058
rect 65782 56006 65834 56058
rect 65846 56006 65898 56058
rect 65910 56006 65962 56058
rect 19574 55462 19626 55514
rect 19638 55462 19690 55514
rect 19702 55462 19754 55514
rect 19766 55462 19818 55514
rect 19830 55462 19882 55514
rect 50294 55462 50346 55514
rect 50358 55462 50410 55514
rect 50422 55462 50474 55514
rect 50486 55462 50538 55514
rect 50550 55462 50602 55514
rect 4214 54918 4266 54970
rect 4278 54918 4330 54970
rect 4342 54918 4394 54970
rect 4406 54918 4458 54970
rect 4470 54918 4522 54970
rect 34934 54918 34986 54970
rect 34998 54918 35050 54970
rect 35062 54918 35114 54970
rect 35126 54918 35178 54970
rect 35190 54918 35242 54970
rect 65654 54918 65706 54970
rect 65718 54918 65770 54970
rect 65782 54918 65834 54970
rect 65846 54918 65898 54970
rect 65910 54918 65962 54970
rect 68100 54655 68152 54664
rect 68100 54621 68109 54655
rect 68109 54621 68143 54655
rect 68143 54621 68152 54655
rect 68100 54612 68152 54621
rect 19574 54374 19626 54426
rect 19638 54374 19690 54426
rect 19702 54374 19754 54426
rect 19766 54374 19818 54426
rect 19830 54374 19882 54426
rect 50294 54374 50346 54426
rect 50358 54374 50410 54426
rect 50422 54374 50474 54426
rect 50486 54374 50538 54426
rect 50550 54374 50602 54426
rect 4214 53830 4266 53882
rect 4278 53830 4330 53882
rect 4342 53830 4394 53882
rect 4406 53830 4458 53882
rect 4470 53830 4522 53882
rect 34934 53830 34986 53882
rect 34998 53830 35050 53882
rect 35062 53830 35114 53882
rect 35126 53830 35178 53882
rect 35190 53830 35242 53882
rect 65654 53830 65706 53882
rect 65718 53830 65770 53882
rect 65782 53830 65834 53882
rect 65846 53830 65898 53882
rect 65910 53830 65962 53882
rect 68100 53567 68152 53576
rect 68100 53533 68109 53567
rect 68109 53533 68143 53567
rect 68143 53533 68152 53567
rect 68100 53524 68152 53533
rect 19574 53286 19626 53338
rect 19638 53286 19690 53338
rect 19702 53286 19754 53338
rect 19766 53286 19818 53338
rect 19830 53286 19882 53338
rect 50294 53286 50346 53338
rect 50358 53286 50410 53338
rect 50422 53286 50474 53338
rect 50486 53286 50538 53338
rect 50550 53286 50602 53338
rect 4214 52742 4266 52794
rect 4278 52742 4330 52794
rect 4342 52742 4394 52794
rect 4406 52742 4458 52794
rect 4470 52742 4522 52794
rect 34934 52742 34986 52794
rect 34998 52742 35050 52794
rect 35062 52742 35114 52794
rect 35126 52742 35178 52794
rect 35190 52742 35242 52794
rect 65654 52742 65706 52794
rect 65718 52742 65770 52794
rect 65782 52742 65834 52794
rect 65846 52742 65898 52794
rect 65910 52742 65962 52794
rect 19574 52198 19626 52250
rect 19638 52198 19690 52250
rect 19702 52198 19754 52250
rect 19766 52198 19818 52250
rect 19830 52198 19882 52250
rect 50294 52198 50346 52250
rect 50358 52198 50410 52250
rect 50422 52198 50474 52250
rect 50486 52198 50538 52250
rect 50550 52198 50602 52250
rect 67640 51799 67692 51808
rect 67640 51765 67649 51799
rect 67649 51765 67683 51799
rect 67683 51765 67692 51799
rect 67640 51756 67692 51765
rect 4214 51654 4266 51706
rect 4278 51654 4330 51706
rect 4342 51654 4394 51706
rect 4406 51654 4458 51706
rect 4470 51654 4522 51706
rect 34934 51654 34986 51706
rect 34998 51654 35050 51706
rect 35062 51654 35114 51706
rect 35126 51654 35178 51706
rect 35190 51654 35242 51706
rect 65654 51654 65706 51706
rect 65718 51654 65770 51706
rect 65782 51654 65834 51706
rect 65846 51654 65898 51706
rect 65910 51654 65962 51706
rect 19574 51110 19626 51162
rect 19638 51110 19690 51162
rect 19702 51110 19754 51162
rect 19766 51110 19818 51162
rect 19830 51110 19882 51162
rect 50294 51110 50346 51162
rect 50358 51110 50410 51162
rect 50422 51110 50474 51162
rect 50486 51110 50538 51162
rect 50550 51110 50602 51162
rect 4214 50566 4266 50618
rect 4278 50566 4330 50618
rect 4342 50566 4394 50618
rect 4406 50566 4458 50618
rect 4470 50566 4522 50618
rect 34934 50566 34986 50618
rect 34998 50566 35050 50618
rect 35062 50566 35114 50618
rect 35126 50566 35178 50618
rect 35190 50566 35242 50618
rect 65654 50566 65706 50618
rect 65718 50566 65770 50618
rect 65782 50566 65834 50618
rect 65846 50566 65898 50618
rect 65910 50566 65962 50618
rect 68100 50303 68152 50312
rect 68100 50269 68109 50303
rect 68109 50269 68143 50303
rect 68143 50269 68152 50303
rect 68100 50260 68152 50269
rect 19574 50022 19626 50074
rect 19638 50022 19690 50074
rect 19702 50022 19754 50074
rect 19766 50022 19818 50074
rect 19830 50022 19882 50074
rect 50294 50022 50346 50074
rect 50358 50022 50410 50074
rect 50422 50022 50474 50074
rect 50486 50022 50538 50074
rect 50550 50022 50602 50074
rect 4214 49478 4266 49530
rect 4278 49478 4330 49530
rect 4342 49478 4394 49530
rect 4406 49478 4458 49530
rect 4470 49478 4522 49530
rect 34934 49478 34986 49530
rect 34998 49478 35050 49530
rect 35062 49478 35114 49530
rect 35126 49478 35178 49530
rect 35190 49478 35242 49530
rect 65654 49478 65706 49530
rect 65718 49478 65770 49530
rect 65782 49478 65834 49530
rect 65846 49478 65898 49530
rect 65910 49478 65962 49530
rect 19574 48934 19626 48986
rect 19638 48934 19690 48986
rect 19702 48934 19754 48986
rect 19766 48934 19818 48986
rect 19830 48934 19882 48986
rect 50294 48934 50346 48986
rect 50358 48934 50410 48986
rect 50422 48934 50474 48986
rect 50486 48934 50538 48986
rect 50550 48934 50602 48986
rect 67640 48603 67692 48612
rect 67640 48569 67649 48603
rect 67649 48569 67683 48603
rect 67683 48569 67692 48603
rect 67640 48560 67692 48569
rect 4214 48390 4266 48442
rect 4278 48390 4330 48442
rect 4342 48390 4394 48442
rect 4406 48390 4458 48442
rect 4470 48390 4522 48442
rect 34934 48390 34986 48442
rect 34998 48390 35050 48442
rect 35062 48390 35114 48442
rect 35126 48390 35178 48442
rect 35190 48390 35242 48442
rect 65654 48390 65706 48442
rect 65718 48390 65770 48442
rect 65782 48390 65834 48442
rect 65846 48390 65898 48442
rect 65910 48390 65962 48442
rect 19574 47846 19626 47898
rect 19638 47846 19690 47898
rect 19702 47846 19754 47898
rect 19766 47846 19818 47898
rect 19830 47846 19882 47898
rect 50294 47846 50346 47898
rect 50358 47846 50410 47898
rect 50422 47846 50474 47898
rect 50486 47846 50538 47898
rect 50550 47846 50602 47898
rect 67640 47447 67692 47456
rect 67640 47413 67649 47447
rect 67649 47413 67683 47447
rect 67683 47413 67692 47447
rect 67640 47404 67692 47413
rect 4214 47302 4266 47354
rect 4278 47302 4330 47354
rect 4342 47302 4394 47354
rect 4406 47302 4458 47354
rect 4470 47302 4522 47354
rect 34934 47302 34986 47354
rect 34998 47302 35050 47354
rect 35062 47302 35114 47354
rect 35126 47302 35178 47354
rect 35190 47302 35242 47354
rect 65654 47302 65706 47354
rect 65718 47302 65770 47354
rect 65782 47302 65834 47354
rect 65846 47302 65898 47354
rect 65910 47302 65962 47354
rect 19574 46758 19626 46810
rect 19638 46758 19690 46810
rect 19702 46758 19754 46810
rect 19766 46758 19818 46810
rect 19830 46758 19882 46810
rect 50294 46758 50346 46810
rect 50358 46758 50410 46810
rect 50422 46758 50474 46810
rect 50486 46758 50538 46810
rect 50550 46758 50602 46810
rect 4214 46214 4266 46266
rect 4278 46214 4330 46266
rect 4342 46214 4394 46266
rect 4406 46214 4458 46266
rect 4470 46214 4522 46266
rect 34934 46214 34986 46266
rect 34998 46214 35050 46266
rect 35062 46214 35114 46266
rect 35126 46214 35178 46266
rect 35190 46214 35242 46266
rect 65654 46214 65706 46266
rect 65718 46214 65770 46266
rect 65782 46214 65834 46266
rect 65846 46214 65898 46266
rect 65910 46214 65962 46266
rect 68100 45951 68152 45960
rect 68100 45917 68109 45951
rect 68109 45917 68143 45951
rect 68143 45917 68152 45951
rect 68100 45908 68152 45917
rect 19574 45670 19626 45722
rect 19638 45670 19690 45722
rect 19702 45670 19754 45722
rect 19766 45670 19818 45722
rect 19830 45670 19882 45722
rect 50294 45670 50346 45722
rect 50358 45670 50410 45722
rect 50422 45670 50474 45722
rect 50486 45670 50538 45722
rect 50550 45670 50602 45722
rect 4214 45126 4266 45178
rect 4278 45126 4330 45178
rect 4342 45126 4394 45178
rect 4406 45126 4458 45178
rect 4470 45126 4522 45178
rect 34934 45126 34986 45178
rect 34998 45126 35050 45178
rect 35062 45126 35114 45178
rect 35126 45126 35178 45178
rect 35190 45126 35242 45178
rect 65654 45126 65706 45178
rect 65718 45126 65770 45178
rect 65782 45126 65834 45178
rect 65846 45126 65898 45178
rect 65910 45126 65962 45178
rect 19574 44582 19626 44634
rect 19638 44582 19690 44634
rect 19702 44582 19754 44634
rect 19766 44582 19818 44634
rect 19830 44582 19882 44634
rect 50294 44582 50346 44634
rect 50358 44582 50410 44634
rect 50422 44582 50474 44634
rect 50486 44582 50538 44634
rect 50550 44582 50602 44634
rect 67548 44140 67600 44192
rect 4214 44038 4266 44090
rect 4278 44038 4330 44090
rect 4342 44038 4394 44090
rect 4406 44038 4458 44090
rect 4470 44038 4522 44090
rect 34934 44038 34986 44090
rect 34998 44038 35050 44090
rect 35062 44038 35114 44090
rect 35126 44038 35178 44090
rect 35190 44038 35242 44090
rect 65654 44038 65706 44090
rect 65718 44038 65770 44090
rect 65782 44038 65834 44090
rect 65846 44038 65898 44090
rect 65910 44038 65962 44090
rect 19574 43494 19626 43546
rect 19638 43494 19690 43546
rect 19702 43494 19754 43546
rect 19766 43494 19818 43546
rect 19830 43494 19882 43546
rect 50294 43494 50346 43546
rect 50358 43494 50410 43546
rect 50422 43494 50474 43546
rect 50486 43494 50538 43546
rect 50550 43494 50602 43546
rect 4214 42950 4266 43002
rect 4278 42950 4330 43002
rect 4342 42950 4394 43002
rect 4406 42950 4458 43002
rect 4470 42950 4522 43002
rect 34934 42950 34986 43002
rect 34998 42950 35050 43002
rect 35062 42950 35114 43002
rect 35126 42950 35178 43002
rect 35190 42950 35242 43002
rect 65654 42950 65706 43002
rect 65718 42950 65770 43002
rect 65782 42950 65834 43002
rect 65846 42950 65898 43002
rect 65910 42950 65962 43002
rect 68100 42687 68152 42696
rect 68100 42653 68109 42687
rect 68109 42653 68143 42687
rect 68143 42653 68152 42687
rect 68100 42644 68152 42653
rect 19574 42406 19626 42458
rect 19638 42406 19690 42458
rect 19702 42406 19754 42458
rect 19766 42406 19818 42458
rect 19830 42406 19882 42458
rect 50294 42406 50346 42458
rect 50358 42406 50410 42458
rect 50422 42406 50474 42458
rect 50486 42406 50538 42458
rect 50550 42406 50602 42458
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 34934 41862 34986 41914
rect 34998 41862 35050 41914
rect 35062 41862 35114 41914
rect 35126 41862 35178 41914
rect 35190 41862 35242 41914
rect 65654 41862 65706 41914
rect 65718 41862 65770 41914
rect 65782 41862 65834 41914
rect 65846 41862 65898 41914
rect 65910 41862 65962 41914
rect 68100 41599 68152 41608
rect 68100 41565 68109 41599
rect 68109 41565 68143 41599
rect 68143 41565 68152 41599
rect 68100 41556 68152 41565
rect 19574 41318 19626 41370
rect 19638 41318 19690 41370
rect 19702 41318 19754 41370
rect 19766 41318 19818 41370
rect 19830 41318 19882 41370
rect 50294 41318 50346 41370
rect 50358 41318 50410 41370
rect 50422 41318 50474 41370
rect 50486 41318 50538 41370
rect 50550 41318 50602 41370
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 34934 40774 34986 40826
rect 34998 40774 35050 40826
rect 35062 40774 35114 40826
rect 35126 40774 35178 40826
rect 35190 40774 35242 40826
rect 65654 40774 65706 40826
rect 65718 40774 65770 40826
rect 65782 40774 65834 40826
rect 65846 40774 65898 40826
rect 65910 40774 65962 40826
rect 19574 40230 19626 40282
rect 19638 40230 19690 40282
rect 19702 40230 19754 40282
rect 19766 40230 19818 40282
rect 19830 40230 19882 40282
rect 50294 40230 50346 40282
rect 50358 40230 50410 40282
rect 50422 40230 50474 40282
rect 50486 40230 50538 40282
rect 50550 40230 50602 40282
rect 67640 39831 67692 39840
rect 67640 39797 67649 39831
rect 67649 39797 67683 39831
rect 67683 39797 67692 39831
rect 67640 39788 67692 39797
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 65654 39686 65706 39738
rect 65718 39686 65770 39738
rect 65782 39686 65834 39738
rect 65846 39686 65898 39738
rect 65910 39686 65962 39738
rect 19574 39142 19626 39194
rect 19638 39142 19690 39194
rect 19702 39142 19754 39194
rect 19766 39142 19818 39194
rect 19830 39142 19882 39194
rect 50294 39142 50346 39194
rect 50358 39142 50410 39194
rect 50422 39142 50474 39194
rect 50486 39142 50538 39194
rect 50550 39142 50602 39194
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 65654 38598 65706 38650
rect 65718 38598 65770 38650
rect 65782 38598 65834 38650
rect 65846 38598 65898 38650
rect 65910 38598 65962 38650
rect 68100 38335 68152 38344
rect 68100 38301 68109 38335
rect 68109 38301 68143 38335
rect 68143 38301 68152 38335
rect 68100 38292 68152 38301
rect 19574 38054 19626 38106
rect 19638 38054 19690 38106
rect 19702 38054 19754 38106
rect 19766 38054 19818 38106
rect 19830 38054 19882 38106
rect 50294 38054 50346 38106
rect 50358 38054 50410 38106
rect 50422 38054 50474 38106
rect 50486 38054 50538 38106
rect 50550 38054 50602 38106
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 65654 37510 65706 37562
rect 65718 37510 65770 37562
rect 65782 37510 65834 37562
rect 65846 37510 65898 37562
rect 65910 37510 65962 37562
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 50294 36966 50346 37018
rect 50358 36966 50410 37018
rect 50422 36966 50474 37018
rect 50486 36966 50538 37018
rect 50550 36966 50602 37018
rect 67640 36635 67692 36644
rect 67640 36601 67649 36635
rect 67649 36601 67683 36635
rect 67683 36601 67692 36635
rect 67640 36592 67692 36601
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 65654 36422 65706 36474
rect 65718 36422 65770 36474
rect 65782 36422 65834 36474
rect 65846 36422 65898 36474
rect 65910 36422 65962 36474
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 50294 35878 50346 35930
rect 50358 35878 50410 35930
rect 50422 35878 50474 35930
rect 50486 35878 50538 35930
rect 50550 35878 50602 35930
rect 67640 35479 67692 35488
rect 67640 35445 67649 35479
rect 67649 35445 67683 35479
rect 67683 35445 67692 35479
rect 67640 35436 67692 35445
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 65654 35334 65706 35386
rect 65718 35334 65770 35386
rect 65782 35334 65834 35386
rect 65846 35334 65898 35386
rect 65910 35334 65962 35386
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 50294 34790 50346 34842
rect 50358 34790 50410 34842
rect 50422 34790 50474 34842
rect 50486 34790 50538 34842
rect 50550 34790 50602 34842
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 65654 34246 65706 34298
rect 65718 34246 65770 34298
rect 65782 34246 65834 34298
rect 65846 34246 65898 34298
rect 65910 34246 65962 34298
rect 68100 33983 68152 33992
rect 68100 33949 68109 33983
rect 68109 33949 68143 33983
rect 68143 33949 68152 33983
rect 68100 33940 68152 33949
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 50294 33702 50346 33754
rect 50358 33702 50410 33754
rect 50422 33702 50474 33754
rect 50486 33702 50538 33754
rect 50550 33702 50602 33754
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 65654 33158 65706 33210
rect 65718 33158 65770 33210
rect 65782 33158 65834 33210
rect 65846 33158 65898 33210
rect 65910 33158 65962 33210
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 50294 32614 50346 32666
rect 50358 32614 50410 32666
rect 50422 32614 50474 32666
rect 50486 32614 50538 32666
rect 50550 32614 50602 32666
rect 67640 32215 67692 32224
rect 67640 32181 67649 32215
rect 67649 32181 67683 32215
rect 67683 32181 67692 32215
rect 67640 32172 67692 32181
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 65654 32070 65706 32122
rect 65718 32070 65770 32122
rect 65782 32070 65834 32122
rect 65846 32070 65898 32122
rect 65910 32070 65962 32122
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 50294 31526 50346 31578
rect 50358 31526 50410 31578
rect 50422 31526 50474 31578
rect 50486 31526 50538 31578
rect 50550 31526 50602 31578
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 65654 30982 65706 31034
rect 65718 30982 65770 31034
rect 65782 30982 65834 31034
rect 65846 30982 65898 31034
rect 65910 30982 65962 31034
rect 68100 30719 68152 30728
rect 68100 30685 68109 30719
rect 68109 30685 68143 30719
rect 68143 30685 68152 30719
rect 68100 30676 68152 30685
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 50294 30438 50346 30490
rect 50358 30438 50410 30490
rect 50422 30438 50474 30490
rect 50486 30438 50538 30490
rect 50550 30438 50602 30490
rect 7564 30200 7616 30252
rect 30104 30200 30156 30252
rect 6736 30132 6788 30184
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 65654 29894 65706 29946
rect 65718 29894 65770 29946
rect 65782 29894 65834 29946
rect 65846 29894 65898 29946
rect 65910 29894 65962 29946
rect 27160 29835 27212 29844
rect 27160 29801 27169 29835
rect 27169 29801 27203 29835
rect 27203 29801 27212 29835
rect 27160 29792 27212 29801
rect 8024 29588 8076 29640
rect 25780 29588 25832 29640
rect 26424 29631 26476 29640
rect 26424 29597 26433 29631
rect 26433 29597 26467 29631
rect 26467 29597 26476 29631
rect 26424 29588 26476 29597
rect 68100 29631 68152 29640
rect 68100 29597 68109 29631
rect 68109 29597 68143 29631
rect 68143 29597 68152 29631
rect 68100 29588 68152 29597
rect 7932 29520 7984 29572
rect 7564 29452 7616 29504
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 50294 29350 50346 29402
rect 50358 29350 50410 29402
rect 50422 29350 50474 29402
rect 50486 29350 50538 29402
rect 50550 29350 50602 29402
rect 5080 29155 5132 29164
rect 5080 29121 5089 29155
rect 5089 29121 5123 29155
rect 5123 29121 5132 29155
rect 5080 29112 5132 29121
rect 7932 29180 7984 29232
rect 7012 29044 7064 29096
rect 19892 29112 19944 29164
rect 25044 29112 25096 29164
rect 8116 29044 8168 29096
rect 19432 29087 19484 29096
rect 19432 29053 19441 29087
rect 19441 29053 19475 29087
rect 19475 29053 19484 29087
rect 19432 29044 19484 29053
rect 5816 29019 5868 29028
rect 5816 28985 5825 29019
rect 5825 28985 5859 29019
rect 5859 28985 5868 29019
rect 5816 28976 5868 28985
rect 8024 28976 8076 29028
rect 18972 29019 19024 29028
rect 4804 28908 4856 28960
rect 6736 28908 6788 28960
rect 6920 28951 6972 28960
rect 6920 28917 6929 28951
rect 6929 28917 6963 28951
rect 6963 28917 6972 28951
rect 6920 28908 6972 28917
rect 7656 28908 7708 28960
rect 18972 28985 18981 29019
rect 18981 28985 19015 29019
rect 19015 28985 19024 29019
rect 18972 28976 19024 28985
rect 9404 28908 9456 28960
rect 24400 28951 24452 28960
rect 24400 28917 24409 28951
rect 24409 28917 24443 28951
rect 24443 28917 24452 28951
rect 24400 28908 24452 28917
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 65654 28806 65706 28858
rect 65718 28806 65770 28858
rect 65782 28806 65834 28858
rect 65846 28806 65898 28858
rect 65910 28806 65962 28858
rect 6736 28747 6788 28756
rect 6736 28713 6745 28747
rect 6745 28713 6779 28747
rect 6779 28713 6788 28747
rect 6736 28704 6788 28713
rect 8300 28747 8352 28756
rect 8300 28713 8309 28747
rect 8309 28713 8343 28747
rect 8343 28713 8352 28747
rect 8300 28704 8352 28713
rect 4804 28611 4856 28620
rect 4804 28577 4813 28611
rect 4813 28577 4847 28611
rect 4847 28577 4856 28611
rect 4804 28568 4856 28577
rect 5080 28500 5132 28552
rect 9680 28636 9732 28688
rect 6276 28543 6328 28552
rect 6276 28509 6285 28543
rect 6285 28509 6319 28543
rect 6319 28509 6328 28543
rect 6276 28500 6328 28509
rect 6920 28543 6972 28552
rect 6920 28509 6929 28543
rect 6929 28509 6963 28543
rect 6963 28509 6972 28543
rect 6920 28500 6972 28509
rect 7656 28500 7708 28552
rect 8116 28543 8168 28552
rect 8116 28509 8125 28543
rect 8125 28509 8159 28543
rect 8159 28509 8168 28543
rect 8116 28500 8168 28509
rect 9404 28500 9456 28552
rect 18972 28636 19024 28688
rect 18604 28568 18656 28620
rect 19248 28704 19300 28756
rect 9128 28432 9180 28484
rect 3792 28407 3844 28416
rect 3792 28373 3801 28407
rect 3801 28373 3835 28407
rect 3835 28373 3844 28407
rect 3792 28364 3844 28373
rect 7840 28364 7892 28416
rect 7932 28364 7984 28416
rect 10232 28500 10284 28552
rect 14004 28500 14056 28552
rect 18052 28543 18104 28552
rect 15384 28475 15436 28484
rect 15384 28441 15393 28475
rect 15393 28441 15427 28475
rect 15427 28441 15436 28475
rect 15384 28432 15436 28441
rect 18052 28509 18061 28543
rect 18061 28509 18095 28543
rect 18095 28509 18104 28543
rect 18052 28500 18104 28509
rect 19340 28500 19392 28552
rect 19892 28543 19944 28552
rect 19892 28509 19901 28543
rect 19901 28509 19935 28543
rect 19935 28509 19944 28543
rect 19892 28500 19944 28509
rect 20076 28500 20128 28552
rect 26056 28704 26108 28756
rect 16764 28432 16816 28484
rect 17776 28475 17828 28484
rect 17776 28441 17785 28475
rect 17785 28441 17819 28475
rect 17819 28441 17828 28475
rect 17776 28432 17828 28441
rect 19432 28364 19484 28416
rect 20076 28364 20128 28416
rect 25688 28568 25740 28620
rect 22008 28543 22060 28552
rect 22008 28509 22017 28543
rect 22017 28509 22051 28543
rect 22051 28509 22060 28543
rect 22008 28500 22060 28509
rect 23204 28543 23256 28552
rect 23204 28509 23213 28543
rect 23213 28509 23247 28543
rect 23247 28509 23256 28543
rect 23204 28500 23256 28509
rect 23296 28543 23348 28552
rect 23296 28509 23305 28543
rect 23305 28509 23339 28543
rect 23339 28509 23348 28543
rect 23296 28500 23348 28509
rect 24400 28500 24452 28552
rect 25044 28543 25096 28552
rect 25044 28509 25053 28543
rect 25053 28509 25087 28543
rect 25087 28509 25096 28543
rect 25044 28500 25096 28509
rect 25136 28543 25188 28552
rect 25136 28509 25145 28543
rect 25145 28509 25179 28543
rect 25179 28509 25188 28543
rect 26056 28543 26108 28552
rect 25136 28500 25188 28509
rect 26056 28509 26065 28543
rect 26065 28509 26099 28543
rect 26099 28509 26108 28543
rect 26056 28500 26108 28509
rect 25688 28432 25740 28484
rect 22008 28364 22060 28416
rect 23572 28364 23624 28416
rect 25136 28364 25188 28416
rect 25596 28364 25648 28416
rect 26792 28407 26844 28416
rect 26792 28373 26801 28407
rect 26801 28373 26835 28407
rect 26835 28373 26844 28407
rect 26792 28364 26844 28373
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 50294 28262 50346 28314
rect 50358 28262 50410 28314
rect 50422 28262 50474 28314
rect 50486 28262 50538 28314
rect 50550 28262 50602 28314
rect 6276 28160 6328 28212
rect 9128 28203 9180 28212
rect 9128 28169 9137 28203
rect 9137 28169 9171 28203
rect 9171 28169 9180 28203
rect 9128 28160 9180 28169
rect 9680 28160 9732 28212
rect 23204 28160 23256 28212
rect 23296 28160 23348 28212
rect 25688 28160 25740 28212
rect 7564 28067 7616 28076
rect 7564 28033 7573 28067
rect 7573 28033 7607 28067
rect 7607 28033 7616 28067
rect 7564 28024 7616 28033
rect 7840 28067 7892 28076
rect 7840 28033 7849 28067
rect 7849 28033 7883 28067
rect 7883 28033 7892 28067
rect 7840 28024 7892 28033
rect 8576 28024 8628 28076
rect 9404 28067 9456 28076
rect 9404 28033 9413 28067
rect 9413 28033 9447 28067
rect 9447 28033 9456 28067
rect 9404 28024 9456 28033
rect 11612 28024 11664 28076
rect 12164 28024 12216 28076
rect 9588 27956 9640 28008
rect 14004 27956 14056 28008
rect 8300 27888 8352 27940
rect 9496 27888 9548 27940
rect 18052 28092 18104 28144
rect 22376 28092 22428 28144
rect 18236 28024 18288 28076
rect 19340 28067 19392 28076
rect 19340 28033 19349 28067
rect 19349 28033 19383 28067
rect 19383 28033 19392 28067
rect 19340 28024 19392 28033
rect 19524 28067 19576 28076
rect 19524 28033 19533 28067
rect 19533 28033 19567 28067
rect 19567 28033 19576 28067
rect 19524 28024 19576 28033
rect 20076 28024 20128 28076
rect 23480 28067 23532 28076
rect 23480 28033 23489 28067
rect 23489 28033 23523 28067
rect 23523 28033 23532 28067
rect 23480 28024 23532 28033
rect 24400 28067 24452 28076
rect 24400 28033 24409 28067
rect 24409 28033 24443 28067
rect 24443 28033 24452 28067
rect 24400 28024 24452 28033
rect 19984 27956 20036 28008
rect 15384 27888 15436 27940
rect 17224 27888 17276 27940
rect 18328 27888 18380 27940
rect 19248 27888 19300 27940
rect 25136 28024 25188 28076
rect 25596 28067 25648 28076
rect 25596 28033 25605 28067
rect 25605 28033 25639 28067
rect 25639 28033 25648 28067
rect 25596 28024 25648 28033
rect 9220 27863 9272 27872
rect 9220 27829 9229 27863
rect 9229 27829 9263 27863
rect 9263 27829 9272 27863
rect 9220 27820 9272 27829
rect 9312 27863 9364 27872
rect 9312 27829 9321 27863
rect 9321 27829 9355 27863
rect 9355 27829 9364 27863
rect 9312 27820 9364 27829
rect 10876 27820 10928 27872
rect 13912 27820 13964 27872
rect 14556 27820 14608 27872
rect 17408 27863 17460 27872
rect 17408 27829 17417 27863
rect 17417 27829 17451 27863
rect 17451 27829 17460 27863
rect 17408 27820 17460 27829
rect 17960 27863 18012 27872
rect 17960 27829 17969 27863
rect 17969 27829 18003 27863
rect 18003 27829 18012 27863
rect 17960 27820 18012 27829
rect 19524 27820 19576 27872
rect 22468 27820 22520 27872
rect 24308 27820 24360 27872
rect 26424 27820 26476 27872
rect 67640 27863 67692 27872
rect 67640 27829 67649 27863
rect 67649 27829 67683 27863
rect 67683 27829 67692 27863
rect 67640 27820 67692 27829
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 65654 27718 65706 27770
rect 65718 27718 65770 27770
rect 65782 27718 65834 27770
rect 65846 27718 65898 27770
rect 65910 27718 65962 27770
rect 3792 27616 3844 27668
rect 9312 27616 9364 27668
rect 10232 27659 10284 27668
rect 10232 27625 10241 27659
rect 10241 27625 10275 27659
rect 10275 27625 10284 27659
rect 10232 27616 10284 27625
rect 1952 27523 2004 27532
rect 1952 27489 1961 27523
rect 1961 27489 1995 27523
rect 1995 27489 2004 27523
rect 1952 27480 2004 27489
rect 7012 27548 7064 27600
rect 9588 27548 9640 27600
rect 10876 27523 10928 27532
rect 10876 27489 10885 27523
rect 10885 27489 10919 27523
rect 10919 27489 10928 27523
rect 10876 27480 10928 27489
rect 2964 27412 3016 27464
rect 7748 27455 7800 27464
rect 7748 27421 7757 27455
rect 7757 27421 7791 27455
rect 7791 27421 7800 27455
rect 7748 27412 7800 27421
rect 7932 27455 7984 27464
rect 7932 27421 7939 27455
rect 7939 27421 7984 27455
rect 7932 27412 7984 27421
rect 8024 27455 8076 27464
rect 8024 27421 8033 27455
rect 8033 27421 8067 27455
rect 8067 27421 8076 27455
rect 8024 27412 8076 27421
rect 9404 27412 9456 27464
rect 9772 27455 9824 27464
rect 9772 27421 9781 27455
rect 9781 27421 9815 27455
rect 9815 27421 9824 27455
rect 13820 27480 13872 27532
rect 9772 27412 9824 27421
rect 5172 27344 5224 27396
rect 10692 27387 10744 27396
rect 5724 27276 5776 27328
rect 7196 27319 7248 27328
rect 7196 27285 7205 27319
rect 7205 27285 7239 27319
rect 7239 27285 7248 27319
rect 7196 27276 7248 27285
rect 8024 27276 8076 27328
rect 8576 27276 8628 27328
rect 10692 27353 10701 27387
rect 10701 27353 10735 27387
rect 10735 27353 10744 27387
rect 10692 27344 10744 27353
rect 9956 27276 10008 27328
rect 11520 27412 11572 27464
rect 14556 27455 14608 27464
rect 13452 27344 13504 27396
rect 13084 27276 13136 27328
rect 14004 27276 14056 27328
rect 14096 27276 14148 27328
rect 14556 27421 14565 27455
rect 14565 27421 14599 27455
rect 14599 27421 14608 27455
rect 14556 27412 14608 27421
rect 19340 27616 19392 27668
rect 21272 27616 21324 27668
rect 25044 27616 25096 27668
rect 26792 27616 26844 27668
rect 20352 27548 20404 27600
rect 14740 27455 14792 27464
rect 14740 27421 14749 27455
rect 14749 27421 14783 27455
rect 14783 27421 14792 27455
rect 14740 27412 14792 27421
rect 16580 27412 16632 27464
rect 17408 27412 17460 27464
rect 19800 27480 19852 27532
rect 17960 27455 18012 27464
rect 17960 27421 17969 27455
rect 17969 27421 18003 27455
rect 18003 27421 18012 27455
rect 17960 27412 18012 27421
rect 19892 27455 19944 27464
rect 19892 27421 19901 27455
rect 19901 27421 19935 27455
rect 19935 27421 19944 27455
rect 19892 27412 19944 27421
rect 19984 27412 20036 27464
rect 17224 27276 17276 27328
rect 17500 27319 17552 27328
rect 17500 27285 17509 27319
rect 17509 27285 17543 27319
rect 17543 27285 17552 27319
rect 17500 27276 17552 27285
rect 17684 27276 17736 27328
rect 19800 27344 19852 27396
rect 20260 27455 20312 27464
rect 20260 27421 20269 27455
rect 20269 27421 20303 27455
rect 20303 27421 20312 27455
rect 20260 27412 20312 27421
rect 27896 27412 27948 27464
rect 20352 27344 20404 27396
rect 26976 27344 27028 27396
rect 20260 27276 20312 27328
rect 22468 27319 22520 27328
rect 22468 27285 22477 27319
rect 22477 27285 22511 27319
rect 22511 27285 22520 27319
rect 22468 27276 22520 27285
rect 23204 27276 23256 27328
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 50294 27174 50346 27226
rect 50358 27174 50410 27226
rect 50422 27174 50474 27226
rect 50486 27174 50538 27226
rect 50550 27174 50602 27226
rect 1952 27072 2004 27124
rect 4620 27072 4672 27124
rect 5172 27072 5224 27124
rect 5816 27004 5868 27056
rect 7104 27004 7156 27056
rect 9404 27072 9456 27124
rect 9680 27072 9732 27124
rect 10692 27072 10744 27124
rect 11612 27072 11664 27124
rect 13452 27115 13504 27124
rect 13452 27081 13461 27115
rect 13461 27081 13495 27115
rect 13495 27081 13504 27115
rect 13452 27072 13504 27081
rect 14372 27072 14424 27124
rect 18236 27072 18288 27124
rect 3148 26936 3200 26988
rect 5724 26936 5776 26988
rect 2964 26868 3016 26920
rect 6276 26868 6328 26920
rect 4712 26732 4764 26784
rect 7932 26800 7984 26852
rect 7656 26732 7708 26784
rect 10048 26936 10100 26988
rect 14740 27004 14792 27056
rect 17500 27004 17552 27056
rect 12164 26800 12216 26852
rect 13820 26979 13872 26988
rect 13820 26945 13829 26979
rect 13829 26945 13863 26979
rect 13863 26945 13872 26979
rect 13820 26936 13872 26945
rect 13912 26979 13964 26988
rect 13912 26945 13921 26979
rect 13921 26945 13955 26979
rect 13955 26945 13964 26979
rect 13912 26936 13964 26945
rect 14096 26979 14148 26988
rect 14096 26945 14105 26979
rect 14105 26945 14139 26979
rect 14139 26945 14148 26979
rect 17684 26979 17736 26988
rect 14096 26936 14148 26945
rect 17684 26945 17693 26979
rect 17693 26945 17727 26979
rect 17727 26945 17736 26979
rect 17684 26936 17736 26945
rect 19984 27072 20036 27124
rect 25136 27072 25188 27124
rect 26976 27072 27028 27124
rect 23572 27004 23624 27056
rect 25320 27004 25372 27056
rect 12992 26911 13044 26920
rect 12992 26877 13001 26911
rect 13001 26877 13035 26911
rect 13035 26877 13044 26911
rect 12992 26868 13044 26877
rect 13084 26868 13136 26920
rect 14556 26868 14608 26920
rect 17132 26868 17184 26920
rect 20168 26979 20220 26988
rect 20168 26945 20177 26979
rect 20177 26945 20211 26979
rect 20211 26945 20220 26979
rect 20168 26936 20220 26945
rect 21272 26979 21324 26988
rect 20352 26868 20404 26920
rect 21272 26945 21281 26979
rect 21281 26945 21315 26979
rect 21315 26945 21324 26979
rect 21272 26936 21324 26945
rect 25780 26936 25832 26988
rect 23572 26911 23624 26920
rect 16304 26800 16356 26852
rect 10876 26775 10928 26784
rect 10876 26741 10885 26775
rect 10885 26741 10919 26775
rect 10919 26741 10928 26775
rect 10876 26732 10928 26741
rect 14372 26732 14424 26784
rect 18328 26732 18380 26784
rect 18972 26732 19024 26784
rect 23572 26877 23581 26911
rect 23581 26877 23615 26911
rect 23615 26877 23624 26911
rect 23572 26868 23624 26877
rect 23756 26732 23808 26784
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 65654 26630 65706 26682
rect 65718 26630 65770 26682
rect 65782 26630 65834 26682
rect 65846 26630 65898 26682
rect 65910 26630 65962 26682
rect 7104 26571 7156 26580
rect 7104 26537 7113 26571
rect 7113 26537 7147 26571
rect 7147 26537 7156 26571
rect 7104 26528 7156 26537
rect 7196 26528 7248 26580
rect 10876 26528 10928 26580
rect 14280 26528 14332 26580
rect 4712 26460 4764 26512
rect 7564 26460 7616 26512
rect 9588 26460 9640 26512
rect 17408 26528 17460 26580
rect 21272 26528 21324 26580
rect 25320 26528 25372 26580
rect 36820 26571 36872 26580
rect 36820 26537 36829 26571
rect 36829 26537 36863 26571
rect 36863 26537 36872 26571
rect 36820 26528 36872 26537
rect 17132 26503 17184 26512
rect 5724 26256 5776 26308
rect 7656 26324 7708 26376
rect 10784 26367 10836 26376
rect 10784 26333 10793 26367
rect 10793 26333 10827 26367
rect 10827 26333 10836 26367
rect 10784 26324 10836 26333
rect 11244 26392 11296 26444
rect 17132 26469 17141 26503
rect 17141 26469 17175 26503
rect 17175 26469 17184 26503
rect 17132 26460 17184 26469
rect 10048 26231 10100 26240
rect 10048 26197 10057 26231
rect 10057 26197 10091 26231
rect 10091 26197 10100 26231
rect 10048 26188 10100 26197
rect 12900 26324 12952 26376
rect 13268 26324 13320 26376
rect 12164 26256 12216 26308
rect 14096 26392 14148 26444
rect 14188 26324 14240 26376
rect 15568 26324 15620 26376
rect 16580 26324 16632 26376
rect 17684 26324 17736 26376
rect 21456 26324 21508 26376
rect 25320 26367 25372 26376
rect 25320 26333 25329 26367
rect 25329 26333 25363 26367
rect 25363 26333 25372 26367
rect 25780 26367 25832 26376
rect 25320 26324 25372 26333
rect 25780 26333 25789 26367
rect 25789 26333 25823 26367
rect 25823 26333 25832 26367
rect 25780 26324 25832 26333
rect 32220 26367 32272 26376
rect 32220 26333 32229 26367
rect 32229 26333 32263 26367
rect 32263 26333 32272 26367
rect 32220 26324 32272 26333
rect 32404 26324 32456 26376
rect 35164 26367 35216 26376
rect 11060 26188 11112 26240
rect 11428 26231 11480 26240
rect 11428 26197 11437 26231
rect 11437 26197 11471 26231
rect 11471 26197 11480 26231
rect 11428 26188 11480 26197
rect 15844 26256 15896 26308
rect 17040 26256 17092 26308
rect 19248 26256 19300 26308
rect 20168 26256 20220 26308
rect 20536 26256 20588 26308
rect 35164 26333 35173 26367
rect 35173 26333 35207 26367
rect 35207 26333 35216 26367
rect 35164 26324 35216 26333
rect 35440 26256 35492 26308
rect 35808 26367 35860 26376
rect 35808 26333 35817 26367
rect 35817 26333 35851 26367
rect 35851 26333 35860 26367
rect 35808 26324 35860 26333
rect 36084 26367 36136 26376
rect 36084 26333 36093 26367
rect 36093 26333 36127 26367
rect 36127 26333 36136 26367
rect 36084 26324 36136 26333
rect 68100 26367 68152 26376
rect 68100 26333 68109 26367
rect 68109 26333 68143 26367
rect 68143 26333 68152 26367
rect 68100 26324 68152 26333
rect 37740 26256 37792 26308
rect 33232 26231 33284 26240
rect 33232 26197 33241 26231
rect 33241 26197 33275 26231
rect 33275 26197 33284 26231
rect 33232 26188 33284 26197
rect 34060 26231 34112 26240
rect 34060 26197 34069 26231
rect 34069 26197 34103 26231
rect 34103 26197 34112 26231
rect 34060 26188 34112 26197
rect 35348 26231 35400 26240
rect 35348 26197 35357 26231
rect 35357 26197 35391 26231
rect 35391 26197 35400 26231
rect 35348 26188 35400 26197
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 50294 26086 50346 26138
rect 50358 26086 50410 26138
rect 50422 26086 50474 26138
rect 50486 26086 50538 26138
rect 50550 26086 50602 26138
rect 3148 26027 3200 26036
rect 3148 25993 3157 26027
rect 3157 25993 3191 26027
rect 3191 25993 3200 26027
rect 3148 25984 3200 25993
rect 3424 25984 3476 26036
rect 7656 25984 7708 26036
rect 10692 25984 10744 26036
rect 14188 25984 14240 26036
rect 19248 26027 19300 26036
rect 19248 25993 19257 26027
rect 19257 25993 19291 26027
rect 19291 25993 19300 26027
rect 19248 25984 19300 25993
rect 34796 26027 34848 26036
rect 34796 25993 34805 26027
rect 34805 25993 34839 26027
rect 34839 25993 34848 26027
rect 34796 25984 34848 25993
rect 35164 25984 35216 26036
rect 2320 25891 2372 25900
rect 2320 25857 2329 25891
rect 2329 25857 2363 25891
rect 2363 25857 2372 25891
rect 2320 25848 2372 25857
rect 2504 25891 2556 25900
rect 2504 25857 2513 25891
rect 2513 25857 2547 25891
rect 2547 25857 2556 25891
rect 2504 25848 2556 25857
rect 3403 25891 3455 25900
rect 3403 25857 3421 25891
rect 3421 25857 3455 25891
rect 3403 25848 3455 25857
rect 3608 25891 3660 25900
rect 3608 25857 3617 25891
rect 3617 25857 3651 25891
rect 3651 25857 3660 25891
rect 3608 25848 3660 25857
rect 3332 25712 3384 25764
rect 3240 25644 3292 25696
rect 6276 25780 6328 25832
rect 6644 25891 6696 25900
rect 6644 25857 6678 25891
rect 6678 25857 6696 25891
rect 11428 25916 11480 25968
rect 33232 25916 33284 25968
rect 34060 25916 34112 25968
rect 6644 25848 6696 25857
rect 8760 25848 8812 25900
rect 11520 25891 11572 25900
rect 11520 25857 11529 25891
rect 11529 25857 11563 25891
rect 11563 25857 11572 25891
rect 11520 25848 11572 25857
rect 15384 25848 15436 25900
rect 16580 25848 16632 25900
rect 16672 25891 16724 25900
rect 16672 25857 16681 25891
rect 16681 25857 16715 25891
rect 16715 25857 16724 25891
rect 16672 25848 16724 25857
rect 17684 25848 17736 25900
rect 17960 25848 18012 25900
rect 20352 25848 20404 25900
rect 22468 25848 22520 25900
rect 23480 25848 23532 25900
rect 23848 25891 23900 25900
rect 23848 25857 23857 25891
rect 23857 25857 23891 25891
rect 23891 25857 23900 25891
rect 23848 25848 23900 25857
rect 25136 25848 25188 25900
rect 35348 25891 35400 25900
rect 35348 25857 35357 25891
rect 35357 25857 35391 25891
rect 35391 25857 35400 25891
rect 35348 25848 35400 25857
rect 19984 25780 20036 25832
rect 23572 25780 23624 25832
rect 24768 25780 24820 25832
rect 33048 25823 33100 25832
rect 33048 25789 33057 25823
rect 33057 25789 33091 25823
rect 33091 25789 33100 25823
rect 33048 25780 33100 25789
rect 3884 25712 3936 25764
rect 4988 25712 5040 25764
rect 19248 25712 19300 25764
rect 7656 25644 7708 25696
rect 10048 25687 10100 25696
rect 10048 25653 10057 25687
rect 10057 25653 10091 25687
rect 10091 25653 10100 25687
rect 10048 25644 10100 25653
rect 13268 25644 13320 25696
rect 14280 25644 14332 25696
rect 15936 25644 15988 25696
rect 16856 25687 16908 25696
rect 16856 25653 16865 25687
rect 16865 25653 16899 25687
rect 16899 25653 16908 25687
rect 16856 25644 16908 25653
rect 21916 25644 21968 25696
rect 22284 25644 22336 25696
rect 24400 25644 24452 25696
rect 24584 25687 24636 25696
rect 24584 25653 24593 25687
rect 24593 25653 24627 25687
rect 24627 25653 24636 25687
rect 24584 25644 24636 25653
rect 26056 25644 26108 25696
rect 32220 25644 32272 25696
rect 34704 25644 34756 25696
rect 35808 25644 35860 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 65654 25542 65706 25594
rect 65718 25542 65770 25594
rect 65782 25542 65834 25594
rect 65846 25542 65898 25594
rect 65910 25542 65962 25594
rect 2504 25440 2556 25492
rect 3332 25440 3384 25492
rect 6644 25440 6696 25492
rect 8760 25440 8812 25492
rect 15384 25440 15436 25492
rect 17960 25440 18012 25492
rect 23848 25440 23900 25492
rect 25136 25483 25188 25492
rect 10784 25372 10836 25424
rect 2964 25236 3016 25288
rect 4712 25236 4764 25288
rect 4160 25211 4212 25220
rect 4160 25177 4194 25211
rect 4194 25177 4212 25211
rect 4160 25168 4212 25177
rect 7012 25276 7064 25288
rect 7012 25242 7021 25276
rect 7021 25242 7055 25276
rect 7055 25242 7064 25276
rect 7012 25236 7064 25242
rect 7472 25236 7524 25288
rect 7656 25236 7708 25288
rect 7932 25279 7984 25288
rect 7932 25245 7941 25279
rect 7941 25245 7975 25279
rect 7975 25245 7984 25279
rect 7932 25236 7984 25245
rect 11244 25304 11296 25356
rect 8116 25279 8168 25288
rect 8116 25245 8125 25279
rect 8125 25245 8159 25279
rect 8159 25245 8168 25279
rect 8116 25236 8168 25245
rect 10140 25236 10192 25288
rect 10692 25279 10744 25288
rect 10692 25245 10701 25279
rect 10701 25245 10735 25279
rect 10735 25245 10744 25279
rect 10692 25236 10744 25245
rect 10784 25168 10836 25220
rect 14924 25236 14976 25288
rect 24676 25372 24728 25424
rect 25136 25449 25145 25483
rect 25145 25449 25179 25483
rect 25179 25449 25188 25483
rect 25136 25440 25188 25449
rect 15660 25304 15712 25356
rect 15292 25168 15344 25220
rect 5264 25143 5316 25152
rect 5264 25109 5273 25143
rect 5273 25109 5307 25143
rect 5307 25109 5316 25143
rect 6000 25143 6052 25152
rect 5264 25100 5316 25109
rect 6000 25109 6009 25143
rect 6009 25109 6043 25143
rect 6043 25109 6052 25143
rect 6000 25100 6052 25109
rect 6828 25100 6880 25152
rect 7472 25100 7524 25152
rect 8300 25100 8352 25152
rect 13820 25100 13872 25152
rect 15936 25279 15988 25288
rect 15936 25245 15945 25279
rect 15945 25245 15979 25279
rect 15979 25245 15988 25279
rect 17132 25279 17184 25288
rect 15936 25236 15988 25245
rect 17132 25245 17141 25279
rect 17141 25245 17175 25279
rect 17175 25245 17184 25279
rect 17132 25236 17184 25245
rect 17316 25279 17368 25288
rect 17316 25245 17325 25279
rect 17325 25245 17359 25279
rect 17359 25245 17368 25279
rect 17316 25236 17368 25245
rect 19984 25304 20036 25356
rect 20720 25279 20772 25288
rect 20720 25245 20729 25279
rect 20729 25245 20763 25279
rect 20763 25245 20772 25279
rect 20720 25236 20772 25245
rect 21456 25236 21508 25288
rect 24216 25236 24268 25288
rect 34796 25372 34848 25424
rect 32220 25304 32272 25356
rect 27896 25279 27948 25288
rect 23480 25211 23532 25220
rect 19340 25100 19392 25152
rect 21272 25100 21324 25152
rect 23480 25177 23489 25211
rect 23489 25177 23523 25211
rect 23523 25177 23532 25211
rect 23480 25168 23532 25177
rect 23664 25211 23716 25220
rect 23664 25177 23673 25211
rect 23673 25177 23707 25211
rect 23707 25177 23716 25211
rect 23664 25168 23716 25177
rect 23848 25168 23900 25220
rect 24584 25168 24636 25220
rect 27896 25245 27905 25279
rect 27905 25245 27939 25279
rect 27939 25245 27948 25279
rect 27896 25236 27948 25245
rect 28356 25236 28408 25288
rect 30656 25236 30708 25288
rect 34244 25304 34296 25356
rect 36084 25440 36136 25492
rect 35348 25279 35400 25288
rect 26240 25168 26292 25220
rect 22560 25143 22612 25152
rect 22560 25109 22569 25143
rect 22569 25109 22603 25143
rect 22603 25109 22612 25143
rect 22560 25100 22612 25109
rect 35348 25245 35357 25279
rect 35357 25245 35391 25279
rect 35391 25245 35400 25279
rect 35348 25236 35400 25245
rect 35900 25236 35952 25288
rect 33508 25168 33560 25220
rect 36728 25211 36780 25220
rect 36728 25177 36737 25211
rect 36737 25177 36771 25211
rect 36771 25177 36780 25211
rect 36728 25168 36780 25177
rect 37464 25168 37516 25220
rect 35440 25100 35492 25152
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 50294 24998 50346 25050
rect 50358 24998 50410 25050
rect 50422 24998 50474 25050
rect 50486 24998 50538 25050
rect 50550 24998 50602 25050
rect 3332 24896 3384 24948
rect 7012 24939 7064 24948
rect 2320 24828 2372 24880
rect 7012 24905 7021 24939
rect 7021 24905 7055 24939
rect 7055 24905 7064 24939
rect 7012 24896 7064 24905
rect 7932 24896 7984 24948
rect 6000 24828 6052 24880
rect 8116 24828 8168 24880
rect 3240 24803 3292 24812
rect 3240 24769 3249 24803
rect 3249 24769 3283 24803
rect 3283 24769 3292 24803
rect 3240 24760 3292 24769
rect 3700 24760 3752 24812
rect 7196 24803 7248 24812
rect 7196 24769 7205 24803
rect 7205 24769 7239 24803
rect 7239 24769 7248 24803
rect 7196 24760 7248 24769
rect 15476 24896 15528 24948
rect 15936 24896 15988 24948
rect 17316 24939 17368 24948
rect 17316 24905 17325 24939
rect 17325 24905 17359 24939
rect 17359 24905 17368 24939
rect 17316 24896 17368 24905
rect 20444 24896 20496 24948
rect 15292 24828 15344 24880
rect 14556 24803 14608 24812
rect 4160 24692 4212 24744
rect 4620 24624 4672 24676
rect 5264 24624 5316 24676
rect 2320 24556 2372 24608
rect 7196 24624 7248 24676
rect 6828 24556 6880 24608
rect 8668 24556 8720 24608
rect 13268 24692 13320 24744
rect 11060 24624 11112 24676
rect 10048 24556 10100 24608
rect 10968 24556 11020 24608
rect 14556 24769 14565 24803
rect 14565 24769 14599 24803
rect 14599 24769 14608 24803
rect 14556 24760 14608 24769
rect 15016 24760 15068 24812
rect 15200 24803 15252 24812
rect 15200 24769 15209 24803
rect 15209 24769 15243 24803
rect 15243 24769 15252 24803
rect 15200 24760 15252 24769
rect 15660 24828 15712 24880
rect 16856 24828 16908 24880
rect 17684 24828 17736 24880
rect 16028 24760 16080 24812
rect 17040 24760 17092 24812
rect 18328 24803 18380 24812
rect 18328 24769 18337 24803
rect 18337 24769 18371 24803
rect 18371 24769 18380 24803
rect 18328 24760 18380 24769
rect 18420 24760 18472 24812
rect 20168 24803 20220 24812
rect 20168 24769 20177 24803
rect 20177 24769 20211 24803
rect 20211 24769 20220 24803
rect 20168 24760 20220 24769
rect 20352 24803 20404 24812
rect 20352 24769 20361 24803
rect 20361 24769 20395 24803
rect 20395 24769 20404 24803
rect 20352 24760 20404 24769
rect 24492 24896 24544 24948
rect 20720 24828 20772 24880
rect 24676 24896 24728 24948
rect 34244 24939 34296 24948
rect 34244 24905 34253 24939
rect 34253 24905 34287 24939
rect 34287 24905 34296 24939
rect 34244 24896 34296 24905
rect 36728 24896 36780 24948
rect 21824 24803 21876 24812
rect 15844 24735 15896 24744
rect 15844 24701 15853 24735
rect 15853 24701 15887 24735
rect 15887 24701 15896 24735
rect 15844 24692 15896 24701
rect 15936 24692 15988 24744
rect 17684 24692 17736 24744
rect 21824 24769 21833 24803
rect 21833 24769 21867 24803
rect 21867 24769 21876 24803
rect 21824 24760 21876 24769
rect 22008 24803 22060 24812
rect 22008 24769 22017 24803
rect 22017 24769 22051 24803
rect 22051 24769 22060 24803
rect 22008 24760 22060 24769
rect 22192 24803 22244 24812
rect 22192 24769 22201 24803
rect 22201 24769 22235 24803
rect 22235 24769 22244 24803
rect 22192 24760 22244 24769
rect 22560 24760 22612 24812
rect 23756 24803 23808 24812
rect 23756 24769 23765 24803
rect 23765 24769 23799 24803
rect 23799 24769 23808 24803
rect 23756 24760 23808 24769
rect 24216 24760 24268 24812
rect 24400 24760 24452 24812
rect 20720 24692 20772 24744
rect 22468 24692 22520 24744
rect 23940 24692 23992 24744
rect 28448 24760 28500 24812
rect 26240 24692 26292 24744
rect 28356 24735 28408 24744
rect 28356 24701 28365 24735
rect 28365 24701 28399 24735
rect 28399 24701 28408 24735
rect 28356 24692 28408 24701
rect 33140 24760 33192 24812
rect 34796 24828 34848 24880
rect 39948 24828 40000 24880
rect 33692 24760 33744 24812
rect 34428 24803 34480 24812
rect 34428 24769 34437 24803
rect 34437 24769 34471 24803
rect 34471 24769 34480 24803
rect 34428 24760 34480 24769
rect 37464 24760 37516 24812
rect 37740 24803 37792 24812
rect 37740 24769 37749 24803
rect 37749 24769 37783 24803
rect 37783 24769 37792 24803
rect 37740 24760 37792 24769
rect 38936 24760 38988 24812
rect 43260 24760 43312 24812
rect 32680 24692 32732 24744
rect 34704 24692 34756 24744
rect 36268 24692 36320 24744
rect 38660 24692 38712 24744
rect 41788 24692 41840 24744
rect 42892 24735 42944 24744
rect 42892 24701 42901 24735
rect 42901 24701 42935 24735
rect 42935 24701 42944 24735
rect 42892 24692 42944 24701
rect 16212 24624 16264 24676
rect 17040 24624 17092 24676
rect 19340 24624 19392 24676
rect 24676 24624 24728 24676
rect 32404 24667 32456 24676
rect 32404 24633 32413 24667
rect 32413 24633 32447 24667
rect 32447 24633 32456 24667
rect 32404 24624 32456 24633
rect 67640 24667 67692 24676
rect 67640 24633 67649 24667
rect 67649 24633 67683 24667
rect 67683 24633 67692 24667
rect 67640 24624 67692 24633
rect 16672 24556 16724 24608
rect 19432 24556 19484 24608
rect 20168 24556 20220 24608
rect 21824 24556 21876 24608
rect 22468 24599 22520 24608
rect 22468 24565 22477 24599
rect 22477 24565 22511 24599
rect 22511 24565 22520 24599
rect 22468 24556 22520 24565
rect 22744 24556 22796 24608
rect 23388 24599 23440 24608
rect 23388 24565 23397 24599
rect 23397 24565 23431 24599
rect 23431 24565 23440 24599
rect 23388 24556 23440 24565
rect 23664 24556 23716 24608
rect 26056 24556 26108 24608
rect 29736 24599 29788 24608
rect 29736 24565 29745 24599
rect 29745 24565 29779 24599
rect 29779 24565 29788 24599
rect 29736 24556 29788 24565
rect 32772 24556 32824 24608
rect 33508 24599 33560 24608
rect 33508 24565 33517 24599
rect 33517 24565 33551 24599
rect 33551 24565 33560 24599
rect 33508 24556 33560 24565
rect 35440 24556 35492 24608
rect 41144 24556 41196 24608
rect 56324 24556 56376 24608
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 65654 24454 65706 24506
rect 65718 24454 65770 24506
rect 65782 24454 65834 24506
rect 65846 24454 65898 24506
rect 65910 24454 65962 24506
rect 5632 24352 5684 24404
rect 8024 24395 8076 24404
rect 8024 24361 8033 24395
rect 8033 24361 8067 24395
rect 8067 24361 8076 24395
rect 8024 24352 8076 24361
rect 13084 24395 13136 24404
rect 13084 24361 13093 24395
rect 13093 24361 13127 24395
rect 13127 24361 13136 24395
rect 13084 24352 13136 24361
rect 15292 24352 15344 24404
rect 15936 24352 15988 24404
rect 16028 24395 16080 24404
rect 16028 24361 16037 24395
rect 16037 24361 16071 24395
rect 16071 24361 16080 24395
rect 16028 24352 16080 24361
rect 17408 24352 17460 24404
rect 2964 24216 3016 24268
rect 6276 24148 6328 24200
rect 5540 24123 5592 24132
rect 5540 24089 5574 24123
rect 5574 24089 5592 24123
rect 5540 24080 5592 24089
rect 3700 24012 3752 24064
rect 5264 24012 5316 24064
rect 9772 24284 9824 24336
rect 15660 24284 15712 24336
rect 16488 24284 16540 24336
rect 11520 24216 11572 24268
rect 7932 24148 7984 24200
rect 8116 24191 8168 24200
rect 8116 24157 8125 24191
rect 8125 24157 8159 24191
rect 8159 24157 8168 24191
rect 8116 24148 8168 24157
rect 7472 24055 7524 24064
rect 7472 24021 7481 24055
rect 7481 24021 7515 24055
rect 7515 24021 7524 24055
rect 7472 24012 7524 24021
rect 8852 24012 8904 24064
rect 9128 24191 9180 24200
rect 9128 24157 9137 24191
rect 9137 24157 9171 24191
rect 9171 24157 9180 24191
rect 9128 24148 9180 24157
rect 9588 24148 9640 24200
rect 14648 24148 14700 24200
rect 16212 24148 16264 24200
rect 16764 24148 16816 24200
rect 17224 24148 17276 24200
rect 17684 24284 17736 24336
rect 18420 24352 18472 24404
rect 20352 24352 20404 24404
rect 20444 24395 20496 24404
rect 20444 24361 20453 24395
rect 20453 24361 20487 24395
rect 20487 24361 20496 24395
rect 20444 24352 20496 24361
rect 22008 24352 22060 24404
rect 24676 24352 24728 24404
rect 32680 24352 32732 24404
rect 34428 24352 34480 24404
rect 35348 24395 35400 24404
rect 35348 24361 35357 24395
rect 35357 24361 35391 24395
rect 35391 24361 35400 24395
rect 35348 24352 35400 24361
rect 39948 24395 40000 24404
rect 39948 24361 39957 24395
rect 39957 24361 39991 24395
rect 39991 24361 40000 24395
rect 39948 24352 40000 24361
rect 41788 24395 41840 24404
rect 41788 24361 41797 24395
rect 41797 24361 41831 24395
rect 41831 24361 41840 24395
rect 41788 24352 41840 24361
rect 43260 24395 43312 24404
rect 43260 24361 43269 24395
rect 43269 24361 43303 24395
rect 43303 24361 43312 24395
rect 43260 24352 43312 24361
rect 20076 24216 20128 24268
rect 17684 24191 17736 24200
rect 17684 24157 17693 24191
rect 17693 24157 17727 24191
rect 17727 24157 17736 24191
rect 17684 24148 17736 24157
rect 17868 24148 17920 24200
rect 19984 24191 20036 24200
rect 19984 24157 19993 24191
rect 19993 24157 20027 24191
rect 20027 24157 20036 24191
rect 19984 24148 20036 24157
rect 20168 24148 20220 24200
rect 9404 24080 9456 24132
rect 11796 24080 11848 24132
rect 13544 24080 13596 24132
rect 19432 24080 19484 24132
rect 9680 24012 9732 24064
rect 11152 24055 11204 24064
rect 11152 24021 11161 24055
rect 11161 24021 11195 24055
rect 11195 24021 11204 24055
rect 11152 24012 11204 24021
rect 16580 24012 16632 24064
rect 17224 24012 17276 24064
rect 17684 24012 17736 24064
rect 22192 24284 22244 24336
rect 35440 24284 35492 24336
rect 20628 24216 20680 24268
rect 21272 24191 21324 24200
rect 21272 24157 21281 24191
rect 21281 24157 21315 24191
rect 21315 24157 21324 24191
rect 21272 24148 21324 24157
rect 34796 24216 34848 24268
rect 22468 24148 22520 24200
rect 24768 24148 24820 24200
rect 28356 24148 28408 24200
rect 29368 24148 29420 24200
rect 31024 24148 31076 24200
rect 32772 24191 32824 24200
rect 32772 24157 32781 24191
rect 32781 24157 32815 24191
rect 32815 24157 32824 24191
rect 38660 24191 38712 24200
rect 32772 24148 32824 24157
rect 38660 24157 38669 24191
rect 38669 24157 38703 24191
rect 38703 24157 38712 24191
rect 38660 24148 38712 24157
rect 38936 24148 38988 24200
rect 40040 24148 40092 24200
rect 41144 24191 41196 24200
rect 41144 24157 41153 24191
rect 41153 24157 41187 24191
rect 41187 24157 41196 24191
rect 41144 24148 41196 24157
rect 42524 24191 42576 24200
rect 42524 24157 42533 24191
rect 42533 24157 42567 24191
rect 42567 24157 42576 24191
rect 42524 24148 42576 24157
rect 42892 24148 42944 24200
rect 43260 24191 43312 24200
rect 43260 24157 43269 24191
rect 43269 24157 43303 24191
rect 43303 24157 43312 24191
rect 43260 24148 43312 24157
rect 24124 24080 24176 24132
rect 24676 24080 24728 24132
rect 24860 24080 24912 24132
rect 27068 24123 27120 24132
rect 27068 24089 27102 24123
rect 27102 24089 27120 24123
rect 27068 24080 27120 24089
rect 30288 24080 30340 24132
rect 32220 24080 32272 24132
rect 37924 24080 37976 24132
rect 21732 24012 21784 24064
rect 25964 24012 26016 24064
rect 27804 24012 27856 24064
rect 29920 24012 29972 24064
rect 36452 24012 36504 24064
rect 42432 24012 42484 24064
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 50294 23910 50346 23962
rect 50358 23910 50410 23962
rect 50422 23910 50474 23962
rect 50486 23910 50538 23962
rect 50550 23910 50602 23962
rect 3424 23808 3476 23860
rect 4344 23851 4396 23860
rect 4344 23817 4353 23851
rect 4353 23817 4387 23851
rect 4387 23817 4396 23851
rect 4344 23808 4396 23817
rect 5540 23851 5592 23860
rect 5540 23817 5549 23851
rect 5549 23817 5583 23851
rect 5583 23817 5592 23851
rect 5540 23808 5592 23817
rect 9404 23851 9456 23860
rect 7472 23740 7524 23792
rect 2136 23715 2188 23724
rect 2136 23681 2145 23715
rect 2145 23681 2179 23715
rect 2179 23681 2188 23715
rect 2136 23672 2188 23681
rect 2320 23715 2372 23724
rect 2320 23681 2329 23715
rect 2329 23681 2363 23715
rect 2363 23681 2372 23715
rect 2320 23672 2372 23681
rect 2504 23715 2556 23724
rect 2504 23681 2513 23715
rect 2513 23681 2547 23715
rect 2547 23681 2556 23715
rect 4896 23715 4948 23724
rect 2504 23672 2556 23681
rect 4896 23681 4905 23715
rect 4905 23681 4939 23715
rect 4939 23681 4948 23715
rect 4896 23672 4948 23681
rect 5080 23715 5132 23724
rect 5080 23681 5089 23715
rect 5089 23681 5123 23715
rect 5123 23681 5132 23715
rect 5080 23672 5132 23681
rect 2688 23604 2740 23656
rect 2964 23647 3016 23656
rect 2964 23613 2973 23647
rect 2973 23613 3007 23647
rect 3007 23613 3016 23647
rect 2964 23604 3016 23613
rect 5264 23715 5316 23724
rect 5264 23681 5273 23715
rect 5273 23681 5307 23715
rect 5307 23681 5316 23715
rect 5264 23672 5316 23681
rect 7840 23672 7892 23724
rect 8300 23715 8352 23724
rect 8300 23681 8309 23715
rect 8309 23681 8343 23715
rect 8343 23681 8352 23715
rect 8300 23672 8352 23681
rect 8484 23672 8536 23724
rect 9404 23817 9413 23851
rect 9413 23817 9447 23851
rect 9447 23817 9456 23851
rect 9404 23808 9456 23817
rect 9680 23808 9732 23860
rect 13820 23808 13872 23860
rect 9864 23740 9916 23792
rect 16488 23740 16540 23792
rect 8852 23672 8904 23724
rect 9039 23715 9091 23724
rect 9039 23681 9064 23715
rect 9064 23681 9091 23715
rect 9039 23672 9091 23681
rect 5264 23536 5316 23588
rect 7656 23511 7708 23520
rect 7656 23477 7665 23511
rect 7665 23477 7699 23511
rect 7699 23477 7708 23511
rect 7656 23468 7708 23477
rect 8668 23604 8720 23656
rect 11152 23672 11204 23724
rect 9772 23604 9824 23656
rect 12992 23604 13044 23656
rect 13360 23604 13412 23656
rect 16212 23672 16264 23724
rect 16580 23672 16632 23724
rect 16856 23715 16908 23724
rect 16856 23681 16865 23715
rect 16865 23681 16899 23715
rect 16899 23681 16908 23715
rect 16856 23672 16908 23681
rect 20628 23808 20680 23860
rect 22376 23851 22428 23860
rect 22376 23817 22385 23851
rect 22385 23817 22419 23851
rect 22419 23817 22428 23851
rect 22376 23808 22428 23817
rect 24860 23851 24912 23860
rect 24860 23817 24869 23851
rect 24869 23817 24903 23851
rect 24903 23817 24912 23851
rect 24860 23808 24912 23817
rect 21640 23740 21692 23792
rect 21916 23783 21968 23792
rect 21916 23749 21925 23783
rect 21925 23749 21959 23783
rect 21959 23749 21968 23783
rect 21916 23740 21968 23749
rect 23480 23740 23532 23792
rect 18788 23715 18840 23724
rect 14280 23604 14332 23656
rect 15200 23604 15252 23656
rect 15568 23604 15620 23656
rect 8760 23468 8812 23520
rect 16580 23536 16632 23588
rect 16672 23536 16724 23588
rect 16948 23536 17000 23588
rect 18788 23681 18797 23715
rect 18797 23681 18831 23715
rect 18831 23681 18840 23715
rect 18788 23672 18840 23681
rect 19340 23672 19392 23724
rect 12072 23468 12124 23520
rect 14372 23511 14424 23520
rect 14372 23477 14381 23511
rect 14381 23477 14415 23511
rect 14415 23477 14424 23511
rect 14372 23468 14424 23477
rect 15936 23468 15988 23520
rect 17684 23536 17736 23588
rect 20628 23672 20680 23724
rect 22192 23715 22244 23724
rect 22192 23681 22201 23715
rect 22201 23681 22235 23715
rect 22235 23681 22244 23715
rect 22192 23672 22244 23681
rect 23296 23672 23348 23724
rect 24216 23715 24268 23724
rect 20168 23604 20220 23656
rect 24216 23681 24225 23715
rect 24225 23681 24259 23715
rect 24259 23681 24268 23715
rect 24216 23672 24268 23681
rect 24492 23715 24544 23724
rect 24492 23681 24501 23715
rect 24501 23681 24535 23715
rect 24535 23681 24544 23715
rect 24492 23672 24544 23681
rect 24676 23672 24728 23724
rect 29644 23715 29696 23724
rect 29644 23681 29653 23715
rect 29653 23681 29687 23715
rect 29687 23681 29696 23715
rect 29644 23672 29696 23681
rect 29828 23715 29880 23724
rect 29828 23681 29837 23715
rect 29837 23681 29871 23715
rect 29871 23681 29880 23715
rect 29828 23672 29880 23681
rect 30104 23808 30156 23860
rect 30288 23851 30340 23860
rect 30288 23817 30297 23851
rect 30297 23817 30331 23851
rect 30331 23817 30340 23851
rect 30288 23808 30340 23817
rect 37924 23851 37976 23860
rect 37924 23817 37933 23851
rect 37933 23817 37967 23851
rect 37967 23817 37976 23851
rect 37924 23808 37976 23817
rect 42800 23808 42852 23860
rect 43260 23808 43312 23860
rect 34060 23715 34112 23724
rect 25964 23604 26016 23656
rect 34060 23681 34069 23715
rect 34069 23681 34103 23715
rect 34103 23681 34112 23715
rect 34060 23672 34112 23681
rect 36452 23715 36504 23724
rect 23112 23536 23164 23588
rect 33876 23604 33928 23656
rect 36452 23681 36461 23715
rect 36461 23681 36495 23715
rect 36495 23681 36504 23715
rect 36452 23672 36504 23681
rect 37280 23715 37332 23724
rect 37280 23681 37289 23715
rect 37289 23681 37323 23715
rect 37323 23681 37332 23715
rect 37280 23672 37332 23681
rect 37648 23715 37700 23724
rect 37648 23681 37657 23715
rect 37657 23681 37691 23715
rect 37691 23681 37700 23715
rect 37648 23672 37700 23681
rect 42432 23715 42484 23724
rect 41604 23604 41656 23656
rect 42432 23681 42441 23715
rect 42441 23681 42475 23715
rect 42475 23681 42484 23715
rect 42432 23672 42484 23681
rect 37464 23536 37516 23588
rect 17592 23468 17644 23520
rect 17868 23468 17920 23520
rect 20076 23511 20128 23520
rect 20076 23477 20085 23511
rect 20085 23477 20119 23511
rect 20119 23477 20128 23511
rect 20076 23468 20128 23477
rect 21732 23468 21784 23520
rect 28264 23468 28316 23520
rect 29460 23468 29512 23520
rect 33784 23468 33836 23520
rect 33968 23468 34020 23520
rect 41696 23468 41748 23520
rect 67548 23468 67600 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 65654 23366 65706 23418
rect 65718 23366 65770 23418
rect 65782 23366 65834 23418
rect 65846 23366 65898 23418
rect 65910 23366 65962 23418
rect 2320 23264 2372 23316
rect 5080 23264 5132 23316
rect 5632 23307 5684 23316
rect 5632 23273 5641 23307
rect 5641 23273 5675 23307
rect 5675 23273 5684 23307
rect 5632 23264 5684 23273
rect 5264 23196 5316 23248
rect 9036 23264 9088 23316
rect 11796 23307 11848 23316
rect 6276 23171 6328 23180
rect 6276 23137 6285 23171
rect 6285 23137 6319 23171
rect 6319 23137 6328 23171
rect 6276 23128 6328 23137
rect 8944 23171 8996 23180
rect 8944 23137 8953 23171
rect 8953 23137 8987 23171
rect 8987 23137 8996 23171
rect 8944 23128 8996 23137
rect 9128 23128 9180 23180
rect 11796 23273 11805 23307
rect 11805 23273 11839 23307
rect 11839 23273 11848 23307
rect 11796 23264 11848 23273
rect 13544 23307 13596 23316
rect 13544 23273 13553 23307
rect 13553 23273 13587 23307
rect 13587 23273 13596 23307
rect 13544 23264 13596 23273
rect 16856 23264 16908 23316
rect 3424 23060 3476 23112
rect 2228 22992 2280 23044
rect 6368 23060 6420 23112
rect 7656 23060 7708 23112
rect 8208 23060 8260 23112
rect 11336 23103 11388 23112
rect 11336 23069 11345 23103
rect 11345 23069 11379 23103
rect 11379 23069 11388 23103
rect 11336 23060 11388 23069
rect 12348 23128 12400 23180
rect 12624 23128 12676 23180
rect 12808 23128 12860 23180
rect 19340 23264 19392 23316
rect 21916 23264 21968 23316
rect 22192 23264 22244 23316
rect 23112 23307 23164 23316
rect 23112 23273 23121 23307
rect 23121 23273 23155 23307
rect 23155 23273 23164 23307
rect 23112 23264 23164 23273
rect 27068 23264 27120 23316
rect 29828 23264 29880 23316
rect 26332 23196 26384 23248
rect 34060 23264 34112 23316
rect 33508 23196 33560 23248
rect 36084 23264 36136 23316
rect 37648 23307 37700 23316
rect 37648 23273 37657 23307
rect 37657 23273 37691 23307
rect 37691 23273 37700 23307
rect 37648 23264 37700 23273
rect 41604 23307 41656 23316
rect 41604 23273 41613 23307
rect 41613 23273 41647 23307
rect 41647 23273 41656 23307
rect 41604 23264 41656 23273
rect 5632 22992 5684 23044
rect 5816 22992 5868 23044
rect 7840 22992 7892 23044
rect 12256 23103 12308 23112
rect 12256 23069 12270 23103
rect 12270 23069 12304 23103
rect 12304 23069 12308 23103
rect 12256 23060 12308 23069
rect 12440 23103 12492 23112
rect 12440 23069 12449 23103
rect 12449 23069 12483 23103
rect 12483 23069 12492 23103
rect 12440 23060 12492 23069
rect 13084 23103 13136 23112
rect 13084 23069 13093 23103
rect 13093 23069 13127 23103
rect 13127 23069 13136 23103
rect 13084 23060 13136 23069
rect 13360 23060 13412 23112
rect 18328 23128 18380 23180
rect 21824 23128 21876 23180
rect 24216 23128 24268 23180
rect 33048 23128 33100 23180
rect 14372 23060 14424 23112
rect 14648 23060 14700 23112
rect 15108 23060 15160 23112
rect 20076 23060 20128 23112
rect 27252 23103 27304 23112
rect 16212 23035 16264 23044
rect 2136 22924 2188 22976
rect 3332 22924 3384 22976
rect 6000 22924 6052 22976
rect 7380 22924 7432 22976
rect 8116 22924 8168 22976
rect 16212 23001 16221 23035
rect 16221 23001 16255 23035
rect 16255 23001 16264 23035
rect 16212 22992 16264 23001
rect 17592 23035 17644 23044
rect 17592 23001 17626 23035
rect 17626 23001 17644 23035
rect 8668 22924 8720 22976
rect 17592 22992 17644 23001
rect 19984 22992 20036 23044
rect 20444 22992 20496 23044
rect 27252 23069 27261 23103
rect 27261 23069 27295 23103
rect 27295 23069 27304 23103
rect 27252 23060 27304 23069
rect 27436 23100 27488 23112
rect 27436 23066 27445 23100
rect 27445 23066 27479 23100
rect 27479 23066 27488 23100
rect 27436 23060 27488 23066
rect 27620 23103 27672 23112
rect 27620 23069 27629 23103
rect 27629 23069 27663 23103
rect 27663 23069 27672 23103
rect 27620 23060 27672 23069
rect 28632 23060 28684 23112
rect 29092 23060 29144 23112
rect 29920 23060 29972 23112
rect 33784 23103 33836 23112
rect 33784 23069 33793 23103
rect 33793 23069 33827 23103
rect 33827 23069 33836 23103
rect 33784 23060 33836 23069
rect 23296 23035 23348 23044
rect 23296 23001 23305 23035
rect 23305 23001 23339 23035
rect 23339 23001 23348 23035
rect 23296 22992 23348 23001
rect 23480 23035 23532 23044
rect 23480 23001 23489 23035
rect 23489 23001 23523 23035
rect 23523 23001 23532 23035
rect 23480 22992 23532 23001
rect 25044 23035 25096 23044
rect 25044 23001 25053 23035
rect 25053 23001 25087 23035
rect 25087 23001 25096 23035
rect 25044 22992 25096 23001
rect 17960 22924 18012 22976
rect 23388 22924 23440 22976
rect 27160 22924 27212 22976
rect 28264 22992 28316 23044
rect 29368 22992 29420 23044
rect 30472 22992 30524 23044
rect 33968 23103 34020 23112
rect 33968 23069 33977 23103
rect 33977 23069 34011 23103
rect 34011 23069 34020 23103
rect 33968 23060 34020 23069
rect 34152 23103 34204 23112
rect 34152 23069 34161 23103
rect 34161 23069 34195 23103
rect 34195 23069 34204 23103
rect 34152 23060 34204 23069
rect 35900 23060 35952 23112
rect 38660 23060 38712 23112
rect 39856 23103 39908 23112
rect 39856 23069 39865 23103
rect 39865 23069 39899 23103
rect 39899 23069 39908 23103
rect 39856 23060 39908 23069
rect 43352 23103 43404 23112
rect 43352 23069 43361 23103
rect 43361 23069 43395 23103
rect 43395 23069 43404 23103
rect 43352 23060 43404 23069
rect 43628 23103 43680 23112
rect 43628 23069 43637 23103
rect 43637 23069 43671 23103
rect 43671 23069 43680 23103
rect 43628 23060 43680 23069
rect 34428 22992 34480 23044
rect 34796 22992 34848 23044
rect 35624 22992 35676 23044
rect 36912 23035 36964 23044
rect 36912 23001 36921 23035
rect 36921 23001 36955 23035
rect 36955 23001 36964 23035
rect 36912 22992 36964 23001
rect 40132 22992 40184 23044
rect 27988 22924 28040 22976
rect 29920 22924 29972 22976
rect 30012 22924 30064 22976
rect 33600 22924 33652 22976
rect 34152 22924 34204 22976
rect 37372 22924 37424 22976
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 50294 22822 50346 22874
rect 50358 22822 50410 22874
rect 50422 22822 50474 22874
rect 50486 22822 50538 22874
rect 50550 22822 50602 22874
rect 3424 22720 3476 22772
rect 12256 22720 12308 22772
rect 2228 22695 2280 22704
rect 2228 22661 2237 22695
rect 2237 22661 2271 22695
rect 2271 22661 2280 22695
rect 2228 22652 2280 22661
rect 2688 22652 2740 22704
rect 5264 22652 5316 22704
rect 2596 22423 2648 22432
rect 2596 22389 2605 22423
rect 2605 22389 2639 22423
rect 2639 22389 2648 22423
rect 2596 22380 2648 22389
rect 5080 22584 5132 22636
rect 6276 22652 6328 22704
rect 9588 22652 9640 22704
rect 12716 22720 12768 22772
rect 12992 22720 13044 22772
rect 13084 22720 13136 22772
rect 14280 22720 14332 22772
rect 17776 22763 17828 22772
rect 5632 22627 5684 22636
rect 5632 22593 5641 22627
rect 5641 22593 5675 22627
rect 5675 22593 5684 22627
rect 5632 22584 5684 22593
rect 5908 22584 5960 22636
rect 7472 22584 7524 22636
rect 9404 22584 9456 22636
rect 10876 22584 10928 22636
rect 17776 22729 17785 22763
rect 17785 22729 17819 22763
rect 17819 22729 17828 22763
rect 17776 22720 17828 22729
rect 12532 22627 12584 22636
rect 12532 22593 12541 22627
rect 12541 22593 12575 22627
rect 12575 22593 12584 22627
rect 12532 22584 12584 22593
rect 15200 22584 15252 22636
rect 15568 22584 15620 22636
rect 15844 22584 15896 22636
rect 17132 22627 17184 22636
rect 17132 22593 17141 22627
rect 17141 22593 17175 22627
rect 17175 22593 17184 22627
rect 17132 22584 17184 22593
rect 17224 22627 17276 22636
rect 17224 22593 17234 22627
rect 17234 22593 17268 22627
rect 17268 22593 17276 22627
rect 17224 22584 17276 22593
rect 17500 22627 17552 22636
rect 17500 22593 17509 22627
rect 17509 22593 17543 22627
rect 17543 22593 17552 22627
rect 17500 22584 17552 22593
rect 17868 22584 17920 22636
rect 19340 22584 19392 22636
rect 19984 22627 20036 22636
rect 19984 22593 19993 22627
rect 19993 22593 20027 22627
rect 20027 22593 20036 22627
rect 19984 22584 20036 22593
rect 15292 22516 15344 22568
rect 22836 22720 22888 22772
rect 24032 22720 24084 22772
rect 22284 22652 22336 22704
rect 22652 22627 22704 22636
rect 22652 22593 22656 22627
rect 22656 22593 22690 22627
rect 22690 22593 22704 22627
rect 22652 22584 22704 22593
rect 22836 22627 22888 22636
rect 22836 22593 22845 22627
rect 22845 22593 22879 22627
rect 22879 22593 22888 22627
rect 22836 22584 22888 22593
rect 23940 22695 23992 22704
rect 23940 22661 23949 22695
rect 23949 22661 23983 22695
rect 23983 22661 23992 22695
rect 23940 22652 23992 22661
rect 4620 22380 4672 22432
rect 5172 22423 5224 22432
rect 5172 22389 5181 22423
rect 5181 22389 5215 22423
rect 5215 22389 5224 22423
rect 5172 22380 5224 22389
rect 9312 22380 9364 22432
rect 11336 22448 11388 22500
rect 20260 22448 20312 22500
rect 11060 22380 11112 22432
rect 12808 22380 12860 22432
rect 22836 22380 22888 22432
rect 23480 22584 23532 22636
rect 24860 22652 24912 22704
rect 24768 22584 24820 22636
rect 27436 22720 27488 22772
rect 28448 22720 28500 22772
rect 28908 22720 28960 22772
rect 29552 22720 29604 22772
rect 34796 22763 34848 22772
rect 34796 22729 34805 22763
rect 34805 22729 34839 22763
rect 34839 22729 34848 22763
rect 34796 22720 34848 22729
rect 35808 22720 35860 22772
rect 36912 22720 36964 22772
rect 40132 22763 40184 22772
rect 40132 22729 40141 22763
rect 40141 22729 40175 22763
rect 40175 22729 40184 22763
rect 40132 22720 40184 22729
rect 42892 22720 42944 22772
rect 43628 22720 43680 22772
rect 26056 22695 26108 22704
rect 26056 22661 26065 22695
rect 26065 22661 26099 22695
rect 26099 22661 26108 22695
rect 26056 22652 26108 22661
rect 27160 22695 27212 22704
rect 27160 22661 27169 22695
rect 27169 22661 27203 22695
rect 27203 22661 27212 22695
rect 27160 22652 27212 22661
rect 27804 22652 27856 22704
rect 27988 22652 28040 22704
rect 25136 22627 25188 22636
rect 25136 22593 25145 22627
rect 25145 22593 25179 22627
rect 25179 22593 25188 22627
rect 25136 22584 25188 22593
rect 25780 22584 25832 22636
rect 25872 22584 25924 22636
rect 26148 22627 26200 22636
rect 26148 22593 26157 22627
rect 26157 22593 26191 22627
rect 26191 22593 26200 22627
rect 26148 22584 26200 22593
rect 26332 22627 26384 22636
rect 26332 22593 26341 22627
rect 26341 22593 26375 22627
rect 26375 22593 26384 22627
rect 26976 22627 27028 22636
rect 26332 22584 26384 22593
rect 26976 22593 26985 22627
rect 26985 22593 27019 22627
rect 27019 22593 27028 22627
rect 26976 22584 27028 22593
rect 29184 22652 29236 22704
rect 35900 22652 35952 22704
rect 38660 22652 38712 22704
rect 29000 22627 29052 22636
rect 23388 22380 23440 22432
rect 23572 22423 23624 22432
rect 23572 22389 23581 22423
rect 23581 22389 23615 22423
rect 23615 22389 23624 22423
rect 23572 22380 23624 22389
rect 29000 22593 29009 22627
rect 29009 22593 29043 22627
rect 29043 22593 29052 22627
rect 29000 22584 29052 22593
rect 30012 22627 30064 22636
rect 29552 22516 29604 22568
rect 29644 22516 29696 22568
rect 30012 22593 30021 22627
rect 30021 22593 30055 22627
rect 30055 22593 30064 22627
rect 30012 22584 30064 22593
rect 30104 22627 30156 22636
rect 30104 22593 30113 22627
rect 30113 22593 30147 22627
rect 30147 22593 30156 22627
rect 30104 22584 30156 22593
rect 30288 22584 30340 22636
rect 33508 22627 33560 22636
rect 33508 22593 33517 22627
rect 33517 22593 33551 22627
rect 33551 22593 33560 22627
rect 33508 22584 33560 22593
rect 33876 22584 33928 22636
rect 34152 22627 34204 22636
rect 34152 22593 34161 22627
rect 34161 22593 34195 22627
rect 34195 22593 34204 22627
rect 34152 22584 34204 22593
rect 34428 22627 34480 22636
rect 34428 22593 34437 22627
rect 34437 22593 34471 22627
rect 34471 22593 34480 22627
rect 34428 22584 34480 22593
rect 34796 22584 34848 22636
rect 35348 22584 35400 22636
rect 38752 22627 38804 22636
rect 38752 22593 38770 22627
rect 38770 22593 38804 22627
rect 38752 22584 38804 22593
rect 40040 22627 40092 22636
rect 40040 22593 40049 22627
rect 40049 22593 40083 22627
rect 40083 22593 40092 22627
rect 40040 22584 40092 22593
rect 41696 22627 41748 22636
rect 41696 22593 41705 22627
rect 41705 22593 41739 22627
rect 41739 22593 41748 22627
rect 41696 22584 41748 22593
rect 41880 22627 41932 22636
rect 41880 22593 41889 22627
rect 41889 22593 41923 22627
rect 41923 22593 41932 22627
rect 41880 22584 41932 22593
rect 42432 22584 42484 22636
rect 42616 22627 42668 22636
rect 42616 22593 42625 22627
rect 42625 22593 42659 22627
rect 42659 22593 42668 22627
rect 42616 22584 42668 22593
rect 42800 22627 42852 22636
rect 42800 22593 42809 22627
rect 42809 22593 42843 22627
rect 42843 22593 42852 22627
rect 42800 22584 42852 22593
rect 33876 22448 33928 22500
rect 35624 22448 35676 22500
rect 32128 22380 32180 22432
rect 33784 22380 33836 22432
rect 36636 22380 36688 22432
rect 42064 22380 42116 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 65654 22278 65706 22330
rect 65718 22278 65770 22330
rect 65782 22278 65834 22330
rect 65846 22278 65898 22330
rect 65910 22278 65962 22330
rect 5632 22176 5684 22228
rect 8300 22176 8352 22228
rect 9036 22176 9088 22228
rect 10876 22219 10928 22228
rect 2596 22108 2648 22160
rect 2688 22108 2740 22160
rect 2412 22015 2464 22024
rect 2412 21981 2421 22015
rect 2421 21981 2455 22015
rect 2455 21981 2464 22015
rect 2412 21972 2464 21981
rect 2964 22040 3016 22092
rect 3240 21972 3292 22024
rect 5172 21972 5224 22024
rect 7932 22040 7984 22092
rect 8944 22083 8996 22092
rect 8944 22049 8953 22083
rect 8953 22049 8987 22083
rect 8987 22049 8996 22083
rect 10876 22185 10885 22219
rect 10885 22185 10919 22219
rect 10919 22185 10928 22219
rect 10876 22176 10928 22185
rect 11060 22176 11112 22228
rect 13452 22176 13504 22228
rect 12808 22108 12860 22160
rect 8944 22040 8996 22049
rect 3148 21836 3200 21888
rect 8300 21972 8352 22024
rect 8760 21972 8812 22024
rect 6368 21947 6420 21956
rect 6368 21913 6377 21947
rect 6377 21913 6411 21947
rect 6411 21913 6420 21947
rect 6368 21904 6420 21913
rect 8116 21904 8168 21956
rect 7196 21879 7248 21888
rect 7196 21845 7205 21879
rect 7205 21845 7239 21879
rect 7239 21845 7248 21879
rect 7196 21836 7248 21845
rect 8484 21836 8536 21888
rect 8944 21836 8996 21888
rect 10600 22015 10652 22024
rect 10600 21981 10609 22015
rect 10609 21981 10643 22015
rect 10643 21981 10652 22015
rect 10600 21972 10652 21981
rect 12440 21972 12492 22024
rect 13176 22040 13228 22092
rect 14740 22176 14792 22228
rect 15016 22176 15068 22228
rect 19432 22176 19484 22228
rect 20076 22176 20128 22228
rect 22652 22176 22704 22228
rect 23480 22176 23532 22228
rect 35808 22219 35860 22228
rect 35808 22185 35817 22219
rect 35817 22185 35851 22219
rect 35851 22185 35860 22219
rect 35808 22176 35860 22185
rect 12072 21947 12124 21956
rect 12072 21913 12081 21947
rect 12081 21913 12115 21947
rect 12115 21913 12124 21947
rect 12072 21904 12124 21913
rect 12348 21904 12400 21956
rect 15108 21972 15160 22024
rect 16212 22015 16264 22024
rect 16212 21981 16221 22015
rect 16221 21981 16255 22015
rect 16255 21981 16264 22015
rect 16212 21972 16264 21981
rect 14924 21904 14976 21956
rect 16396 22015 16448 22024
rect 16396 21981 16405 22015
rect 16405 21981 16439 22015
rect 16439 21981 16448 22015
rect 16580 22015 16632 22024
rect 16396 21972 16448 21981
rect 16580 21981 16589 22015
rect 16589 21981 16623 22015
rect 16623 21981 16632 22015
rect 16580 21972 16632 21981
rect 17592 21972 17644 22024
rect 15200 21836 15252 21888
rect 15752 21836 15804 21888
rect 15936 21879 15988 21888
rect 15936 21845 15945 21879
rect 15945 21845 15979 21879
rect 15979 21845 15988 21879
rect 15936 21836 15988 21845
rect 17592 21879 17644 21888
rect 17592 21845 17601 21879
rect 17601 21845 17635 21879
rect 17635 21845 17644 21879
rect 17592 21836 17644 21845
rect 17960 22040 18012 22092
rect 18880 21972 18932 22024
rect 19432 22015 19484 22024
rect 19432 21981 19436 22015
rect 19436 21981 19470 22015
rect 19470 21981 19484 22015
rect 19432 21972 19484 21981
rect 26976 22108 27028 22160
rect 29920 22108 29972 22160
rect 28172 22040 28224 22092
rect 29552 22083 29604 22092
rect 29552 22049 29561 22083
rect 29561 22049 29595 22083
rect 29595 22049 29604 22083
rect 29552 22040 29604 22049
rect 34796 22040 34848 22092
rect 35440 22040 35492 22092
rect 35992 22108 36044 22160
rect 19340 21904 19392 21956
rect 19984 21972 20036 22024
rect 20536 21972 20588 22024
rect 21824 22015 21876 22024
rect 21824 21981 21833 22015
rect 21833 21981 21867 22015
rect 21867 21981 21876 22015
rect 21824 21972 21876 21981
rect 21916 22015 21968 22024
rect 21916 21981 21925 22015
rect 21925 21981 21959 22015
rect 21959 21981 21968 22015
rect 22192 22015 22244 22024
rect 21916 21972 21968 21981
rect 22192 21981 22201 22015
rect 22201 21981 22235 22015
rect 22235 21981 22244 22015
rect 22192 21972 22244 21981
rect 22928 21972 22980 22024
rect 23020 22015 23072 22024
rect 23020 21981 23029 22015
rect 23029 21981 23063 22015
rect 23063 21981 23072 22015
rect 23020 21972 23072 21981
rect 18512 21836 18564 21888
rect 20996 21904 21048 21956
rect 22468 21904 22520 21956
rect 24768 21972 24820 22024
rect 25872 22015 25924 22024
rect 25872 21981 25881 22015
rect 25881 21981 25915 22015
rect 25915 21981 25924 22015
rect 25872 21972 25924 21981
rect 25964 22015 26016 22024
rect 25964 21981 25973 22015
rect 25973 21981 26007 22015
rect 26007 21981 26016 22015
rect 25964 21972 26016 21981
rect 27988 22015 28040 22024
rect 20260 21836 20312 21888
rect 21548 21836 21600 21888
rect 25136 21904 25188 21956
rect 26148 21904 26200 21956
rect 23204 21836 23256 21888
rect 23664 21836 23716 21888
rect 24492 21879 24544 21888
rect 24492 21845 24501 21879
rect 24501 21845 24535 21879
rect 24535 21845 24544 21879
rect 24492 21836 24544 21845
rect 27988 21981 27997 22015
rect 27997 21981 28031 22015
rect 28031 21981 28040 22015
rect 27988 21972 28040 21981
rect 29920 22015 29972 22024
rect 29920 21981 29929 22015
rect 29929 21981 29963 22015
rect 29963 21981 29972 22015
rect 29920 21972 29972 21981
rect 30288 21972 30340 22024
rect 31668 21972 31720 22024
rect 32128 22015 32180 22024
rect 32128 21981 32146 22015
rect 32146 21981 32180 22015
rect 32128 21972 32180 21981
rect 32404 22015 32456 22024
rect 32404 21981 32413 22015
rect 32413 21981 32447 22015
rect 32447 21981 32456 22015
rect 32404 21972 32456 21981
rect 68100 22151 68152 22160
rect 68100 22117 68109 22151
rect 68109 22117 68143 22151
rect 68143 22117 68152 22151
rect 68100 22108 68152 22117
rect 36452 22040 36504 22092
rect 38752 22040 38804 22092
rect 39856 22083 39908 22092
rect 39856 22049 39865 22083
rect 39865 22049 39899 22083
rect 39899 22049 39908 22083
rect 39856 22040 39908 22049
rect 27620 21904 27672 21956
rect 29736 21947 29788 21956
rect 29736 21913 29745 21947
rect 29745 21913 29779 21947
rect 29779 21913 29788 21947
rect 29736 21904 29788 21913
rect 37372 22015 37424 22024
rect 35532 21904 35584 21956
rect 37372 21981 37381 22015
rect 37381 21981 37415 22015
rect 37415 21981 37424 22015
rect 37372 21972 37424 21981
rect 37464 22015 37516 22024
rect 37464 21981 37473 22015
rect 37473 21981 37507 22015
rect 37507 21981 37516 22015
rect 37464 21972 37516 21981
rect 38384 21972 38436 22024
rect 42064 22015 42116 22024
rect 42064 21981 42073 22015
rect 42073 21981 42107 22015
rect 42107 21981 42116 22015
rect 42064 21972 42116 21981
rect 37280 21904 37332 21956
rect 38200 21904 38252 21956
rect 30472 21836 30524 21888
rect 35348 21836 35400 21888
rect 36544 21836 36596 21888
rect 41788 21836 41840 21888
rect 42524 21836 42576 21888
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 50294 21734 50346 21786
rect 50358 21734 50410 21786
rect 50422 21734 50474 21786
rect 50486 21734 50538 21786
rect 50550 21734 50602 21786
rect 5816 21632 5868 21684
rect 10508 21632 10560 21684
rect 10600 21632 10652 21684
rect 12624 21632 12676 21684
rect 16212 21632 16264 21684
rect 16396 21632 16448 21684
rect 17684 21632 17736 21684
rect 20168 21632 20220 21684
rect 20996 21632 21048 21684
rect 2964 21496 3016 21548
rect 3148 21539 3200 21548
rect 3148 21505 3182 21539
rect 3182 21505 3200 21539
rect 3148 21496 3200 21505
rect 6644 21539 6696 21548
rect 6644 21505 6678 21539
rect 6678 21505 6696 21539
rect 8208 21539 8260 21548
rect 6644 21496 6696 21505
rect 8208 21505 8217 21539
rect 8217 21505 8251 21539
rect 8251 21505 8260 21539
rect 8208 21496 8260 21505
rect 8300 21496 8352 21548
rect 9036 21539 9088 21548
rect 9036 21505 9045 21539
rect 9045 21505 9079 21539
rect 9079 21505 9088 21539
rect 9036 21496 9088 21505
rect 12256 21564 12308 21616
rect 5540 21428 5592 21480
rect 7840 21428 7892 21480
rect 8760 21428 8812 21480
rect 10232 21496 10284 21548
rect 11704 21496 11756 21548
rect 9680 21428 9732 21480
rect 12440 21496 12492 21548
rect 12900 21564 12952 21616
rect 17224 21564 17276 21616
rect 19800 21564 19852 21616
rect 20076 21607 20128 21616
rect 20076 21573 20085 21607
rect 20085 21573 20119 21607
rect 20119 21573 20128 21607
rect 20076 21564 20128 21573
rect 13176 21496 13228 21548
rect 15568 21539 15620 21548
rect 15568 21505 15577 21539
rect 15577 21505 15611 21539
rect 15611 21505 15620 21539
rect 15568 21496 15620 21505
rect 15752 21539 15804 21548
rect 15752 21505 15761 21539
rect 15761 21505 15795 21539
rect 15795 21505 15804 21539
rect 15752 21496 15804 21505
rect 16028 21496 16080 21548
rect 16764 21496 16816 21548
rect 17868 21539 17920 21548
rect 12256 21428 12308 21480
rect 17868 21505 17877 21539
rect 17877 21505 17911 21539
rect 17911 21505 17920 21539
rect 17868 21496 17920 21505
rect 19064 21496 19116 21548
rect 19432 21496 19484 21548
rect 20260 21496 20312 21548
rect 23388 21564 23440 21616
rect 23480 21564 23532 21616
rect 23940 21564 23992 21616
rect 20444 21539 20496 21548
rect 20444 21505 20453 21539
rect 20453 21505 20487 21539
rect 20487 21505 20496 21539
rect 20904 21539 20956 21548
rect 20444 21496 20496 21505
rect 20904 21505 20913 21539
rect 20913 21505 20947 21539
rect 20947 21505 20956 21539
rect 20904 21496 20956 21505
rect 16580 21428 16632 21480
rect 17224 21428 17276 21480
rect 19156 21428 19208 21480
rect 22376 21496 22428 21548
rect 23020 21496 23072 21548
rect 23572 21496 23624 21548
rect 24308 21539 24360 21548
rect 24308 21505 24317 21539
rect 24317 21505 24351 21539
rect 24351 21505 24360 21539
rect 24308 21496 24360 21505
rect 25596 21564 25648 21616
rect 27896 21564 27948 21616
rect 24676 21539 24728 21548
rect 24676 21505 24685 21539
rect 24685 21505 24719 21539
rect 24719 21505 24728 21539
rect 24676 21496 24728 21505
rect 24860 21496 24912 21548
rect 27712 21539 27764 21548
rect 22468 21428 22520 21480
rect 27712 21505 27721 21539
rect 27721 21505 27755 21539
rect 27755 21505 27764 21539
rect 27712 21496 27764 21505
rect 29092 21632 29144 21684
rect 32496 21632 32548 21684
rect 35992 21632 36044 21684
rect 38200 21675 38252 21684
rect 38200 21641 38209 21675
rect 38209 21641 38243 21675
rect 38243 21641 38252 21675
rect 38200 21632 38252 21641
rect 42616 21632 42668 21684
rect 43352 21632 43404 21684
rect 32956 21564 33008 21616
rect 28632 21539 28684 21548
rect 28632 21505 28641 21539
rect 28641 21505 28675 21539
rect 28675 21505 28684 21539
rect 28632 21496 28684 21505
rect 28724 21496 28776 21548
rect 27620 21428 27672 21480
rect 29000 21496 29052 21548
rect 29368 21496 29420 21548
rect 30288 21496 30340 21548
rect 32312 21496 32364 21548
rect 32404 21496 32456 21548
rect 33048 21496 33100 21548
rect 34428 21496 34480 21548
rect 37464 21496 37516 21548
rect 37740 21539 37792 21548
rect 29184 21428 29236 21480
rect 34704 21428 34756 21480
rect 9588 21360 9640 21412
rect 4620 21292 4672 21344
rect 7288 21292 7340 21344
rect 8392 21292 8444 21344
rect 9680 21335 9732 21344
rect 9680 21301 9689 21335
rect 9689 21301 9723 21335
rect 9723 21301 9732 21335
rect 9680 21292 9732 21301
rect 10232 21335 10284 21344
rect 10232 21301 10241 21335
rect 10241 21301 10275 21335
rect 10275 21301 10284 21335
rect 10232 21292 10284 21301
rect 11704 21292 11756 21344
rect 17592 21360 17644 21412
rect 19340 21360 19392 21412
rect 20260 21360 20312 21412
rect 22192 21360 22244 21412
rect 30104 21360 30156 21412
rect 14832 21292 14884 21344
rect 15844 21292 15896 21344
rect 16580 21292 16632 21344
rect 17316 21292 17368 21344
rect 20076 21292 20128 21344
rect 21916 21292 21968 21344
rect 24032 21335 24084 21344
rect 24032 21301 24041 21335
rect 24041 21301 24075 21335
rect 24075 21301 24084 21335
rect 24032 21292 24084 21301
rect 27804 21335 27856 21344
rect 27804 21301 27813 21335
rect 27813 21301 27847 21335
rect 27847 21301 27856 21335
rect 27804 21292 27856 21301
rect 30840 21292 30892 21344
rect 30932 21292 30984 21344
rect 32772 21292 32824 21344
rect 33600 21292 33652 21344
rect 37280 21428 37332 21480
rect 37740 21505 37749 21539
rect 37749 21505 37783 21539
rect 37783 21505 37792 21539
rect 37740 21496 37792 21505
rect 42524 21564 42576 21616
rect 41236 21539 41288 21548
rect 41236 21505 41245 21539
rect 41245 21505 41279 21539
rect 41279 21505 41288 21539
rect 41236 21496 41288 21505
rect 41604 21496 41656 21548
rect 42432 21539 42484 21548
rect 42432 21505 42441 21539
rect 42441 21505 42475 21539
rect 42475 21505 42484 21539
rect 42432 21496 42484 21505
rect 42800 21496 42852 21548
rect 41420 21471 41472 21480
rect 41420 21437 41429 21471
rect 41429 21437 41463 21471
rect 41463 21437 41472 21471
rect 41420 21428 41472 21437
rect 36360 21292 36412 21344
rect 37832 21292 37884 21344
rect 41604 21292 41656 21344
rect 41880 21292 41932 21344
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 65654 21190 65706 21242
rect 65718 21190 65770 21242
rect 65782 21190 65834 21242
rect 65846 21190 65898 21242
rect 65910 21190 65962 21242
rect 6552 21088 6604 21140
rect 6644 21088 6696 21140
rect 7748 21088 7800 21140
rect 3240 21063 3292 21072
rect 3240 21029 3249 21063
rect 3249 21029 3283 21063
rect 3283 21029 3292 21063
rect 3240 21020 3292 21029
rect 3424 21020 3476 21072
rect 7288 21020 7340 21072
rect 8760 21088 8812 21140
rect 8484 21020 8536 21072
rect 9312 21020 9364 21072
rect 16856 21088 16908 21140
rect 17132 21088 17184 21140
rect 20444 21088 20496 21140
rect 27712 21131 27764 21140
rect 21364 21020 21416 21072
rect 21916 21020 21968 21072
rect 24676 21020 24728 21072
rect 27712 21097 27721 21131
rect 27721 21097 27755 21131
rect 27755 21097 27764 21131
rect 27712 21088 27764 21097
rect 28724 21088 28776 21140
rect 28908 21131 28960 21140
rect 28908 21097 28917 21131
rect 28917 21097 28951 21131
rect 28951 21097 28960 21131
rect 28908 21088 28960 21097
rect 29920 21088 29972 21140
rect 33692 21088 33744 21140
rect 34060 21088 34112 21140
rect 37740 21088 37792 21140
rect 38016 21088 38068 21140
rect 42432 21088 42484 21140
rect 35532 21020 35584 21072
rect 4620 20952 4672 21004
rect 6920 20952 6972 21004
rect 1492 20884 1544 20936
rect 1860 20927 1912 20936
rect 1860 20893 1869 20927
rect 1869 20893 1903 20927
rect 1903 20893 1912 20927
rect 1860 20884 1912 20893
rect 5540 20748 5592 20800
rect 5724 20748 5776 20800
rect 7288 20927 7340 20936
rect 9036 20952 9088 21004
rect 7288 20893 7302 20927
rect 7302 20893 7336 20927
rect 7336 20893 7340 20927
rect 7288 20884 7340 20893
rect 8116 20927 8168 20936
rect 8116 20893 8125 20927
rect 8125 20893 8159 20927
rect 8159 20893 8168 20927
rect 8116 20884 8168 20893
rect 7840 20816 7892 20868
rect 7748 20748 7800 20800
rect 8300 20884 8352 20936
rect 8668 20884 8720 20936
rect 9680 20884 9732 20936
rect 11612 20927 11664 20936
rect 11612 20893 11621 20927
rect 11621 20893 11655 20927
rect 11655 20893 11664 20927
rect 11612 20884 11664 20893
rect 11704 20884 11756 20936
rect 14004 20884 14056 20936
rect 8392 20859 8444 20868
rect 8392 20825 8401 20859
rect 8401 20825 8435 20859
rect 8435 20825 8444 20859
rect 8392 20816 8444 20825
rect 8852 20816 8904 20868
rect 10508 20816 10560 20868
rect 14648 20884 14700 20936
rect 15292 20927 15344 20936
rect 15292 20893 15301 20927
rect 15301 20893 15335 20927
rect 15335 20893 15344 20927
rect 15292 20884 15344 20893
rect 15936 20884 15988 20936
rect 18788 20952 18840 21004
rect 18880 20952 18932 21004
rect 17960 20927 18012 20936
rect 17960 20893 17969 20927
rect 17969 20893 18003 20927
rect 18003 20893 18012 20927
rect 18144 20927 18196 20936
rect 17960 20884 18012 20893
rect 18144 20893 18153 20927
rect 18153 20893 18187 20927
rect 18187 20893 18196 20927
rect 18144 20884 18196 20893
rect 18236 20927 18288 20936
rect 18236 20893 18245 20927
rect 18245 20893 18279 20927
rect 18279 20893 18288 20927
rect 19432 20927 19484 20936
rect 18236 20884 18288 20893
rect 19432 20893 19436 20927
rect 19436 20893 19470 20927
rect 19470 20893 19484 20927
rect 19432 20884 19484 20893
rect 20168 20952 20220 21004
rect 20628 20952 20680 21004
rect 19156 20816 19208 20868
rect 19340 20816 19392 20868
rect 21548 20884 21600 20936
rect 21824 20952 21876 21004
rect 20628 20816 20680 20868
rect 9404 20748 9456 20800
rect 10416 20748 10468 20800
rect 12992 20791 13044 20800
rect 12992 20757 13001 20791
rect 13001 20757 13035 20791
rect 13035 20757 13044 20791
rect 12992 20748 13044 20757
rect 15016 20748 15068 20800
rect 17132 20791 17184 20800
rect 17132 20757 17141 20791
rect 17141 20757 17175 20791
rect 17175 20757 17184 20791
rect 17132 20748 17184 20757
rect 18420 20748 18472 20800
rect 19800 20748 19852 20800
rect 20904 20748 20956 20800
rect 21732 20927 21784 20936
rect 21732 20893 21741 20927
rect 21741 20893 21775 20927
rect 21775 20893 21784 20927
rect 22008 20927 22060 20936
rect 21732 20884 21784 20893
rect 22008 20893 22017 20927
rect 22017 20893 22051 20927
rect 22051 20893 22060 20927
rect 22008 20884 22060 20893
rect 24768 20952 24820 21004
rect 27344 20952 27396 21004
rect 26240 20884 26292 20936
rect 28172 20927 28224 20936
rect 22468 20816 22520 20868
rect 23756 20816 23808 20868
rect 21732 20748 21784 20800
rect 23020 20748 23072 20800
rect 25136 20816 25188 20868
rect 25412 20859 25464 20868
rect 25412 20825 25421 20859
rect 25421 20825 25455 20859
rect 25455 20825 25464 20859
rect 25412 20816 25464 20825
rect 25596 20859 25648 20868
rect 25596 20825 25605 20859
rect 25605 20825 25639 20859
rect 25639 20825 25648 20859
rect 25596 20816 25648 20825
rect 26148 20816 26200 20868
rect 28172 20893 28181 20927
rect 28181 20893 28215 20927
rect 28215 20893 28224 20927
rect 28172 20884 28224 20893
rect 28908 20884 28960 20936
rect 29092 20884 29144 20936
rect 29552 20927 29604 20936
rect 29552 20893 29561 20927
rect 29561 20893 29595 20927
rect 29595 20893 29604 20927
rect 29552 20884 29604 20893
rect 30472 20952 30524 21004
rect 30748 20995 30800 21004
rect 30748 20961 30757 20995
rect 30757 20961 30791 20995
rect 30791 20961 30800 20995
rect 30748 20952 30800 20961
rect 28448 20816 28500 20868
rect 29920 20927 29972 20936
rect 29920 20893 29929 20927
rect 29929 20893 29963 20927
rect 29963 20893 29972 20927
rect 29920 20884 29972 20893
rect 30104 20884 30156 20936
rect 30840 20927 30892 20936
rect 30380 20816 30432 20868
rect 30564 20859 30616 20868
rect 30564 20825 30573 20859
rect 30573 20825 30607 20859
rect 30607 20825 30616 20859
rect 30564 20816 30616 20825
rect 30840 20893 30849 20927
rect 30849 20893 30883 20927
rect 30883 20893 30892 20927
rect 30840 20884 30892 20893
rect 32128 20884 32180 20936
rect 34336 20952 34388 21004
rect 35716 20952 35768 21004
rect 41420 21020 41472 21072
rect 32496 20884 32548 20936
rect 33324 20927 33376 20936
rect 33324 20893 33333 20927
rect 33333 20893 33367 20927
rect 33367 20893 33376 20927
rect 33324 20884 33376 20893
rect 33600 20927 33652 20936
rect 33600 20893 33609 20927
rect 33609 20893 33643 20927
rect 33643 20893 33652 20927
rect 33600 20884 33652 20893
rect 33692 20884 33744 20936
rect 36084 20884 36136 20936
rect 36544 20952 36596 21004
rect 40132 20952 40184 21004
rect 41696 20952 41748 21004
rect 38292 20927 38344 20936
rect 35808 20816 35860 20868
rect 25688 20748 25740 20800
rect 31760 20748 31812 20800
rect 32496 20748 32548 20800
rect 35624 20748 35676 20800
rect 38292 20893 38301 20927
rect 38301 20893 38335 20927
rect 38335 20893 38344 20927
rect 38292 20884 38344 20893
rect 41512 20927 41564 20936
rect 41512 20893 41521 20927
rect 41521 20893 41555 20927
rect 41555 20893 41564 20927
rect 41512 20884 41564 20893
rect 41604 20927 41656 20936
rect 41604 20893 41613 20927
rect 41613 20893 41647 20927
rect 41647 20893 41656 20927
rect 41604 20884 41656 20893
rect 41788 20816 41840 20868
rect 35992 20748 36044 20800
rect 41328 20791 41380 20800
rect 41328 20757 41337 20791
rect 41337 20757 41371 20791
rect 41371 20757 41380 20791
rect 41328 20748 41380 20757
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 50294 20646 50346 20698
rect 50358 20646 50410 20698
rect 50422 20646 50474 20698
rect 50486 20646 50538 20698
rect 50550 20646 50602 20698
rect 7564 20544 7616 20596
rect 8116 20544 8168 20596
rect 12256 20544 12308 20596
rect 9404 20476 9456 20528
rect 12992 20544 13044 20596
rect 12532 20519 12584 20528
rect 12532 20485 12541 20519
rect 12541 20485 12575 20519
rect 12575 20485 12584 20519
rect 12532 20476 12584 20485
rect 15200 20476 15252 20528
rect 1400 20408 1452 20460
rect 5540 20451 5592 20460
rect 5540 20417 5549 20451
rect 5549 20417 5583 20451
rect 5583 20417 5592 20451
rect 5540 20408 5592 20417
rect 8208 20408 8260 20460
rect 10140 20451 10192 20460
rect 10140 20417 10149 20451
rect 10149 20417 10183 20451
rect 10183 20417 10192 20451
rect 10140 20408 10192 20417
rect 15384 20476 15436 20528
rect 16672 20519 16724 20528
rect 16672 20485 16681 20519
rect 16681 20485 16715 20519
rect 16715 20485 16724 20519
rect 16672 20476 16724 20485
rect 17960 20544 18012 20596
rect 19064 20544 19116 20596
rect 21824 20544 21876 20596
rect 22284 20544 22336 20596
rect 18604 20476 18656 20528
rect 19340 20476 19392 20528
rect 20352 20519 20404 20528
rect 20352 20485 20361 20519
rect 20361 20485 20395 20519
rect 20395 20485 20404 20519
rect 20352 20476 20404 20485
rect 21640 20476 21692 20528
rect 15476 20451 15528 20460
rect 15476 20417 15485 20451
rect 15485 20417 15519 20451
rect 15519 20417 15528 20451
rect 15476 20408 15528 20417
rect 15752 20451 15804 20460
rect 15752 20417 15761 20451
rect 15761 20417 15795 20451
rect 15795 20417 15804 20451
rect 15752 20408 15804 20417
rect 17132 20408 17184 20460
rect 17224 20408 17276 20460
rect 17500 20408 17552 20460
rect 19432 20408 19484 20460
rect 20260 20451 20312 20460
rect 20260 20417 20269 20451
rect 20269 20417 20303 20451
rect 20303 20417 20312 20451
rect 20536 20451 20588 20460
rect 20260 20408 20312 20417
rect 20536 20417 20545 20451
rect 20545 20417 20579 20451
rect 20579 20417 20588 20451
rect 20536 20408 20588 20417
rect 1492 20340 1544 20392
rect 4896 20383 4948 20392
rect 4896 20349 4905 20383
rect 4905 20349 4939 20383
rect 4939 20349 4948 20383
rect 4896 20340 4948 20349
rect 5448 20340 5500 20392
rect 6920 20340 6972 20392
rect 7932 20340 7984 20392
rect 8668 20383 8720 20392
rect 8668 20349 8677 20383
rect 8677 20349 8711 20383
rect 8711 20349 8720 20383
rect 8668 20340 8720 20349
rect 8484 20272 8536 20324
rect 12992 20340 13044 20392
rect 15660 20383 15712 20392
rect 15660 20349 15669 20383
rect 15669 20349 15703 20383
rect 15703 20349 15712 20383
rect 15660 20340 15712 20349
rect 16304 20340 16356 20392
rect 21916 20451 21968 20460
rect 21916 20417 21925 20451
rect 21925 20417 21959 20451
rect 21959 20417 21968 20451
rect 21916 20408 21968 20417
rect 22100 20451 22152 20460
rect 22100 20417 22109 20451
rect 22109 20417 22143 20451
rect 22143 20417 22152 20451
rect 22100 20408 22152 20417
rect 22376 20408 22428 20460
rect 22928 20408 22980 20460
rect 23572 20544 23624 20596
rect 25412 20544 25464 20596
rect 26240 20544 26292 20596
rect 32956 20587 33008 20596
rect 26976 20476 27028 20528
rect 29552 20476 29604 20528
rect 32404 20476 32456 20528
rect 32956 20553 32965 20587
rect 32965 20553 32999 20587
rect 32999 20553 33008 20587
rect 32956 20544 33008 20553
rect 35716 20544 35768 20596
rect 38292 20544 38344 20596
rect 41328 20544 41380 20596
rect 42800 20544 42852 20596
rect 34336 20519 34388 20528
rect 23388 20451 23440 20460
rect 23388 20417 23397 20451
rect 23397 20417 23431 20451
rect 23431 20417 23440 20451
rect 23388 20408 23440 20417
rect 23664 20451 23716 20460
rect 23664 20417 23673 20451
rect 23673 20417 23707 20451
rect 23707 20417 23716 20451
rect 24400 20451 24452 20460
rect 23664 20408 23716 20417
rect 24400 20417 24409 20451
rect 24409 20417 24443 20451
rect 24443 20417 24452 20451
rect 24400 20408 24452 20417
rect 26608 20408 26660 20460
rect 27436 20451 27488 20460
rect 27436 20417 27445 20451
rect 27445 20417 27479 20451
rect 27479 20417 27488 20451
rect 27436 20408 27488 20417
rect 28264 20451 28316 20460
rect 28264 20417 28273 20451
rect 28273 20417 28307 20451
rect 28307 20417 28316 20451
rect 28264 20408 28316 20417
rect 25136 20340 25188 20392
rect 25320 20383 25372 20392
rect 25320 20349 25329 20383
rect 25329 20349 25363 20383
rect 25363 20349 25372 20383
rect 25320 20340 25372 20349
rect 28080 20340 28132 20392
rect 28448 20340 28500 20392
rect 32036 20408 32088 20460
rect 32496 20451 32548 20460
rect 32496 20417 32500 20451
rect 32500 20417 32534 20451
rect 32534 20417 32548 20451
rect 32496 20408 32548 20417
rect 34336 20485 34345 20519
rect 34345 20485 34379 20519
rect 34379 20485 34388 20519
rect 34336 20476 34388 20485
rect 3148 20247 3200 20256
rect 3148 20213 3157 20247
rect 3157 20213 3191 20247
rect 3191 20213 3200 20247
rect 3148 20204 3200 20213
rect 6368 20247 6420 20256
rect 6368 20213 6377 20247
rect 6377 20213 6411 20247
rect 6411 20213 6420 20247
rect 6368 20204 6420 20213
rect 14556 20204 14608 20256
rect 15384 20204 15436 20256
rect 18052 20204 18104 20256
rect 22100 20272 22152 20324
rect 29736 20272 29788 20324
rect 33692 20408 33744 20460
rect 35900 20476 35952 20528
rect 38108 20476 38160 20528
rect 41420 20476 41472 20528
rect 33784 20340 33836 20392
rect 34244 20340 34296 20392
rect 37648 20383 37700 20392
rect 37648 20349 37657 20383
rect 37657 20349 37691 20383
rect 37691 20349 37700 20383
rect 37648 20340 37700 20349
rect 21824 20204 21876 20256
rect 22928 20204 22980 20256
rect 23296 20204 23348 20256
rect 25228 20204 25280 20256
rect 25872 20204 25924 20256
rect 27896 20204 27948 20256
rect 30196 20204 30248 20256
rect 37372 20272 37424 20324
rect 37924 20408 37976 20460
rect 41788 20408 41840 20460
rect 42432 20451 42484 20460
rect 42432 20417 42441 20451
rect 42441 20417 42475 20451
rect 42475 20417 42484 20451
rect 42432 20408 42484 20417
rect 38844 20383 38896 20392
rect 38844 20349 38853 20383
rect 38853 20349 38887 20383
rect 38887 20349 38896 20383
rect 38844 20340 38896 20349
rect 40224 20340 40276 20392
rect 41696 20383 41748 20392
rect 41696 20349 41705 20383
rect 41705 20349 41739 20383
rect 41739 20349 41748 20383
rect 41696 20340 41748 20349
rect 32220 20204 32272 20256
rect 34152 20247 34204 20256
rect 34152 20213 34161 20247
rect 34161 20213 34195 20247
rect 34195 20213 34204 20247
rect 34152 20204 34204 20213
rect 37740 20247 37792 20256
rect 37740 20213 37749 20247
rect 37749 20213 37783 20247
rect 37783 20213 37792 20247
rect 37740 20204 37792 20213
rect 39488 20204 39540 20256
rect 41788 20204 41840 20256
rect 67640 20247 67692 20256
rect 67640 20213 67649 20247
rect 67649 20213 67683 20247
rect 67683 20213 67692 20247
rect 67640 20204 67692 20213
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 65654 20102 65706 20154
rect 65718 20102 65770 20154
rect 65782 20102 65834 20154
rect 65846 20102 65898 20154
rect 65910 20102 65962 20154
rect 7288 20000 7340 20052
rect 8116 20043 8168 20052
rect 8116 20009 8125 20043
rect 8125 20009 8159 20043
rect 8159 20009 8168 20043
rect 8116 20000 8168 20009
rect 9220 20000 9272 20052
rect 11060 20000 11112 20052
rect 18052 20000 18104 20052
rect 7840 19932 7892 19984
rect 8024 19907 8076 19916
rect 2228 19796 2280 19848
rect 4620 19796 4672 19848
rect 4896 19796 4948 19848
rect 7104 19839 7156 19848
rect 7104 19805 7113 19839
rect 7113 19805 7147 19839
rect 7147 19805 7156 19839
rect 7104 19796 7156 19805
rect 8024 19873 8033 19907
rect 8033 19873 8067 19907
rect 8067 19873 8076 19907
rect 8024 19864 8076 19873
rect 7472 19839 7524 19848
rect 1492 19660 1544 19712
rect 6920 19660 6972 19712
rect 7472 19805 7481 19839
rect 7481 19805 7515 19839
rect 7515 19805 7524 19839
rect 8484 19864 8536 19916
rect 9772 19864 9824 19916
rect 13268 19864 13320 19916
rect 7472 19796 7524 19805
rect 9107 19836 9159 19845
rect 7932 19771 7984 19780
rect 7932 19737 7941 19771
rect 7941 19737 7975 19771
rect 7975 19737 7984 19771
rect 7932 19728 7984 19737
rect 7840 19660 7892 19712
rect 9107 19802 9116 19836
rect 9116 19802 9150 19836
rect 9150 19802 9159 19836
rect 9107 19793 9159 19802
rect 9404 19796 9456 19848
rect 11612 19796 11664 19848
rect 12164 19796 12216 19848
rect 15660 19796 15712 19848
rect 16672 19864 16724 19916
rect 17040 19796 17092 19848
rect 22192 20000 22244 20052
rect 24400 20000 24452 20052
rect 24676 20043 24728 20052
rect 24676 20009 24685 20043
rect 24685 20009 24719 20043
rect 24719 20009 24728 20043
rect 24676 20000 24728 20009
rect 26148 20043 26200 20052
rect 26148 20009 26157 20043
rect 26157 20009 26191 20043
rect 26191 20009 26200 20043
rect 26148 20000 26200 20009
rect 26976 20000 27028 20052
rect 30564 20000 30616 20052
rect 32128 20043 32180 20052
rect 32128 20009 32137 20043
rect 32137 20009 32171 20043
rect 32171 20009 32180 20043
rect 32128 20000 32180 20009
rect 34244 20000 34296 20052
rect 37924 20043 37976 20052
rect 37924 20009 37933 20043
rect 37933 20009 37967 20043
rect 37967 20009 37976 20043
rect 37924 20000 37976 20009
rect 14464 19771 14516 19780
rect 14464 19737 14473 19771
rect 14473 19737 14507 19771
rect 14507 19737 14516 19771
rect 14464 19728 14516 19737
rect 15108 19728 15160 19780
rect 15292 19771 15344 19780
rect 15292 19737 15301 19771
rect 15301 19737 15335 19771
rect 15335 19737 15344 19771
rect 15292 19728 15344 19737
rect 15568 19728 15620 19780
rect 15752 19728 15804 19780
rect 16304 19728 16356 19780
rect 10140 19660 10192 19712
rect 14372 19660 14424 19712
rect 16488 19660 16540 19712
rect 17500 19660 17552 19712
rect 17684 19703 17736 19712
rect 17684 19669 17693 19703
rect 17693 19669 17727 19703
rect 17727 19669 17736 19703
rect 17684 19660 17736 19669
rect 19340 19932 19392 19984
rect 20628 19932 20680 19984
rect 27436 19932 27488 19984
rect 27712 19932 27764 19984
rect 28356 19932 28408 19984
rect 29644 19932 29696 19984
rect 29736 19932 29788 19984
rect 18328 19864 18380 19916
rect 19432 19864 19484 19916
rect 18880 19796 18932 19848
rect 20352 19796 20404 19848
rect 23388 19864 23440 19916
rect 25320 19864 25372 19916
rect 21824 19728 21876 19780
rect 23480 19796 23532 19848
rect 24584 19796 24636 19848
rect 25044 19796 25096 19848
rect 25688 19839 25740 19848
rect 25688 19805 25697 19839
rect 25697 19805 25731 19839
rect 25731 19805 25740 19839
rect 25688 19796 25740 19805
rect 24952 19771 25004 19780
rect 24952 19737 24961 19771
rect 24961 19737 24995 19771
rect 24995 19737 25004 19771
rect 24952 19728 25004 19737
rect 25964 19796 26016 19848
rect 26608 19839 26660 19848
rect 26608 19805 26617 19839
rect 26617 19805 26651 19839
rect 26651 19805 26660 19839
rect 26608 19796 26660 19805
rect 27712 19839 27764 19848
rect 27712 19805 27721 19839
rect 27721 19805 27755 19839
rect 27755 19805 27764 19839
rect 27712 19796 27764 19805
rect 27896 19839 27948 19848
rect 27896 19805 27905 19839
rect 27905 19805 27939 19839
rect 27939 19805 27948 19839
rect 27896 19796 27948 19805
rect 28172 19864 28224 19916
rect 30288 19864 30340 19916
rect 31024 19864 31076 19916
rect 31760 19907 31812 19916
rect 31760 19873 31769 19907
rect 31769 19873 31803 19907
rect 31803 19873 31812 19907
rect 31760 19864 31812 19873
rect 28080 19839 28132 19848
rect 28080 19805 28089 19839
rect 28089 19805 28123 19839
rect 28123 19805 28132 19839
rect 28080 19796 28132 19805
rect 29736 19796 29788 19848
rect 30196 19796 30248 19848
rect 30656 19839 30708 19848
rect 30656 19805 30665 19839
rect 30665 19805 30699 19839
rect 30699 19805 30708 19839
rect 30656 19796 30708 19805
rect 30932 19839 30984 19848
rect 30932 19805 30941 19839
rect 30941 19805 30975 19839
rect 30975 19805 30984 19839
rect 30932 19796 30984 19805
rect 37740 19932 37792 19984
rect 40224 20000 40276 20052
rect 41236 20000 41288 20052
rect 41880 20000 41932 20052
rect 32772 19839 32824 19848
rect 32772 19805 32781 19839
rect 32781 19805 32815 19839
rect 32815 19805 32824 19839
rect 32772 19796 32824 19805
rect 33508 19839 33560 19848
rect 33508 19805 33517 19839
rect 33517 19805 33551 19839
rect 33551 19805 33560 19839
rect 33508 19796 33560 19805
rect 34152 19864 34204 19916
rect 36084 19864 36136 19916
rect 38844 19864 38896 19916
rect 27620 19728 27672 19780
rect 28264 19728 28316 19780
rect 28816 19771 28868 19780
rect 28816 19737 28825 19771
rect 28825 19737 28859 19771
rect 28859 19737 28868 19771
rect 28816 19728 28868 19737
rect 33876 19839 33928 19848
rect 33876 19805 33885 19839
rect 33885 19805 33919 19839
rect 33919 19805 33928 19839
rect 33876 19796 33928 19805
rect 36728 19796 36780 19848
rect 34796 19728 34848 19780
rect 35348 19728 35400 19780
rect 37096 19728 37148 19780
rect 37556 19839 37608 19848
rect 37556 19805 37565 19839
rect 37565 19805 37599 19839
rect 37599 19805 37608 19839
rect 37556 19796 37608 19805
rect 38200 19796 38252 19848
rect 38292 19728 38344 19780
rect 40132 19839 40184 19848
rect 40132 19805 40141 19839
rect 40141 19805 40175 19839
rect 40175 19805 40184 19839
rect 40132 19796 40184 19805
rect 39488 19728 39540 19780
rect 20352 19660 20404 19712
rect 25872 19660 25924 19712
rect 28632 19660 28684 19712
rect 31116 19660 31168 19712
rect 32404 19660 32456 19712
rect 34704 19660 34756 19712
rect 34888 19703 34940 19712
rect 34888 19669 34897 19703
rect 34897 19669 34931 19703
rect 34931 19669 34940 19703
rect 34888 19660 34940 19669
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 50294 19558 50346 19610
rect 50358 19558 50410 19610
rect 50422 19558 50474 19610
rect 50486 19558 50538 19610
rect 50550 19558 50602 19610
rect 2228 19499 2280 19508
rect 2228 19465 2237 19499
rect 2237 19465 2271 19499
rect 2271 19465 2280 19499
rect 2228 19456 2280 19465
rect 8024 19456 8076 19508
rect 6368 19431 6420 19440
rect 6368 19397 6377 19431
rect 6377 19397 6411 19431
rect 6411 19397 6420 19431
rect 6368 19388 6420 19397
rect 7840 19388 7892 19440
rect 8208 19388 8260 19440
rect 9128 19456 9180 19508
rect 10048 19388 10100 19440
rect 14372 19388 14424 19440
rect 15200 19456 15252 19508
rect 16764 19456 16816 19508
rect 15292 19388 15344 19440
rect 18328 19456 18380 19508
rect 25320 19456 25372 19508
rect 29552 19456 29604 19508
rect 2872 19320 2924 19372
rect 6920 19320 6972 19372
rect 8116 19320 8168 19372
rect 10140 19320 10192 19372
rect 12164 19363 12216 19372
rect 12164 19329 12173 19363
rect 12173 19329 12207 19363
rect 12207 19329 12216 19363
rect 12164 19320 12216 19329
rect 14096 19320 14148 19372
rect 16948 19388 17000 19440
rect 15660 19363 15712 19372
rect 2780 19252 2832 19304
rect 3148 19252 3200 19304
rect 7288 19252 7340 19304
rect 9772 19295 9824 19304
rect 9772 19261 9781 19295
rect 9781 19261 9815 19295
rect 9815 19261 9824 19295
rect 9772 19252 9824 19261
rect 11980 19252 12032 19304
rect 13176 19252 13228 19304
rect 14464 19252 14516 19304
rect 15660 19329 15669 19363
rect 15669 19329 15703 19363
rect 15703 19329 15712 19363
rect 15660 19320 15712 19329
rect 16672 19320 16724 19372
rect 17960 19320 18012 19372
rect 18788 19320 18840 19372
rect 22376 19320 22428 19372
rect 23480 19363 23532 19372
rect 23480 19329 23489 19363
rect 23489 19329 23523 19363
rect 23523 19329 23532 19363
rect 23480 19320 23532 19329
rect 24584 19363 24636 19372
rect 24584 19329 24593 19363
rect 24593 19329 24627 19363
rect 24627 19329 24636 19363
rect 24584 19320 24636 19329
rect 25596 19388 25648 19440
rect 28632 19431 28684 19440
rect 28632 19397 28666 19431
rect 28666 19397 28684 19431
rect 28632 19388 28684 19397
rect 25688 19363 25740 19372
rect 16764 19252 16816 19304
rect 17132 19252 17184 19304
rect 18880 19295 18932 19304
rect 7288 19159 7340 19168
rect 7288 19125 7297 19159
rect 7297 19125 7331 19159
rect 7331 19125 7340 19159
rect 7288 19116 7340 19125
rect 7932 19116 7984 19168
rect 13912 19116 13964 19168
rect 15844 19116 15896 19168
rect 16672 19116 16724 19168
rect 17132 19116 17184 19168
rect 18880 19261 18889 19295
rect 18889 19261 18923 19295
rect 18923 19261 18932 19295
rect 18880 19252 18932 19261
rect 19064 19252 19116 19304
rect 20996 19252 21048 19304
rect 21732 19252 21784 19304
rect 20444 19184 20496 19236
rect 23572 19252 23624 19304
rect 25688 19329 25697 19363
rect 25697 19329 25731 19363
rect 25731 19329 25740 19363
rect 25688 19320 25740 19329
rect 25228 19252 25280 19304
rect 28448 19320 28500 19372
rect 30472 19320 30524 19372
rect 31852 19388 31904 19440
rect 33784 19388 33836 19440
rect 35992 19388 36044 19440
rect 36820 19388 36872 19440
rect 37096 19456 37148 19508
rect 31116 19363 31168 19372
rect 31116 19329 31125 19363
rect 31125 19329 31159 19363
rect 31159 19329 31168 19363
rect 32588 19363 32640 19372
rect 31116 19320 31168 19329
rect 32588 19329 32597 19363
rect 32597 19329 32631 19363
rect 32631 19329 32640 19363
rect 32588 19320 32640 19329
rect 33508 19320 33560 19372
rect 34612 19320 34664 19372
rect 34796 19320 34848 19372
rect 36268 19363 36320 19372
rect 36268 19329 36277 19363
rect 36277 19329 36311 19363
rect 36311 19329 36320 19363
rect 36268 19320 36320 19329
rect 37372 19320 37424 19372
rect 39488 19431 39540 19440
rect 39488 19397 39497 19431
rect 39497 19397 39531 19431
rect 39531 19397 39540 19431
rect 39488 19388 39540 19397
rect 40224 19388 40276 19440
rect 38292 19363 38344 19372
rect 38292 19329 38301 19363
rect 38301 19329 38335 19363
rect 38335 19329 38344 19363
rect 38292 19320 38344 19329
rect 31300 19252 31352 19304
rect 31760 19252 31812 19304
rect 33324 19252 33376 19304
rect 34704 19295 34756 19304
rect 34704 19261 34713 19295
rect 34713 19261 34747 19295
rect 34747 19261 34756 19295
rect 34704 19252 34756 19261
rect 20536 19116 20588 19168
rect 22560 19116 22612 19168
rect 26424 19116 26476 19168
rect 27344 19116 27396 19168
rect 27804 19116 27856 19168
rect 30104 19184 30156 19236
rect 38200 19184 38252 19236
rect 32036 19116 32088 19168
rect 32496 19116 32548 19168
rect 34704 19116 34756 19168
rect 36268 19116 36320 19168
rect 37004 19116 37056 19168
rect 41328 19116 41380 19168
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 65654 19014 65706 19066
rect 65718 19014 65770 19066
rect 65782 19014 65834 19066
rect 65846 19014 65898 19066
rect 65910 19014 65962 19066
rect 7288 18955 7340 18964
rect 7288 18921 7297 18955
rect 7297 18921 7331 18955
rect 7331 18921 7340 18955
rect 7288 18912 7340 18921
rect 13912 18912 13964 18964
rect 14096 18955 14148 18964
rect 14096 18921 14105 18955
rect 14105 18921 14139 18955
rect 14139 18921 14148 18955
rect 14096 18912 14148 18921
rect 15660 18912 15712 18964
rect 15384 18844 15436 18896
rect 15752 18844 15804 18896
rect 1492 18819 1544 18828
rect 1492 18785 1501 18819
rect 1501 18785 1535 18819
rect 1535 18785 1544 18819
rect 1492 18776 1544 18785
rect 8668 18776 8720 18828
rect 18880 18844 18932 18896
rect 25504 18912 25556 18964
rect 25688 18912 25740 18964
rect 24952 18844 25004 18896
rect 26056 18844 26108 18896
rect 1768 18751 1820 18760
rect 1768 18717 1777 18751
rect 1777 18717 1811 18751
rect 1811 18717 1820 18751
rect 1768 18708 1820 18717
rect 5816 18708 5868 18760
rect 19984 18776 20036 18828
rect 20444 18776 20496 18828
rect 13452 18708 13504 18760
rect 14188 18708 14240 18760
rect 14464 18751 14516 18760
rect 14464 18717 14473 18751
rect 14473 18717 14507 18751
rect 14507 18717 14516 18751
rect 14464 18708 14516 18717
rect 14556 18751 14608 18760
rect 14556 18717 14565 18751
rect 14565 18717 14599 18751
rect 14599 18717 14608 18751
rect 14556 18708 14608 18717
rect 10324 18640 10376 18692
rect 14924 18708 14976 18760
rect 15384 18751 15436 18760
rect 15384 18717 15393 18751
rect 15393 18717 15427 18751
rect 15427 18717 15436 18751
rect 15384 18708 15436 18717
rect 15660 18708 15712 18760
rect 17316 18708 17368 18760
rect 16120 18640 16172 18692
rect 17592 18640 17644 18692
rect 20168 18708 20220 18760
rect 20628 18708 20680 18760
rect 22376 18776 22428 18828
rect 21916 18751 21968 18760
rect 21916 18717 21925 18751
rect 21925 18717 21959 18751
rect 21959 18717 21968 18751
rect 21916 18708 21968 18717
rect 22560 18708 22612 18760
rect 25412 18776 25464 18828
rect 25504 18776 25556 18828
rect 25964 18776 26016 18828
rect 29644 18912 29696 18964
rect 30288 18955 30340 18964
rect 30288 18921 30297 18955
rect 30297 18921 30331 18955
rect 30331 18921 30340 18955
rect 30288 18912 30340 18921
rect 30380 18912 30432 18964
rect 37648 18912 37700 18964
rect 38292 18912 38344 18964
rect 40224 18955 40276 18964
rect 40224 18921 40233 18955
rect 40233 18921 40267 18955
rect 40267 18921 40276 18955
rect 40224 18912 40276 18921
rect 27344 18844 27396 18896
rect 30564 18844 30616 18896
rect 34796 18844 34848 18896
rect 30012 18819 30064 18828
rect 30012 18785 30021 18819
rect 30021 18785 30055 18819
rect 30055 18785 30064 18819
rect 30012 18776 30064 18785
rect 36268 18844 36320 18896
rect 41788 18887 41840 18896
rect 22100 18640 22152 18692
rect 25136 18640 25188 18692
rect 26424 18708 26476 18760
rect 28448 18708 28500 18760
rect 29828 18708 29880 18760
rect 4344 18572 4396 18624
rect 4988 18615 5040 18624
rect 4988 18581 4997 18615
rect 4997 18581 5031 18615
rect 5031 18581 5040 18615
rect 4988 18572 5040 18581
rect 11704 18615 11756 18624
rect 11704 18581 11713 18615
rect 11713 18581 11747 18615
rect 11747 18581 11756 18615
rect 11704 18572 11756 18581
rect 15384 18572 15436 18624
rect 15936 18572 15988 18624
rect 16764 18615 16816 18624
rect 16764 18581 16773 18615
rect 16773 18581 16807 18615
rect 16807 18581 16816 18615
rect 16764 18572 16816 18581
rect 17040 18572 17092 18624
rect 17224 18615 17276 18624
rect 17224 18581 17233 18615
rect 17233 18581 17267 18615
rect 17267 18581 17276 18615
rect 17224 18572 17276 18581
rect 20628 18572 20680 18624
rect 27620 18640 27672 18692
rect 32404 18708 32456 18760
rect 33048 18708 33100 18760
rect 33508 18708 33560 18760
rect 33784 18751 33836 18760
rect 33784 18717 33793 18751
rect 33793 18717 33827 18751
rect 33827 18717 33836 18751
rect 33784 18708 33836 18717
rect 34612 18708 34664 18760
rect 32680 18640 32732 18692
rect 33968 18683 34020 18692
rect 33968 18649 33977 18683
rect 33977 18649 34011 18683
rect 34011 18649 34020 18683
rect 33968 18640 34020 18649
rect 35072 18751 35124 18760
rect 35072 18717 35081 18751
rect 35081 18717 35115 18751
rect 35115 18717 35124 18751
rect 35072 18708 35124 18717
rect 36728 18708 36780 18760
rect 37004 18751 37056 18760
rect 37004 18717 37013 18751
rect 37013 18717 37047 18751
rect 37047 18717 37056 18751
rect 37004 18708 37056 18717
rect 41788 18853 41797 18887
rect 41797 18853 41831 18887
rect 41831 18853 41840 18887
rect 41788 18844 41840 18853
rect 41328 18819 41380 18828
rect 41328 18785 41337 18819
rect 41337 18785 41371 18819
rect 41371 18785 41380 18819
rect 41328 18776 41380 18785
rect 35992 18683 36044 18692
rect 35992 18649 36001 18683
rect 36001 18649 36035 18683
rect 36035 18649 36044 18683
rect 35992 18640 36044 18649
rect 36452 18640 36504 18692
rect 37556 18708 37608 18760
rect 38752 18708 38804 18760
rect 41420 18751 41472 18760
rect 41420 18717 41429 18751
rect 41429 18717 41463 18751
rect 41463 18717 41472 18751
rect 41420 18708 41472 18717
rect 68100 18751 68152 18760
rect 68100 18717 68109 18751
rect 68109 18717 68143 18751
rect 68143 18717 68152 18751
rect 68100 18708 68152 18717
rect 27712 18615 27764 18624
rect 27712 18581 27721 18615
rect 27721 18581 27755 18615
rect 27755 18581 27764 18615
rect 27712 18572 27764 18581
rect 28080 18572 28132 18624
rect 29552 18572 29604 18624
rect 31852 18572 31904 18624
rect 33324 18572 33376 18624
rect 34612 18572 34664 18624
rect 35072 18572 35124 18624
rect 35348 18615 35400 18624
rect 35348 18581 35357 18615
rect 35357 18581 35391 18615
rect 35391 18581 35400 18615
rect 35348 18572 35400 18581
rect 37648 18572 37700 18624
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 50294 18470 50346 18522
rect 50358 18470 50410 18522
rect 50422 18470 50474 18522
rect 50486 18470 50538 18522
rect 50550 18470 50602 18522
rect 2872 18411 2924 18420
rect 2872 18377 2881 18411
rect 2881 18377 2915 18411
rect 2915 18377 2924 18411
rect 2872 18368 2924 18377
rect 8484 18368 8536 18420
rect 8760 18368 8812 18420
rect 9864 18368 9916 18420
rect 10324 18411 10376 18420
rect 10324 18377 10333 18411
rect 10333 18377 10367 18411
rect 10367 18377 10376 18411
rect 10324 18368 10376 18377
rect 4988 18300 5040 18352
rect 2780 18232 2832 18284
rect 7288 18300 7340 18352
rect 4344 18207 4396 18216
rect 4344 18173 4353 18207
rect 4353 18173 4387 18207
rect 4387 18173 4396 18207
rect 4344 18164 4396 18173
rect 4620 18207 4672 18216
rect 4620 18173 4629 18207
rect 4629 18173 4663 18207
rect 4663 18173 4672 18207
rect 4620 18164 4672 18173
rect 2320 18071 2372 18080
rect 2320 18037 2329 18071
rect 2329 18037 2363 18071
rect 2363 18037 2372 18071
rect 2320 18028 2372 18037
rect 6460 18071 6512 18080
rect 6460 18037 6469 18071
rect 6469 18037 6503 18071
rect 6503 18037 6512 18071
rect 6460 18028 6512 18037
rect 6920 18275 6972 18284
rect 6920 18241 6929 18275
rect 6929 18241 6963 18275
rect 6963 18241 6972 18275
rect 6920 18232 6972 18241
rect 7104 18275 7156 18284
rect 7104 18241 7113 18275
rect 7113 18241 7147 18275
rect 7147 18241 7156 18275
rect 7104 18232 7156 18241
rect 7656 18164 7708 18216
rect 8668 18300 8720 18352
rect 8024 18275 8076 18284
rect 8024 18241 8058 18275
rect 8058 18241 8076 18275
rect 10232 18300 10284 18352
rect 14832 18368 14884 18420
rect 15200 18300 15252 18352
rect 8024 18232 8076 18241
rect 9864 18275 9916 18284
rect 9864 18241 9873 18275
rect 9873 18241 9907 18275
rect 9907 18241 9916 18275
rect 9864 18232 9916 18241
rect 8760 18164 8812 18216
rect 11060 18164 11112 18216
rect 14096 18164 14148 18216
rect 14648 18164 14700 18216
rect 15384 18232 15436 18284
rect 15660 18232 15712 18284
rect 16212 18300 16264 18352
rect 15476 18164 15528 18216
rect 16120 18275 16172 18284
rect 16120 18241 16129 18275
rect 16129 18241 16163 18275
rect 16163 18241 16172 18275
rect 16120 18232 16172 18241
rect 17132 18368 17184 18420
rect 17592 18411 17644 18420
rect 17592 18377 17601 18411
rect 17601 18377 17635 18411
rect 17635 18377 17644 18411
rect 17592 18368 17644 18377
rect 18696 18368 18748 18420
rect 19248 18368 19300 18420
rect 21916 18368 21968 18420
rect 30380 18368 30432 18420
rect 23572 18300 23624 18352
rect 16212 18164 16264 18216
rect 17408 18232 17460 18284
rect 18788 18275 18840 18284
rect 18788 18241 18797 18275
rect 18797 18241 18831 18275
rect 18831 18241 18840 18275
rect 18788 18232 18840 18241
rect 19064 18275 19116 18284
rect 19064 18241 19073 18275
rect 19073 18241 19107 18275
rect 19107 18241 19116 18275
rect 19064 18232 19116 18241
rect 19248 18232 19300 18284
rect 19984 18232 20036 18284
rect 21732 18232 21784 18284
rect 22008 18232 22060 18284
rect 25136 18300 25188 18352
rect 25412 18300 25464 18352
rect 27620 18343 27672 18352
rect 27620 18309 27629 18343
rect 27629 18309 27663 18343
rect 27663 18309 27672 18343
rect 27620 18300 27672 18309
rect 23940 18207 23992 18216
rect 23940 18173 23949 18207
rect 23949 18173 23983 18207
rect 23983 18173 23992 18207
rect 23940 18164 23992 18173
rect 24860 18275 24912 18284
rect 24860 18241 24869 18275
rect 24869 18241 24903 18275
rect 24903 18241 24912 18275
rect 24860 18232 24912 18241
rect 25044 18275 25096 18284
rect 25044 18241 25053 18275
rect 25053 18241 25087 18275
rect 25087 18241 25096 18275
rect 25044 18232 25096 18241
rect 25688 18232 25740 18284
rect 25228 18164 25280 18216
rect 26056 18232 26108 18284
rect 29000 18300 29052 18352
rect 29644 18300 29696 18352
rect 30196 18300 30248 18352
rect 33968 18368 34020 18420
rect 35900 18368 35952 18420
rect 40224 18368 40276 18420
rect 33600 18300 33652 18352
rect 35348 18300 35400 18352
rect 37556 18300 37608 18352
rect 27620 18164 27672 18216
rect 19616 18096 19668 18148
rect 22008 18139 22060 18148
rect 22008 18105 22017 18139
rect 22017 18105 22051 18139
rect 22051 18105 22060 18139
rect 22008 18096 22060 18105
rect 24584 18096 24636 18148
rect 36084 18232 36136 18284
rect 36728 18232 36780 18284
rect 37648 18275 37700 18284
rect 37648 18241 37657 18275
rect 37657 18241 37691 18275
rect 37691 18241 37700 18275
rect 37648 18232 37700 18241
rect 37832 18275 37884 18284
rect 37832 18241 37841 18275
rect 37841 18241 37875 18275
rect 37875 18241 37884 18275
rect 37832 18232 37884 18241
rect 38844 18232 38896 18284
rect 28448 18164 28500 18216
rect 29552 18164 29604 18216
rect 33968 18164 34020 18216
rect 8760 18028 8812 18080
rect 9128 18071 9180 18080
rect 9128 18037 9137 18071
rect 9137 18037 9171 18071
rect 9171 18037 9180 18071
rect 9128 18028 9180 18037
rect 14004 18028 14056 18080
rect 14924 18028 14976 18080
rect 15384 18028 15436 18080
rect 21272 18071 21324 18080
rect 21272 18037 21281 18071
rect 21281 18037 21315 18071
rect 21315 18037 21324 18071
rect 21272 18028 21324 18037
rect 23664 18028 23716 18080
rect 26056 18028 26108 18080
rect 27712 18071 27764 18080
rect 27712 18037 27721 18071
rect 27721 18037 27755 18071
rect 27755 18037 27764 18071
rect 27712 18028 27764 18037
rect 30748 18096 30800 18148
rect 29828 18028 29880 18080
rect 30196 18028 30248 18080
rect 33876 18096 33928 18148
rect 34704 18028 34756 18080
rect 36452 18028 36504 18080
rect 37740 18028 37792 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 65654 17926 65706 17978
rect 65718 17926 65770 17978
rect 65782 17926 65834 17978
rect 65846 17926 65898 17978
rect 65910 17926 65962 17978
rect 1860 17824 1912 17876
rect 4620 17824 4672 17876
rect 2872 17688 2924 17740
rect 2320 17620 2372 17672
rect 7656 17824 7708 17876
rect 8024 17867 8076 17876
rect 8024 17833 8033 17867
rect 8033 17833 8067 17867
rect 8067 17833 8076 17867
rect 8024 17824 8076 17833
rect 9864 17824 9916 17876
rect 14096 17867 14148 17876
rect 14096 17833 14105 17867
rect 14105 17833 14139 17867
rect 14139 17833 14148 17867
rect 14096 17824 14148 17833
rect 14832 17824 14884 17876
rect 18788 17824 18840 17876
rect 19616 17867 19668 17876
rect 19616 17833 19625 17867
rect 19625 17833 19659 17867
rect 19659 17833 19668 17867
rect 19616 17824 19668 17833
rect 21456 17867 21508 17876
rect 21456 17833 21465 17867
rect 21465 17833 21499 17867
rect 21499 17833 21508 17867
rect 21456 17824 21508 17833
rect 22560 17824 22612 17876
rect 23112 17824 23164 17876
rect 23572 17824 23624 17876
rect 24860 17824 24912 17876
rect 27620 17824 27672 17876
rect 32680 17867 32732 17876
rect 32680 17833 32689 17867
rect 32689 17833 32723 17867
rect 32723 17833 32732 17867
rect 32680 17824 32732 17833
rect 9956 17756 10008 17808
rect 15660 17756 15712 17808
rect 16672 17756 16724 17808
rect 20904 17756 20956 17808
rect 21916 17756 21968 17808
rect 23940 17756 23992 17808
rect 25688 17756 25740 17808
rect 8760 17688 8812 17740
rect 12164 17731 12216 17740
rect 12164 17697 12173 17731
rect 12173 17697 12207 17731
rect 12207 17697 12216 17731
rect 12164 17688 12216 17697
rect 16212 17731 16264 17740
rect 16212 17697 16221 17731
rect 16221 17697 16255 17731
rect 16255 17697 16264 17731
rect 16212 17688 16264 17697
rect 19064 17688 19116 17740
rect 25228 17688 25280 17740
rect 1860 17552 1912 17604
rect 5264 17527 5316 17536
rect 5264 17493 5273 17527
rect 5273 17493 5307 17527
rect 5307 17493 5316 17527
rect 5264 17484 5316 17493
rect 6460 17552 6512 17604
rect 7748 17663 7800 17672
rect 7748 17629 7757 17663
rect 7757 17629 7791 17663
rect 7791 17629 7800 17663
rect 7748 17620 7800 17629
rect 9220 17620 9272 17672
rect 9128 17595 9180 17604
rect 9128 17561 9137 17595
rect 9137 17561 9171 17595
rect 9171 17561 9180 17595
rect 11704 17620 11756 17672
rect 15384 17620 15436 17672
rect 15476 17663 15528 17672
rect 15476 17629 15485 17663
rect 15485 17629 15519 17663
rect 15519 17629 15528 17663
rect 15476 17620 15528 17629
rect 16304 17620 16356 17672
rect 16948 17620 17000 17672
rect 17776 17620 17828 17672
rect 21272 17620 21324 17672
rect 9128 17552 9180 17561
rect 11612 17552 11664 17604
rect 7012 17484 7064 17536
rect 11244 17484 11296 17536
rect 11796 17484 11848 17536
rect 12256 17552 12308 17604
rect 14924 17552 14976 17604
rect 16580 17484 16632 17536
rect 17224 17527 17276 17536
rect 17224 17493 17233 17527
rect 17233 17493 17267 17527
rect 17267 17493 17276 17527
rect 17224 17484 17276 17493
rect 19156 17552 19208 17604
rect 21732 17663 21784 17672
rect 21732 17629 21741 17663
rect 21741 17629 21775 17663
rect 21775 17629 21784 17663
rect 21732 17620 21784 17629
rect 22376 17552 22428 17604
rect 21732 17484 21784 17536
rect 24860 17620 24912 17672
rect 25320 17620 25372 17672
rect 25504 17663 25556 17672
rect 26332 17688 26384 17740
rect 25504 17629 25519 17663
rect 25519 17629 25553 17663
rect 25553 17629 25556 17663
rect 25504 17620 25556 17629
rect 32220 17688 32272 17740
rect 24584 17595 24636 17604
rect 24584 17561 24593 17595
rect 24593 17561 24627 17595
rect 24627 17561 24636 17595
rect 24584 17552 24636 17561
rect 28448 17620 28500 17672
rect 31116 17620 31168 17672
rect 31484 17663 31536 17672
rect 31484 17629 31493 17663
rect 31493 17629 31527 17663
rect 31527 17629 31536 17663
rect 31484 17620 31536 17629
rect 33232 17756 33284 17808
rect 33416 17620 33468 17672
rect 26056 17552 26108 17604
rect 40040 17688 40092 17740
rect 37740 17620 37792 17672
rect 68100 17663 68152 17672
rect 68100 17629 68109 17663
rect 68109 17629 68143 17663
rect 68143 17629 68152 17663
rect 68100 17620 68152 17629
rect 26240 17484 26292 17536
rect 32220 17527 32272 17536
rect 32220 17493 32229 17527
rect 32229 17493 32263 17527
rect 32263 17493 32272 17527
rect 32220 17484 32272 17493
rect 32864 17484 32916 17536
rect 37648 17595 37700 17604
rect 37648 17561 37657 17595
rect 37657 17561 37691 17595
rect 37691 17561 37700 17595
rect 37648 17552 37700 17561
rect 37832 17595 37884 17604
rect 37832 17561 37841 17595
rect 37841 17561 37875 17595
rect 37875 17561 37884 17595
rect 37832 17552 37884 17561
rect 35440 17484 35492 17536
rect 35624 17484 35676 17536
rect 35716 17484 35768 17536
rect 36268 17527 36320 17536
rect 36268 17493 36277 17527
rect 36277 17493 36311 17527
rect 36311 17493 36320 17527
rect 36268 17484 36320 17493
rect 37188 17527 37240 17536
rect 37188 17493 37197 17527
rect 37197 17493 37231 17527
rect 37231 17493 37240 17527
rect 37188 17484 37240 17493
rect 37464 17484 37516 17536
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 50294 17382 50346 17434
rect 50358 17382 50410 17434
rect 50422 17382 50474 17434
rect 50486 17382 50538 17434
rect 50550 17382 50602 17434
rect 1400 17323 1452 17332
rect 1400 17289 1409 17323
rect 1409 17289 1443 17323
rect 1443 17289 1452 17323
rect 1400 17280 1452 17289
rect 2872 17280 2924 17332
rect 6920 17280 6972 17332
rect 12256 17323 12308 17332
rect 2320 17144 2372 17196
rect 2596 17144 2648 17196
rect 3240 17212 3292 17264
rect 2964 17187 3016 17196
rect 2964 17153 2973 17187
rect 2973 17153 3007 17187
rect 3007 17153 3016 17187
rect 2964 17144 3016 17153
rect 3148 17187 3200 17196
rect 3148 17153 3157 17187
rect 3157 17153 3191 17187
rect 3191 17153 3200 17187
rect 4620 17212 4672 17264
rect 5264 17212 5316 17264
rect 3148 17144 3200 17153
rect 2412 17076 2464 17128
rect 4712 17144 4764 17196
rect 1952 16983 2004 16992
rect 1952 16949 1961 16983
rect 1961 16949 1995 16983
rect 1995 16949 2004 16983
rect 1952 16940 2004 16949
rect 7472 17076 7524 17128
rect 3148 16940 3200 16992
rect 7104 17008 7156 17060
rect 8208 17144 8260 17196
rect 8760 17212 8812 17264
rect 8484 17187 8536 17196
rect 8484 17153 8493 17187
rect 8493 17153 8527 17187
rect 8527 17153 8536 17187
rect 8484 17144 8536 17153
rect 9588 17144 9640 17196
rect 12256 17289 12265 17323
rect 12265 17289 12299 17323
rect 12299 17289 12308 17323
rect 12256 17280 12308 17289
rect 9956 17212 10008 17264
rect 10692 17255 10744 17264
rect 10692 17221 10701 17255
rect 10701 17221 10735 17255
rect 10735 17221 10744 17255
rect 10692 17212 10744 17221
rect 11060 17212 11112 17264
rect 11520 17144 11572 17196
rect 11796 17187 11848 17196
rect 11428 17076 11480 17128
rect 11796 17153 11805 17187
rect 11805 17153 11839 17187
rect 11839 17153 11848 17187
rect 11796 17144 11848 17153
rect 11980 17187 12032 17196
rect 11980 17153 11989 17187
rect 11989 17153 12023 17187
rect 12023 17153 12032 17187
rect 16120 17280 16172 17332
rect 16212 17280 16264 17332
rect 18696 17280 18748 17332
rect 11980 17144 12032 17153
rect 15660 17187 15712 17196
rect 15660 17153 15669 17187
rect 15669 17153 15703 17187
rect 15703 17153 15712 17187
rect 15660 17144 15712 17153
rect 16396 17212 16448 17264
rect 16212 17144 16264 17196
rect 19984 17212 20036 17264
rect 20904 17212 20956 17264
rect 23848 17280 23900 17332
rect 25228 17280 25280 17332
rect 25320 17280 25372 17332
rect 25504 17280 25556 17332
rect 12072 17076 12124 17128
rect 19248 17187 19300 17196
rect 19248 17153 19257 17187
rect 19257 17153 19291 17187
rect 19291 17153 19300 17187
rect 19248 17144 19300 17153
rect 19432 17187 19484 17196
rect 19432 17153 19441 17187
rect 19441 17153 19475 17187
rect 19475 17153 19484 17187
rect 19432 17144 19484 17153
rect 19064 17076 19116 17128
rect 19708 17144 19760 17196
rect 20260 17144 20312 17196
rect 21272 17187 21324 17196
rect 21272 17153 21281 17187
rect 21281 17153 21315 17187
rect 21315 17153 21324 17187
rect 21272 17144 21324 17153
rect 22836 17144 22888 17196
rect 23940 17187 23992 17196
rect 23940 17153 23949 17187
rect 23949 17153 23983 17187
rect 23983 17153 23992 17187
rect 23940 17144 23992 17153
rect 28356 17187 28408 17196
rect 4988 16983 5040 16992
rect 4988 16949 4997 16983
rect 4997 16949 5031 16983
rect 5031 16949 5040 16983
rect 8760 16983 8812 16992
rect 4988 16940 5040 16949
rect 8760 16949 8769 16983
rect 8769 16949 8803 16983
rect 8803 16949 8812 16983
rect 8760 16940 8812 16949
rect 13636 17008 13688 17060
rect 18788 17051 18840 17060
rect 18788 17017 18797 17051
rect 18797 17017 18831 17051
rect 18831 17017 18840 17051
rect 22192 17076 22244 17128
rect 28356 17153 28365 17187
rect 28365 17153 28399 17187
rect 28399 17153 28408 17187
rect 28356 17144 28408 17153
rect 28540 17280 28592 17332
rect 28632 17280 28684 17332
rect 29000 17323 29052 17332
rect 29000 17289 29009 17323
rect 29009 17289 29043 17323
rect 29043 17289 29052 17323
rect 29000 17280 29052 17289
rect 28908 17212 28960 17264
rect 37740 17280 37792 17332
rect 37832 17280 37884 17332
rect 35716 17212 35768 17264
rect 26516 17076 26568 17128
rect 29920 17144 29972 17196
rect 33232 17187 33284 17196
rect 33232 17153 33241 17187
rect 33241 17153 33275 17187
rect 33275 17153 33284 17187
rect 33232 17144 33284 17153
rect 35348 17144 35400 17196
rect 36084 17187 36136 17196
rect 36084 17153 36093 17187
rect 36093 17153 36127 17187
rect 36127 17153 36136 17187
rect 36084 17144 36136 17153
rect 37280 17187 37332 17196
rect 37280 17153 37289 17187
rect 37289 17153 37323 17187
rect 37323 17153 37332 17187
rect 37280 17144 37332 17153
rect 37464 17187 37516 17196
rect 37464 17153 37473 17187
rect 37473 17153 37507 17187
rect 37507 17153 37516 17187
rect 37464 17144 37516 17153
rect 37556 17187 37608 17196
rect 37556 17153 37565 17187
rect 37565 17153 37599 17187
rect 37599 17153 37608 17187
rect 37556 17144 37608 17153
rect 18788 17008 18840 17017
rect 20904 17008 20956 17060
rect 11428 16940 11480 16992
rect 17960 16940 18012 16992
rect 20260 16940 20312 16992
rect 20444 16983 20496 16992
rect 20444 16949 20453 16983
rect 20453 16949 20487 16983
rect 20487 16949 20496 16983
rect 20444 16940 20496 16949
rect 22100 16940 22152 16992
rect 25044 16940 25096 16992
rect 26332 16983 26384 16992
rect 26332 16949 26341 16983
rect 26341 16949 26375 16983
rect 26375 16949 26384 16983
rect 26332 16940 26384 16949
rect 27988 16940 28040 16992
rect 28448 16940 28500 16992
rect 31484 17076 31536 17128
rect 31208 16940 31260 16992
rect 34520 16940 34572 16992
rect 36084 16940 36136 16992
rect 38844 17144 38896 17196
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 65654 16838 65706 16890
rect 65718 16838 65770 16890
rect 65782 16838 65834 16890
rect 65846 16838 65898 16890
rect 65910 16838 65962 16890
rect 1952 16736 2004 16788
rect 2872 16736 2924 16788
rect 2964 16736 3016 16788
rect 8208 16736 8260 16788
rect 15660 16779 15712 16788
rect 2596 16668 2648 16720
rect 5080 16668 5132 16720
rect 7748 16668 7800 16720
rect 15660 16745 15669 16779
rect 15669 16745 15703 16779
rect 15703 16745 15712 16779
rect 15660 16736 15712 16745
rect 19248 16736 19300 16788
rect 16212 16668 16264 16720
rect 16856 16668 16908 16720
rect 2964 16600 3016 16652
rect 3240 16600 3292 16652
rect 2320 16532 2372 16584
rect 4988 16532 5040 16584
rect 5448 16532 5500 16584
rect 8668 16600 8720 16652
rect 10692 16600 10744 16652
rect 12164 16643 12216 16652
rect 7472 16575 7524 16584
rect 7472 16541 7481 16575
rect 7481 16541 7515 16575
rect 7515 16541 7524 16575
rect 7472 16532 7524 16541
rect 7656 16575 7708 16584
rect 7656 16541 7665 16575
rect 7665 16541 7699 16575
rect 7699 16541 7708 16575
rect 7656 16532 7708 16541
rect 8760 16532 8812 16584
rect 12164 16609 12173 16643
rect 12173 16609 12207 16643
rect 12207 16609 12216 16643
rect 12164 16600 12216 16609
rect 14924 16600 14976 16652
rect 16304 16600 16356 16652
rect 11244 16575 11296 16584
rect 11244 16541 11253 16575
rect 11253 16541 11287 16575
rect 11287 16541 11296 16575
rect 11244 16532 11296 16541
rect 4712 16507 4764 16516
rect 4712 16473 4721 16507
rect 4721 16473 4755 16507
rect 4755 16473 4764 16507
rect 4712 16464 4764 16473
rect 10968 16464 11020 16516
rect 11428 16575 11480 16584
rect 11428 16541 11437 16575
rect 11437 16541 11471 16575
rect 11471 16541 11480 16575
rect 11428 16532 11480 16541
rect 5356 16396 5408 16448
rect 7012 16439 7064 16448
rect 7012 16405 7021 16439
rect 7021 16405 7055 16439
rect 7055 16405 7064 16439
rect 7012 16396 7064 16405
rect 9496 16396 9548 16448
rect 14096 16532 14148 16584
rect 13084 16464 13136 16516
rect 17960 16532 18012 16584
rect 23480 16736 23532 16788
rect 25320 16736 25372 16788
rect 26516 16779 26568 16788
rect 26516 16745 26525 16779
rect 26525 16745 26559 16779
rect 26559 16745 26568 16779
rect 26516 16736 26568 16745
rect 28540 16736 28592 16788
rect 29920 16779 29972 16788
rect 29920 16745 29929 16779
rect 29929 16745 29963 16779
rect 29963 16745 29972 16779
rect 29920 16736 29972 16745
rect 22192 16711 22244 16720
rect 22192 16677 22201 16711
rect 22201 16677 22235 16711
rect 22235 16677 22244 16711
rect 22192 16668 22244 16677
rect 23572 16668 23624 16720
rect 31392 16736 31444 16788
rect 31944 16736 31996 16788
rect 32864 16779 32916 16788
rect 32864 16745 32873 16779
rect 32873 16745 32907 16779
rect 32907 16745 32916 16779
rect 32864 16736 32916 16745
rect 30196 16668 30248 16720
rect 34704 16736 34756 16788
rect 35348 16779 35400 16788
rect 35348 16745 35357 16779
rect 35357 16745 35391 16779
rect 35391 16745 35400 16779
rect 35348 16736 35400 16745
rect 35716 16736 35768 16788
rect 35992 16736 36044 16788
rect 19984 16600 20036 16652
rect 23756 16600 23808 16652
rect 15936 16464 15988 16516
rect 18972 16464 19024 16516
rect 19156 16464 19208 16516
rect 11796 16396 11848 16448
rect 17132 16396 17184 16448
rect 19248 16439 19300 16448
rect 19248 16405 19257 16439
rect 19257 16405 19291 16439
rect 19291 16405 19300 16439
rect 19248 16396 19300 16405
rect 20260 16532 20312 16584
rect 22008 16532 22060 16584
rect 22100 16532 22152 16584
rect 24860 16575 24912 16584
rect 24860 16541 24869 16575
rect 24869 16541 24903 16575
rect 24903 16541 24912 16575
rect 24860 16532 24912 16541
rect 25044 16575 25096 16584
rect 25044 16541 25053 16575
rect 25053 16541 25087 16575
rect 25087 16541 25096 16575
rect 25044 16532 25096 16541
rect 25320 16532 25372 16584
rect 27988 16600 28040 16652
rect 28908 16600 28960 16652
rect 28356 16532 28408 16584
rect 28816 16532 28868 16584
rect 30104 16532 30156 16584
rect 30293 16569 30345 16584
rect 31576 16600 31628 16652
rect 37832 16668 37884 16720
rect 30293 16535 30310 16569
rect 30310 16535 30344 16569
rect 30344 16535 30345 16569
rect 30293 16532 30345 16535
rect 19984 16464 20036 16516
rect 22376 16507 22428 16516
rect 22376 16473 22385 16507
rect 22385 16473 22419 16507
rect 22419 16473 22428 16507
rect 22376 16464 22428 16473
rect 25228 16464 25280 16516
rect 28264 16507 28316 16516
rect 28264 16473 28273 16507
rect 28273 16473 28307 16507
rect 28307 16473 28316 16507
rect 28264 16464 28316 16473
rect 29920 16464 29972 16516
rect 19616 16396 19668 16448
rect 21732 16439 21784 16448
rect 21732 16405 21741 16439
rect 21741 16405 21775 16439
rect 21775 16405 21784 16439
rect 21732 16396 21784 16405
rect 25872 16439 25924 16448
rect 25872 16405 25881 16439
rect 25881 16405 25915 16439
rect 25915 16405 25924 16439
rect 25872 16396 25924 16405
rect 31208 16575 31260 16584
rect 31208 16541 31217 16575
rect 31217 16541 31251 16575
rect 31251 16541 31260 16575
rect 31208 16532 31260 16541
rect 33600 16532 33652 16584
rect 34704 16575 34756 16584
rect 34704 16541 34713 16575
rect 34713 16541 34747 16575
rect 34747 16541 34756 16575
rect 34704 16532 34756 16541
rect 35624 16600 35676 16652
rect 30840 16464 30892 16516
rect 33324 16464 33376 16516
rect 33784 16507 33836 16516
rect 33784 16473 33793 16507
rect 33793 16473 33827 16507
rect 33827 16473 33836 16507
rect 33784 16464 33836 16473
rect 34520 16464 34572 16516
rect 32404 16396 32456 16448
rect 33232 16396 33284 16448
rect 35532 16532 35584 16584
rect 37280 16575 37332 16584
rect 37280 16541 37289 16575
rect 37289 16541 37323 16575
rect 37323 16541 37332 16575
rect 37280 16532 37332 16541
rect 38292 16736 38344 16788
rect 37188 16464 37240 16516
rect 37372 16396 37424 16448
rect 37556 16396 37608 16448
rect 37924 16439 37976 16448
rect 37924 16405 37933 16439
rect 37933 16405 37967 16439
rect 37967 16405 37976 16439
rect 37924 16396 37976 16405
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 50294 16294 50346 16346
rect 50358 16294 50410 16346
rect 50422 16294 50474 16346
rect 50486 16294 50538 16346
rect 50550 16294 50602 16346
rect 3148 16192 3200 16244
rect 7656 16192 7708 16244
rect 11244 16192 11296 16244
rect 18236 16235 18288 16244
rect 18236 16201 18245 16235
rect 18245 16201 18279 16235
rect 18279 16201 18288 16235
rect 18236 16192 18288 16201
rect 19432 16192 19484 16244
rect 22376 16192 22428 16244
rect 3240 16099 3292 16108
rect 3240 16065 3249 16099
rect 3249 16065 3283 16099
rect 3283 16065 3292 16099
rect 3240 16056 3292 16065
rect 3424 16056 3476 16108
rect 9220 16124 9272 16176
rect 3148 15920 3200 15972
rect 6920 16056 6972 16108
rect 9312 16056 9364 16108
rect 9496 16099 9548 16108
rect 9496 16065 9505 16099
rect 9505 16065 9539 16099
rect 9539 16065 9548 16099
rect 9496 16056 9548 16065
rect 7196 15988 7248 16040
rect 7012 15920 7064 15972
rect 11796 16124 11848 16176
rect 13636 16124 13688 16176
rect 17776 16167 17828 16176
rect 17776 16133 17785 16167
rect 17785 16133 17819 16167
rect 17819 16133 17828 16167
rect 17776 16124 17828 16133
rect 18972 16167 19024 16176
rect 18972 16133 18981 16167
rect 18981 16133 19015 16167
rect 19015 16133 19024 16167
rect 18972 16124 19024 16133
rect 11520 16099 11572 16108
rect 11520 16065 11529 16099
rect 11529 16065 11563 16099
rect 11563 16065 11572 16099
rect 11520 16056 11572 16065
rect 11704 16056 11756 16108
rect 14648 16099 14700 16108
rect 14648 16065 14658 16099
rect 14658 16065 14692 16099
rect 14692 16065 14700 16099
rect 14648 16056 14700 16065
rect 14832 16099 14884 16108
rect 14832 16065 14841 16099
rect 14841 16065 14875 16099
rect 14875 16065 14884 16099
rect 14832 16056 14884 16065
rect 15016 16099 15068 16108
rect 15016 16065 15030 16099
rect 15030 16065 15064 16099
rect 15064 16065 15068 16099
rect 17960 16099 18012 16108
rect 15016 16056 15068 16065
rect 17960 16065 17969 16099
rect 17969 16065 18003 16099
rect 18003 16065 18012 16099
rect 17960 16056 18012 16065
rect 18052 16099 18104 16108
rect 18052 16065 18061 16099
rect 18061 16065 18095 16099
rect 18095 16065 18104 16099
rect 18052 16056 18104 16065
rect 12072 15988 12124 16040
rect 21732 16124 21784 16176
rect 24124 16192 24176 16244
rect 23204 16124 23256 16176
rect 36452 16192 36504 16244
rect 40040 16235 40092 16244
rect 40040 16201 40049 16235
rect 40049 16201 40083 16235
rect 40083 16201 40092 16235
rect 40040 16192 40092 16201
rect 22376 16056 22428 16108
rect 22560 16099 22612 16108
rect 22560 16065 22569 16099
rect 22569 16065 22603 16099
rect 22603 16065 22612 16099
rect 22560 16056 22612 16065
rect 23756 16099 23808 16108
rect 11980 15920 12032 15972
rect 3884 15852 3936 15904
rect 4712 15852 4764 15904
rect 6552 15895 6604 15904
rect 6552 15861 6561 15895
rect 6561 15861 6595 15895
rect 6595 15861 6604 15895
rect 6552 15852 6604 15861
rect 15568 15852 15620 15904
rect 17040 15852 17092 15904
rect 22100 15988 22152 16040
rect 23756 16065 23765 16099
rect 23765 16065 23799 16099
rect 23799 16065 23808 16099
rect 23756 16056 23808 16065
rect 24584 16056 24636 16108
rect 25688 16099 25740 16108
rect 25688 16065 25697 16099
rect 25697 16065 25731 16099
rect 25731 16065 25740 16099
rect 25688 16056 25740 16065
rect 27712 16056 27764 16108
rect 27988 16056 28040 16108
rect 28540 16099 28592 16108
rect 28540 16065 28549 16099
rect 28549 16065 28583 16099
rect 28583 16065 28592 16099
rect 28540 16056 28592 16065
rect 28724 16056 28776 16108
rect 28816 16099 28868 16108
rect 28816 16065 28825 16099
rect 28825 16065 28859 16099
rect 28859 16065 28868 16099
rect 28816 16056 28868 16065
rect 30472 15988 30524 16040
rect 35072 16124 35124 16176
rect 37924 16124 37976 16176
rect 32864 16056 32916 16108
rect 33508 16099 33560 16108
rect 33508 16065 33517 16099
rect 33517 16065 33551 16099
rect 33551 16065 33560 16099
rect 33508 16056 33560 16065
rect 34888 16056 34940 16108
rect 35532 16099 35584 16108
rect 35532 16065 35541 16099
rect 35541 16065 35575 16099
rect 35575 16065 35584 16099
rect 35532 16056 35584 16065
rect 33692 15988 33744 16040
rect 34704 15988 34756 16040
rect 35072 16031 35124 16040
rect 35072 15997 35081 16031
rect 35081 15997 35115 16031
rect 35115 15997 35124 16031
rect 35072 15988 35124 15997
rect 35348 15988 35400 16040
rect 35440 15988 35492 16040
rect 35808 16099 35860 16108
rect 35808 16065 35817 16099
rect 35817 16065 35851 16099
rect 35851 16065 35860 16099
rect 35808 16056 35860 16065
rect 35992 16056 36044 16108
rect 37648 16099 37700 16108
rect 37648 16065 37657 16099
rect 37657 16065 37691 16099
rect 37691 16065 37700 16099
rect 37648 16056 37700 16065
rect 38752 16056 38804 16108
rect 37924 15988 37976 16040
rect 18144 15920 18196 15972
rect 24676 15920 24728 15972
rect 22744 15895 22796 15904
rect 22744 15861 22753 15895
rect 22753 15861 22787 15895
rect 22787 15861 22796 15895
rect 22744 15852 22796 15861
rect 23480 15852 23532 15904
rect 29000 15920 29052 15972
rect 27160 15895 27212 15904
rect 27160 15861 27169 15895
rect 27169 15861 27203 15895
rect 27203 15861 27212 15895
rect 27160 15852 27212 15861
rect 28356 15852 28408 15904
rect 30012 15852 30064 15904
rect 30104 15852 30156 15904
rect 33600 15852 33652 15904
rect 36176 15895 36228 15904
rect 36176 15861 36185 15895
rect 36185 15861 36219 15895
rect 36219 15861 36228 15895
rect 36176 15852 36228 15861
rect 37464 15852 37516 15904
rect 67640 15895 67692 15904
rect 67640 15861 67649 15895
rect 67649 15861 67683 15895
rect 67683 15861 67692 15895
rect 67640 15852 67692 15861
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 65654 15750 65706 15802
rect 65718 15750 65770 15802
rect 65782 15750 65834 15802
rect 65846 15750 65898 15802
rect 65910 15750 65962 15802
rect 1768 15648 1820 15700
rect 2780 15691 2832 15700
rect 2780 15657 2789 15691
rect 2789 15657 2823 15691
rect 2823 15657 2832 15691
rect 2780 15648 2832 15657
rect 6460 15648 6512 15700
rect 9312 15648 9364 15700
rect 11888 15648 11940 15700
rect 11980 15691 12032 15700
rect 11980 15657 11989 15691
rect 11989 15657 12023 15691
rect 12023 15657 12032 15691
rect 11980 15648 12032 15657
rect 14924 15648 14976 15700
rect 18328 15648 18380 15700
rect 19984 15648 20036 15700
rect 27804 15648 27856 15700
rect 28724 15648 28776 15700
rect 32864 15691 32916 15700
rect 32864 15657 32873 15691
rect 32873 15657 32907 15691
rect 32907 15657 32916 15691
rect 32864 15648 32916 15657
rect 36912 15691 36964 15700
rect 36912 15657 36921 15691
rect 36921 15657 36955 15691
rect 36955 15657 36964 15691
rect 36912 15648 36964 15657
rect 38108 15648 38160 15700
rect 1400 15444 1452 15496
rect 2136 15487 2188 15496
rect 2136 15453 2145 15487
rect 2145 15453 2179 15487
rect 2179 15453 2188 15487
rect 2136 15444 2188 15453
rect 2964 15512 3016 15564
rect 3424 15512 3476 15564
rect 3608 15444 3660 15496
rect 3884 15444 3936 15496
rect 7196 15555 7248 15564
rect 7196 15521 7205 15555
rect 7205 15521 7239 15555
rect 7239 15521 7248 15555
rect 7196 15512 7248 15521
rect 7932 15512 7984 15564
rect 6460 15487 6512 15496
rect 6460 15453 6469 15487
rect 6469 15453 6503 15487
rect 6503 15453 6512 15487
rect 6460 15444 6512 15453
rect 6552 15487 6604 15496
rect 6552 15453 6561 15487
rect 6561 15453 6595 15487
rect 6595 15453 6604 15487
rect 6552 15444 6604 15453
rect 7656 15444 7708 15496
rect 7012 15419 7064 15428
rect 7012 15385 7021 15419
rect 7021 15385 7055 15419
rect 7055 15385 7064 15419
rect 7012 15376 7064 15385
rect 4896 15308 4948 15360
rect 5264 15308 5316 15360
rect 6644 15308 6696 15360
rect 8392 15444 8444 15496
rect 8484 15444 8536 15496
rect 9588 15512 9640 15564
rect 9772 15444 9824 15496
rect 10324 15487 10376 15496
rect 10324 15453 10333 15487
rect 10333 15453 10367 15487
rect 10367 15453 10376 15487
rect 10324 15444 10376 15453
rect 10692 15444 10744 15496
rect 11796 15512 11848 15564
rect 11336 15487 11388 15496
rect 11336 15453 11345 15487
rect 11345 15453 11379 15487
rect 11379 15453 11388 15487
rect 11336 15444 11388 15453
rect 11612 15444 11664 15496
rect 8116 15419 8168 15428
rect 8116 15385 8125 15419
rect 8125 15385 8159 15419
rect 8159 15385 8168 15419
rect 8116 15376 8168 15385
rect 8852 15376 8904 15428
rect 9588 15376 9640 15428
rect 11704 15376 11756 15428
rect 12624 15444 12676 15496
rect 12992 15580 13044 15632
rect 13084 15487 13136 15496
rect 13084 15453 13091 15487
rect 13091 15453 13136 15487
rect 13084 15444 13136 15453
rect 15016 15512 15068 15564
rect 14280 15444 14332 15496
rect 14832 15444 14884 15496
rect 14924 15487 14976 15496
rect 14924 15453 14933 15487
rect 14933 15453 14967 15487
rect 14967 15453 14976 15487
rect 17868 15580 17920 15632
rect 15200 15512 15252 15564
rect 25964 15580 26016 15632
rect 29736 15580 29788 15632
rect 34520 15580 34572 15632
rect 14924 15444 14976 15453
rect 15752 15444 15804 15496
rect 16856 15487 16908 15496
rect 10600 15351 10652 15360
rect 10600 15317 10609 15351
rect 10609 15317 10643 15351
rect 10643 15317 10652 15351
rect 10600 15308 10652 15317
rect 11336 15308 11388 15360
rect 12808 15376 12860 15428
rect 13176 15419 13228 15428
rect 13176 15385 13185 15419
rect 13185 15385 13219 15419
rect 13219 15385 13228 15419
rect 13176 15376 13228 15385
rect 16856 15453 16865 15487
rect 16865 15453 16899 15487
rect 16899 15453 16908 15487
rect 16856 15444 16908 15453
rect 17040 15487 17092 15496
rect 17040 15453 17047 15487
rect 17047 15453 17092 15487
rect 17040 15444 17092 15453
rect 17224 15487 17276 15496
rect 17224 15453 17233 15487
rect 17233 15453 17267 15487
rect 17267 15453 17276 15487
rect 17224 15444 17276 15453
rect 17316 15487 17368 15496
rect 17316 15453 17330 15487
rect 17330 15453 17364 15487
rect 17364 15453 17368 15487
rect 17316 15444 17368 15453
rect 18052 15444 18104 15496
rect 20260 15444 20312 15496
rect 24400 15487 24452 15496
rect 24400 15453 24409 15487
rect 24409 15453 24443 15487
rect 24443 15453 24452 15487
rect 24400 15444 24452 15453
rect 25228 15487 25280 15496
rect 25228 15453 25237 15487
rect 25237 15453 25271 15487
rect 25271 15453 25280 15487
rect 25228 15444 25280 15453
rect 26884 15444 26936 15496
rect 27528 15512 27580 15564
rect 27804 15512 27856 15564
rect 30564 15512 30616 15564
rect 31116 15512 31168 15564
rect 31484 15555 31536 15564
rect 31484 15521 31493 15555
rect 31493 15521 31527 15555
rect 31527 15521 31536 15555
rect 31484 15512 31536 15521
rect 27620 15444 27672 15496
rect 28540 15444 28592 15496
rect 15936 15376 15988 15428
rect 18420 15376 18472 15428
rect 18972 15376 19024 15428
rect 21272 15376 21324 15428
rect 21824 15376 21876 15428
rect 22008 15419 22060 15428
rect 22008 15385 22017 15419
rect 22017 15385 22051 15419
rect 22051 15385 22060 15419
rect 22008 15376 22060 15385
rect 13544 15351 13596 15360
rect 13544 15317 13553 15351
rect 13553 15317 13587 15351
rect 13587 15317 13596 15351
rect 13544 15308 13596 15317
rect 14372 15308 14424 15360
rect 14924 15308 14976 15360
rect 18236 15308 18288 15360
rect 22836 15308 22888 15360
rect 25320 15376 25372 15428
rect 25688 15308 25740 15360
rect 28264 15419 28316 15428
rect 28264 15385 28273 15419
rect 28273 15385 28307 15419
rect 28307 15385 28316 15419
rect 28264 15376 28316 15385
rect 29000 15376 29052 15428
rect 29644 15444 29696 15496
rect 29828 15487 29880 15496
rect 29828 15453 29837 15487
rect 29837 15453 29871 15487
rect 29871 15453 29880 15487
rect 29828 15444 29880 15453
rect 30012 15487 30064 15496
rect 30012 15453 30021 15487
rect 30021 15453 30055 15487
rect 30055 15453 30064 15487
rect 30012 15444 30064 15453
rect 30196 15487 30248 15496
rect 30196 15453 30205 15487
rect 30205 15453 30239 15487
rect 30239 15453 30248 15487
rect 31760 15487 31812 15496
rect 30196 15444 30248 15453
rect 30288 15376 30340 15428
rect 31760 15453 31769 15487
rect 31769 15453 31803 15487
rect 31803 15453 31812 15487
rect 31760 15444 31812 15453
rect 31116 15376 31168 15428
rect 33416 15444 33468 15496
rect 33600 15444 33652 15496
rect 35348 15444 35400 15496
rect 36176 15444 36228 15496
rect 39304 15487 39356 15496
rect 39304 15453 39313 15487
rect 39313 15453 39347 15487
rect 39347 15453 39356 15487
rect 39304 15444 39356 15453
rect 34796 15376 34848 15428
rect 30380 15308 30432 15360
rect 30840 15308 30892 15360
rect 32128 15308 32180 15360
rect 33692 15308 33744 15360
rect 33784 15308 33836 15360
rect 37648 15376 37700 15428
rect 38660 15376 38712 15428
rect 37924 15351 37976 15360
rect 37924 15317 37933 15351
rect 37933 15317 37967 15351
rect 37967 15317 37976 15351
rect 37924 15308 37976 15317
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 50294 15206 50346 15258
rect 50358 15206 50410 15258
rect 50422 15206 50474 15258
rect 50486 15206 50538 15258
rect 50550 15206 50602 15258
rect 3148 15104 3200 15156
rect 4896 15147 4948 15156
rect 4896 15113 4905 15147
rect 4905 15113 4939 15147
rect 4939 15113 4948 15147
rect 4896 15104 4948 15113
rect 7840 15104 7892 15156
rect 8944 15104 8996 15156
rect 2596 14968 2648 15020
rect 4712 15036 4764 15088
rect 7472 15036 7524 15088
rect 11060 15104 11112 15156
rect 12624 15104 12676 15156
rect 11704 15036 11756 15088
rect 13176 15036 13228 15088
rect 5172 14968 5224 15020
rect 5356 15011 5408 15020
rect 5356 14977 5365 15011
rect 5365 14977 5399 15011
rect 5399 14977 5408 15011
rect 5356 14968 5408 14977
rect 7564 14968 7616 15020
rect 8392 15011 8444 15020
rect 8392 14977 8401 15011
rect 8401 14977 8435 15011
rect 8435 14977 8444 15011
rect 8392 14968 8444 14977
rect 8852 14968 8904 15020
rect 10232 14968 10284 15020
rect 11796 15011 11848 15020
rect 11796 14977 11805 15011
rect 11805 14977 11839 15011
rect 11839 14977 11848 15011
rect 11796 14968 11848 14977
rect 11980 15011 12032 15020
rect 11980 14977 11989 15011
rect 11989 14977 12023 15011
rect 12023 14977 12032 15011
rect 12532 15011 12584 15020
rect 11980 14968 12032 14977
rect 12532 14977 12541 15011
rect 12541 14977 12575 15011
rect 12575 14977 12584 15011
rect 12532 14968 12584 14977
rect 12716 15011 12768 15020
rect 12716 14977 12723 15011
rect 12723 14977 12768 15011
rect 12716 14968 12768 14977
rect 5264 14943 5316 14952
rect 5264 14909 5273 14943
rect 5273 14909 5307 14943
rect 5307 14909 5316 14943
rect 5264 14900 5316 14909
rect 8392 14832 8444 14884
rect 11704 14900 11756 14952
rect 12992 15011 13044 15020
rect 12992 14977 13006 15011
rect 13006 14977 13040 15011
rect 13040 14977 13044 15011
rect 12992 14968 13044 14977
rect 13728 14968 13780 15020
rect 16948 15104 17000 15156
rect 17224 15104 17276 15156
rect 18052 15104 18104 15156
rect 19064 15104 19116 15156
rect 20260 15147 20312 15156
rect 20260 15113 20269 15147
rect 20269 15113 20303 15147
rect 20303 15113 20312 15147
rect 20260 15104 20312 15113
rect 22744 15104 22796 15156
rect 14188 15036 14240 15088
rect 14648 15036 14700 15088
rect 16580 15036 16632 15088
rect 17684 15079 17736 15088
rect 17684 15045 17693 15079
rect 17693 15045 17727 15079
rect 17727 15045 17736 15079
rect 18420 15079 18472 15088
rect 17684 15036 17736 15045
rect 18420 15045 18429 15079
rect 18429 15045 18463 15079
rect 18463 15045 18472 15079
rect 18420 15036 18472 15045
rect 14280 15011 14332 15020
rect 14280 14977 14289 15011
rect 14289 14977 14323 15011
rect 14323 14977 14332 15011
rect 14280 14968 14332 14977
rect 15016 14968 15068 15020
rect 15292 14968 15344 15020
rect 15752 15011 15804 15020
rect 15752 14977 15761 15011
rect 15761 14977 15795 15011
rect 15795 14977 15804 15011
rect 15752 14968 15804 14977
rect 17408 14900 17460 14952
rect 17776 14968 17828 15020
rect 28264 15104 28316 15156
rect 19248 15036 19300 15088
rect 22928 15036 22980 15088
rect 24768 15036 24820 15088
rect 26240 15036 26292 15088
rect 30012 15104 30064 15156
rect 30656 15147 30708 15156
rect 30656 15113 30665 15147
rect 30665 15113 30699 15147
rect 30699 15113 30708 15147
rect 30656 15104 30708 15113
rect 31484 15104 31536 15156
rect 31760 15104 31812 15156
rect 20904 15011 20956 15020
rect 20904 14977 20913 15011
rect 20913 14977 20947 15011
rect 20947 14977 20956 15011
rect 20904 14968 20956 14977
rect 18880 14943 18932 14952
rect 5448 14764 5500 14816
rect 6184 14764 6236 14816
rect 7012 14764 7064 14816
rect 7104 14764 7156 14816
rect 15752 14832 15804 14884
rect 16304 14832 16356 14884
rect 17684 14832 17736 14884
rect 11980 14764 12032 14816
rect 12992 14764 13044 14816
rect 15292 14764 15344 14816
rect 15936 14764 15988 14816
rect 17776 14764 17828 14816
rect 18880 14909 18889 14943
rect 18889 14909 18923 14943
rect 18923 14909 18932 14943
rect 18880 14900 18932 14909
rect 20812 14900 20864 14952
rect 19984 14832 20036 14884
rect 22284 14968 22336 15020
rect 23480 14968 23532 15020
rect 24952 14968 25004 15020
rect 25044 15011 25096 15020
rect 25044 14977 25053 15011
rect 25053 14977 25087 15011
rect 25087 14977 25096 15011
rect 25044 14968 25096 14977
rect 25688 14968 25740 15020
rect 24216 14943 24268 14952
rect 24216 14909 24225 14943
rect 24225 14909 24259 14943
rect 24259 14909 24268 14943
rect 24216 14900 24268 14909
rect 28172 14968 28224 15020
rect 30196 15036 30248 15088
rect 28632 15011 28684 15020
rect 28632 14977 28641 15011
rect 28641 14977 28675 15011
rect 28675 14977 28684 15011
rect 28632 14968 28684 14977
rect 30288 15011 30340 15020
rect 30288 14977 30297 15011
rect 30297 14977 30331 15011
rect 30331 14977 30340 15011
rect 30288 14968 30340 14977
rect 17960 14764 18012 14816
rect 21272 14807 21324 14816
rect 21272 14773 21281 14807
rect 21281 14773 21315 14807
rect 21315 14773 21324 14807
rect 21272 14764 21324 14773
rect 22560 14764 22612 14816
rect 24860 14832 24912 14884
rect 25228 14832 25280 14884
rect 25412 14807 25464 14816
rect 25412 14773 25421 14807
rect 25421 14773 25455 14807
rect 25455 14773 25464 14807
rect 25412 14764 25464 14773
rect 28080 14764 28132 14816
rect 28172 14764 28224 14816
rect 28816 14807 28868 14816
rect 28816 14773 28825 14807
rect 28825 14773 28859 14807
rect 28859 14773 28868 14807
rect 28816 14764 28868 14773
rect 30012 14900 30064 14952
rect 30656 14968 30708 15020
rect 31024 14968 31076 15020
rect 31392 15011 31444 15020
rect 31392 14977 31401 15011
rect 31401 14977 31435 15011
rect 31435 14977 31444 15011
rect 31392 14968 31444 14977
rect 32128 15011 32180 15020
rect 32128 14977 32137 15011
rect 32137 14977 32171 15011
rect 32171 14977 32180 15011
rect 32128 14968 32180 14977
rect 32312 15011 32364 15020
rect 32312 14977 32321 15011
rect 32321 14977 32355 15011
rect 32355 14977 32364 15011
rect 32312 14968 32364 14977
rect 35440 15104 35492 15156
rect 36636 15147 36688 15156
rect 36636 15113 36645 15147
rect 36645 15113 36679 15147
rect 36679 15113 36688 15147
rect 36636 15104 36688 15113
rect 33508 15079 33560 15088
rect 33508 15045 33517 15079
rect 33517 15045 33551 15079
rect 33551 15045 33560 15079
rect 33508 15036 33560 15045
rect 33968 15036 34020 15088
rect 36912 15036 36964 15088
rect 37372 15036 37424 15088
rect 32864 14968 32916 15020
rect 34796 14968 34848 15020
rect 34704 14900 34756 14952
rect 37464 15011 37516 15020
rect 37464 14977 37473 15011
rect 37473 14977 37507 15011
rect 37507 14977 37516 15011
rect 37464 14968 37516 14977
rect 38660 15104 38712 15156
rect 41420 15104 41472 15156
rect 35256 14900 35308 14952
rect 35532 14900 35584 14952
rect 30196 14832 30248 14884
rect 31208 14832 31260 14884
rect 32680 14832 32732 14884
rect 37924 14832 37976 14884
rect 32772 14807 32824 14816
rect 32772 14773 32781 14807
rect 32781 14773 32815 14807
rect 32815 14773 32824 14807
rect 32772 14764 32824 14773
rect 37096 14764 37148 14816
rect 38384 14968 38436 15020
rect 39304 14764 39356 14816
rect 39856 14764 39908 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 65654 14662 65706 14714
rect 65718 14662 65770 14714
rect 65782 14662 65834 14714
rect 65846 14662 65898 14714
rect 65910 14662 65962 14714
rect 2872 14560 2924 14612
rect 3332 14560 3384 14612
rect 8576 14560 8628 14612
rect 8760 14560 8812 14612
rect 9036 14560 9088 14612
rect 12532 14560 12584 14612
rect 14004 14560 14056 14612
rect 14648 14560 14700 14612
rect 15844 14560 15896 14612
rect 7472 14424 7524 14476
rect 7196 14399 7248 14408
rect 7196 14365 7205 14399
rect 7205 14365 7239 14399
rect 7239 14365 7248 14399
rect 7196 14356 7248 14365
rect 7748 14356 7800 14408
rect 10968 14424 11020 14476
rect 5264 14288 5316 14340
rect 2320 14220 2372 14272
rect 5632 14220 5684 14272
rect 9404 14288 9456 14340
rect 10416 14356 10468 14408
rect 10508 14356 10560 14408
rect 11152 14399 11204 14408
rect 11152 14365 11161 14399
rect 11161 14365 11195 14399
rect 11195 14365 11204 14399
rect 11152 14356 11204 14365
rect 11244 14399 11296 14408
rect 11244 14365 11253 14399
rect 11253 14365 11287 14399
rect 11287 14365 11296 14399
rect 11244 14356 11296 14365
rect 12348 14356 12400 14408
rect 12716 14399 12768 14408
rect 12716 14365 12725 14399
rect 12725 14365 12759 14399
rect 12759 14365 12768 14399
rect 12716 14356 12768 14365
rect 16028 14492 16080 14544
rect 16580 14492 16632 14544
rect 16304 14467 16356 14476
rect 16304 14433 16313 14467
rect 16313 14433 16347 14467
rect 16347 14433 16356 14467
rect 16304 14424 16356 14433
rect 17868 14560 17920 14612
rect 20444 14560 20496 14612
rect 23204 14603 23256 14612
rect 23204 14569 23213 14603
rect 23213 14569 23247 14603
rect 23247 14569 23256 14603
rect 23204 14560 23256 14569
rect 24400 14603 24452 14612
rect 24400 14569 24409 14603
rect 24409 14569 24443 14603
rect 24443 14569 24452 14603
rect 24400 14560 24452 14569
rect 28356 14603 28408 14612
rect 19156 14492 19208 14544
rect 19340 14535 19392 14544
rect 19340 14501 19349 14535
rect 19349 14501 19383 14535
rect 19383 14501 19392 14535
rect 19340 14492 19392 14501
rect 9128 14220 9180 14272
rect 11428 14288 11480 14340
rect 14648 14331 14700 14340
rect 14648 14297 14657 14331
rect 14657 14297 14691 14331
rect 14691 14297 14700 14331
rect 14648 14288 14700 14297
rect 14740 14331 14792 14340
rect 14740 14297 14749 14331
rect 14749 14297 14783 14331
rect 14783 14297 14792 14331
rect 14740 14288 14792 14297
rect 10416 14263 10468 14272
rect 10416 14229 10425 14263
rect 10425 14229 10459 14263
rect 10459 14229 10468 14263
rect 10416 14220 10468 14229
rect 11796 14220 11848 14272
rect 13452 14220 13504 14272
rect 13636 14220 13688 14272
rect 15844 14356 15896 14408
rect 17960 14424 18012 14476
rect 16580 14356 16632 14408
rect 17316 14356 17368 14408
rect 23020 14492 23072 14544
rect 20628 14424 20680 14476
rect 22008 14424 22060 14476
rect 20444 14356 20496 14408
rect 21916 14356 21968 14408
rect 25320 14399 25372 14408
rect 17592 14288 17644 14340
rect 20812 14288 20864 14340
rect 22192 14288 22244 14340
rect 25320 14365 25329 14399
rect 25329 14365 25363 14399
rect 25363 14365 25372 14399
rect 25320 14356 25372 14365
rect 25780 14424 25832 14476
rect 28356 14569 28365 14603
rect 28365 14569 28399 14603
rect 28399 14569 28408 14603
rect 28356 14560 28408 14569
rect 30196 14603 30248 14612
rect 30196 14569 30205 14603
rect 30205 14569 30239 14603
rect 30239 14569 30248 14603
rect 30196 14560 30248 14569
rect 30288 14560 30340 14612
rect 32312 14560 32364 14612
rect 33784 14560 33836 14612
rect 38384 14603 38436 14612
rect 38384 14569 38393 14603
rect 38393 14569 38427 14603
rect 38427 14569 38436 14603
rect 38384 14560 38436 14569
rect 28816 14492 28868 14544
rect 29000 14424 29052 14476
rect 26056 14356 26108 14408
rect 26240 14399 26292 14408
rect 26240 14365 26249 14399
rect 26249 14365 26283 14399
rect 26283 14365 26292 14399
rect 26240 14356 26292 14365
rect 21088 14263 21140 14272
rect 21088 14229 21097 14263
rect 21097 14229 21131 14263
rect 21131 14229 21140 14263
rect 21088 14220 21140 14229
rect 22376 14263 22428 14272
rect 22376 14229 22385 14263
rect 22385 14229 22419 14263
rect 22419 14229 22428 14263
rect 22376 14220 22428 14229
rect 25596 14220 25648 14272
rect 26332 14220 26384 14272
rect 31024 14399 31076 14408
rect 31024 14365 31033 14399
rect 31033 14365 31067 14399
rect 31067 14365 31076 14399
rect 31024 14356 31076 14365
rect 31392 14424 31444 14476
rect 32680 14424 32732 14476
rect 32496 14356 32548 14408
rect 37740 14492 37792 14544
rect 35440 14424 35492 14476
rect 35532 14399 35584 14408
rect 35532 14365 35541 14399
rect 35541 14365 35575 14399
rect 35575 14365 35584 14399
rect 35532 14356 35584 14365
rect 37648 14356 37700 14408
rect 68100 14399 68152 14408
rect 27804 14288 27856 14340
rect 29920 14331 29972 14340
rect 29920 14297 29929 14331
rect 29929 14297 29963 14331
rect 29963 14297 29972 14331
rect 29920 14288 29972 14297
rect 30840 14331 30892 14340
rect 30840 14297 30849 14331
rect 30849 14297 30883 14331
rect 30883 14297 30892 14331
rect 30840 14288 30892 14297
rect 33140 14288 33192 14340
rect 33324 14288 33376 14340
rect 34520 14288 34572 14340
rect 36912 14331 36964 14340
rect 36912 14297 36921 14331
rect 36921 14297 36955 14331
rect 36955 14297 36964 14331
rect 36912 14288 36964 14297
rect 37096 14331 37148 14340
rect 37096 14297 37105 14331
rect 37105 14297 37139 14331
rect 37139 14297 37148 14331
rect 37096 14288 37148 14297
rect 27528 14220 27580 14272
rect 28908 14263 28960 14272
rect 28908 14229 28917 14263
rect 28917 14229 28951 14263
rect 28951 14229 28960 14263
rect 28908 14220 28960 14229
rect 37832 14220 37884 14272
rect 68100 14365 68109 14399
rect 68109 14365 68143 14399
rect 68143 14365 68152 14399
rect 68100 14356 68152 14365
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 50294 14118 50346 14170
rect 50358 14118 50410 14170
rect 50422 14118 50474 14170
rect 50486 14118 50538 14170
rect 50550 14118 50602 14170
rect 2688 14016 2740 14068
rect 7104 14016 7156 14068
rect 7748 14059 7800 14068
rect 7748 14025 7757 14059
rect 7757 14025 7791 14059
rect 7791 14025 7800 14059
rect 7748 14016 7800 14025
rect 9036 14059 9088 14068
rect 9036 14025 9045 14059
rect 9045 14025 9079 14059
rect 9079 14025 9088 14059
rect 9036 14016 9088 14025
rect 9128 14016 9180 14068
rect 17592 14016 17644 14068
rect 18328 14016 18380 14068
rect 19892 14059 19944 14068
rect 19892 14025 19901 14059
rect 19901 14025 19935 14059
rect 19935 14025 19944 14059
rect 19892 14016 19944 14025
rect 22192 14016 22244 14068
rect 22560 14016 22612 14068
rect 24952 14059 25004 14068
rect 24952 14025 24961 14059
rect 24961 14025 24995 14059
rect 24995 14025 25004 14059
rect 24952 14016 25004 14025
rect 25320 14016 25372 14068
rect 29092 14016 29144 14068
rect 31024 14016 31076 14068
rect 31668 14016 31720 14068
rect 2504 13923 2556 13932
rect 2504 13889 2513 13923
rect 2513 13889 2547 13923
rect 2547 13889 2556 13923
rect 2504 13880 2556 13889
rect 3056 13948 3108 14000
rect 8760 13991 8812 14000
rect 8760 13957 8769 13991
rect 8769 13957 8803 13991
rect 8803 13957 8812 13991
rect 8760 13948 8812 13957
rect 9588 13948 9640 14000
rect 1492 13855 1544 13864
rect 1492 13821 1501 13855
rect 1501 13821 1535 13855
rect 1535 13821 1544 13855
rect 1492 13812 1544 13821
rect 2872 13923 2924 13932
rect 2872 13889 2881 13923
rect 2881 13889 2915 13923
rect 2915 13889 2924 13923
rect 3608 13923 3660 13932
rect 2872 13880 2924 13889
rect 3608 13889 3617 13923
rect 3617 13889 3651 13923
rect 3651 13889 3660 13923
rect 3608 13880 3660 13889
rect 6092 13880 6144 13932
rect 8300 13880 8352 13932
rect 8668 13880 8720 13932
rect 8852 13923 8904 13932
rect 8852 13889 8861 13923
rect 8861 13889 8895 13923
rect 8895 13889 8904 13923
rect 8852 13880 8904 13889
rect 9404 13880 9456 13932
rect 15844 13948 15896 14000
rect 19156 13948 19208 14000
rect 12992 13880 13044 13932
rect 13452 13880 13504 13932
rect 15476 13923 15528 13932
rect 15476 13889 15485 13923
rect 15485 13889 15519 13923
rect 15519 13889 15528 13923
rect 15476 13880 15528 13889
rect 17040 13923 17092 13932
rect 6368 13855 6420 13864
rect 6368 13821 6377 13855
rect 6377 13821 6411 13855
rect 6411 13821 6420 13855
rect 6368 13812 6420 13821
rect 10324 13855 10376 13864
rect 10324 13821 10333 13855
rect 10333 13821 10367 13855
rect 10367 13821 10376 13855
rect 10324 13812 10376 13821
rect 11244 13812 11296 13864
rect 11520 13855 11572 13864
rect 11520 13821 11529 13855
rect 11529 13821 11563 13855
rect 11563 13821 11572 13855
rect 11520 13812 11572 13821
rect 12808 13812 12860 13864
rect 13636 13855 13688 13864
rect 13636 13821 13645 13855
rect 13645 13821 13679 13855
rect 13679 13821 13688 13855
rect 13636 13812 13688 13821
rect 16396 13812 16448 13864
rect 17040 13889 17049 13923
rect 17049 13889 17083 13923
rect 17083 13889 17092 13923
rect 17040 13880 17092 13889
rect 17224 13923 17276 13932
rect 17224 13889 17231 13923
rect 17231 13889 17276 13923
rect 17224 13880 17276 13889
rect 17408 13923 17460 13932
rect 17408 13889 17417 13923
rect 17417 13889 17451 13923
rect 17451 13889 17460 13923
rect 17408 13880 17460 13889
rect 17500 13923 17552 13932
rect 17500 13889 17514 13923
rect 17514 13889 17548 13923
rect 17548 13889 17552 13923
rect 17500 13880 17552 13889
rect 17684 13880 17736 13932
rect 20904 13948 20956 14000
rect 19708 13923 19760 13932
rect 19708 13889 19717 13923
rect 19717 13889 19751 13923
rect 19751 13889 19760 13923
rect 19708 13880 19760 13889
rect 20260 13880 20312 13932
rect 20720 13880 20772 13932
rect 2872 13744 2924 13796
rect 13268 13744 13320 13796
rect 18052 13744 18104 13796
rect 2780 13676 2832 13728
rect 3608 13676 3660 13728
rect 3792 13676 3844 13728
rect 10692 13676 10744 13728
rect 13820 13676 13872 13728
rect 14372 13676 14424 13728
rect 19432 13812 19484 13864
rect 20536 13812 20588 13864
rect 18972 13744 19024 13796
rect 22836 13812 22888 13864
rect 25136 13880 25188 13932
rect 25780 13948 25832 14000
rect 26056 13991 26108 14000
rect 26056 13957 26065 13991
rect 26065 13957 26099 13991
rect 26099 13957 26108 13991
rect 26056 13948 26108 13957
rect 29276 13991 29328 14000
rect 29276 13957 29285 13991
rect 29285 13957 29319 13991
rect 29319 13957 29328 13991
rect 29276 13948 29328 13957
rect 32772 13948 32824 14000
rect 33508 13948 33560 14000
rect 34520 13991 34572 14000
rect 34520 13957 34529 13991
rect 34529 13957 34563 13991
rect 34563 13957 34572 13991
rect 34520 13948 34572 13957
rect 37372 14016 37424 14068
rect 25412 13923 25464 13932
rect 25412 13889 25426 13923
rect 25426 13889 25460 13923
rect 25460 13889 25464 13923
rect 25412 13880 25464 13889
rect 25596 13923 25648 13932
rect 25596 13889 25605 13923
rect 25605 13889 25639 13923
rect 25639 13889 25648 13923
rect 25596 13880 25648 13889
rect 26148 13880 26200 13932
rect 27528 13880 27580 13932
rect 27804 13880 27856 13932
rect 29184 13923 29236 13932
rect 29184 13889 29193 13923
rect 29193 13889 29227 13923
rect 29227 13889 29236 13923
rect 29184 13880 29236 13889
rect 29552 13923 29604 13932
rect 25780 13812 25832 13864
rect 26792 13812 26844 13864
rect 27620 13812 27672 13864
rect 28172 13812 28224 13864
rect 28540 13812 28592 13864
rect 29552 13889 29561 13923
rect 29561 13889 29595 13923
rect 29595 13889 29604 13923
rect 29552 13880 29604 13889
rect 34704 13923 34756 13932
rect 34704 13889 34713 13923
rect 34713 13889 34747 13923
rect 34747 13889 34756 13923
rect 34704 13880 34756 13889
rect 35348 13923 35400 13932
rect 35348 13889 35357 13923
rect 35357 13889 35391 13923
rect 35391 13889 35400 13923
rect 35348 13880 35400 13889
rect 35624 13923 35676 13932
rect 35624 13889 35658 13923
rect 35658 13889 35676 13923
rect 37648 13923 37700 13932
rect 35624 13880 35676 13889
rect 37648 13889 37657 13923
rect 37657 13889 37691 13923
rect 37691 13889 37700 13923
rect 37648 13880 37700 13889
rect 26240 13744 26292 13796
rect 27252 13744 27304 13796
rect 37924 13923 37976 13932
rect 37924 13889 37936 13923
rect 37936 13889 37970 13923
rect 37970 13889 37976 13923
rect 37924 13880 37976 13889
rect 38200 13880 38252 13932
rect 39948 13812 40000 13864
rect 29092 13744 29144 13796
rect 29828 13744 29880 13796
rect 37740 13744 37792 13796
rect 19616 13676 19668 13728
rect 20260 13676 20312 13728
rect 27528 13676 27580 13728
rect 29644 13676 29696 13728
rect 34796 13676 34848 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 65654 13574 65706 13626
rect 65718 13574 65770 13626
rect 65782 13574 65834 13626
rect 65846 13574 65898 13626
rect 65910 13574 65962 13626
rect 2872 13515 2924 13524
rect 2872 13481 2881 13515
rect 2881 13481 2915 13515
rect 2915 13481 2924 13515
rect 2872 13472 2924 13481
rect 2964 13472 3016 13524
rect 6092 13515 6144 13524
rect 6092 13481 6101 13515
rect 6101 13481 6135 13515
rect 6135 13481 6144 13515
rect 6092 13472 6144 13481
rect 13728 13472 13780 13524
rect 13820 13472 13872 13524
rect 14556 13515 14608 13524
rect 14556 13481 14565 13515
rect 14565 13481 14599 13515
rect 14599 13481 14608 13515
rect 14556 13472 14608 13481
rect 15476 13472 15528 13524
rect 15844 13472 15896 13524
rect 16488 13472 16540 13524
rect 2504 13336 2556 13388
rect 11336 13404 11388 13456
rect 2688 13311 2740 13320
rect 2688 13277 2697 13311
rect 2697 13277 2731 13311
rect 2731 13277 2740 13311
rect 2688 13268 2740 13277
rect 5632 13311 5684 13320
rect 5632 13277 5641 13311
rect 5641 13277 5675 13311
rect 5675 13277 5684 13311
rect 5632 13268 5684 13277
rect 6552 13311 6604 13320
rect 2596 13200 2648 13252
rect 3056 13200 3108 13252
rect 6552 13277 6561 13311
rect 6561 13277 6595 13311
rect 6595 13277 6604 13311
rect 6552 13268 6604 13277
rect 8668 13336 8720 13388
rect 9588 13336 9640 13388
rect 11520 13336 11572 13388
rect 19984 13472 20036 13524
rect 22468 13472 22520 13524
rect 24032 13472 24084 13524
rect 28540 13472 28592 13524
rect 28724 13515 28776 13524
rect 28724 13481 28733 13515
rect 28733 13481 28767 13515
rect 28767 13481 28776 13515
rect 28724 13472 28776 13481
rect 29828 13472 29880 13524
rect 12440 13336 12492 13388
rect 13452 13336 13504 13388
rect 8392 13268 8444 13320
rect 8944 13311 8996 13320
rect 8944 13277 8953 13311
rect 8953 13277 8987 13311
rect 8987 13277 8996 13311
rect 8944 13268 8996 13277
rect 7380 13200 7432 13252
rect 9404 13268 9456 13320
rect 11428 13311 11480 13320
rect 11428 13277 11437 13311
rect 11437 13277 11471 13311
rect 11471 13277 11480 13311
rect 11428 13268 11480 13277
rect 12900 13311 12952 13320
rect 12900 13277 12909 13311
rect 12909 13277 12943 13311
rect 12943 13277 12952 13311
rect 12900 13268 12952 13277
rect 15660 13336 15712 13388
rect 16488 13336 16540 13388
rect 16580 13336 16632 13388
rect 6828 13132 6880 13184
rect 8852 13132 8904 13184
rect 14648 13243 14700 13252
rect 14648 13209 14657 13243
rect 14657 13209 14691 13243
rect 14691 13209 14700 13243
rect 14648 13200 14700 13209
rect 10876 13132 10928 13184
rect 15844 13311 15896 13320
rect 15844 13277 15853 13311
rect 15853 13277 15887 13311
rect 15887 13277 15896 13311
rect 15844 13268 15896 13277
rect 16028 13268 16080 13320
rect 18972 13336 19024 13388
rect 19064 13336 19116 13388
rect 20352 13336 20404 13388
rect 16764 13200 16816 13252
rect 17500 13200 17552 13252
rect 19340 13268 19392 13320
rect 19432 13311 19484 13320
rect 19432 13277 19441 13311
rect 19441 13277 19475 13311
rect 19475 13277 19484 13311
rect 19432 13268 19484 13277
rect 19984 13268 20036 13320
rect 20720 13311 20772 13320
rect 20720 13277 20729 13311
rect 20729 13277 20763 13311
rect 20763 13277 20772 13311
rect 24308 13404 24360 13456
rect 26516 13447 26568 13456
rect 26516 13413 26525 13447
rect 26525 13413 26559 13447
rect 26559 13413 26568 13447
rect 26516 13404 26568 13413
rect 31392 13447 31444 13456
rect 21272 13336 21324 13388
rect 20720 13268 20772 13277
rect 21640 13311 21692 13320
rect 21640 13277 21649 13311
rect 21649 13277 21683 13311
rect 21683 13277 21692 13311
rect 21640 13268 21692 13277
rect 22008 13268 22060 13320
rect 22560 13311 22612 13320
rect 22560 13277 22569 13311
rect 22569 13277 22603 13311
rect 22603 13277 22612 13311
rect 22560 13268 22612 13277
rect 23388 13311 23440 13320
rect 23388 13277 23397 13311
rect 23397 13277 23431 13311
rect 23431 13277 23440 13311
rect 23388 13268 23440 13277
rect 25136 13336 25188 13388
rect 23756 13311 23808 13320
rect 23756 13277 23765 13311
rect 23765 13277 23799 13311
rect 23799 13277 23808 13311
rect 23756 13268 23808 13277
rect 25596 13268 25648 13320
rect 27436 13311 27488 13320
rect 27436 13277 27445 13311
rect 27445 13277 27479 13311
rect 27479 13277 27488 13311
rect 27436 13268 27488 13277
rect 31392 13413 31401 13447
rect 31401 13413 31435 13447
rect 31435 13413 31444 13447
rect 31392 13404 31444 13413
rect 34980 13472 35032 13524
rect 35440 13472 35492 13524
rect 35624 13515 35676 13524
rect 35624 13481 35633 13515
rect 35633 13481 35667 13515
rect 35667 13481 35676 13515
rect 35624 13472 35676 13481
rect 36636 13472 36688 13524
rect 37004 13472 37056 13524
rect 37740 13515 37792 13524
rect 37740 13481 37749 13515
rect 37749 13481 37783 13515
rect 37783 13481 37792 13515
rect 37740 13472 37792 13481
rect 38200 13515 38252 13524
rect 38200 13481 38209 13515
rect 38209 13481 38243 13515
rect 38243 13481 38252 13515
rect 38200 13472 38252 13481
rect 30196 13336 30248 13388
rect 28264 13311 28316 13320
rect 28264 13277 28271 13311
rect 28271 13277 28316 13311
rect 28264 13268 28316 13277
rect 28356 13311 28408 13320
rect 28356 13277 28365 13311
rect 28365 13277 28399 13311
rect 28399 13277 28408 13311
rect 28356 13268 28408 13277
rect 29460 13268 29512 13320
rect 29644 13268 29696 13320
rect 34796 13336 34848 13388
rect 35808 13404 35860 13456
rect 31392 13268 31444 13320
rect 31668 13311 31720 13320
rect 31668 13277 31677 13311
rect 31677 13277 31711 13311
rect 31711 13277 31720 13311
rect 31668 13268 31720 13277
rect 33508 13268 33560 13320
rect 34152 13268 34204 13320
rect 34980 13311 35032 13320
rect 34980 13277 34989 13311
rect 34989 13277 35023 13311
rect 35023 13277 35032 13311
rect 34980 13268 35032 13277
rect 36912 13268 36964 13320
rect 39856 13311 39908 13320
rect 39856 13277 39865 13311
rect 39865 13277 39899 13311
rect 39899 13277 39908 13311
rect 39856 13268 39908 13277
rect 39948 13268 40000 13320
rect 20444 13200 20496 13252
rect 20812 13243 20864 13252
rect 20812 13209 20821 13243
rect 20821 13209 20855 13243
rect 20855 13209 20864 13243
rect 20812 13200 20864 13209
rect 15844 13132 15896 13184
rect 16304 13132 16356 13184
rect 18144 13132 18196 13184
rect 19616 13132 19668 13184
rect 23664 13200 23716 13252
rect 25044 13200 25096 13252
rect 26148 13200 26200 13252
rect 26332 13243 26384 13252
rect 26332 13209 26341 13243
rect 26341 13209 26375 13243
rect 26375 13209 26384 13243
rect 26332 13200 26384 13209
rect 24676 13175 24728 13184
rect 24676 13141 24685 13175
rect 24685 13141 24719 13175
rect 24719 13141 24728 13175
rect 24676 13132 24728 13141
rect 25964 13132 26016 13184
rect 27436 13132 27488 13184
rect 27988 13132 28040 13184
rect 29920 13132 29972 13184
rect 30196 13243 30248 13252
rect 30196 13209 30205 13243
rect 30205 13209 30239 13243
rect 30239 13209 30248 13243
rect 30196 13200 30248 13209
rect 30656 13132 30708 13184
rect 33876 13200 33928 13252
rect 37648 13200 37700 13252
rect 33968 13132 34020 13184
rect 35256 13132 35308 13184
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 50294 13030 50346 13082
rect 50358 13030 50410 13082
rect 50422 13030 50474 13082
rect 50486 13030 50538 13082
rect 50550 13030 50602 13082
rect 2044 12792 2096 12844
rect 4620 12928 4672 12980
rect 2596 12860 2648 12912
rect 3792 12860 3844 12912
rect 8944 12860 8996 12912
rect 10048 12928 10100 12980
rect 10876 12971 10928 12980
rect 10876 12937 10885 12971
rect 10885 12937 10919 12971
rect 10919 12937 10928 12971
rect 10876 12928 10928 12937
rect 11336 12928 11388 12980
rect 11704 12971 11756 12980
rect 11704 12937 11713 12971
rect 11713 12937 11747 12971
rect 11747 12937 11756 12971
rect 11704 12928 11756 12937
rect 12072 12928 12124 12980
rect 13268 12928 13320 12980
rect 17224 12928 17276 12980
rect 18052 12928 18104 12980
rect 18788 12928 18840 12980
rect 18972 12971 19024 12980
rect 18972 12937 18981 12971
rect 18981 12937 19015 12971
rect 19015 12937 19024 12971
rect 18972 12928 19024 12937
rect 20996 12928 21048 12980
rect 21640 12928 21692 12980
rect 22284 12928 22336 12980
rect 22560 12928 22612 12980
rect 11612 12903 11664 12912
rect 11612 12869 11621 12903
rect 11621 12869 11655 12903
rect 11655 12869 11664 12903
rect 11612 12860 11664 12869
rect 3148 12792 3200 12844
rect 7748 12835 7800 12844
rect 7748 12801 7757 12835
rect 7757 12801 7791 12835
rect 7791 12801 7800 12835
rect 7748 12792 7800 12801
rect 9680 12835 9732 12844
rect 9680 12801 9689 12835
rect 9689 12801 9723 12835
rect 9723 12801 9732 12835
rect 9680 12792 9732 12801
rect 10692 12792 10744 12844
rect 11428 12792 11480 12844
rect 12532 12835 12584 12844
rect 12532 12801 12541 12835
rect 12541 12801 12575 12835
rect 12575 12801 12584 12835
rect 12532 12792 12584 12801
rect 13360 12835 13412 12844
rect 13360 12801 13394 12835
rect 13394 12801 13412 12835
rect 13360 12792 13412 12801
rect 16120 12835 16172 12844
rect 4620 12656 4672 12708
rect 6552 12656 6604 12708
rect 2688 12588 2740 12640
rect 7472 12588 7524 12640
rect 8392 12588 8444 12640
rect 10048 12656 10100 12708
rect 16120 12801 16129 12835
rect 16129 12801 16163 12835
rect 16163 12801 16172 12835
rect 16120 12792 16172 12801
rect 16212 12792 16264 12844
rect 18880 12860 18932 12912
rect 22192 12903 22244 12912
rect 22192 12869 22201 12903
rect 22201 12869 22235 12903
rect 22235 12869 22244 12903
rect 22192 12860 22244 12869
rect 25412 12928 25464 12980
rect 25780 12928 25832 12980
rect 26148 12928 26200 12980
rect 34704 12928 34756 12980
rect 23480 12903 23532 12912
rect 23480 12869 23489 12903
rect 23489 12869 23523 12903
rect 23523 12869 23532 12903
rect 23480 12860 23532 12869
rect 17132 12792 17184 12844
rect 19340 12792 19392 12844
rect 20904 12792 20956 12844
rect 12256 12588 12308 12640
rect 14464 12631 14516 12640
rect 14464 12597 14473 12631
rect 14473 12597 14507 12631
rect 14507 12597 14516 12631
rect 14464 12588 14516 12597
rect 14924 12588 14976 12640
rect 15936 12631 15988 12640
rect 15936 12597 15945 12631
rect 15945 12597 15979 12631
rect 15979 12597 15988 12631
rect 15936 12588 15988 12597
rect 25964 12860 26016 12912
rect 27528 12860 27580 12912
rect 29368 12860 29420 12912
rect 30932 12903 30984 12912
rect 30932 12869 30941 12903
rect 30941 12869 30975 12903
rect 30975 12869 30984 12903
rect 30932 12860 30984 12869
rect 23756 12792 23808 12844
rect 24032 12792 24084 12844
rect 24124 12767 24176 12776
rect 24124 12733 24133 12767
rect 24133 12733 24167 12767
rect 24167 12733 24176 12767
rect 24124 12724 24176 12733
rect 26240 12792 26292 12844
rect 26424 12792 26476 12844
rect 27988 12835 28040 12844
rect 26516 12724 26568 12776
rect 27068 12767 27120 12776
rect 27068 12733 27077 12767
rect 27077 12733 27111 12767
rect 27111 12733 27120 12767
rect 27068 12724 27120 12733
rect 27988 12801 27997 12835
rect 27997 12801 28031 12835
rect 28031 12801 28040 12835
rect 27988 12792 28040 12801
rect 28356 12792 28408 12844
rect 28632 12792 28684 12844
rect 29184 12792 29236 12844
rect 29460 12792 29512 12844
rect 30656 12835 30708 12844
rect 30656 12801 30665 12835
rect 30665 12801 30699 12835
rect 30699 12801 30708 12835
rect 30656 12792 30708 12801
rect 30748 12835 30800 12844
rect 30748 12801 30758 12835
rect 30758 12801 30792 12835
rect 30792 12801 30800 12835
rect 30748 12792 30800 12801
rect 31116 12835 31168 12844
rect 31116 12801 31130 12835
rect 31130 12801 31164 12835
rect 31164 12801 31168 12835
rect 33324 12835 33376 12844
rect 31116 12792 31168 12801
rect 33324 12801 33333 12835
rect 33333 12801 33367 12835
rect 33367 12801 33376 12835
rect 33324 12792 33376 12801
rect 29644 12724 29696 12776
rect 23940 12656 23992 12708
rect 33508 12835 33560 12844
rect 33508 12801 33517 12835
rect 33517 12801 33551 12835
rect 33551 12801 33560 12835
rect 34152 12835 34204 12844
rect 33508 12792 33560 12801
rect 34152 12801 34161 12835
rect 34161 12801 34195 12835
rect 34195 12801 34204 12835
rect 34152 12792 34204 12801
rect 35256 12860 35308 12912
rect 35900 12860 35952 12912
rect 37832 12928 37884 12980
rect 38016 12928 38068 12980
rect 41696 12928 41748 12980
rect 34612 12792 34664 12844
rect 36728 12835 36780 12844
rect 36728 12801 36737 12835
rect 36737 12801 36771 12835
rect 36771 12801 36780 12835
rect 36728 12792 36780 12801
rect 37648 12792 37700 12844
rect 37832 12792 37884 12844
rect 41236 12835 41288 12844
rect 41236 12801 41245 12835
rect 41245 12801 41279 12835
rect 41279 12801 41288 12835
rect 41236 12792 41288 12801
rect 36084 12724 36136 12776
rect 67640 12699 67692 12708
rect 67640 12665 67649 12699
rect 67649 12665 67683 12699
rect 67683 12665 67692 12699
rect 67640 12656 67692 12665
rect 19432 12588 19484 12640
rect 20720 12588 20772 12640
rect 22008 12631 22060 12640
rect 22008 12597 22017 12631
rect 22017 12597 22051 12631
rect 22051 12597 22060 12631
rect 22008 12588 22060 12597
rect 24492 12588 24544 12640
rect 25964 12588 26016 12640
rect 27344 12588 27396 12640
rect 29460 12588 29512 12640
rect 29736 12588 29788 12640
rect 31300 12631 31352 12640
rect 31300 12597 31309 12631
rect 31309 12597 31343 12631
rect 31343 12597 31352 12631
rect 31300 12588 31352 12597
rect 34796 12631 34848 12640
rect 34796 12597 34805 12631
rect 34805 12597 34839 12631
rect 34839 12597 34848 12631
rect 34796 12588 34848 12597
rect 37372 12588 37424 12640
rect 38384 12631 38436 12640
rect 38384 12597 38393 12631
rect 38393 12597 38427 12631
rect 38427 12597 38436 12631
rect 38384 12588 38436 12597
rect 38660 12588 38712 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 65654 12486 65706 12538
rect 65718 12486 65770 12538
rect 65782 12486 65834 12538
rect 65846 12486 65898 12538
rect 65910 12486 65962 12538
rect 3148 12427 3200 12436
rect 3148 12393 3157 12427
rect 3157 12393 3191 12427
rect 3191 12393 3200 12427
rect 3148 12384 3200 12393
rect 3700 12384 3752 12436
rect 6368 12384 6420 12436
rect 7104 12384 7156 12436
rect 13268 12427 13320 12436
rect 13268 12393 13277 12427
rect 13277 12393 13311 12427
rect 13311 12393 13320 12427
rect 13268 12384 13320 12393
rect 16672 12384 16724 12436
rect 17776 12427 17828 12436
rect 17776 12393 17785 12427
rect 17785 12393 17819 12427
rect 17819 12393 17828 12427
rect 17776 12384 17828 12393
rect 20812 12384 20864 12436
rect 20996 12384 21048 12436
rect 2504 12223 2556 12232
rect 2504 12189 2513 12223
rect 2513 12189 2547 12223
rect 2547 12189 2556 12223
rect 2504 12180 2556 12189
rect 2688 12223 2740 12232
rect 2688 12189 2697 12223
rect 2697 12189 2731 12223
rect 2731 12189 2740 12223
rect 2688 12180 2740 12189
rect 3056 12248 3108 12300
rect 5816 12316 5868 12368
rect 6828 12316 6880 12368
rect 7656 12316 7708 12368
rect 8392 12316 8444 12368
rect 24676 12384 24728 12436
rect 25136 12384 25188 12436
rect 25872 12384 25924 12436
rect 26516 12427 26568 12436
rect 26516 12393 26525 12427
rect 26525 12393 26559 12427
rect 26559 12393 26568 12427
rect 26516 12384 26568 12393
rect 26884 12384 26936 12436
rect 3700 12180 3752 12232
rect 3792 12180 3844 12232
rect 6368 12180 6420 12232
rect 6920 12248 6972 12300
rect 3148 12044 3200 12096
rect 5724 12087 5776 12096
rect 5724 12053 5733 12087
rect 5733 12053 5767 12087
rect 5767 12053 5776 12087
rect 5724 12044 5776 12053
rect 6736 12180 6788 12232
rect 6828 12223 6880 12232
rect 6828 12189 6837 12223
rect 6837 12189 6871 12223
rect 6871 12189 6880 12223
rect 6828 12180 6880 12189
rect 7472 12223 7524 12232
rect 7472 12189 7481 12223
rect 7481 12189 7515 12223
rect 7515 12189 7524 12223
rect 7472 12180 7524 12189
rect 17132 12248 17184 12300
rect 7656 12223 7708 12232
rect 7656 12189 7665 12223
rect 7665 12189 7699 12223
rect 7699 12189 7708 12223
rect 9864 12223 9916 12232
rect 7656 12180 7708 12189
rect 9864 12189 9873 12223
rect 9873 12189 9907 12223
rect 9907 12189 9916 12223
rect 9864 12180 9916 12189
rect 10048 12223 10100 12232
rect 10048 12189 10057 12223
rect 10057 12189 10091 12223
rect 10091 12189 10100 12223
rect 10048 12180 10100 12189
rect 10324 12180 10376 12232
rect 11336 12180 11388 12232
rect 11704 12223 11756 12232
rect 11704 12189 11713 12223
rect 11713 12189 11747 12223
rect 11747 12189 11756 12223
rect 11704 12180 11756 12189
rect 10140 12155 10192 12164
rect 10140 12121 10149 12155
rect 10149 12121 10183 12155
rect 10183 12121 10192 12155
rect 10140 12112 10192 12121
rect 11060 12155 11112 12164
rect 11060 12121 11069 12155
rect 11069 12121 11103 12155
rect 11103 12121 11112 12155
rect 11060 12112 11112 12121
rect 12072 12223 12124 12232
rect 12072 12189 12081 12223
rect 12081 12189 12115 12223
rect 12115 12189 12124 12223
rect 12072 12180 12124 12189
rect 12256 12112 12308 12164
rect 13820 12180 13872 12232
rect 14464 12180 14516 12232
rect 14740 12180 14792 12232
rect 14924 12223 14976 12232
rect 14924 12189 14933 12223
rect 14933 12189 14967 12223
rect 14967 12189 14976 12223
rect 14924 12180 14976 12189
rect 15108 12180 15160 12232
rect 15476 12223 15528 12232
rect 15476 12189 15485 12223
rect 15485 12189 15519 12223
rect 15519 12189 15528 12223
rect 15660 12223 15712 12232
rect 15476 12180 15528 12189
rect 15660 12189 15669 12223
rect 15669 12189 15703 12223
rect 15703 12189 15712 12223
rect 15660 12180 15712 12189
rect 15752 12223 15804 12232
rect 15752 12189 15761 12223
rect 15761 12189 15795 12223
rect 15795 12189 15804 12223
rect 15752 12180 15804 12189
rect 16764 12180 16816 12232
rect 17684 12223 17736 12232
rect 17684 12189 17693 12223
rect 17693 12189 17727 12223
rect 17727 12189 17736 12223
rect 19432 12248 19484 12300
rect 19984 12248 20036 12300
rect 22928 12248 22980 12300
rect 23480 12248 23532 12300
rect 17684 12180 17736 12189
rect 20260 12180 20312 12232
rect 22192 12180 22244 12232
rect 24584 12316 24636 12368
rect 24768 12316 24820 12368
rect 25412 12359 25464 12368
rect 25412 12325 25421 12359
rect 25421 12325 25455 12359
rect 25455 12325 25464 12359
rect 25412 12316 25464 12325
rect 26608 12316 26660 12368
rect 26240 12248 26292 12300
rect 27988 12316 28040 12368
rect 7196 12044 7248 12096
rect 8024 12044 8076 12096
rect 8300 12044 8352 12096
rect 9956 12044 10008 12096
rect 12808 12087 12860 12096
rect 12808 12053 12817 12087
rect 12817 12053 12851 12087
rect 12851 12053 12860 12087
rect 12808 12044 12860 12053
rect 13636 12112 13688 12164
rect 14556 12112 14608 12164
rect 20996 12112 21048 12164
rect 22100 12155 22152 12164
rect 22100 12121 22109 12155
rect 22109 12121 22143 12155
rect 22143 12121 22152 12155
rect 22100 12112 22152 12121
rect 24584 12223 24636 12232
rect 24584 12189 24593 12223
rect 24593 12189 24627 12223
rect 24627 12189 24636 12223
rect 24584 12180 24636 12189
rect 25136 12180 25188 12232
rect 25688 12223 25740 12232
rect 25688 12189 25697 12223
rect 25697 12189 25731 12223
rect 25731 12189 25740 12223
rect 25688 12180 25740 12189
rect 26056 12180 26108 12232
rect 29460 12248 29512 12300
rect 29828 12248 29880 12300
rect 31392 12384 31444 12436
rect 36084 12427 36136 12436
rect 31116 12316 31168 12368
rect 29644 12223 29696 12232
rect 14832 12044 14884 12096
rect 15752 12044 15804 12096
rect 16672 12044 16724 12096
rect 17868 12044 17920 12096
rect 20444 12044 20496 12096
rect 20720 12044 20772 12096
rect 22928 12044 22980 12096
rect 24400 12087 24452 12096
rect 24400 12053 24409 12087
rect 24409 12053 24443 12087
rect 24443 12053 24452 12087
rect 24400 12044 24452 12053
rect 25412 12112 25464 12164
rect 25872 12112 25924 12164
rect 27988 12112 28040 12164
rect 28632 12155 28684 12164
rect 28632 12121 28641 12155
rect 28641 12121 28675 12155
rect 28675 12121 28684 12155
rect 28632 12112 28684 12121
rect 29644 12189 29653 12223
rect 29653 12189 29687 12223
rect 29687 12189 29696 12223
rect 29644 12180 29696 12189
rect 29920 12223 29972 12232
rect 29920 12189 29929 12223
rect 29929 12189 29963 12223
rect 29963 12189 29972 12223
rect 29920 12180 29972 12189
rect 30932 12248 30984 12300
rect 32496 12248 32548 12300
rect 30196 12180 30248 12232
rect 31300 12223 31352 12232
rect 31300 12189 31309 12223
rect 31309 12189 31343 12223
rect 31343 12189 31352 12223
rect 31300 12180 31352 12189
rect 31392 12180 31444 12232
rect 32128 12180 32180 12232
rect 32680 12180 32732 12232
rect 33600 12248 33652 12300
rect 36084 12393 36093 12427
rect 36093 12393 36127 12427
rect 36127 12393 36136 12427
rect 36084 12384 36136 12393
rect 41236 12427 41288 12436
rect 41236 12393 41245 12427
rect 41245 12393 41279 12427
rect 41279 12393 41288 12427
rect 41236 12384 41288 12393
rect 35348 12180 35400 12232
rect 35808 12180 35860 12232
rect 36820 12223 36872 12232
rect 36820 12189 36829 12223
rect 36829 12189 36863 12223
rect 36863 12189 36872 12223
rect 36820 12180 36872 12189
rect 29552 12112 29604 12164
rect 28724 12087 28776 12096
rect 28724 12053 28733 12087
rect 28733 12053 28767 12087
rect 28767 12053 28776 12087
rect 28724 12044 28776 12053
rect 29000 12044 29052 12096
rect 31576 12155 31628 12164
rect 31576 12121 31585 12155
rect 31585 12121 31619 12155
rect 31619 12121 31628 12155
rect 32404 12155 32456 12164
rect 31576 12112 31628 12121
rect 32404 12121 32413 12155
rect 32413 12121 32447 12155
rect 32447 12121 32456 12155
rect 32404 12112 32456 12121
rect 33508 12112 33560 12164
rect 33876 12112 33928 12164
rect 34796 12112 34848 12164
rect 37004 12223 37056 12232
rect 37004 12189 37013 12223
rect 37013 12189 37047 12223
rect 37047 12189 37056 12223
rect 37004 12180 37056 12189
rect 37556 12180 37608 12232
rect 38660 12248 38712 12300
rect 37924 12112 37976 12164
rect 38384 12180 38436 12232
rect 39028 12180 39080 12232
rect 39856 12223 39908 12232
rect 39856 12189 39865 12223
rect 39865 12189 39899 12223
rect 39899 12189 39908 12223
rect 39856 12180 39908 12189
rect 30380 12044 30432 12096
rect 32220 12044 32272 12096
rect 37280 12087 37332 12096
rect 37280 12053 37289 12087
rect 37289 12053 37323 12087
rect 37323 12053 37332 12087
rect 37280 12044 37332 12053
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 50294 11942 50346 11994
rect 50358 11942 50410 11994
rect 50422 11942 50474 11994
rect 50486 11942 50538 11994
rect 50550 11942 50602 11994
rect 2136 11840 2188 11892
rect 2412 11840 2464 11892
rect 4620 11840 4672 11892
rect 6736 11883 6788 11892
rect 6736 11849 6745 11883
rect 6745 11849 6779 11883
rect 6779 11849 6788 11883
rect 6736 11840 6788 11849
rect 7196 11883 7248 11892
rect 7196 11849 7205 11883
rect 7205 11849 7239 11883
rect 7239 11849 7248 11883
rect 7196 11840 7248 11849
rect 1952 11772 2004 11824
rect 2044 11747 2096 11756
rect 2044 11713 2053 11747
rect 2053 11713 2087 11747
rect 2087 11713 2096 11747
rect 2044 11704 2096 11713
rect 5724 11772 5776 11824
rect 8484 11772 8536 11824
rect 5816 11704 5868 11756
rect 6000 11704 6052 11756
rect 8024 11747 8076 11756
rect 8024 11713 8058 11747
rect 8058 11713 8076 11747
rect 8024 11704 8076 11713
rect 2504 11636 2556 11688
rect 7104 11636 7156 11688
rect 3240 11568 3292 11620
rect 8944 11840 8996 11892
rect 17132 11840 17184 11892
rect 18788 11883 18840 11892
rect 18788 11849 18797 11883
rect 18797 11849 18831 11883
rect 18831 11849 18840 11883
rect 18788 11840 18840 11849
rect 23296 11883 23348 11892
rect 23296 11849 23305 11883
rect 23305 11849 23339 11883
rect 23339 11849 23348 11883
rect 23296 11840 23348 11849
rect 10048 11772 10100 11824
rect 11336 11704 11388 11756
rect 13176 11772 13228 11824
rect 16212 11772 16264 11824
rect 15200 11704 15252 11756
rect 15752 11747 15804 11756
rect 15752 11713 15761 11747
rect 15761 11713 15795 11747
rect 15795 11713 15804 11747
rect 15752 11704 15804 11713
rect 16304 11704 16356 11756
rect 23204 11772 23256 11824
rect 25504 11840 25556 11892
rect 23940 11772 23992 11824
rect 24124 11772 24176 11824
rect 24768 11772 24820 11824
rect 25136 11815 25188 11824
rect 25136 11781 25145 11815
rect 25145 11781 25179 11815
rect 25179 11781 25188 11815
rect 25136 11772 25188 11781
rect 25412 11772 25464 11824
rect 29000 11840 29052 11892
rect 29460 11840 29512 11892
rect 29644 11840 29696 11892
rect 33048 11840 33100 11892
rect 34520 11840 34572 11892
rect 35624 11840 35676 11892
rect 17132 11704 17184 11756
rect 15292 11636 15344 11688
rect 18512 11704 18564 11756
rect 20076 11704 20128 11756
rect 18236 11636 18288 11688
rect 11520 11568 11572 11620
rect 17040 11568 17092 11620
rect 17408 11568 17460 11620
rect 19248 11568 19300 11620
rect 2504 11500 2556 11552
rect 6000 11500 6052 11552
rect 10876 11500 10928 11552
rect 11060 11500 11112 11552
rect 12072 11500 12124 11552
rect 12624 11500 12676 11552
rect 15936 11500 15988 11552
rect 16580 11500 16632 11552
rect 18972 11543 19024 11552
rect 18972 11509 18981 11543
rect 18981 11509 19015 11543
rect 19015 11509 19024 11543
rect 18972 11500 19024 11509
rect 19524 11500 19576 11552
rect 20076 11500 20128 11552
rect 20536 11747 20588 11756
rect 20536 11713 20545 11747
rect 20545 11713 20579 11747
rect 20579 11713 20588 11747
rect 20536 11704 20588 11713
rect 22376 11747 22428 11756
rect 20260 11636 20312 11688
rect 20996 11636 21048 11688
rect 22376 11713 22385 11747
rect 22385 11713 22419 11747
rect 22419 11713 22428 11747
rect 22376 11704 22428 11713
rect 22284 11568 22336 11620
rect 20720 11500 20772 11552
rect 22928 11704 22980 11756
rect 23480 11747 23532 11756
rect 23480 11713 23489 11747
rect 23489 11713 23523 11747
rect 23523 11713 23532 11747
rect 23480 11704 23532 11713
rect 24584 11747 24636 11756
rect 24584 11713 24593 11747
rect 24593 11713 24627 11747
rect 24627 11713 24636 11747
rect 29276 11772 29328 11824
rect 35348 11772 35400 11824
rect 35808 11772 35860 11824
rect 24584 11704 24636 11713
rect 26240 11747 26292 11756
rect 26240 11713 26249 11747
rect 26249 11713 26283 11747
rect 26283 11713 26292 11747
rect 26240 11704 26292 11713
rect 26424 11704 26476 11756
rect 27436 11704 27488 11756
rect 23756 11568 23808 11620
rect 23940 11568 23992 11620
rect 25412 11568 25464 11620
rect 26700 11636 26752 11688
rect 26792 11636 26844 11688
rect 27712 11747 27764 11756
rect 27712 11713 27721 11747
rect 27721 11713 27755 11747
rect 27755 11713 27764 11747
rect 27712 11704 27764 11713
rect 29828 11704 29880 11756
rect 30196 11747 30248 11756
rect 30196 11713 30241 11747
rect 30241 11713 30248 11747
rect 30196 11704 30248 11713
rect 30380 11747 30432 11756
rect 30380 11713 30389 11747
rect 30389 11713 30423 11747
rect 30423 11713 30432 11747
rect 30380 11704 30432 11713
rect 32864 11704 32916 11756
rect 33600 11747 33652 11756
rect 33600 11713 33609 11747
rect 33609 11713 33643 11747
rect 33643 11713 33652 11747
rect 33600 11704 33652 11713
rect 34796 11704 34848 11756
rect 37556 11747 37608 11756
rect 34520 11679 34572 11688
rect 34520 11645 34529 11679
rect 34529 11645 34563 11679
rect 34563 11645 34572 11679
rect 37556 11713 37565 11747
rect 37565 11713 37599 11747
rect 37599 11713 37608 11747
rect 37556 11704 37608 11713
rect 34520 11636 34572 11645
rect 27712 11500 27764 11552
rect 27804 11500 27856 11552
rect 28080 11500 28132 11552
rect 28632 11500 28684 11552
rect 29736 11543 29788 11552
rect 29736 11509 29745 11543
rect 29745 11509 29779 11543
rect 29779 11509 29788 11543
rect 29736 11500 29788 11509
rect 30012 11500 30064 11552
rect 30196 11500 30248 11552
rect 32864 11543 32916 11552
rect 32864 11509 32873 11543
rect 32873 11509 32907 11543
rect 32907 11509 32916 11543
rect 32864 11500 32916 11509
rect 36636 11568 36688 11620
rect 36912 11500 36964 11552
rect 37832 11500 37884 11552
rect 67640 11543 67692 11552
rect 67640 11509 67649 11543
rect 67649 11509 67683 11543
rect 67683 11509 67692 11543
rect 67640 11500 67692 11509
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 65654 11398 65706 11450
rect 65718 11398 65770 11450
rect 65782 11398 65834 11450
rect 65846 11398 65898 11450
rect 65910 11398 65962 11450
rect 9956 11296 10008 11348
rect 13360 11296 13412 11348
rect 13544 11296 13596 11348
rect 15108 11339 15160 11348
rect 15108 11305 15117 11339
rect 15117 11305 15151 11339
rect 15151 11305 15160 11339
rect 15108 11296 15160 11305
rect 15568 11296 15620 11348
rect 18420 11296 18472 11348
rect 20168 11296 20220 11348
rect 22100 11296 22152 11348
rect 22376 11339 22428 11348
rect 22376 11305 22385 11339
rect 22385 11305 22419 11339
rect 22419 11305 22428 11339
rect 22376 11296 22428 11305
rect 23756 11339 23808 11348
rect 23756 11305 23765 11339
rect 23765 11305 23799 11339
rect 23799 11305 23808 11339
rect 23756 11296 23808 11305
rect 24676 11296 24728 11348
rect 28724 11296 28776 11348
rect 3148 11092 3200 11144
rect 3792 11135 3844 11144
rect 3792 11101 3801 11135
rect 3801 11101 3835 11135
rect 3835 11101 3844 11135
rect 3792 11092 3844 11101
rect 11428 11228 11480 11280
rect 11612 11228 11664 11280
rect 14740 11228 14792 11280
rect 14832 11228 14884 11280
rect 6092 11160 6144 11212
rect 7104 11160 7156 11212
rect 16488 11160 16540 11212
rect 17316 11160 17368 11212
rect 17684 11228 17736 11280
rect 29828 11271 29880 11280
rect 29828 11237 29837 11271
rect 29837 11237 29871 11271
rect 29871 11237 29880 11271
rect 29828 11228 29880 11237
rect 32864 11271 32916 11280
rect 9772 11092 9824 11144
rect 11612 11092 11664 11144
rect 11888 11092 11940 11144
rect 5080 11024 5132 11076
rect 6000 11067 6052 11076
rect 6000 11033 6009 11067
rect 6009 11033 6043 11067
rect 6043 11033 6052 11067
rect 6000 11024 6052 11033
rect 6644 11067 6696 11076
rect 6644 11033 6653 11067
rect 6653 11033 6687 11067
rect 6687 11033 6696 11067
rect 6644 11024 6696 11033
rect 8300 11067 8352 11076
rect 2504 10956 2556 11008
rect 5632 10999 5684 11008
rect 5632 10965 5641 10999
rect 5641 10965 5675 10999
rect 5675 10965 5684 10999
rect 5632 10956 5684 10965
rect 8300 11033 8309 11067
rect 8309 11033 8343 11067
rect 8343 11033 8352 11067
rect 8300 11024 8352 11033
rect 10232 11024 10284 11076
rect 10508 11024 10560 11076
rect 11336 11067 11388 11076
rect 11336 11033 11345 11067
rect 11345 11033 11379 11067
rect 11379 11033 11388 11067
rect 11336 11024 11388 11033
rect 11520 11067 11572 11076
rect 11520 11033 11529 11067
rect 11529 11033 11563 11067
rect 11563 11033 11572 11067
rect 11520 11024 11572 11033
rect 7748 10956 7800 11008
rect 8944 10956 8996 11008
rect 12440 11135 12492 11144
rect 12440 11101 12449 11135
rect 12449 11101 12483 11135
rect 12483 11101 12492 11135
rect 12440 11092 12492 11101
rect 13820 11092 13872 11144
rect 13544 11024 13596 11076
rect 14648 11024 14700 11076
rect 15476 11135 15528 11144
rect 15476 11101 15485 11135
rect 15485 11101 15519 11135
rect 15519 11101 15528 11135
rect 15476 11092 15528 11101
rect 16304 11067 16356 11076
rect 16304 11033 16313 11067
rect 16313 11033 16347 11067
rect 16347 11033 16356 11067
rect 16304 11024 16356 11033
rect 16764 11135 16816 11144
rect 16764 11101 16773 11135
rect 16773 11101 16807 11135
rect 16807 11101 16816 11135
rect 17040 11135 17092 11144
rect 16764 11092 16816 11101
rect 17040 11101 17049 11135
rect 17049 11101 17083 11135
rect 17083 11101 17092 11135
rect 17040 11092 17092 11101
rect 18328 11160 18380 11212
rect 19432 11160 19484 11212
rect 20536 11160 20588 11212
rect 20812 11160 20864 11212
rect 23940 11160 23992 11212
rect 27988 11160 28040 11212
rect 28172 11203 28224 11212
rect 28172 11169 28181 11203
rect 28181 11169 28215 11203
rect 28215 11169 28224 11203
rect 28172 11160 28224 11169
rect 28632 11160 28684 11212
rect 30472 11160 30524 11212
rect 32864 11237 32873 11271
rect 32873 11237 32907 11271
rect 32907 11237 32916 11271
rect 32864 11228 32916 11237
rect 18236 11135 18288 11144
rect 18236 11101 18245 11135
rect 18245 11101 18279 11135
rect 18279 11101 18288 11135
rect 18236 11092 18288 11101
rect 20076 11135 20128 11144
rect 18328 11024 18380 11076
rect 18604 11024 18656 11076
rect 20076 11101 20085 11135
rect 20085 11101 20119 11135
rect 20119 11101 20128 11135
rect 20076 11092 20128 11101
rect 22192 11135 22244 11144
rect 20260 11024 20312 11076
rect 20812 11024 20864 11076
rect 22192 11101 22201 11135
rect 22201 11101 22235 11135
rect 22235 11101 22244 11135
rect 22192 11092 22244 11101
rect 23848 11092 23900 11144
rect 24768 11135 24820 11144
rect 22560 11024 22612 11076
rect 16948 10999 17000 11008
rect 16948 10965 16957 10999
rect 16957 10965 16991 10999
rect 16991 10965 17000 10999
rect 16948 10956 17000 10965
rect 24768 11101 24777 11135
rect 24777 11101 24811 11135
rect 24811 11101 24820 11135
rect 24768 11092 24820 11101
rect 24952 11135 25004 11144
rect 24952 11101 24961 11135
rect 24961 11101 24995 11135
rect 24995 11101 25004 11135
rect 24952 11092 25004 11101
rect 25044 11092 25096 11144
rect 26056 11092 26108 11144
rect 27160 11092 27212 11144
rect 30196 11092 30248 11144
rect 32220 11135 32272 11144
rect 32220 11101 32229 11135
rect 32229 11101 32263 11135
rect 32263 11101 32272 11135
rect 32220 11092 32272 11101
rect 32496 11135 32548 11144
rect 32496 11101 32505 11135
rect 32505 11101 32539 11135
rect 32539 11101 32548 11135
rect 32496 11092 32548 11101
rect 33600 11160 33652 11212
rect 33232 11092 33284 11144
rect 33968 11092 34020 11144
rect 36820 11296 36872 11348
rect 36084 11228 36136 11280
rect 40408 11296 40460 11348
rect 34428 11160 34480 11212
rect 34980 11135 35032 11144
rect 34980 11101 34989 11135
rect 34989 11101 35023 11135
rect 35023 11101 35032 11135
rect 34980 11092 35032 11101
rect 25136 11024 25188 11076
rect 25964 11067 26016 11076
rect 25964 11033 25973 11067
rect 25973 11033 26007 11067
rect 26007 11033 26016 11067
rect 25964 11024 26016 11033
rect 26240 11024 26292 11076
rect 26884 11024 26936 11076
rect 27528 11024 27580 11076
rect 33416 11067 33468 11076
rect 29184 10956 29236 11008
rect 29368 10956 29420 11008
rect 29920 10956 29972 11008
rect 33416 11033 33425 11067
rect 33425 11033 33459 11067
rect 33459 11033 33468 11067
rect 33416 11024 33468 11033
rect 34612 11024 34664 11076
rect 35164 11135 35216 11144
rect 35164 11101 35173 11135
rect 35173 11101 35207 11135
rect 35207 11101 35216 11135
rect 37372 11160 37424 11212
rect 35164 11092 35216 11101
rect 35808 11092 35860 11144
rect 39028 11092 39080 11144
rect 35440 11024 35492 11076
rect 36084 11067 36136 11076
rect 36084 11033 36093 11067
rect 36093 11033 36127 11067
rect 36127 11033 36136 11067
rect 36084 11024 36136 11033
rect 36360 11024 36412 11076
rect 36912 11067 36964 11076
rect 36912 11033 36921 11067
rect 36921 11033 36955 11067
rect 36955 11033 36964 11067
rect 36912 11024 36964 11033
rect 34704 10999 34756 11008
rect 34704 10965 34713 10999
rect 34713 10965 34747 10999
rect 34747 10965 34756 10999
rect 34704 10956 34756 10965
rect 37280 11024 37332 11076
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 50294 10854 50346 10906
rect 50358 10854 50410 10906
rect 50422 10854 50474 10906
rect 50486 10854 50538 10906
rect 50550 10854 50602 10906
rect 1492 10752 1544 10804
rect 5080 10752 5132 10804
rect 6828 10752 6880 10804
rect 9864 10752 9916 10804
rect 10232 10795 10284 10804
rect 10232 10761 10241 10795
rect 10241 10761 10275 10795
rect 10275 10761 10284 10795
rect 10232 10752 10284 10761
rect 2504 10616 2556 10668
rect 4712 10659 4764 10668
rect 4712 10625 4721 10659
rect 4721 10625 4755 10659
rect 4755 10625 4764 10659
rect 4712 10616 4764 10625
rect 5540 10659 5592 10668
rect 5540 10625 5549 10659
rect 5549 10625 5583 10659
rect 5583 10625 5592 10659
rect 5540 10616 5592 10625
rect 5632 10659 5684 10668
rect 5632 10625 5641 10659
rect 5641 10625 5675 10659
rect 5675 10625 5684 10659
rect 5632 10616 5684 10625
rect 5908 10616 5960 10668
rect 6828 10616 6880 10668
rect 7104 10659 7156 10668
rect 7104 10625 7113 10659
rect 7113 10625 7147 10659
rect 7147 10625 7156 10659
rect 7104 10616 7156 10625
rect 7380 10659 7432 10668
rect 7380 10625 7414 10659
rect 7414 10625 7432 10659
rect 7380 10616 7432 10625
rect 8484 10616 8536 10668
rect 8852 10616 8904 10668
rect 9496 10616 9548 10668
rect 11704 10684 11756 10736
rect 11796 10684 11848 10736
rect 9680 10616 9732 10668
rect 1952 10548 2004 10600
rect 9956 10659 10008 10668
rect 9956 10625 9965 10659
rect 9965 10625 9999 10659
rect 9999 10625 10008 10659
rect 10784 10659 10836 10668
rect 9956 10616 10008 10625
rect 10784 10625 10793 10659
rect 10793 10625 10827 10659
rect 10827 10625 10836 10659
rect 10784 10616 10836 10625
rect 11152 10616 11204 10668
rect 11888 10659 11940 10668
rect 11888 10625 11897 10659
rect 11897 10625 11931 10659
rect 11931 10625 11940 10659
rect 11888 10616 11940 10625
rect 12072 10659 12124 10668
rect 12072 10625 12081 10659
rect 12081 10625 12115 10659
rect 12115 10625 12124 10659
rect 12072 10616 12124 10625
rect 12348 10684 12400 10736
rect 12256 10659 12308 10668
rect 12256 10625 12265 10659
rect 12265 10625 12299 10659
rect 12299 10625 12308 10659
rect 16948 10752 17000 10804
rect 17316 10752 17368 10804
rect 22192 10752 22244 10804
rect 25964 10752 26016 10804
rect 26056 10752 26108 10804
rect 27436 10795 27488 10804
rect 27436 10761 27445 10795
rect 27445 10761 27479 10795
rect 27479 10761 27488 10795
rect 27436 10752 27488 10761
rect 28356 10752 28408 10804
rect 27712 10684 27764 10736
rect 28908 10684 28960 10736
rect 13176 10659 13228 10668
rect 12256 10616 12308 10625
rect 13176 10625 13185 10659
rect 13185 10625 13219 10659
rect 13219 10625 13228 10659
rect 13176 10616 13228 10625
rect 18512 10616 18564 10668
rect 22284 10616 22336 10668
rect 25320 10616 25372 10668
rect 25596 10616 25648 10668
rect 11612 10548 11664 10600
rect 18328 10548 18380 10600
rect 20536 10548 20588 10600
rect 23388 10548 23440 10600
rect 26240 10659 26292 10668
rect 26240 10625 26249 10659
rect 26249 10625 26283 10659
rect 26283 10625 26292 10659
rect 26240 10616 26292 10625
rect 26424 10659 26476 10668
rect 26424 10625 26433 10659
rect 26433 10625 26467 10659
rect 26467 10625 26476 10659
rect 26424 10616 26476 10625
rect 27988 10616 28040 10668
rect 30104 10684 30156 10736
rect 29368 10659 29420 10668
rect 9956 10480 10008 10532
rect 2504 10455 2556 10464
rect 2504 10421 2513 10455
rect 2513 10421 2547 10455
rect 2547 10421 2556 10455
rect 2504 10412 2556 10421
rect 5448 10412 5500 10464
rect 7288 10412 7340 10464
rect 9128 10412 9180 10464
rect 10876 10412 10928 10464
rect 15200 10455 15252 10464
rect 15200 10421 15209 10455
rect 15209 10421 15243 10455
rect 15243 10421 15252 10455
rect 15200 10412 15252 10421
rect 17316 10412 17368 10464
rect 22652 10412 22704 10464
rect 23020 10412 23072 10464
rect 23296 10412 23348 10464
rect 26792 10548 26844 10600
rect 29368 10625 29376 10659
rect 29376 10625 29410 10659
rect 29410 10625 29420 10659
rect 29368 10616 29420 10625
rect 29460 10659 29512 10668
rect 29460 10625 29469 10659
rect 29469 10625 29503 10659
rect 29503 10625 29512 10659
rect 29460 10616 29512 10625
rect 30380 10659 30432 10668
rect 30380 10625 30389 10659
rect 30389 10625 30423 10659
rect 30423 10625 30432 10659
rect 30380 10616 30432 10625
rect 31944 10684 31996 10736
rect 31484 10659 31536 10668
rect 31484 10625 31493 10659
rect 31493 10625 31527 10659
rect 31527 10625 31536 10659
rect 33048 10752 33100 10804
rect 33140 10684 33192 10736
rect 35164 10752 35216 10804
rect 40408 10795 40460 10804
rect 40408 10761 40417 10795
rect 40417 10761 40451 10795
rect 40451 10761 40460 10795
rect 40408 10752 40460 10761
rect 42432 10752 42484 10804
rect 31484 10616 31536 10625
rect 27160 10480 27212 10532
rect 30840 10523 30892 10532
rect 30840 10489 30849 10523
rect 30849 10489 30883 10523
rect 30883 10489 30892 10523
rect 30840 10480 30892 10489
rect 31760 10548 31812 10600
rect 33600 10616 33652 10668
rect 32128 10523 32180 10532
rect 32128 10489 32137 10523
rect 32137 10489 32171 10523
rect 32171 10489 32180 10523
rect 32128 10480 32180 10489
rect 24216 10412 24268 10464
rect 28080 10455 28132 10464
rect 28080 10421 28089 10455
rect 28089 10421 28123 10455
rect 28123 10421 28132 10455
rect 28080 10412 28132 10421
rect 28816 10455 28868 10464
rect 28816 10421 28825 10455
rect 28825 10421 28859 10455
rect 28859 10421 28868 10455
rect 28816 10412 28868 10421
rect 30288 10455 30340 10464
rect 30288 10421 30297 10455
rect 30297 10421 30331 10455
rect 30331 10421 30340 10455
rect 30288 10412 30340 10421
rect 31116 10412 31168 10464
rect 33784 10548 33836 10600
rect 34704 10684 34756 10736
rect 34796 10616 34848 10668
rect 35900 10616 35952 10668
rect 36636 10616 36688 10668
rect 37188 10616 37240 10668
rect 37924 10616 37976 10668
rect 39028 10659 39080 10668
rect 39028 10625 39037 10659
rect 39037 10625 39071 10659
rect 39071 10625 39080 10659
rect 39028 10616 39080 10625
rect 39120 10616 39172 10668
rect 39856 10616 39908 10668
rect 40960 10591 41012 10600
rect 40960 10557 40969 10591
rect 40969 10557 41003 10591
rect 41003 10557 41012 10591
rect 40960 10548 41012 10557
rect 34244 10412 34296 10464
rect 35348 10412 35400 10464
rect 36360 10412 36412 10464
rect 40868 10455 40920 10464
rect 40868 10421 40877 10455
rect 40877 10421 40911 10455
rect 40911 10421 40920 10455
rect 40868 10412 40920 10421
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 65654 10310 65706 10362
rect 65718 10310 65770 10362
rect 65782 10310 65834 10362
rect 65846 10310 65898 10362
rect 65910 10310 65962 10362
rect 6644 10208 6696 10260
rect 7380 10208 7432 10260
rect 7564 10208 7616 10260
rect 12256 10251 12308 10260
rect 12256 10217 12265 10251
rect 12265 10217 12299 10251
rect 12299 10217 12308 10251
rect 12256 10208 12308 10217
rect 6920 10140 6972 10192
rect 3792 10115 3844 10124
rect 3792 10081 3801 10115
rect 3801 10081 3835 10115
rect 3835 10081 3844 10115
rect 3792 10072 3844 10081
rect 5540 10072 5592 10124
rect 6092 10047 6144 10056
rect 6092 10013 6101 10047
rect 6101 10013 6135 10047
rect 6135 10013 6144 10047
rect 6092 10004 6144 10013
rect 6276 10047 6328 10056
rect 6276 10013 6285 10047
rect 6285 10013 6319 10047
rect 6319 10013 6328 10047
rect 6828 10047 6880 10056
rect 6276 10004 6328 10013
rect 6828 10013 6837 10047
rect 6837 10013 6871 10047
rect 6871 10013 6880 10047
rect 7728 10047 7780 10056
rect 6828 10004 6880 10013
rect 6920 9936 6972 9988
rect 6092 9868 6144 9920
rect 7104 9868 7156 9920
rect 7728 10013 7745 10047
rect 7745 10013 7780 10047
rect 7728 10004 7780 10013
rect 8116 10047 8168 10056
rect 8116 10013 8125 10047
rect 8125 10013 8159 10047
rect 8159 10013 8168 10047
rect 8944 10047 8996 10056
rect 8116 10004 8168 10013
rect 8944 10013 8953 10047
rect 8953 10013 8987 10047
rect 8987 10013 8996 10047
rect 8944 10004 8996 10013
rect 9864 10004 9916 10056
rect 10324 10072 10376 10124
rect 10692 10072 10744 10124
rect 11428 10115 11480 10124
rect 11428 10081 11437 10115
rect 11437 10081 11471 10115
rect 11471 10081 11480 10115
rect 11428 10072 11480 10081
rect 13268 10208 13320 10260
rect 13636 10140 13688 10192
rect 10140 10047 10192 10056
rect 10140 10013 10149 10047
rect 10149 10013 10183 10047
rect 10183 10013 10192 10047
rect 10140 10004 10192 10013
rect 11152 10047 11204 10056
rect 11152 10013 11161 10047
rect 11161 10013 11195 10047
rect 11195 10013 11204 10047
rect 11152 10004 11204 10013
rect 11888 10004 11940 10056
rect 12256 10047 12308 10056
rect 12256 10013 12265 10047
rect 12265 10013 12299 10047
rect 12299 10013 12308 10047
rect 14096 10047 14148 10056
rect 12256 10004 12308 10013
rect 10324 9936 10376 9988
rect 14096 10013 14105 10047
rect 14105 10013 14139 10047
rect 14139 10013 14148 10047
rect 14096 10004 14148 10013
rect 14188 10047 14240 10056
rect 14188 10013 14197 10047
rect 14197 10013 14231 10047
rect 14231 10013 14240 10047
rect 17316 10208 17368 10260
rect 20076 10208 20128 10260
rect 20352 10208 20404 10260
rect 25596 10251 25648 10260
rect 25596 10217 25605 10251
rect 25605 10217 25639 10251
rect 25639 10217 25648 10251
rect 25596 10208 25648 10217
rect 26056 10208 26108 10260
rect 29460 10208 29512 10260
rect 31484 10208 31536 10260
rect 34796 10208 34848 10260
rect 35808 10208 35860 10260
rect 39120 10208 39172 10260
rect 23848 10140 23900 10192
rect 26424 10140 26476 10192
rect 20076 10115 20128 10124
rect 14188 10004 14240 10013
rect 15476 10004 15528 10056
rect 20076 10081 20085 10115
rect 20085 10081 20119 10115
rect 20119 10081 20128 10115
rect 20076 10072 20128 10081
rect 20352 10072 20404 10124
rect 20720 10115 20772 10124
rect 20720 10081 20729 10115
rect 20729 10081 20763 10115
rect 20763 10081 20772 10115
rect 20720 10072 20772 10081
rect 27436 10072 27488 10124
rect 29920 10140 29972 10192
rect 32036 10115 32088 10124
rect 14556 9936 14608 9988
rect 9864 9868 9916 9920
rect 14832 9868 14884 9920
rect 15200 9911 15252 9920
rect 15200 9877 15209 9911
rect 15209 9877 15243 9911
rect 15243 9877 15252 9911
rect 15200 9868 15252 9877
rect 16028 9911 16080 9920
rect 16028 9877 16037 9911
rect 16037 9877 16071 9911
rect 16071 9877 16080 9911
rect 16028 9868 16080 9877
rect 16672 10004 16724 10056
rect 16856 9868 16908 9920
rect 18420 10047 18472 10056
rect 18420 10013 18429 10047
rect 18429 10013 18463 10047
rect 18463 10013 18472 10047
rect 18420 10004 18472 10013
rect 20168 10004 20220 10056
rect 20536 10004 20588 10056
rect 20812 10004 20864 10056
rect 20904 10004 20956 10056
rect 19340 9936 19392 9988
rect 20352 9936 20404 9988
rect 19984 9911 20036 9920
rect 19984 9877 19993 9911
rect 19993 9877 20027 9911
rect 20027 9877 20036 9911
rect 19984 9868 20036 9877
rect 20168 9868 20220 9920
rect 23296 10047 23348 10056
rect 22284 9936 22336 9988
rect 23296 10013 23305 10047
rect 23305 10013 23339 10047
rect 23339 10013 23348 10047
rect 23296 10004 23348 10013
rect 27160 10047 27212 10056
rect 27160 10013 27169 10047
rect 27169 10013 27203 10047
rect 27203 10013 27212 10047
rect 27160 10004 27212 10013
rect 28448 10047 28500 10056
rect 28448 10013 28457 10047
rect 28457 10013 28491 10047
rect 28491 10013 28500 10047
rect 28448 10004 28500 10013
rect 28540 10004 28592 10056
rect 28724 9979 28776 9988
rect 28724 9945 28733 9979
rect 28733 9945 28767 9979
rect 28767 9945 28776 9979
rect 28724 9936 28776 9945
rect 29000 10004 29052 10056
rect 29920 10047 29972 10056
rect 29920 10013 29929 10047
rect 29929 10013 29963 10047
rect 29963 10013 29972 10047
rect 29920 10004 29972 10013
rect 31208 10004 31260 10056
rect 31760 10004 31812 10056
rect 32036 10081 32045 10115
rect 32045 10081 32079 10115
rect 32079 10081 32088 10115
rect 32036 10072 32088 10081
rect 32588 10072 32640 10124
rect 33324 10115 33376 10124
rect 33324 10081 33333 10115
rect 33333 10081 33367 10115
rect 33367 10081 33376 10115
rect 33324 10072 33376 10081
rect 33692 10072 33744 10124
rect 33508 10047 33560 10056
rect 29184 9936 29236 9988
rect 29828 9979 29880 9988
rect 29828 9945 29837 9979
rect 29837 9945 29871 9979
rect 29871 9945 29880 9979
rect 31116 9979 31168 9988
rect 29828 9936 29880 9945
rect 31116 9945 31125 9979
rect 31125 9945 31159 9979
rect 31159 9945 31168 9979
rect 31116 9936 31168 9945
rect 25136 9911 25188 9920
rect 25136 9877 25145 9911
rect 25145 9877 25179 9911
rect 25179 9877 25188 9911
rect 25136 9868 25188 9877
rect 25320 9868 25372 9920
rect 29920 9868 29972 9920
rect 31944 9868 31996 9920
rect 33508 10013 33517 10047
rect 33517 10013 33551 10047
rect 33551 10013 33560 10047
rect 33508 10004 33560 10013
rect 33784 10004 33836 10056
rect 34704 10047 34756 10056
rect 34704 10013 34713 10047
rect 34713 10013 34747 10047
rect 34747 10013 34756 10047
rect 34704 10004 34756 10013
rect 37556 10072 37608 10124
rect 37280 10047 37332 10056
rect 37280 10013 37289 10047
rect 37289 10013 37323 10047
rect 37323 10013 37332 10047
rect 37280 10004 37332 10013
rect 68100 10047 68152 10056
rect 34796 9936 34848 9988
rect 37188 9936 37240 9988
rect 68100 10013 68109 10047
rect 68109 10013 68143 10047
rect 68143 10013 68152 10047
rect 68100 10004 68152 10013
rect 33876 9868 33928 9920
rect 35072 9911 35124 9920
rect 35072 9877 35081 9911
rect 35081 9877 35115 9911
rect 35115 9877 35124 9911
rect 35072 9868 35124 9877
rect 38200 9911 38252 9920
rect 38200 9877 38209 9911
rect 38209 9877 38243 9911
rect 38243 9877 38252 9911
rect 38200 9868 38252 9877
rect 39304 9868 39356 9920
rect 39856 9868 39908 9920
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 50294 9766 50346 9818
rect 50358 9766 50410 9818
rect 50422 9766 50474 9818
rect 50486 9766 50538 9818
rect 50550 9766 50602 9818
rect 5172 9664 5224 9716
rect 12256 9664 12308 9716
rect 14556 9664 14608 9716
rect 20536 9707 20588 9716
rect 6092 9596 6144 9648
rect 8300 9596 8352 9648
rect 11428 9596 11480 9648
rect 5448 9571 5500 9580
rect 5448 9537 5457 9571
rect 5457 9537 5491 9571
rect 5491 9537 5500 9571
rect 5448 9528 5500 9537
rect 5724 9528 5776 9580
rect 6920 9571 6972 9580
rect 6920 9537 6929 9571
rect 6929 9537 6963 9571
rect 6963 9537 6972 9571
rect 6920 9528 6972 9537
rect 9680 9528 9732 9580
rect 9772 9571 9824 9580
rect 9772 9537 9781 9571
rect 9781 9537 9815 9571
rect 9815 9537 9824 9571
rect 9772 9528 9824 9537
rect 10324 9528 10376 9580
rect 6552 9460 6604 9512
rect 7288 9460 7340 9512
rect 8760 9460 8812 9512
rect 7104 9392 7156 9444
rect 10508 9528 10560 9580
rect 10784 9571 10836 9580
rect 10784 9537 10793 9571
rect 10793 9537 10827 9571
rect 10827 9537 10836 9571
rect 10784 9528 10836 9537
rect 5632 9324 5684 9376
rect 7748 9324 7800 9376
rect 11152 9528 11204 9580
rect 11980 9528 12032 9580
rect 15200 9596 15252 9648
rect 14740 9571 14792 9580
rect 14740 9537 14749 9571
rect 14749 9537 14783 9571
rect 14783 9537 14792 9571
rect 14740 9528 14792 9537
rect 11796 9392 11848 9444
rect 11428 9324 11480 9376
rect 12716 9460 12768 9512
rect 14832 9460 14884 9512
rect 15476 9528 15528 9580
rect 16856 9571 16908 9580
rect 16856 9537 16865 9571
rect 16865 9537 16899 9571
rect 16899 9537 16908 9571
rect 16856 9528 16908 9537
rect 20536 9673 20545 9707
rect 20545 9673 20579 9707
rect 20579 9673 20588 9707
rect 20536 9664 20588 9673
rect 20812 9664 20864 9716
rect 25688 9664 25740 9716
rect 18420 9596 18472 9648
rect 17132 9571 17184 9580
rect 17132 9537 17141 9571
rect 17141 9537 17175 9571
rect 17175 9537 17184 9571
rect 17132 9528 17184 9537
rect 17224 9571 17276 9580
rect 17224 9537 17233 9571
rect 17233 9537 17267 9571
rect 17267 9537 17276 9571
rect 17224 9528 17276 9537
rect 12532 9392 12584 9444
rect 15384 9392 15436 9444
rect 18236 9435 18288 9444
rect 18236 9401 18245 9435
rect 18245 9401 18279 9435
rect 18279 9401 18288 9435
rect 18236 9392 18288 9401
rect 12164 9367 12216 9376
rect 12164 9333 12173 9367
rect 12173 9333 12207 9367
rect 12207 9333 12216 9367
rect 12164 9324 12216 9333
rect 15660 9324 15712 9376
rect 18788 9571 18840 9580
rect 18788 9537 18797 9571
rect 18797 9537 18831 9571
rect 18831 9537 18840 9571
rect 18788 9528 18840 9537
rect 19340 9460 19392 9512
rect 19984 9528 20036 9580
rect 21272 9596 21324 9648
rect 22560 9639 22612 9648
rect 22560 9605 22569 9639
rect 22569 9605 22603 9639
rect 22603 9605 22612 9639
rect 22560 9596 22612 9605
rect 24492 9639 24544 9648
rect 20812 9571 20864 9580
rect 20812 9537 20821 9571
rect 20821 9537 20855 9571
rect 20855 9537 20864 9571
rect 20812 9528 20864 9537
rect 22284 9528 22336 9580
rect 23388 9571 23440 9580
rect 23388 9537 23397 9571
rect 23397 9537 23431 9571
rect 23431 9537 23440 9571
rect 23388 9528 23440 9537
rect 24032 9528 24084 9580
rect 24492 9605 24526 9639
rect 24526 9605 24544 9639
rect 24492 9596 24544 9605
rect 27436 9664 27488 9716
rect 26792 9528 26844 9580
rect 29092 9571 29144 9580
rect 29092 9537 29101 9571
rect 29101 9537 29135 9571
rect 29135 9537 29144 9571
rect 29092 9528 29144 9537
rect 29276 9571 29328 9580
rect 29276 9537 29285 9571
rect 29285 9537 29319 9571
rect 29319 9537 29328 9571
rect 29276 9528 29328 9537
rect 30288 9596 30340 9648
rect 30564 9596 30616 9648
rect 33692 9596 33744 9648
rect 34428 9664 34480 9716
rect 30748 9571 30800 9580
rect 18512 9392 18564 9444
rect 20996 9460 21048 9512
rect 24216 9503 24268 9512
rect 24216 9469 24225 9503
rect 24225 9469 24259 9503
rect 24259 9469 24268 9503
rect 24216 9460 24268 9469
rect 30748 9537 30757 9571
rect 30757 9537 30791 9571
rect 30791 9537 30800 9571
rect 30748 9528 30800 9537
rect 29092 9392 29144 9444
rect 31116 9460 31168 9512
rect 33508 9528 33560 9580
rect 32036 9460 32088 9512
rect 33876 9571 33928 9580
rect 33876 9537 33885 9571
rect 33885 9537 33919 9571
rect 33919 9537 33928 9571
rect 35072 9596 35124 9648
rect 33876 9528 33928 9537
rect 34244 9571 34296 9580
rect 34244 9537 34253 9571
rect 34253 9537 34287 9571
rect 34287 9537 34296 9571
rect 34244 9528 34296 9537
rect 34428 9528 34480 9580
rect 35164 9571 35216 9580
rect 35164 9537 35173 9571
rect 35173 9537 35207 9571
rect 35207 9537 35216 9571
rect 35164 9528 35216 9537
rect 35440 9596 35492 9648
rect 35808 9528 35860 9580
rect 36360 9571 36412 9580
rect 36360 9537 36369 9571
rect 36369 9537 36403 9571
rect 36403 9537 36412 9571
rect 36360 9528 36412 9537
rect 30288 9392 30340 9444
rect 33232 9392 33284 9444
rect 35716 9460 35768 9512
rect 37188 9528 37240 9580
rect 37556 9528 37608 9580
rect 37927 9574 37979 9580
rect 37927 9540 37936 9574
rect 37936 9540 37970 9574
rect 37970 9540 37979 9574
rect 37927 9528 37979 9540
rect 38200 9528 38252 9580
rect 38568 9460 38620 9512
rect 21088 9324 21140 9376
rect 24584 9324 24636 9376
rect 29736 9367 29788 9376
rect 29736 9333 29745 9367
rect 29745 9333 29779 9367
rect 29779 9333 29788 9367
rect 29736 9324 29788 9333
rect 35532 9324 35584 9376
rect 37096 9324 37148 9376
rect 40868 9324 40920 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 65654 9222 65706 9274
rect 65718 9222 65770 9274
rect 65782 9222 65834 9274
rect 65846 9222 65898 9274
rect 65910 9222 65962 9274
rect 1952 9163 2004 9172
rect 1952 9129 1961 9163
rect 1961 9129 1995 9163
rect 1995 9129 2004 9163
rect 1952 9120 2004 9129
rect 5172 9163 5224 9172
rect 5172 9129 5181 9163
rect 5181 9129 5215 9163
rect 5215 9129 5224 9163
rect 5172 9120 5224 9129
rect 10324 9163 10376 9172
rect 10324 9129 10333 9163
rect 10333 9129 10367 9163
rect 10367 9129 10376 9163
rect 10324 9120 10376 9129
rect 13268 9163 13320 9172
rect 13268 9129 13277 9163
rect 13277 9129 13311 9163
rect 13311 9129 13320 9163
rect 13268 9120 13320 9129
rect 14188 9120 14240 9172
rect 9864 8984 9916 9036
rect 2780 8916 2832 8968
rect 3516 8916 3568 8968
rect 5264 8916 5316 8968
rect 6920 8916 6972 8968
rect 7748 8959 7800 8968
rect 7748 8925 7757 8959
rect 7757 8925 7791 8959
rect 7791 8925 7800 8959
rect 7748 8916 7800 8925
rect 7932 8959 7984 8968
rect 7932 8925 7941 8959
rect 7941 8925 7975 8959
rect 7975 8925 7984 8959
rect 7932 8916 7984 8925
rect 2228 8848 2280 8900
rect 2412 8848 2464 8900
rect 2780 8780 2832 8832
rect 3056 8780 3108 8832
rect 5080 8848 5132 8900
rect 8116 8959 8168 8968
rect 8116 8925 8125 8959
rect 8125 8925 8159 8959
rect 8159 8925 8168 8959
rect 8116 8916 8168 8925
rect 11796 9052 11848 9104
rect 17132 9120 17184 9172
rect 17500 9120 17552 9172
rect 18512 9120 18564 9172
rect 20076 9163 20128 9172
rect 20076 9129 20085 9163
rect 20085 9129 20119 9163
rect 20119 9129 20128 9163
rect 20076 9120 20128 9129
rect 23388 9120 23440 9172
rect 11612 8984 11664 9036
rect 16212 8984 16264 9036
rect 10140 8916 10192 8968
rect 10692 8916 10744 8968
rect 12164 8959 12216 8968
rect 12164 8925 12198 8959
rect 12198 8925 12216 8959
rect 12164 8916 12216 8925
rect 15660 8959 15712 8968
rect 15660 8925 15678 8959
rect 15678 8925 15712 8959
rect 15660 8916 15712 8925
rect 7012 8780 7064 8832
rect 7288 8823 7340 8832
rect 7288 8789 7297 8823
rect 7297 8789 7331 8823
rect 7331 8789 7340 8823
rect 7288 8780 7340 8789
rect 8392 8823 8444 8832
rect 8392 8789 8401 8823
rect 8401 8789 8435 8823
rect 8435 8789 8444 8823
rect 8392 8780 8444 8789
rect 10784 8780 10836 8832
rect 11152 8823 11204 8832
rect 11152 8789 11161 8823
rect 11161 8789 11195 8823
rect 11195 8789 11204 8823
rect 11152 8780 11204 8789
rect 13360 8780 13412 8832
rect 15476 8780 15528 8832
rect 19340 8916 19392 8968
rect 20168 8916 20220 8968
rect 20812 8984 20864 9036
rect 20352 8916 20404 8968
rect 20628 8916 20680 8968
rect 23112 8916 23164 8968
rect 18788 8848 18840 8900
rect 21180 8891 21232 8900
rect 21180 8857 21189 8891
rect 21189 8857 21223 8891
rect 21223 8857 21232 8891
rect 21180 8848 21232 8857
rect 21640 8848 21692 8900
rect 24216 8984 24268 9036
rect 27712 9120 27764 9172
rect 29000 9120 29052 9172
rect 29276 9120 29328 9172
rect 36360 9120 36412 9172
rect 29828 9052 29880 9104
rect 35716 9052 35768 9104
rect 35808 9052 35860 9104
rect 30748 9027 30800 9036
rect 19156 8780 19208 8832
rect 20076 8780 20128 8832
rect 22100 8780 22152 8832
rect 27252 8916 27304 8968
rect 30748 8993 30757 9027
rect 30757 8993 30791 9027
rect 30791 8993 30800 9027
rect 30748 8984 30800 8993
rect 30840 8984 30892 9036
rect 31852 8984 31904 9036
rect 29368 8916 29420 8968
rect 29920 8959 29972 8968
rect 23848 8823 23900 8832
rect 23848 8789 23857 8823
rect 23857 8789 23891 8823
rect 23891 8789 23900 8823
rect 23848 8780 23900 8789
rect 24308 8780 24360 8832
rect 24492 8780 24544 8832
rect 24676 8848 24728 8900
rect 25780 8848 25832 8900
rect 27804 8891 27856 8900
rect 27804 8857 27838 8891
rect 27838 8857 27856 8891
rect 29920 8925 29929 8959
rect 29929 8925 29963 8959
rect 29963 8925 29972 8959
rect 29920 8916 29972 8925
rect 30196 8916 30248 8968
rect 31116 8916 31168 8968
rect 31944 8959 31996 8968
rect 31944 8925 31953 8959
rect 31953 8925 31987 8959
rect 31987 8925 31996 8959
rect 31944 8916 31996 8925
rect 33232 8959 33284 8968
rect 27804 8848 27856 8857
rect 31024 8848 31076 8900
rect 31484 8848 31536 8900
rect 33232 8925 33241 8959
rect 33241 8925 33275 8959
rect 33275 8925 33284 8959
rect 33232 8916 33284 8925
rect 33508 8984 33560 9036
rect 33416 8959 33468 8968
rect 33416 8925 33425 8959
rect 33425 8925 33459 8959
rect 33459 8925 33468 8959
rect 33416 8916 33468 8925
rect 33876 8916 33928 8968
rect 28448 8780 28500 8832
rect 28816 8780 28868 8832
rect 31852 8780 31904 8832
rect 34520 8848 34572 8900
rect 35716 8848 35768 8900
rect 37188 8959 37240 8968
rect 37188 8925 37197 8959
rect 37197 8925 37231 8959
rect 37231 8925 37240 8959
rect 37372 8959 37424 8968
rect 37188 8916 37240 8925
rect 37372 8925 37381 8959
rect 37381 8925 37415 8959
rect 37415 8925 37424 8959
rect 37372 8916 37424 8925
rect 38200 8984 38252 9036
rect 32404 8823 32456 8832
rect 32404 8789 32413 8823
rect 32413 8789 32447 8823
rect 32447 8789 32456 8823
rect 32404 8780 32456 8789
rect 33048 8780 33100 8832
rect 34060 8823 34112 8832
rect 34060 8789 34069 8823
rect 34069 8789 34103 8823
rect 34103 8789 34112 8823
rect 34060 8780 34112 8789
rect 37924 8848 37976 8900
rect 39304 8848 39356 8900
rect 38660 8823 38712 8832
rect 38660 8789 38669 8823
rect 38669 8789 38703 8823
rect 38703 8789 38712 8823
rect 38660 8780 38712 8789
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 50294 8678 50346 8730
rect 50358 8678 50410 8730
rect 50422 8678 50474 8730
rect 50486 8678 50538 8730
rect 50550 8678 50602 8730
rect 2044 8576 2096 8628
rect 1860 8440 1912 8492
rect 2412 8440 2464 8492
rect 3516 8508 3568 8560
rect 5080 8576 5132 8628
rect 5632 8576 5684 8628
rect 7932 8576 7984 8628
rect 5264 8508 5316 8560
rect 5172 8440 5224 8492
rect 7012 8508 7064 8560
rect 14372 8576 14424 8628
rect 8392 8508 8444 8560
rect 17040 8576 17092 8628
rect 6920 8440 6972 8492
rect 7104 8440 7156 8492
rect 7932 8483 7984 8492
rect 7932 8449 7941 8483
rect 7941 8449 7975 8483
rect 7975 8449 7984 8483
rect 7932 8440 7984 8449
rect 15016 8508 15068 8560
rect 14464 8483 14516 8492
rect 2136 8304 2188 8356
rect 5908 8372 5960 8424
rect 7012 8415 7064 8424
rect 7012 8381 7021 8415
rect 7021 8381 7055 8415
rect 7055 8381 7064 8415
rect 7012 8372 7064 8381
rect 7472 8372 7524 8424
rect 3792 8304 3844 8356
rect 14464 8449 14473 8483
rect 14473 8449 14507 8483
rect 14507 8449 14516 8483
rect 14464 8440 14516 8449
rect 15108 8440 15160 8492
rect 8760 8415 8812 8424
rect 8760 8381 8769 8415
rect 8769 8381 8803 8415
rect 8803 8381 8812 8415
rect 8760 8372 8812 8381
rect 14372 8372 14424 8424
rect 16764 8440 16816 8492
rect 16672 8415 16724 8424
rect 16672 8381 16681 8415
rect 16681 8381 16715 8415
rect 16715 8381 16724 8415
rect 16672 8372 16724 8381
rect 8116 8304 8168 8356
rect 13636 8304 13688 8356
rect 15292 8304 15344 8356
rect 9772 8236 9824 8288
rect 10692 8279 10744 8288
rect 10692 8245 10701 8279
rect 10701 8245 10735 8279
rect 10735 8245 10744 8279
rect 10692 8236 10744 8245
rect 14740 8236 14792 8288
rect 14832 8236 14884 8288
rect 17408 8236 17460 8288
rect 18696 8440 18748 8492
rect 18972 8483 19024 8492
rect 18972 8449 18981 8483
rect 18981 8449 19015 8483
rect 19015 8449 19024 8483
rect 18972 8440 19024 8449
rect 19248 8576 19300 8628
rect 24492 8576 24544 8628
rect 25320 8576 25372 8628
rect 30840 8576 30892 8628
rect 31484 8619 31536 8628
rect 31484 8585 31493 8619
rect 31493 8585 31527 8619
rect 31527 8585 31536 8619
rect 31484 8576 31536 8585
rect 20076 8551 20128 8560
rect 20076 8517 20085 8551
rect 20085 8517 20119 8551
rect 20119 8517 20128 8551
rect 20076 8508 20128 8517
rect 19156 8483 19208 8492
rect 19156 8449 19165 8483
rect 19165 8449 19199 8483
rect 19199 8449 19208 8483
rect 19156 8440 19208 8449
rect 22100 8440 22152 8492
rect 23572 8440 23624 8492
rect 24400 8508 24452 8560
rect 27528 8508 27580 8560
rect 34060 8576 34112 8628
rect 34612 8576 34664 8628
rect 32404 8508 32456 8560
rect 34704 8551 34756 8560
rect 34704 8517 34713 8551
rect 34713 8517 34747 8551
rect 34747 8517 34756 8551
rect 34704 8508 34756 8517
rect 24308 8483 24360 8492
rect 24308 8449 24317 8483
rect 24317 8449 24351 8483
rect 24351 8449 24360 8483
rect 24308 8440 24360 8449
rect 25136 8483 25188 8492
rect 23848 8372 23900 8424
rect 25136 8449 25145 8483
rect 25145 8449 25179 8483
rect 25179 8449 25188 8483
rect 25136 8440 25188 8449
rect 27712 8440 27764 8492
rect 33600 8440 33652 8492
rect 34152 8483 34204 8492
rect 34152 8449 34161 8483
rect 34161 8449 34195 8483
rect 34195 8449 34204 8483
rect 34152 8440 34204 8449
rect 29184 8372 29236 8424
rect 33508 8415 33560 8424
rect 33508 8381 33517 8415
rect 33517 8381 33551 8415
rect 33551 8381 33560 8415
rect 33508 8372 33560 8381
rect 27804 8347 27856 8356
rect 19432 8279 19484 8288
rect 19432 8245 19441 8279
rect 19441 8245 19475 8279
rect 19475 8245 19484 8279
rect 19432 8236 19484 8245
rect 25228 8236 25280 8288
rect 27804 8313 27813 8347
rect 27813 8313 27847 8347
rect 27847 8313 27856 8347
rect 27804 8304 27856 8313
rect 27988 8304 28040 8356
rect 35348 8576 35400 8628
rect 37372 8576 37424 8628
rect 36360 8551 36412 8560
rect 36360 8517 36369 8551
rect 36369 8517 36403 8551
rect 36403 8517 36412 8551
rect 36360 8508 36412 8517
rect 38660 8576 38712 8628
rect 38200 8508 38252 8560
rect 36544 8483 36596 8492
rect 36544 8449 36553 8483
rect 36553 8449 36587 8483
rect 36587 8449 36596 8483
rect 36544 8440 36596 8449
rect 37188 8440 37240 8492
rect 35808 8372 35860 8424
rect 37760 8483 37812 8492
rect 37760 8449 37795 8483
rect 37795 8449 37812 8483
rect 37760 8440 37812 8449
rect 38016 8440 38068 8492
rect 37924 8372 37976 8424
rect 38568 8372 38620 8424
rect 28724 8236 28776 8288
rect 31576 8236 31628 8288
rect 32128 8279 32180 8288
rect 32128 8245 32137 8279
rect 32137 8245 32171 8279
rect 32171 8245 32180 8279
rect 37832 8304 37884 8356
rect 40960 8440 41012 8492
rect 67548 8304 67600 8356
rect 32128 8236 32180 8245
rect 34060 8279 34112 8288
rect 34060 8245 34069 8279
rect 34069 8245 34103 8279
rect 34103 8245 34112 8279
rect 34060 8236 34112 8245
rect 34244 8236 34296 8288
rect 37740 8236 37792 8288
rect 38016 8279 38068 8288
rect 38016 8245 38025 8279
rect 38025 8245 38059 8279
rect 38059 8245 38068 8279
rect 38016 8236 38068 8245
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 65654 8134 65706 8186
rect 65718 8134 65770 8186
rect 65782 8134 65834 8186
rect 65846 8134 65898 8186
rect 65910 8134 65962 8186
rect 1860 8032 1912 8084
rect 2504 8032 2556 8084
rect 3792 8032 3844 8084
rect 8668 8032 8720 8084
rect 15568 8032 15620 8084
rect 16764 8032 16816 8084
rect 18972 8032 19024 8084
rect 25780 8032 25832 8084
rect 28908 8032 28960 8084
rect 31024 8075 31076 8084
rect 31024 8041 31033 8075
rect 31033 8041 31067 8075
rect 31067 8041 31076 8075
rect 31024 8032 31076 8041
rect 31760 8032 31812 8084
rect 32128 8032 32180 8084
rect 6000 7964 6052 8016
rect 2136 7896 2188 7948
rect 6276 7896 6328 7948
rect 8576 7964 8628 8016
rect 11152 8007 11204 8016
rect 11152 7973 11161 8007
rect 11161 7973 11195 8007
rect 11195 7973 11204 8007
rect 11152 7964 11204 7973
rect 14648 7964 14700 8016
rect 9772 7896 9824 7948
rect 1768 7828 1820 7880
rect 5448 7828 5500 7880
rect 7472 7828 7524 7880
rect 12716 7828 12768 7880
rect 15752 7896 15804 7948
rect 21640 7939 21692 7948
rect 21640 7905 21649 7939
rect 21649 7905 21683 7939
rect 21683 7905 21692 7939
rect 21640 7896 21692 7905
rect 2320 7760 2372 7812
rect 5724 7803 5776 7812
rect 5724 7769 5733 7803
rect 5733 7769 5767 7803
rect 5767 7769 5776 7803
rect 5724 7760 5776 7769
rect 6460 7760 6512 7812
rect 7932 7760 7984 7812
rect 12256 7803 12308 7812
rect 12256 7769 12274 7803
rect 12274 7769 12308 7803
rect 12256 7760 12308 7769
rect 6000 7692 6052 7744
rect 8392 7692 8444 7744
rect 9312 7692 9364 7744
rect 13820 7692 13872 7744
rect 14280 7735 14332 7744
rect 14280 7701 14289 7735
rect 14289 7701 14323 7735
rect 14323 7701 14332 7735
rect 14280 7692 14332 7701
rect 14740 7871 14792 7880
rect 14740 7837 14749 7871
rect 14749 7837 14783 7871
rect 14783 7837 14792 7871
rect 14740 7828 14792 7837
rect 15568 7871 15620 7880
rect 15568 7837 15577 7871
rect 15577 7837 15611 7871
rect 15611 7837 15620 7871
rect 15568 7828 15620 7837
rect 16120 7760 16172 7812
rect 16304 7871 16356 7880
rect 16304 7837 16313 7871
rect 16313 7837 16347 7871
rect 16347 7837 16356 7871
rect 16304 7828 16356 7837
rect 16764 7828 16816 7880
rect 17132 7871 17184 7880
rect 17132 7837 17141 7871
rect 17141 7837 17175 7871
rect 17175 7837 17184 7871
rect 17132 7828 17184 7837
rect 17408 7871 17460 7880
rect 17408 7837 17417 7871
rect 17417 7837 17451 7871
rect 17451 7837 17460 7871
rect 17408 7828 17460 7837
rect 18236 7871 18288 7880
rect 18236 7837 18245 7871
rect 18245 7837 18279 7871
rect 18279 7837 18288 7871
rect 18236 7828 18288 7837
rect 18512 7871 18564 7880
rect 18512 7837 18521 7871
rect 18521 7837 18555 7871
rect 18555 7837 18564 7871
rect 18512 7828 18564 7837
rect 19892 7828 19944 7880
rect 21088 7828 21140 7880
rect 25780 7896 25832 7948
rect 28540 7939 28592 7948
rect 28540 7905 28549 7939
rect 28549 7905 28583 7939
rect 28583 7905 28592 7939
rect 28540 7896 28592 7905
rect 31300 7896 31352 7948
rect 31576 7939 31628 7948
rect 31576 7905 31585 7939
rect 31585 7905 31619 7939
rect 31619 7905 31628 7939
rect 31576 7896 31628 7905
rect 25228 7871 25280 7880
rect 25228 7837 25237 7871
rect 25237 7837 25271 7871
rect 25271 7837 25280 7871
rect 25228 7828 25280 7837
rect 19248 7760 19300 7812
rect 19432 7760 19484 7812
rect 22192 7760 22244 7812
rect 23848 7803 23900 7812
rect 23848 7769 23857 7803
rect 23857 7769 23891 7803
rect 23891 7769 23900 7803
rect 23848 7760 23900 7769
rect 24676 7760 24728 7812
rect 25412 7871 25464 7880
rect 25412 7837 25421 7871
rect 25421 7837 25455 7871
rect 25455 7837 25464 7871
rect 25412 7828 25464 7837
rect 28356 7803 28408 7812
rect 28356 7769 28365 7803
rect 28365 7769 28399 7803
rect 28399 7769 28408 7803
rect 28356 7760 28408 7769
rect 28448 7760 28500 7812
rect 29184 7828 29236 7880
rect 29736 7828 29788 7880
rect 31024 7828 31076 7880
rect 33508 8032 33560 8084
rect 34152 8075 34204 8084
rect 34152 8041 34161 8075
rect 34161 8041 34195 8075
rect 34195 8041 34204 8075
rect 34152 8032 34204 8041
rect 35808 8032 35860 8084
rect 39304 8075 39356 8084
rect 39304 8041 39313 8075
rect 39313 8041 39347 8075
rect 39347 8041 39356 8075
rect 39304 8032 39356 8041
rect 34520 7964 34572 8016
rect 33048 7871 33100 7880
rect 33048 7837 33082 7871
rect 33082 7837 33100 7871
rect 33048 7828 33100 7837
rect 35716 7828 35768 7880
rect 37924 7871 37976 7880
rect 37924 7837 37933 7871
rect 37933 7837 37967 7871
rect 37967 7837 37976 7871
rect 37924 7828 37976 7837
rect 38016 7828 38068 7880
rect 29552 7760 29604 7812
rect 14924 7692 14976 7744
rect 15016 7692 15068 7744
rect 18328 7735 18380 7744
rect 18328 7701 18337 7735
rect 18337 7701 18371 7735
rect 18371 7701 18380 7735
rect 18328 7692 18380 7701
rect 18512 7692 18564 7744
rect 23112 7692 23164 7744
rect 23572 7692 23624 7744
rect 24124 7692 24176 7744
rect 24492 7735 24544 7744
rect 24492 7701 24501 7735
rect 24501 7701 24535 7735
rect 24535 7701 24544 7735
rect 24492 7692 24544 7701
rect 26148 7692 26200 7744
rect 29828 7692 29880 7744
rect 31944 7735 31996 7744
rect 31944 7701 31953 7735
rect 31953 7701 31987 7735
rect 31987 7701 31996 7735
rect 31944 7692 31996 7701
rect 37096 7803 37148 7812
rect 37096 7769 37114 7803
rect 37114 7769 37148 7803
rect 37096 7760 37148 7769
rect 34796 7692 34848 7744
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 50294 7590 50346 7642
rect 50358 7590 50410 7642
rect 50422 7590 50474 7642
rect 50486 7590 50538 7642
rect 50550 7590 50602 7642
rect 2412 7531 2464 7540
rect 2412 7497 2421 7531
rect 2421 7497 2455 7531
rect 2455 7497 2464 7531
rect 2412 7488 2464 7497
rect 5724 7488 5776 7540
rect 8668 7531 8720 7540
rect 3516 7352 3568 7404
rect 5540 7352 5592 7404
rect 6460 7395 6512 7404
rect 6460 7361 6469 7395
rect 6469 7361 6503 7395
rect 6503 7361 6512 7395
rect 6460 7352 6512 7361
rect 8668 7497 8677 7531
rect 8677 7497 8711 7531
rect 8711 7497 8720 7531
rect 8668 7488 8720 7497
rect 9772 7531 9824 7540
rect 9772 7497 9781 7531
rect 9781 7497 9815 7531
rect 9815 7497 9824 7531
rect 9772 7488 9824 7497
rect 12256 7531 12308 7540
rect 12256 7497 12265 7531
rect 12265 7497 12299 7531
rect 12299 7497 12308 7531
rect 12256 7488 12308 7497
rect 13084 7488 13136 7540
rect 8760 7420 8812 7472
rect 11152 7420 11204 7472
rect 7564 7395 7616 7404
rect 7564 7361 7598 7395
rect 7598 7361 7616 7395
rect 11520 7395 11572 7404
rect 7564 7352 7616 7361
rect 11520 7361 11529 7395
rect 11529 7361 11563 7395
rect 11563 7361 11572 7395
rect 11520 7352 11572 7361
rect 11704 7395 11756 7404
rect 11704 7361 11713 7395
rect 11713 7361 11747 7395
rect 11747 7361 11756 7395
rect 11704 7352 11756 7361
rect 14280 7420 14332 7472
rect 11612 7284 11664 7336
rect 12532 7284 12584 7336
rect 2320 7148 2372 7200
rect 7104 7148 7156 7200
rect 9036 7216 9088 7268
rect 12716 7327 12768 7336
rect 12716 7293 12725 7327
rect 12725 7293 12759 7327
rect 12759 7293 12768 7327
rect 12716 7284 12768 7293
rect 7932 7148 7984 7200
rect 10232 7191 10284 7200
rect 10232 7157 10241 7191
rect 10241 7157 10275 7191
rect 10275 7157 10284 7191
rect 10232 7148 10284 7157
rect 11336 7148 11388 7200
rect 18328 7488 18380 7540
rect 19432 7488 19484 7540
rect 20076 7488 20128 7540
rect 25596 7488 25648 7540
rect 22192 7420 22244 7472
rect 19156 7352 19208 7404
rect 21088 7395 21140 7404
rect 21088 7361 21097 7395
rect 21097 7361 21131 7395
rect 21131 7361 21140 7395
rect 21088 7352 21140 7361
rect 22560 7420 22612 7472
rect 24308 7420 24360 7472
rect 15016 7327 15068 7336
rect 15016 7293 15025 7327
rect 15025 7293 15059 7327
rect 15059 7293 15068 7327
rect 15016 7284 15068 7293
rect 16764 7284 16816 7336
rect 22468 7395 22520 7404
rect 22468 7361 22477 7395
rect 22477 7361 22511 7395
rect 22511 7361 22520 7395
rect 22468 7352 22520 7361
rect 22652 7395 22704 7404
rect 22652 7361 22661 7395
rect 22661 7361 22695 7395
rect 22695 7361 22704 7395
rect 24400 7395 24452 7404
rect 22652 7352 22704 7361
rect 24400 7361 24409 7395
rect 24409 7361 24443 7395
rect 24443 7361 24452 7395
rect 24400 7352 24452 7361
rect 25780 7395 25832 7404
rect 25780 7361 25789 7395
rect 25789 7361 25823 7395
rect 25823 7361 25832 7395
rect 25780 7352 25832 7361
rect 13728 7148 13780 7200
rect 14464 7148 14516 7200
rect 14740 7148 14792 7200
rect 23296 7284 23348 7336
rect 24676 7327 24728 7336
rect 24676 7293 24685 7327
rect 24685 7293 24719 7327
rect 24719 7293 24728 7327
rect 24676 7284 24728 7293
rect 16488 7216 16540 7268
rect 22376 7216 22428 7268
rect 26148 7395 26200 7404
rect 26148 7361 26157 7395
rect 26157 7361 26191 7395
rect 26191 7361 26200 7395
rect 26148 7352 26200 7361
rect 33232 7488 33284 7540
rect 34796 7488 34848 7540
rect 37740 7488 37792 7540
rect 34520 7420 34572 7472
rect 35716 7420 35768 7472
rect 26240 7284 26292 7336
rect 26976 7327 27028 7336
rect 26976 7293 26985 7327
rect 26985 7293 27019 7327
rect 27019 7293 27028 7327
rect 26976 7284 27028 7293
rect 28264 7284 28316 7336
rect 28908 7284 28960 7336
rect 29828 7395 29880 7404
rect 29828 7361 29837 7395
rect 29837 7361 29871 7395
rect 29871 7361 29880 7395
rect 29828 7352 29880 7361
rect 35532 7352 35584 7404
rect 30656 7284 30708 7336
rect 26608 7216 26660 7268
rect 15844 7148 15896 7200
rect 16948 7148 17000 7200
rect 22192 7148 22244 7200
rect 23756 7148 23808 7200
rect 24860 7148 24912 7200
rect 25412 7148 25464 7200
rect 27344 7148 27396 7200
rect 28540 7148 28592 7200
rect 29644 7148 29696 7200
rect 30932 7148 30984 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 65654 7046 65706 7098
rect 65718 7046 65770 7098
rect 65782 7046 65834 7098
rect 65846 7046 65898 7098
rect 65910 7046 65962 7098
rect 7564 6987 7616 6996
rect 7564 6953 7573 6987
rect 7573 6953 7607 6987
rect 7607 6953 7616 6987
rect 7564 6944 7616 6953
rect 4068 6876 4120 6928
rect 6184 6876 6236 6928
rect 11336 6944 11388 6996
rect 11612 6987 11664 6996
rect 11612 6953 11621 6987
rect 11621 6953 11655 6987
rect 11655 6953 11664 6987
rect 11612 6944 11664 6953
rect 12348 6944 12400 6996
rect 12532 6944 12584 6996
rect 11520 6876 11572 6928
rect 12256 6876 12308 6928
rect 18696 6944 18748 6996
rect 26976 6944 27028 6996
rect 29184 6944 29236 6996
rect 29644 6944 29696 6996
rect 31852 6987 31904 6996
rect 31852 6953 31861 6987
rect 31861 6953 31895 6987
rect 31895 6953 31904 6987
rect 31852 6944 31904 6953
rect 5540 6851 5592 6860
rect 5540 6817 5549 6851
rect 5549 6817 5583 6851
rect 5583 6817 5592 6851
rect 5540 6808 5592 6817
rect 1952 6783 2004 6792
rect 1952 6749 1961 6783
rect 1961 6749 1995 6783
rect 1995 6749 2004 6783
rect 1952 6740 2004 6749
rect 2044 6783 2096 6792
rect 2044 6749 2053 6783
rect 2053 6749 2087 6783
rect 2087 6749 2096 6783
rect 2044 6740 2096 6749
rect 3056 6740 3108 6792
rect 4068 6740 4120 6792
rect 5724 6740 5776 6792
rect 2964 6672 3016 6724
rect 6000 6783 6052 6792
rect 6000 6749 6009 6783
rect 6009 6749 6043 6783
rect 6043 6749 6052 6783
rect 6000 6740 6052 6749
rect 6276 6740 6328 6792
rect 8668 6808 8720 6860
rect 8760 6808 8812 6860
rect 15016 6808 15068 6860
rect 7104 6783 7156 6792
rect 7104 6749 7113 6783
rect 7113 6749 7147 6783
rect 7147 6749 7156 6783
rect 7104 6740 7156 6749
rect 6736 6672 6788 6724
rect 7288 6783 7340 6792
rect 7288 6749 7297 6783
rect 7297 6749 7331 6783
rect 7331 6749 7340 6783
rect 7288 6740 7340 6749
rect 7472 6740 7524 6792
rect 11060 6783 11112 6792
rect 9220 6672 9272 6724
rect 2504 6604 2556 6656
rect 3516 6604 3568 6656
rect 8300 6647 8352 6656
rect 8300 6613 8309 6647
rect 8309 6613 8343 6647
rect 8343 6613 8352 6647
rect 8300 6604 8352 6613
rect 10416 6604 10468 6656
rect 11060 6749 11069 6783
rect 11069 6749 11103 6783
rect 11103 6749 11112 6783
rect 11060 6740 11112 6749
rect 11336 6783 11388 6792
rect 11336 6749 11345 6783
rect 11345 6749 11379 6783
rect 11379 6749 11388 6783
rect 11336 6740 11388 6749
rect 11428 6783 11480 6792
rect 11428 6749 11437 6783
rect 11437 6749 11471 6783
rect 11471 6749 11480 6783
rect 11428 6740 11480 6749
rect 14004 6740 14056 6792
rect 14280 6740 14332 6792
rect 12440 6672 12492 6724
rect 12348 6604 12400 6656
rect 12808 6604 12860 6656
rect 15660 6740 15712 6792
rect 16120 6783 16172 6792
rect 16120 6749 16129 6783
rect 16129 6749 16163 6783
rect 16163 6749 16172 6783
rect 16120 6740 16172 6749
rect 16304 6783 16356 6792
rect 16304 6749 16313 6783
rect 16313 6749 16347 6783
rect 16347 6749 16356 6783
rect 16304 6740 16356 6749
rect 16580 6808 16632 6860
rect 16764 6876 16816 6928
rect 28908 6876 28960 6928
rect 19156 6808 19208 6860
rect 19984 6851 20036 6860
rect 19984 6817 19993 6851
rect 19993 6817 20027 6851
rect 20027 6817 20036 6851
rect 19984 6808 20036 6817
rect 22100 6851 22152 6860
rect 22100 6817 22109 6851
rect 22109 6817 22143 6851
rect 22143 6817 22152 6851
rect 22100 6808 22152 6817
rect 24400 6808 24452 6860
rect 26608 6851 26660 6860
rect 26608 6817 26617 6851
rect 26617 6817 26651 6851
rect 26651 6817 26660 6851
rect 26608 6808 26660 6817
rect 30564 6808 30616 6860
rect 30932 6808 30984 6860
rect 14924 6672 14976 6724
rect 17224 6740 17276 6792
rect 17960 6783 18012 6792
rect 17960 6749 17969 6783
rect 17969 6749 18003 6783
rect 18003 6749 18012 6783
rect 17960 6740 18012 6749
rect 19248 6783 19300 6792
rect 19248 6749 19257 6783
rect 19257 6749 19291 6783
rect 19291 6749 19300 6783
rect 19248 6740 19300 6749
rect 19432 6783 19484 6792
rect 19432 6749 19441 6783
rect 19441 6749 19475 6783
rect 19475 6749 19484 6783
rect 19432 6740 19484 6749
rect 21088 6740 21140 6792
rect 22192 6740 22244 6792
rect 24308 6740 24360 6792
rect 20076 6672 20128 6724
rect 16856 6604 16908 6656
rect 18512 6604 18564 6656
rect 20352 6604 20404 6656
rect 23664 6604 23716 6656
rect 25136 6740 25188 6792
rect 29828 6740 29880 6792
rect 30656 6740 30708 6792
rect 32036 6783 32088 6792
rect 32036 6749 32045 6783
rect 32045 6749 32079 6783
rect 32079 6749 32088 6783
rect 32036 6740 32088 6749
rect 32220 6740 32272 6792
rect 34796 6740 34848 6792
rect 68100 6783 68152 6792
rect 28540 6672 28592 6724
rect 31944 6672 31996 6724
rect 68100 6749 68109 6783
rect 68109 6749 68143 6783
rect 68143 6749 68152 6783
rect 68100 6740 68152 6749
rect 28264 6604 28316 6656
rect 31668 6604 31720 6656
rect 33784 6604 33836 6656
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 50294 6502 50346 6554
rect 50358 6502 50410 6554
rect 50422 6502 50474 6554
rect 50486 6502 50538 6554
rect 50550 6502 50602 6554
rect 1952 6400 2004 6452
rect 4068 6443 4120 6452
rect 4068 6409 4077 6443
rect 4077 6409 4111 6443
rect 4111 6409 4120 6443
rect 4068 6400 4120 6409
rect 6460 6443 6512 6452
rect 6460 6409 6469 6443
rect 6469 6409 6503 6443
rect 6503 6409 6512 6443
rect 9220 6443 9272 6452
rect 6460 6400 6512 6409
rect 1768 6375 1820 6384
rect 1768 6341 1777 6375
rect 1777 6341 1811 6375
rect 1811 6341 1820 6375
rect 1768 6332 1820 6341
rect 2780 6332 2832 6384
rect 3424 6332 3476 6384
rect 9220 6409 9229 6443
rect 9229 6409 9263 6443
rect 9263 6409 9272 6443
rect 9220 6400 9272 6409
rect 9772 6400 9824 6452
rect 2964 6307 3016 6316
rect 2964 6273 2998 6307
rect 2998 6273 3016 6307
rect 2964 6264 3016 6273
rect 5816 6264 5868 6316
rect 6644 6307 6696 6316
rect 6644 6273 6653 6307
rect 6653 6273 6687 6307
rect 6687 6273 6696 6307
rect 6644 6264 6696 6273
rect 8668 6264 8720 6316
rect 10416 6332 10468 6384
rect 10600 6400 10652 6452
rect 10876 6375 10928 6384
rect 10876 6341 10885 6375
rect 10885 6341 10919 6375
rect 10919 6341 10928 6375
rect 10876 6332 10928 6341
rect 6736 6196 6788 6248
rect 9128 6264 9180 6316
rect 11060 6264 11112 6316
rect 12440 6332 12492 6384
rect 8300 6128 8352 6180
rect 8668 6128 8720 6180
rect 9220 6196 9272 6248
rect 11244 6196 11296 6248
rect 11428 6128 11480 6180
rect 11980 6264 12032 6316
rect 12164 6264 12216 6316
rect 14924 6400 14976 6452
rect 16120 6400 16172 6452
rect 16028 6332 16080 6384
rect 16672 6332 16724 6384
rect 14372 6307 14424 6316
rect 14372 6273 14381 6307
rect 14381 6273 14415 6307
rect 14415 6273 14424 6307
rect 14372 6264 14424 6273
rect 14096 6196 14148 6248
rect 14924 6264 14976 6316
rect 15384 6307 15436 6316
rect 15384 6273 15393 6307
rect 15393 6273 15427 6307
rect 15427 6273 15436 6307
rect 15384 6264 15436 6273
rect 15476 6307 15528 6316
rect 15476 6273 15485 6307
rect 15485 6273 15519 6307
rect 15519 6273 15528 6307
rect 15476 6264 15528 6273
rect 15660 6307 15712 6316
rect 15660 6273 15669 6307
rect 15669 6273 15703 6307
rect 15703 6273 15712 6307
rect 15660 6264 15712 6273
rect 16856 6264 16908 6316
rect 18604 6332 18656 6384
rect 18696 6307 18748 6316
rect 18696 6273 18705 6307
rect 18705 6273 18739 6307
rect 18739 6273 18748 6307
rect 18696 6264 18748 6273
rect 18880 6307 18932 6316
rect 18880 6273 18889 6307
rect 18889 6273 18923 6307
rect 18923 6273 18932 6307
rect 18880 6264 18932 6273
rect 19156 6264 19208 6316
rect 20076 6400 20128 6452
rect 22468 6400 22520 6452
rect 23480 6400 23532 6452
rect 23664 6332 23716 6384
rect 24216 6332 24268 6384
rect 24584 6332 24636 6384
rect 21088 6264 21140 6316
rect 22192 6264 22244 6316
rect 22652 6264 22704 6316
rect 23480 6307 23532 6316
rect 23480 6273 23489 6307
rect 23489 6273 23523 6307
rect 23523 6273 23532 6307
rect 23480 6264 23532 6273
rect 19984 6196 20036 6248
rect 24768 6307 24820 6316
rect 24768 6273 24777 6307
rect 24777 6273 24811 6307
rect 24811 6273 24820 6307
rect 24768 6264 24820 6273
rect 24952 6264 25004 6316
rect 27712 6400 27764 6452
rect 27896 6400 27948 6452
rect 30656 6400 30708 6452
rect 31852 6400 31904 6452
rect 32036 6400 32088 6452
rect 28080 6196 28132 6248
rect 28264 6196 28316 6248
rect 28540 6307 28592 6316
rect 28540 6273 28554 6307
rect 28554 6273 28588 6307
rect 28588 6273 28592 6307
rect 28540 6264 28592 6273
rect 29000 6264 29052 6316
rect 29184 6307 29236 6316
rect 29184 6273 29193 6307
rect 29193 6273 29227 6307
rect 29227 6273 29236 6307
rect 29184 6264 29236 6273
rect 33692 6332 33744 6384
rect 36728 6332 36780 6384
rect 28816 6196 28868 6248
rect 32680 6307 32732 6316
rect 32680 6273 32689 6307
rect 32689 6273 32723 6307
rect 32723 6273 32732 6307
rect 32680 6264 32732 6273
rect 32956 6264 33008 6316
rect 33784 6307 33836 6316
rect 33784 6273 33793 6307
rect 33793 6273 33827 6307
rect 33827 6273 33836 6307
rect 33784 6264 33836 6273
rect 37740 6264 37792 6316
rect 39396 6264 39448 6316
rect 31116 6239 31168 6248
rect 31116 6205 31125 6239
rect 31125 6205 31159 6239
rect 31159 6205 31168 6239
rect 31116 6196 31168 6205
rect 12348 6128 12400 6180
rect 14280 6128 14332 6180
rect 3056 6060 3108 6112
rect 5816 6103 5868 6112
rect 5816 6069 5825 6103
rect 5825 6069 5859 6103
rect 5859 6069 5868 6103
rect 5816 6060 5868 6069
rect 7288 6103 7340 6112
rect 7288 6069 7297 6103
rect 7297 6069 7331 6103
rect 7331 6069 7340 6103
rect 7288 6060 7340 6069
rect 9956 6060 10008 6112
rect 11612 6060 11664 6112
rect 12072 6103 12124 6112
rect 12072 6069 12081 6103
rect 12081 6069 12115 6103
rect 12115 6069 12124 6103
rect 12072 6060 12124 6069
rect 13912 6103 13964 6112
rect 13912 6069 13921 6103
rect 13921 6069 13955 6103
rect 13955 6069 13964 6103
rect 13912 6060 13964 6069
rect 14004 6060 14056 6112
rect 14648 6060 14700 6112
rect 15200 6060 15252 6112
rect 16396 6060 16448 6112
rect 20444 6103 20496 6112
rect 20444 6069 20453 6103
rect 20453 6069 20487 6103
rect 20487 6069 20496 6103
rect 20444 6060 20496 6069
rect 20904 6060 20956 6112
rect 26056 6128 26108 6180
rect 33048 6239 33100 6248
rect 33048 6205 33057 6239
rect 33057 6205 33091 6239
rect 33091 6205 33100 6239
rect 33048 6196 33100 6205
rect 24952 6103 25004 6112
rect 24952 6069 24961 6103
rect 24961 6069 24995 6103
rect 24995 6069 25004 6103
rect 24952 6060 25004 6069
rect 27620 6060 27672 6112
rect 28356 6060 28408 6112
rect 33232 6060 33284 6112
rect 34520 6196 34572 6248
rect 36268 6196 36320 6248
rect 36268 6060 36320 6112
rect 36728 6103 36780 6112
rect 36728 6069 36737 6103
rect 36737 6069 36771 6103
rect 36771 6069 36780 6103
rect 36728 6060 36780 6069
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 65654 5958 65706 6010
rect 65718 5958 65770 6010
rect 65782 5958 65834 6010
rect 65846 5958 65898 6010
rect 65910 5958 65962 6010
rect 2780 5856 2832 5908
rect 3240 5899 3292 5908
rect 3240 5865 3249 5899
rect 3249 5865 3283 5899
rect 3283 5865 3292 5899
rect 9036 5899 9088 5908
rect 3240 5856 3292 5865
rect 5816 5788 5868 5840
rect 8116 5788 8168 5840
rect 9036 5865 9045 5899
rect 9045 5865 9079 5899
rect 9079 5865 9088 5899
rect 9036 5856 9088 5865
rect 12624 5856 12676 5908
rect 16304 5856 16356 5908
rect 18880 5856 18932 5908
rect 24952 5856 25004 5908
rect 6736 5763 6788 5772
rect 5632 5695 5684 5704
rect 5632 5661 5641 5695
rect 5641 5661 5675 5695
rect 5675 5661 5684 5695
rect 5632 5652 5684 5661
rect 6736 5729 6745 5763
rect 6745 5729 6779 5763
rect 6779 5729 6788 5763
rect 6736 5720 6788 5729
rect 5816 5695 5868 5704
rect 5816 5661 5825 5695
rect 5825 5661 5859 5695
rect 5859 5661 5868 5695
rect 5816 5652 5868 5661
rect 6276 5652 6328 5704
rect 6552 5652 6604 5704
rect 6828 5652 6880 5704
rect 7932 5652 7984 5704
rect 8208 5695 8260 5704
rect 8208 5661 8217 5695
rect 8217 5661 8251 5695
rect 8251 5661 8260 5695
rect 8208 5652 8260 5661
rect 10416 5695 10468 5704
rect 1860 5584 1912 5636
rect 10416 5661 10425 5695
rect 10425 5661 10459 5695
rect 10459 5661 10468 5695
rect 10416 5652 10468 5661
rect 11796 5695 11848 5704
rect 11796 5661 11805 5695
rect 11805 5661 11839 5695
rect 11839 5661 11848 5695
rect 11796 5652 11848 5661
rect 25136 5788 25188 5840
rect 27620 5831 27672 5840
rect 27620 5797 27629 5831
rect 27629 5797 27663 5831
rect 27663 5797 27672 5831
rect 27620 5788 27672 5797
rect 12440 5720 12492 5772
rect 12164 5695 12216 5704
rect 12164 5661 12173 5695
rect 12173 5661 12207 5695
rect 12207 5661 12216 5695
rect 15108 5720 15160 5772
rect 12164 5652 12216 5661
rect 14188 5652 14240 5704
rect 14280 5652 14332 5704
rect 12348 5584 12400 5636
rect 5356 5559 5408 5568
rect 5356 5525 5365 5559
rect 5365 5525 5399 5559
rect 5399 5525 5408 5559
rect 5356 5516 5408 5525
rect 7748 5559 7800 5568
rect 7748 5525 7757 5559
rect 7757 5525 7791 5559
rect 7791 5525 7800 5559
rect 7748 5516 7800 5525
rect 10784 5516 10836 5568
rect 11520 5516 11572 5568
rect 11980 5516 12032 5568
rect 12532 5516 12584 5568
rect 16396 5652 16448 5704
rect 17132 5652 17184 5704
rect 17500 5652 17552 5704
rect 17776 5695 17828 5704
rect 17776 5661 17785 5695
rect 17785 5661 17819 5695
rect 17819 5661 17828 5695
rect 17776 5652 17828 5661
rect 18328 5652 18380 5704
rect 19248 5695 19300 5704
rect 19248 5661 19257 5695
rect 19257 5661 19291 5695
rect 19291 5661 19300 5695
rect 19248 5652 19300 5661
rect 19432 5652 19484 5704
rect 20352 5720 20404 5772
rect 20720 5720 20772 5772
rect 22652 5720 22704 5772
rect 26240 5763 26292 5772
rect 26240 5729 26249 5763
rect 26249 5729 26283 5763
rect 26283 5729 26292 5763
rect 26240 5720 26292 5729
rect 19984 5652 20036 5704
rect 20444 5695 20496 5704
rect 20444 5661 20453 5695
rect 20453 5661 20487 5695
rect 20487 5661 20496 5695
rect 20444 5652 20496 5661
rect 14740 5584 14792 5636
rect 24584 5652 24636 5704
rect 25136 5652 25188 5704
rect 28540 5856 28592 5908
rect 33048 5856 33100 5908
rect 36268 5899 36320 5908
rect 36268 5865 36277 5899
rect 36277 5865 36311 5899
rect 36311 5865 36320 5899
rect 36268 5856 36320 5865
rect 37740 5899 37792 5908
rect 37740 5865 37749 5899
rect 37749 5865 37783 5899
rect 37783 5865 37792 5899
rect 37740 5856 37792 5865
rect 32220 5720 32272 5772
rect 32772 5788 32824 5840
rect 33692 5720 33744 5772
rect 28080 5695 28132 5704
rect 28080 5661 28089 5695
rect 28089 5661 28123 5695
rect 28123 5661 28132 5695
rect 28080 5652 28132 5661
rect 30656 5652 30708 5704
rect 31668 5695 31720 5704
rect 31668 5661 31677 5695
rect 31677 5661 31711 5695
rect 31711 5661 31720 5695
rect 31668 5652 31720 5661
rect 32588 5652 32640 5704
rect 32864 5695 32916 5704
rect 32864 5661 32873 5695
rect 32873 5661 32907 5695
rect 32907 5661 32916 5695
rect 33140 5695 33192 5704
rect 32864 5652 32916 5661
rect 33140 5661 33149 5695
rect 33149 5661 33183 5695
rect 33183 5661 33192 5695
rect 33140 5652 33192 5661
rect 20720 5584 20772 5636
rect 26516 5627 26568 5636
rect 26516 5593 26550 5627
rect 26550 5593 26568 5627
rect 34060 5652 34112 5704
rect 36268 5695 36320 5704
rect 36268 5661 36277 5695
rect 36277 5661 36311 5695
rect 36311 5661 36320 5695
rect 36268 5652 36320 5661
rect 36452 5695 36504 5704
rect 36452 5661 36461 5695
rect 36461 5661 36495 5695
rect 36495 5661 36504 5695
rect 36452 5652 36504 5661
rect 68100 5695 68152 5704
rect 26516 5584 26568 5593
rect 36176 5584 36228 5636
rect 68100 5661 68109 5695
rect 68109 5661 68143 5695
rect 68143 5661 68152 5695
rect 68100 5652 68152 5661
rect 20444 5516 20496 5568
rect 25964 5516 26016 5568
rect 32772 5516 32824 5568
rect 32864 5516 32916 5568
rect 34060 5516 34112 5568
rect 34704 5516 34756 5568
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 50294 5414 50346 5466
rect 50358 5414 50410 5466
rect 50422 5414 50474 5466
rect 50486 5414 50538 5466
rect 50550 5414 50602 5466
rect 1860 5355 1912 5364
rect 1860 5321 1869 5355
rect 1869 5321 1903 5355
rect 1903 5321 1912 5355
rect 1860 5312 1912 5321
rect 3516 5355 3568 5364
rect 3516 5321 3525 5355
rect 3525 5321 3559 5355
rect 3559 5321 3568 5355
rect 3516 5312 3568 5321
rect 5816 5312 5868 5364
rect 8208 5312 8260 5364
rect 3240 5244 3292 5296
rect 2044 5108 2096 5160
rect 2320 5219 2372 5228
rect 2320 5185 2329 5219
rect 2329 5185 2363 5219
rect 2363 5185 2372 5219
rect 2320 5176 2372 5185
rect 2504 5219 2556 5228
rect 2504 5185 2513 5219
rect 2513 5185 2547 5219
rect 2547 5185 2556 5219
rect 5356 5244 5408 5296
rect 6460 5244 6512 5296
rect 9680 5312 9732 5364
rect 9772 5312 9824 5364
rect 10968 5312 11020 5364
rect 11612 5312 11664 5364
rect 13268 5312 13320 5364
rect 14372 5312 14424 5364
rect 14740 5312 14792 5364
rect 15476 5312 15528 5364
rect 19340 5312 19392 5364
rect 20260 5312 20312 5364
rect 20812 5355 20864 5364
rect 20812 5321 20821 5355
rect 20821 5321 20855 5355
rect 20855 5321 20864 5355
rect 20812 5312 20864 5321
rect 22836 5312 22888 5364
rect 24216 5312 24268 5364
rect 26516 5312 26568 5364
rect 31116 5312 31168 5364
rect 34796 5312 34848 5364
rect 36176 5355 36228 5364
rect 36176 5321 36185 5355
rect 36185 5321 36219 5355
rect 36219 5321 36228 5355
rect 36176 5312 36228 5321
rect 2504 5176 2556 5185
rect 2412 5108 2464 5160
rect 3424 5108 3476 5160
rect 7840 5176 7892 5228
rect 8484 5219 8536 5228
rect 8484 5185 8493 5219
rect 8493 5185 8527 5219
rect 8527 5185 8536 5219
rect 8484 5176 8536 5185
rect 9128 5219 9180 5228
rect 8392 5108 8444 5160
rect 9128 5185 9137 5219
rect 9137 5185 9171 5219
rect 9171 5185 9180 5219
rect 9128 5176 9180 5185
rect 11704 5219 11756 5228
rect 11704 5185 11713 5219
rect 11713 5185 11747 5219
rect 11747 5185 11756 5219
rect 11704 5176 11756 5185
rect 11980 5219 12032 5228
rect 11980 5185 11989 5219
rect 11989 5185 12023 5219
rect 12023 5185 12032 5219
rect 11980 5176 12032 5185
rect 12164 5176 12216 5228
rect 12256 5219 12308 5228
rect 12256 5185 12265 5219
rect 12265 5185 12299 5219
rect 12299 5185 12308 5219
rect 14280 5244 14332 5296
rect 16764 5287 16816 5296
rect 16764 5253 16773 5287
rect 16773 5253 16807 5287
rect 16807 5253 16816 5287
rect 16764 5244 16816 5253
rect 12256 5176 12308 5185
rect 13452 5219 13504 5228
rect 13452 5185 13461 5219
rect 13461 5185 13495 5219
rect 13495 5185 13504 5219
rect 13452 5176 13504 5185
rect 14372 5219 14424 5228
rect 14372 5185 14381 5219
rect 14381 5185 14415 5219
rect 14415 5185 14424 5219
rect 14372 5176 14424 5185
rect 15108 5219 15160 5228
rect 15108 5185 15117 5219
rect 15117 5185 15151 5219
rect 15151 5185 15160 5219
rect 15108 5176 15160 5185
rect 9588 5151 9640 5160
rect 3056 5015 3108 5024
rect 3056 4981 3065 5015
rect 3065 4981 3099 5015
rect 3099 4981 3108 5015
rect 3056 4972 3108 4981
rect 6460 4972 6512 5024
rect 9128 5015 9180 5024
rect 9128 4981 9137 5015
rect 9137 4981 9171 5015
rect 9171 4981 9180 5015
rect 9128 4972 9180 4981
rect 9588 5117 9597 5151
rect 9597 5117 9631 5151
rect 9631 5117 9640 5151
rect 9588 5108 9640 5117
rect 11704 5040 11756 5092
rect 12532 5108 12584 5160
rect 12716 5108 12768 5160
rect 13084 5108 13136 5160
rect 14096 5108 14148 5160
rect 17592 5176 17644 5228
rect 17408 5108 17460 5160
rect 9864 4972 9916 5024
rect 10508 4972 10560 5024
rect 16580 5040 16632 5092
rect 14280 4972 14332 5024
rect 18512 5244 18564 5296
rect 19708 5244 19760 5296
rect 20444 5244 20496 5296
rect 24768 5287 24820 5296
rect 19984 5176 20036 5228
rect 24768 5253 24777 5287
rect 24777 5253 24811 5287
rect 24811 5253 24820 5287
rect 24768 5244 24820 5253
rect 28080 5244 28132 5296
rect 28540 5287 28592 5296
rect 28540 5253 28549 5287
rect 28549 5253 28583 5287
rect 28583 5253 28592 5287
rect 28540 5244 28592 5253
rect 29644 5244 29696 5296
rect 30288 5244 30340 5296
rect 19432 5108 19484 5160
rect 22100 5176 22152 5228
rect 22652 5219 22704 5228
rect 22652 5185 22661 5219
rect 22661 5185 22695 5219
rect 22695 5185 22704 5219
rect 22652 5176 22704 5185
rect 22928 5219 22980 5228
rect 22928 5185 22962 5219
rect 22962 5185 22980 5219
rect 22928 5176 22980 5185
rect 25136 5176 25188 5228
rect 25688 5176 25740 5228
rect 25964 5219 26016 5228
rect 25964 5185 25973 5219
rect 25973 5185 26007 5219
rect 26007 5185 26016 5219
rect 25964 5176 26016 5185
rect 18144 5040 18196 5092
rect 18880 4972 18932 5024
rect 19340 5040 19392 5092
rect 21088 5108 21140 5160
rect 26148 5219 26200 5228
rect 26148 5185 26157 5219
rect 26157 5185 26191 5219
rect 26191 5185 26200 5219
rect 26148 5176 26200 5185
rect 27804 5176 27856 5228
rect 33232 5219 33284 5228
rect 33232 5185 33241 5219
rect 33241 5185 33275 5219
rect 33275 5185 33284 5219
rect 33232 5176 33284 5185
rect 36728 5244 36780 5296
rect 34704 5219 34756 5228
rect 34704 5185 34713 5219
rect 34713 5185 34747 5219
rect 34747 5185 34756 5219
rect 34704 5176 34756 5185
rect 36176 5219 36228 5228
rect 36176 5185 36177 5219
rect 36177 5185 36211 5219
rect 36211 5185 36228 5219
rect 36176 5176 36228 5185
rect 36268 5176 36320 5228
rect 26332 5108 26384 5160
rect 29920 5108 29972 5160
rect 30564 5151 30616 5160
rect 30564 5117 30573 5151
rect 30573 5117 30607 5151
rect 30607 5117 30616 5151
rect 30564 5108 30616 5117
rect 58808 5108 58860 5160
rect 20812 5040 20864 5092
rect 25780 5040 25832 5092
rect 59268 5040 59320 5092
rect 19984 4972 20036 5024
rect 24860 4972 24912 5024
rect 28816 4972 28868 5024
rect 34612 4972 34664 5024
rect 58716 4972 58768 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 65654 4870 65706 4922
rect 65718 4870 65770 4922
rect 65782 4870 65834 4922
rect 65846 4870 65898 4922
rect 65910 4870 65962 4922
rect 2320 4768 2372 4820
rect 3976 4768 4028 4820
rect 5632 4768 5684 4820
rect 8392 4811 8444 4820
rect 8392 4777 8401 4811
rect 8401 4777 8435 4811
rect 8435 4777 8444 4811
rect 8392 4768 8444 4777
rect 9772 4768 9824 4820
rect 10600 4768 10652 4820
rect 11244 4768 11296 4820
rect 12164 4768 12216 4820
rect 14096 4811 14148 4820
rect 14096 4777 14105 4811
rect 14105 4777 14139 4811
rect 14139 4777 14148 4811
rect 14096 4768 14148 4777
rect 11612 4700 11664 4752
rect 1768 4607 1820 4616
rect 1768 4573 1777 4607
rect 1777 4573 1811 4607
rect 1811 4573 1820 4607
rect 1768 4564 1820 4573
rect 2228 4632 2280 4684
rect 5724 4632 5776 4684
rect 3148 4496 3200 4548
rect 3976 4496 4028 4548
rect 6644 4496 6696 4548
rect 6920 4564 6972 4616
rect 7748 4564 7800 4616
rect 11152 4632 11204 4684
rect 10324 4607 10376 4616
rect 2320 4428 2372 4480
rect 5540 4428 5592 4480
rect 9772 4471 9824 4480
rect 9772 4437 9781 4471
rect 9781 4437 9815 4471
rect 9815 4437 9824 4471
rect 9772 4428 9824 4437
rect 10324 4573 10333 4607
rect 10333 4573 10367 4607
rect 10367 4573 10376 4607
rect 10324 4564 10376 4573
rect 11244 4564 11296 4616
rect 12256 4700 12308 4752
rect 12072 4675 12124 4684
rect 12072 4641 12081 4675
rect 12081 4641 12115 4675
rect 12115 4641 12124 4675
rect 12072 4632 12124 4641
rect 12532 4632 12584 4684
rect 18052 4700 18104 4752
rect 21272 4768 21324 4820
rect 22192 4768 22244 4820
rect 22928 4811 22980 4820
rect 18604 4700 18656 4752
rect 22560 4700 22612 4752
rect 11980 4607 12032 4616
rect 11980 4573 11989 4607
rect 11989 4573 12023 4607
rect 12023 4573 12032 4607
rect 11980 4564 12032 4573
rect 12348 4607 12400 4616
rect 12348 4573 12357 4607
rect 12357 4573 12391 4607
rect 12391 4573 12400 4607
rect 12348 4564 12400 4573
rect 10140 4496 10192 4548
rect 10876 4496 10928 4548
rect 11888 4496 11940 4548
rect 13728 4564 13780 4616
rect 16672 4632 16724 4684
rect 17408 4632 17460 4684
rect 17868 4607 17920 4616
rect 11336 4428 11388 4480
rect 11980 4428 12032 4480
rect 12532 4471 12584 4480
rect 12532 4437 12541 4471
rect 12541 4437 12575 4471
rect 12575 4437 12584 4471
rect 12532 4428 12584 4437
rect 13268 4428 13320 4480
rect 15200 4539 15252 4548
rect 15200 4505 15218 4539
rect 15218 4505 15252 4539
rect 15200 4496 15252 4505
rect 16580 4496 16632 4548
rect 16764 4428 16816 4480
rect 17040 4428 17092 4480
rect 17592 4496 17644 4548
rect 17868 4573 17877 4607
rect 17877 4573 17911 4607
rect 17911 4573 17920 4607
rect 17868 4564 17920 4573
rect 19156 4632 19208 4684
rect 19064 4564 19116 4616
rect 19340 4607 19392 4616
rect 19340 4573 19349 4607
rect 19349 4573 19383 4607
rect 19383 4573 19392 4607
rect 19340 4564 19392 4573
rect 19432 4564 19484 4616
rect 19708 4564 19760 4616
rect 19984 4607 20036 4616
rect 19984 4573 19993 4607
rect 19993 4573 20027 4607
rect 20027 4573 20036 4607
rect 19984 4564 20036 4573
rect 22192 4564 22244 4616
rect 22928 4777 22937 4811
rect 22937 4777 22971 4811
rect 22971 4777 22980 4811
rect 22928 4768 22980 4777
rect 23848 4811 23900 4820
rect 23848 4777 23857 4811
rect 23857 4777 23891 4811
rect 23891 4777 23900 4811
rect 23848 4768 23900 4777
rect 24584 4768 24636 4820
rect 25044 4768 25096 4820
rect 28724 4768 28776 4820
rect 20536 4496 20588 4548
rect 20168 4428 20220 4480
rect 22192 4428 22244 4480
rect 22836 4564 22888 4616
rect 24584 4564 24636 4616
rect 24860 4607 24912 4616
rect 24860 4573 24869 4607
rect 24869 4573 24903 4607
rect 24903 4573 24912 4607
rect 25596 4632 25648 4684
rect 28172 4700 28224 4752
rect 28264 4700 28316 4752
rect 28632 4700 28684 4752
rect 30288 4768 30340 4820
rect 36452 4768 36504 4820
rect 24860 4564 24912 4573
rect 25688 4607 25740 4616
rect 25688 4573 25697 4607
rect 25697 4573 25731 4607
rect 25731 4573 25740 4607
rect 25688 4564 25740 4573
rect 25872 4607 25924 4616
rect 25872 4573 25881 4607
rect 25881 4573 25915 4607
rect 25915 4573 25924 4607
rect 25872 4564 25924 4573
rect 27804 4607 27856 4616
rect 24400 4471 24452 4480
rect 24400 4437 24409 4471
rect 24409 4437 24443 4471
rect 24443 4437 24452 4471
rect 24400 4428 24452 4437
rect 24676 4428 24728 4480
rect 25780 4496 25832 4548
rect 27804 4573 27813 4607
rect 27813 4573 27847 4607
rect 27847 4573 27856 4607
rect 32128 4700 32180 4752
rect 36268 4700 36320 4752
rect 57244 4700 57296 4752
rect 58256 4700 58308 4752
rect 28908 4632 28960 4684
rect 27804 4564 27856 4573
rect 28816 4607 28868 4616
rect 28816 4573 28825 4607
rect 28825 4573 28859 4607
rect 28859 4573 28868 4607
rect 28816 4564 28868 4573
rect 29000 4607 29052 4616
rect 29000 4573 29009 4607
rect 29009 4573 29043 4607
rect 29043 4573 29052 4607
rect 29000 4564 29052 4573
rect 29736 4607 29788 4616
rect 29736 4573 29745 4607
rect 29745 4573 29779 4607
rect 29779 4573 29788 4607
rect 29736 4564 29788 4573
rect 29920 4607 29972 4616
rect 29920 4573 29929 4607
rect 29929 4573 29963 4607
rect 29963 4573 29972 4607
rect 29920 4564 29972 4573
rect 32588 4564 32640 4616
rect 36176 4632 36228 4684
rect 34520 4564 34572 4616
rect 58900 4632 58952 4684
rect 36912 4607 36964 4616
rect 36912 4573 36921 4607
rect 36921 4573 36955 4607
rect 36955 4573 36964 4607
rect 36912 4564 36964 4573
rect 57152 4564 57204 4616
rect 57612 4564 57664 4616
rect 27252 4496 27304 4548
rect 30288 4428 30340 4480
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 50294 4326 50346 4378
rect 50358 4326 50410 4378
rect 50422 4326 50474 4378
rect 50486 4326 50538 4378
rect 50550 4326 50602 4378
rect 2136 4131 2188 4140
rect 2136 4097 2145 4131
rect 2145 4097 2179 4131
rect 2179 4097 2188 4131
rect 2136 4088 2188 4097
rect 2412 4156 2464 4208
rect 2320 4131 2372 4140
rect 2320 4097 2329 4131
rect 2329 4097 2363 4131
rect 2363 4097 2372 4131
rect 2320 4088 2372 4097
rect 2504 4131 2556 4140
rect 2504 4097 2513 4131
rect 2513 4097 2547 4131
rect 2547 4097 2556 4131
rect 3424 4156 3476 4208
rect 5632 4199 5684 4208
rect 5632 4165 5641 4199
rect 5641 4165 5675 4199
rect 5675 4165 5684 4199
rect 5632 4156 5684 4165
rect 6552 4156 6604 4208
rect 2504 4088 2556 4097
rect 4988 4131 5040 4140
rect 4988 4097 4997 4131
rect 4997 4097 5031 4131
rect 5031 4097 5040 4131
rect 4988 4088 5040 4097
rect 6644 4131 6696 4140
rect 6644 4097 6653 4131
rect 6653 4097 6687 4131
rect 6687 4097 6696 4131
rect 6644 4088 6696 4097
rect 6828 4224 6880 4276
rect 9680 4224 9732 4276
rect 10232 4224 10284 4276
rect 11796 4224 11848 4276
rect 12348 4224 12400 4276
rect 8944 4199 8996 4208
rect 8944 4165 8953 4199
rect 8953 4165 8987 4199
rect 8987 4165 8996 4199
rect 8944 4156 8996 4165
rect 7012 4131 7064 4140
rect 7012 4097 7021 4131
rect 7021 4097 7055 4131
rect 7055 4097 7064 4131
rect 7012 4088 7064 4097
rect 8576 4088 8628 4140
rect 9680 4131 9732 4140
rect 9680 4097 9689 4131
rect 9689 4097 9723 4131
rect 9723 4097 9732 4131
rect 9680 4088 9732 4097
rect 9864 4156 9916 4208
rect 10232 4088 10284 4140
rect 10508 4131 10560 4140
rect 10508 4097 10517 4131
rect 10517 4097 10551 4131
rect 10551 4097 10560 4131
rect 10508 4088 10560 4097
rect 12440 4156 12492 4208
rect 12532 4156 12584 4208
rect 17408 4156 17460 4208
rect 22192 4267 22244 4276
rect 22192 4233 22201 4267
rect 22201 4233 22235 4267
rect 22235 4233 22244 4267
rect 22192 4224 22244 4233
rect 22284 4156 22336 4208
rect 24216 4224 24268 4276
rect 24768 4267 24820 4276
rect 24768 4233 24777 4267
rect 24777 4233 24811 4267
rect 24811 4233 24820 4267
rect 24768 4224 24820 4233
rect 25872 4224 25924 4276
rect 29736 4224 29788 4276
rect 23480 4156 23532 4208
rect 24400 4156 24452 4208
rect 25136 4156 25188 4208
rect 11060 4088 11112 4140
rect 12900 4088 12952 4140
rect 5540 3952 5592 4004
rect 12440 4020 12492 4072
rect 13544 4088 13596 4140
rect 13728 4088 13780 4140
rect 13820 4088 13872 4140
rect 14924 4131 14976 4140
rect 14924 4097 14933 4131
rect 14933 4097 14967 4131
rect 14967 4097 14976 4131
rect 14924 4088 14976 4097
rect 16856 4131 16908 4140
rect 16856 4097 16865 4131
rect 16865 4097 16899 4131
rect 16899 4097 16908 4131
rect 16856 4088 16908 4097
rect 16580 4020 16632 4072
rect 17040 4088 17092 4140
rect 17868 4088 17920 4140
rect 18236 4088 18288 4140
rect 7656 3995 7708 4004
rect 7656 3961 7665 3995
rect 7665 3961 7699 3995
rect 7699 3961 7708 3995
rect 7656 3952 7708 3961
rect 7748 3952 7800 4004
rect 2136 3884 2188 3936
rect 4620 3884 4672 3936
rect 6368 3927 6420 3936
rect 6368 3893 6377 3927
rect 6377 3893 6411 3927
rect 6411 3893 6420 3927
rect 6368 3884 6420 3893
rect 6552 3884 6604 3936
rect 7564 3884 7616 3936
rect 8208 3927 8260 3936
rect 8208 3893 8217 3927
rect 8217 3893 8251 3927
rect 8251 3893 8260 3927
rect 8208 3884 8260 3893
rect 10968 3952 11020 4004
rect 11244 3884 11296 3936
rect 13084 3884 13136 3936
rect 15384 3952 15436 4004
rect 18696 4020 18748 4072
rect 17592 3952 17644 4004
rect 19340 4088 19392 4140
rect 19984 4088 20036 4140
rect 20536 4131 20588 4140
rect 20536 4097 20545 4131
rect 20545 4097 20579 4131
rect 20579 4097 20588 4131
rect 20536 4088 20588 4097
rect 20812 4088 20864 4140
rect 21088 4088 21140 4140
rect 22652 4088 22704 4140
rect 20628 4020 20680 4072
rect 20904 3952 20956 4004
rect 13636 3884 13688 3936
rect 14096 3927 14148 3936
rect 14096 3893 14105 3927
rect 14105 3893 14139 3927
rect 14139 3893 14148 3927
rect 14096 3884 14148 3893
rect 16672 3884 16724 3936
rect 17960 3884 18012 3936
rect 18512 3927 18564 3936
rect 18512 3893 18521 3927
rect 18521 3893 18555 3927
rect 18555 3893 18564 3927
rect 18512 3884 18564 3893
rect 19432 3884 19484 3936
rect 19984 3884 20036 3936
rect 20628 3884 20680 3936
rect 26056 4088 26108 4140
rect 26240 4088 26292 4140
rect 27252 4131 27304 4140
rect 27252 4097 27286 4131
rect 27286 4097 27304 4131
rect 27252 4088 27304 4097
rect 28540 4156 28592 4208
rect 30564 4156 30616 4208
rect 32128 4224 32180 4276
rect 30288 4131 30340 4140
rect 30288 4097 30322 4131
rect 30322 4097 30340 4131
rect 30288 4088 30340 4097
rect 34520 4156 34572 4208
rect 36912 4224 36964 4276
rect 57980 4088 58032 4140
rect 34612 4020 34664 4072
rect 59176 4020 59228 4072
rect 57520 3952 57572 4004
rect 58624 3952 58676 4004
rect 30012 3884 30064 3936
rect 56140 3884 56192 3936
rect 56324 3884 56376 3936
rect 56968 3884 57020 3936
rect 58072 3884 58124 3936
rect 67640 3927 67692 3936
rect 67640 3893 67649 3927
rect 67649 3893 67683 3927
rect 67683 3893 67692 3927
rect 67640 3884 67692 3893
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 65654 3782 65706 3834
rect 65718 3782 65770 3834
rect 65782 3782 65834 3834
rect 65846 3782 65898 3834
rect 65910 3782 65962 3834
rect 2228 3723 2280 3732
rect 2228 3689 2237 3723
rect 2237 3689 2271 3723
rect 2271 3689 2280 3723
rect 2228 3680 2280 3689
rect 2504 3680 2556 3732
rect 8208 3680 8260 3732
rect 11336 3680 11388 3732
rect 11612 3723 11664 3732
rect 11612 3689 11621 3723
rect 11621 3689 11655 3723
rect 11655 3689 11664 3723
rect 11612 3680 11664 3689
rect 12440 3680 12492 3732
rect 3424 3408 3476 3460
rect 4160 3383 4212 3392
rect 4160 3349 4169 3383
rect 4169 3349 4203 3383
rect 4203 3349 4212 3383
rect 4160 3340 4212 3349
rect 5632 3340 5684 3392
rect 6368 3408 6420 3460
rect 6920 3476 6972 3528
rect 7564 3544 7616 3596
rect 7748 3476 7800 3528
rect 7840 3519 7892 3528
rect 7840 3485 7849 3519
rect 7849 3485 7883 3519
rect 7883 3485 7892 3519
rect 7840 3476 7892 3485
rect 9036 3476 9088 3528
rect 6736 3408 6788 3460
rect 8576 3408 8628 3460
rect 13452 3612 13504 3664
rect 15108 3655 15160 3664
rect 15108 3621 15117 3655
rect 15117 3621 15151 3655
rect 15151 3621 15160 3655
rect 15108 3612 15160 3621
rect 18236 3680 18288 3732
rect 18420 3680 18472 3732
rect 18696 3680 18748 3732
rect 22376 3680 22428 3732
rect 57796 3680 57848 3732
rect 58072 3680 58124 3732
rect 18144 3612 18196 3664
rect 18512 3612 18564 3664
rect 11060 3544 11112 3596
rect 9588 3519 9640 3528
rect 9588 3485 9597 3519
rect 9597 3485 9631 3519
rect 9631 3485 9640 3519
rect 9588 3476 9640 3485
rect 9864 3519 9916 3528
rect 9864 3485 9898 3519
rect 9898 3485 9916 3519
rect 9864 3476 9916 3485
rect 10692 3476 10744 3528
rect 10876 3476 10928 3528
rect 11612 3476 11664 3528
rect 11888 3476 11940 3528
rect 16580 3544 16632 3596
rect 19432 3587 19484 3596
rect 12992 3476 13044 3528
rect 13360 3476 13412 3528
rect 12624 3451 12676 3460
rect 12624 3417 12633 3451
rect 12633 3417 12667 3451
rect 12667 3417 12676 3451
rect 12624 3408 12676 3417
rect 13452 3408 13504 3460
rect 15384 3476 15436 3528
rect 15844 3476 15896 3528
rect 16304 3519 16356 3528
rect 16304 3485 16313 3519
rect 16313 3485 16347 3519
rect 16347 3485 16356 3519
rect 16304 3476 16356 3485
rect 19432 3553 19441 3587
rect 19441 3553 19475 3587
rect 19475 3553 19484 3587
rect 19432 3544 19484 3553
rect 20076 3612 20128 3664
rect 41144 3612 41196 3664
rect 56508 3612 56560 3664
rect 58348 3612 58400 3664
rect 55772 3544 55824 3596
rect 56784 3544 56836 3596
rect 58992 3544 59044 3596
rect 16856 3519 16908 3528
rect 15752 3408 15804 3460
rect 16856 3485 16865 3519
rect 16865 3485 16899 3519
rect 16899 3485 16908 3519
rect 16856 3476 16908 3485
rect 17040 3476 17092 3528
rect 17592 3476 17644 3528
rect 16764 3408 16816 3460
rect 20168 3476 20220 3528
rect 20444 3476 20496 3528
rect 21548 3476 21600 3528
rect 22376 3476 22428 3528
rect 23480 3476 23532 3528
rect 24308 3476 24360 3528
rect 25136 3476 25188 3528
rect 25964 3476 26016 3528
rect 26792 3476 26844 3528
rect 27620 3476 27672 3528
rect 28724 3476 28776 3528
rect 29828 3476 29880 3528
rect 30656 3476 30708 3528
rect 31484 3476 31536 3528
rect 32312 3476 32364 3528
rect 33140 3476 33192 3528
rect 39212 3476 39264 3528
rect 40040 3476 40092 3528
rect 40868 3476 40920 3528
rect 42524 3476 42576 3528
rect 43076 3476 43128 3528
rect 45008 3476 45060 3528
rect 45284 3476 45336 3528
rect 46112 3476 46164 3528
rect 46940 3476 46992 3528
rect 47768 3476 47820 3528
rect 48872 3476 48924 3528
rect 50160 3476 50212 3528
rect 50804 3476 50856 3528
rect 51356 3476 51408 3528
rect 52736 3476 52788 3528
rect 53012 3476 53064 3528
rect 54668 3476 54720 3528
rect 55496 3476 55548 3528
rect 56232 3476 56284 3528
rect 57336 3476 57388 3528
rect 60464 3519 60516 3528
rect 60464 3485 60473 3519
rect 60473 3485 60507 3519
rect 60507 3485 60516 3519
rect 60464 3476 60516 3485
rect 19432 3408 19484 3460
rect 19984 3451 20036 3460
rect 19984 3417 19993 3451
rect 19993 3417 20027 3451
rect 20027 3417 20036 3451
rect 19984 3408 20036 3417
rect 7380 3340 7432 3392
rect 7748 3340 7800 3392
rect 10692 3340 10744 3392
rect 11060 3340 11112 3392
rect 11244 3340 11296 3392
rect 12256 3340 12308 3392
rect 13636 3340 13688 3392
rect 14188 3340 14240 3392
rect 19248 3383 19300 3392
rect 19248 3349 19257 3383
rect 19257 3349 19291 3383
rect 19291 3349 19300 3383
rect 19248 3340 19300 3349
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 50294 3238 50346 3290
rect 50358 3238 50410 3290
rect 50422 3238 50474 3290
rect 50486 3238 50538 3290
rect 50550 3238 50602 3290
rect 4160 3000 4212 3052
rect 7748 3136 7800 3188
rect 7840 3136 7892 3188
rect 8576 3136 8628 3188
rect 10416 3179 10468 3188
rect 6736 3000 6788 3052
rect 6920 3000 6972 3052
rect 7840 3000 7892 3052
rect 9588 3068 9640 3120
rect 10416 3145 10425 3179
rect 10425 3145 10459 3179
rect 10459 3145 10468 3179
rect 10416 3136 10468 3145
rect 12440 3136 12492 3188
rect 14924 3179 14976 3188
rect 11244 3068 11296 3120
rect 9128 3000 9180 3052
rect 13268 3068 13320 3120
rect 4896 2932 4948 2984
rect 5632 2864 5684 2916
rect 5908 2864 5960 2916
rect 6460 2907 6512 2916
rect 6460 2873 6469 2907
rect 6469 2873 6503 2907
rect 6503 2873 6512 2907
rect 6460 2864 6512 2873
rect 6736 2864 6788 2916
rect 12256 3043 12308 3052
rect 12256 3009 12265 3043
rect 12265 3009 12299 3043
rect 12299 3009 12308 3043
rect 12256 3000 12308 3009
rect 13544 3043 13596 3052
rect 10416 2932 10468 2984
rect 13544 3009 13553 3043
rect 13553 3009 13587 3043
rect 13587 3009 13596 3043
rect 13544 3000 13596 3009
rect 13912 3068 13964 3120
rect 14924 3145 14933 3179
rect 14933 3145 14967 3179
rect 14967 3145 14976 3179
rect 14924 3136 14976 3145
rect 15660 3136 15712 3188
rect 20076 3136 20128 3188
rect 20536 3136 20588 3188
rect 55956 3136 56008 3188
rect 58072 3136 58124 3188
rect 16396 3068 16448 3120
rect 14372 3000 14424 3052
rect 14924 3000 14976 3052
rect 15200 3000 15252 3052
rect 17316 3000 17368 3052
rect 57704 3068 57756 3120
rect 60464 3068 60516 3120
rect 21732 3000 21784 3052
rect 58164 3000 58216 3052
rect 12716 2932 12768 2984
rect 19984 2932 20036 2984
rect 20168 2932 20220 2984
rect 21824 2932 21876 2984
rect 37280 2932 37332 2984
rect 44732 2932 44784 2984
rect 48596 2932 48648 2984
rect 52460 2932 52512 2984
rect 53564 2932 53616 2984
rect 55220 2932 55272 2984
rect 56692 2932 56744 2984
rect 12072 2796 12124 2848
rect 12532 2796 12584 2848
rect 13912 2796 13964 2848
rect 16764 2864 16816 2916
rect 38384 2864 38436 2916
rect 39764 2864 39816 2916
rect 42248 2864 42300 2916
rect 43628 2864 43680 2916
rect 47492 2864 47544 2916
rect 49424 2864 49476 2916
rect 50620 2864 50672 2916
rect 53288 2864 53340 2916
rect 54392 2864 54444 2916
rect 55680 2864 55732 2916
rect 57060 2864 57112 2916
rect 58440 2932 58492 2984
rect 17040 2796 17092 2848
rect 20260 2796 20312 2848
rect 20996 2796 21048 2848
rect 22652 2796 22704 2848
rect 22928 2796 22980 2848
rect 24032 2796 24084 2848
rect 24860 2796 24912 2848
rect 25412 2796 25464 2848
rect 26240 2796 26292 2848
rect 27068 2796 27120 2848
rect 27896 2796 27948 2848
rect 28448 2796 28500 2848
rect 29276 2796 29328 2848
rect 30104 2796 30156 2848
rect 30380 2796 30432 2848
rect 31208 2796 31260 2848
rect 32036 2796 32088 2848
rect 32864 2839 32916 2848
rect 32864 2805 32873 2839
rect 32873 2805 32907 2839
rect 32907 2805 32916 2839
rect 32864 2796 32916 2805
rect 33692 2796 33744 2848
rect 34244 2796 34296 2848
rect 34520 2796 34572 2848
rect 35348 2796 35400 2848
rect 36176 2796 36228 2848
rect 36728 2796 36780 2848
rect 37832 2796 37884 2848
rect 38936 2796 38988 2848
rect 40316 2796 40368 2848
rect 41696 2796 41748 2848
rect 42800 2796 42852 2848
rect 44180 2796 44232 2848
rect 45560 2796 45612 2848
rect 46664 2796 46716 2848
rect 48044 2796 48096 2848
rect 49976 2796 50028 2848
rect 51908 2796 51960 2848
rect 53840 2796 53892 2848
rect 55404 2796 55456 2848
rect 56048 2796 56100 2848
rect 59360 2864 59412 2916
rect 59452 2796 59504 2848
rect 60464 2839 60516 2848
rect 60464 2805 60473 2839
rect 60473 2805 60507 2839
rect 60507 2805 60516 2839
rect 60464 2796 60516 2805
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 65654 2694 65706 2746
rect 65718 2694 65770 2746
rect 65782 2694 65834 2746
rect 65846 2694 65898 2746
rect 65910 2694 65962 2746
rect 7840 2635 7892 2644
rect 7840 2601 7849 2635
rect 7849 2601 7883 2635
rect 7883 2601 7892 2635
rect 7840 2592 7892 2601
rect 9496 2592 9548 2644
rect 11980 2592 12032 2644
rect 12072 2635 12124 2644
rect 12072 2601 12081 2635
rect 12081 2601 12115 2635
rect 12115 2601 12124 2635
rect 12256 2635 12308 2644
rect 12072 2592 12124 2601
rect 12256 2601 12265 2635
rect 12265 2601 12299 2635
rect 12299 2601 12308 2635
rect 12256 2592 12308 2601
rect 16856 2635 16908 2644
rect 12716 2524 12768 2576
rect 4896 2431 4948 2440
rect 4896 2397 4905 2431
rect 4905 2397 4939 2431
rect 4939 2397 4948 2431
rect 4896 2388 4948 2397
rect 6736 2456 6788 2508
rect 6736 2363 6788 2372
rect 4436 2295 4488 2304
rect 4436 2261 4445 2295
rect 4445 2261 4479 2295
rect 4479 2261 4488 2295
rect 4436 2252 4488 2261
rect 5080 2295 5132 2304
rect 5080 2261 5089 2295
rect 5089 2261 5123 2295
rect 5123 2261 5132 2295
rect 5080 2252 5132 2261
rect 5724 2295 5776 2304
rect 5724 2261 5733 2295
rect 5733 2261 5767 2295
rect 5767 2261 5776 2295
rect 5724 2252 5776 2261
rect 6736 2329 6745 2363
rect 6745 2329 6779 2363
rect 6779 2329 6788 2363
rect 6736 2320 6788 2329
rect 7012 2388 7064 2440
rect 7380 2431 7432 2440
rect 7380 2397 7389 2431
rect 7389 2397 7423 2431
rect 7423 2397 7432 2431
rect 7380 2388 7432 2397
rect 11520 2456 11572 2508
rect 7564 2431 7616 2440
rect 7564 2397 7573 2431
rect 7573 2397 7607 2431
rect 7607 2397 7616 2431
rect 9496 2431 9548 2440
rect 7564 2388 7616 2397
rect 9496 2397 9505 2431
rect 9505 2397 9539 2431
rect 9539 2397 9548 2431
rect 9496 2388 9548 2397
rect 9588 2388 9640 2440
rect 10232 2431 10284 2440
rect 10232 2397 10241 2431
rect 10241 2397 10275 2431
rect 10275 2397 10284 2431
rect 10232 2388 10284 2397
rect 10416 2388 10468 2440
rect 10508 2320 10560 2372
rect 12624 2388 12676 2440
rect 12992 2524 13044 2576
rect 12164 2320 12216 2372
rect 14372 2524 14424 2576
rect 14740 2524 14792 2576
rect 16856 2601 16865 2635
rect 16865 2601 16899 2635
rect 16899 2601 16908 2635
rect 16856 2592 16908 2601
rect 17592 2635 17644 2644
rect 17592 2601 17601 2635
rect 17601 2601 17635 2635
rect 17635 2601 17644 2635
rect 17592 2592 17644 2601
rect 18236 2635 18288 2644
rect 18236 2601 18245 2635
rect 18245 2601 18279 2635
rect 18279 2601 18288 2635
rect 18236 2592 18288 2601
rect 17132 2524 17184 2576
rect 14464 2456 14516 2508
rect 14556 2388 14608 2440
rect 14924 2388 14976 2440
rect 15200 2320 15252 2372
rect 9588 2252 9640 2304
rect 10048 2295 10100 2304
rect 10048 2261 10057 2295
rect 10057 2261 10091 2295
rect 10091 2261 10100 2295
rect 10048 2252 10100 2261
rect 12256 2252 12308 2304
rect 14464 2252 14516 2304
rect 14740 2252 14792 2304
rect 15660 2295 15712 2304
rect 15660 2261 15669 2295
rect 15669 2261 15703 2295
rect 15703 2261 15712 2295
rect 21272 2524 21324 2576
rect 21732 2592 21784 2644
rect 23112 2592 23164 2644
rect 55220 2592 55272 2644
rect 57428 2592 57480 2644
rect 23204 2524 23256 2576
rect 29000 2524 29052 2576
rect 30932 2524 30984 2576
rect 40592 2524 40644 2576
rect 44456 2524 44508 2576
rect 48320 2524 48372 2576
rect 52184 2524 52236 2576
rect 55864 2524 55916 2576
rect 58072 2524 58124 2576
rect 18236 2456 18288 2508
rect 18420 2431 18472 2440
rect 18420 2397 18429 2431
rect 18429 2397 18463 2431
rect 18463 2397 18472 2431
rect 18420 2388 18472 2397
rect 20720 2388 20772 2440
rect 22100 2388 22152 2440
rect 23756 2388 23808 2440
rect 24584 2388 24636 2440
rect 26516 2456 26568 2508
rect 37004 2456 37056 2508
rect 38108 2456 38160 2508
rect 41420 2456 41472 2508
rect 43352 2456 43404 2508
rect 46388 2456 46440 2508
rect 49148 2456 49200 2508
rect 51080 2456 51132 2508
rect 54944 2456 54996 2508
rect 63684 2499 63736 2508
rect 25688 2388 25740 2440
rect 27344 2388 27396 2440
rect 28172 2388 28224 2440
rect 29552 2388 29604 2440
rect 32588 2388 32640 2440
rect 33416 2388 33468 2440
rect 33968 2388 34020 2440
rect 34796 2388 34848 2440
rect 35072 2388 35124 2440
rect 35624 2388 35676 2440
rect 35900 2388 35952 2440
rect 36452 2388 36504 2440
rect 37556 2388 37608 2440
rect 38660 2388 38712 2440
rect 19340 2295 19392 2304
rect 15660 2252 15712 2261
rect 19340 2261 19349 2295
rect 19349 2261 19383 2295
rect 19383 2261 19392 2295
rect 19340 2252 19392 2261
rect 31760 2320 31812 2372
rect 39488 2320 39540 2372
rect 41972 2388 42024 2440
rect 43904 2320 43956 2372
rect 45836 2388 45888 2440
rect 47216 2320 47268 2372
rect 49700 2388 49752 2440
rect 51632 2388 51684 2440
rect 54116 2320 54168 2372
rect 56416 2388 56468 2440
rect 27712 2252 27764 2304
rect 56876 2252 56928 2304
rect 63684 2465 63693 2499
rect 63693 2465 63727 2499
rect 63727 2465 63736 2499
rect 63684 2456 63736 2465
rect 61752 2431 61804 2440
rect 61752 2397 61761 2431
rect 61761 2397 61795 2431
rect 61795 2397 61804 2431
rect 61752 2388 61804 2397
rect 63040 2431 63092 2440
rect 63040 2397 63049 2431
rect 63049 2397 63083 2431
rect 63083 2397 63092 2431
rect 63040 2388 63092 2397
rect 67640 2431 67692 2440
rect 67640 2397 67649 2431
rect 67649 2397 67683 2431
rect 67683 2397 67692 2431
rect 67640 2388 67692 2397
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 50294 2150 50346 2202
rect 50358 2150 50410 2202
rect 50422 2150 50474 2202
rect 50486 2150 50538 2202
rect 50550 2150 50602 2202
rect 4436 2048 4488 2100
rect 12624 2048 12676 2100
rect 14556 2048 14608 2100
rect 20352 2048 20404 2100
rect 58072 2048 58124 2100
rect 61752 2048 61804 2100
rect 5080 1980 5132 2032
rect 10140 1980 10192 2032
rect 12072 1980 12124 2032
rect 5632 1912 5684 1964
rect 10232 1912 10284 1964
rect 12992 1980 13044 2032
rect 59084 1980 59136 2032
rect 63684 1980 63736 2032
rect 12532 1912 12584 1964
rect 15200 1912 15252 1964
rect 58532 1912 58584 1964
rect 63040 1912 63092 1964
rect 12164 1844 12216 1896
rect 19248 1844 19300 1896
rect 13544 1776 13596 1828
rect 15384 1776 15436 1828
rect 4896 1708 4948 1760
rect 10876 1708 10928 1760
rect 11980 1708 12032 1760
rect 18420 1708 18472 1760
rect 19340 1708 19392 1760
rect 19800 1708 19852 1760
rect 7564 1640 7616 1692
rect 12808 1640 12860 1692
rect 5724 1572 5776 1624
rect 14280 1572 14332 1624
rect 12256 1504 12308 1556
rect 13360 1504 13412 1556
rect 19708 1504 19760 1556
rect 20076 1504 20128 1556
rect 12072 1436 12124 1488
rect 17040 1436 17092 1488
rect 10324 1368 10376 1420
rect 10968 1368 11020 1420
rect 11796 1368 11848 1420
rect 12256 1368 12308 1420
rect 12532 1368 12584 1420
rect 11152 1300 11204 1352
rect 11428 1300 11480 1352
rect 18512 1368 18564 1420
rect 19248 1368 19300 1420
rect 19524 1368 19576 1420
rect 20628 1368 20680 1420
rect 9588 1164 9640 1216
rect 11152 1164 11204 1216
rect 12900 1164 12952 1216
rect 56784 1164 56836 1216
rect 57060 1164 57112 1216
rect 57060 1028 57112 1080
rect 59452 1028 59504 1080
<< metal2 >>
rect 4342 59200 4398 60000
rect 13082 59200 13138 60000
rect 21822 59200 21878 60000
rect 30562 59200 30618 60000
rect 39302 59200 39358 60000
rect 48042 59200 48098 60000
rect 56782 59200 56838 60000
rect 65522 59200 65578 60000
rect 4356 57458 4384 59200
rect 13096 57458 13124 59200
rect 21836 57882 21864 59200
rect 21836 57854 22140 57882
rect 19574 57692 19882 57701
rect 19574 57690 19580 57692
rect 19636 57690 19660 57692
rect 19716 57690 19740 57692
rect 19796 57690 19820 57692
rect 19876 57690 19882 57692
rect 19636 57638 19638 57690
rect 19818 57638 19820 57690
rect 19574 57636 19580 57638
rect 19636 57636 19660 57638
rect 19716 57636 19740 57638
rect 19796 57636 19820 57638
rect 19876 57636 19882 57638
rect 19574 57627 19882 57636
rect 22112 57594 22140 57854
rect 30576 57594 30604 59200
rect 39316 57594 39344 59200
rect 48056 57882 48084 59200
rect 48056 57854 48360 57882
rect 48332 57594 48360 57854
rect 50294 57692 50602 57701
rect 50294 57690 50300 57692
rect 50356 57690 50380 57692
rect 50436 57690 50460 57692
rect 50516 57690 50540 57692
rect 50596 57690 50602 57692
rect 50356 57638 50358 57690
rect 50538 57638 50540 57690
rect 50294 57636 50300 57638
rect 50356 57636 50380 57638
rect 50436 57636 50460 57638
rect 50516 57636 50540 57638
rect 50596 57636 50602 57638
rect 50294 57627 50602 57636
rect 56796 57594 56824 59200
rect 65536 57594 65564 59200
rect 67638 57624 67694 57633
rect 22100 57588 22152 57594
rect 22100 57530 22152 57536
rect 30564 57588 30616 57594
rect 30564 57530 30616 57536
rect 39304 57588 39356 57594
rect 39304 57530 39356 57536
rect 48320 57588 48372 57594
rect 48320 57530 48372 57536
rect 56784 57588 56836 57594
rect 56784 57530 56836 57536
rect 65524 57588 65576 57594
rect 67638 57559 67694 57568
rect 65524 57530 65576 57536
rect 36820 57520 36872 57526
rect 36820 57462 36872 57468
rect 4344 57452 4396 57458
rect 4344 57394 4396 57400
rect 13084 57452 13136 57458
rect 13084 57394 13136 57400
rect 21640 57452 21692 57458
rect 21640 57394 21692 57400
rect 30104 57452 30156 57458
rect 30104 57394 30156 57400
rect 4214 57148 4522 57157
rect 4214 57146 4220 57148
rect 4276 57146 4300 57148
rect 4356 57146 4380 57148
rect 4436 57146 4460 57148
rect 4516 57146 4522 57148
rect 4276 57094 4278 57146
rect 4458 57094 4460 57146
rect 4214 57092 4220 57094
rect 4276 57092 4300 57094
rect 4356 57092 4380 57094
rect 4436 57092 4460 57094
rect 4516 57092 4522 57094
rect 4214 57083 4522 57092
rect 21652 56710 21680 57394
rect 30116 57254 30144 57394
rect 30104 57248 30156 57254
rect 30104 57190 30156 57196
rect 27160 57044 27212 57050
rect 27160 56986 27212 56992
rect 21640 56704 21692 56710
rect 21640 56646 21692 56652
rect 19574 56604 19882 56613
rect 19574 56602 19580 56604
rect 19636 56602 19660 56604
rect 19716 56602 19740 56604
rect 19796 56602 19820 56604
rect 19876 56602 19882 56604
rect 19636 56550 19638 56602
rect 19818 56550 19820 56602
rect 19574 56548 19580 56550
rect 19636 56548 19660 56550
rect 19716 56548 19740 56550
rect 19796 56548 19820 56550
rect 19876 56548 19882 56550
rect 19574 56539 19882 56548
rect 4214 56060 4522 56069
rect 4214 56058 4220 56060
rect 4276 56058 4300 56060
rect 4356 56058 4380 56060
rect 4436 56058 4460 56060
rect 4516 56058 4522 56060
rect 4276 56006 4278 56058
rect 4458 56006 4460 56058
rect 4214 56004 4220 56006
rect 4276 56004 4300 56006
rect 4356 56004 4380 56006
rect 4436 56004 4460 56006
rect 4516 56004 4522 56006
rect 4214 55995 4522 56004
rect 19574 55516 19882 55525
rect 19574 55514 19580 55516
rect 19636 55514 19660 55516
rect 19716 55514 19740 55516
rect 19796 55514 19820 55516
rect 19876 55514 19882 55516
rect 19636 55462 19638 55514
rect 19818 55462 19820 55514
rect 19574 55460 19580 55462
rect 19636 55460 19660 55462
rect 19716 55460 19740 55462
rect 19796 55460 19820 55462
rect 19876 55460 19882 55462
rect 19574 55451 19882 55460
rect 4214 54972 4522 54981
rect 4214 54970 4220 54972
rect 4276 54970 4300 54972
rect 4356 54970 4380 54972
rect 4436 54970 4460 54972
rect 4516 54970 4522 54972
rect 4276 54918 4278 54970
rect 4458 54918 4460 54970
rect 4214 54916 4220 54918
rect 4276 54916 4300 54918
rect 4356 54916 4380 54918
rect 4436 54916 4460 54918
rect 4516 54916 4522 54918
rect 4214 54907 4522 54916
rect 19574 54428 19882 54437
rect 19574 54426 19580 54428
rect 19636 54426 19660 54428
rect 19716 54426 19740 54428
rect 19796 54426 19820 54428
rect 19876 54426 19882 54428
rect 19636 54374 19638 54426
rect 19818 54374 19820 54426
rect 19574 54372 19580 54374
rect 19636 54372 19660 54374
rect 19716 54372 19740 54374
rect 19796 54372 19820 54374
rect 19876 54372 19882 54374
rect 19574 54363 19882 54372
rect 4214 53884 4522 53893
rect 4214 53882 4220 53884
rect 4276 53882 4300 53884
rect 4356 53882 4380 53884
rect 4436 53882 4460 53884
rect 4516 53882 4522 53884
rect 4276 53830 4278 53882
rect 4458 53830 4460 53882
rect 4214 53828 4220 53830
rect 4276 53828 4300 53830
rect 4356 53828 4380 53830
rect 4436 53828 4460 53830
rect 4516 53828 4522 53830
rect 4214 53819 4522 53828
rect 19574 53340 19882 53349
rect 19574 53338 19580 53340
rect 19636 53338 19660 53340
rect 19716 53338 19740 53340
rect 19796 53338 19820 53340
rect 19876 53338 19882 53340
rect 19636 53286 19638 53338
rect 19818 53286 19820 53338
rect 19574 53284 19580 53286
rect 19636 53284 19660 53286
rect 19716 53284 19740 53286
rect 19796 53284 19820 53286
rect 19876 53284 19882 53286
rect 19574 53275 19882 53284
rect 4214 52796 4522 52805
rect 4214 52794 4220 52796
rect 4276 52794 4300 52796
rect 4356 52794 4380 52796
rect 4436 52794 4460 52796
rect 4516 52794 4522 52796
rect 4276 52742 4278 52794
rect 4458 52742 4460 52794
rect 4214 52740 4220 52742
rect 4276 52740 4300 52742
rect 4356 52740 4380 52742
rect 4436 52740 4460 52742
rect 4516 52740 4522 52742
rect 4214 52731 4522 52740
rect 19574 52252 19882 52261
rect 19574 52250 19580 52252
rect 19636 52250 19660 52252
rect 19716 52250 19740 52252
rect 19796 52250 19820 52252
rect 19876 52250 19882 52252
rect 19636 52198 19638 52250
rect 19818 52198 19820 52250
rect 19574 52196 19580 52198
rect 19636 52196 19660 52198
rect 19716 52196 19740 52198
rect 19796 52196 19820 52198
rect 19876 52196 19882 52198
rect 19574 52187 19882 52196
rect 4214 51708 4522 51717
rect 4214 51706 4220 51708
rect 4276 51706 4300 51708
rect 4356 51706 4380 51708
rect 4436 51706 4460 51708
rect 4516 51706 4522 51708
rect 4276 51654 4278 51706
rect 4458 51654 4460 51706
rect 4214 51652 4220 51654
rect 4276 51652 4300 51654
rect 4356 51652 4380 51654
rect 4436 51652 4460 51654
rect 4516 51652 4522 51654
rect 4214 51643 4522 51652
rect 19574 51164 19882 51173
rect 19574 51162 19580 51164
rect 19636 51162 19660 51164
rect 19716 51162 19740 51164
rect 19796 51162 19820 51164
rect 19876 51162 19882 51164
rect 19636 51110 19638 51162
rect 19818 51110 19820 51162
rect 19574 51108 19580 51110
rect 19636 51108 19660 51110
rect 19716 51108 19740 51110
rect 19796 51108 19820 51110
rect 19876 51108 19882 51110
rect 19574 51099 19882 51108
rect 4214 50620 4522 50629
rect 4214 50618 4220 50620
rect 4276 50618 4300 50620
rect 4356 50618 4380 50620
rect 4436 50618 4460 50620
rect 4516 50618 4522 50620
rect 4276 50566 4278 50618
rect 4458 50566 4460 50618
rect 4214 50564 4220 50566
rect 4276 50564 4300 50566
rect 4356 50564 4380 50566
rect 4436 50564 4460 50566
rect 4516 50564 4522 50566
rect 4214 50555 4522 50564
rect 19574 50076 19882 50085
rect 19574 50074 19580 50076
rect 19636 50074 19660 50076
rect 19716 50074 19740 50076
rect 19796 50074 19820 50076
rect 19876 50074 19882 50076
rect 19636 50022 19638 50074
rect 19818 50022 19820 50074
rect 19574 50020 19580 50022
rect 19636 50020 19660 50022
rect 19716 50020 19740 50022
rect 19796 50020 19820 50022
rect 19876 50020 19882 50022
rect 19574 50011 19882 50020
rect 4214 49532 4522 49541
rect 4214 49530 4220 49532
rect 4276 49530 4300 49532
rect 4356 49530 4380 49532
rect 4436 49530 4460 49532
rect 4516 49530 4522 49532
rect 4276 49478 4278 49530
rect 4458 49478 4460 49530
rect 4214 49476 4220 49478
rect 4276 49476 4300 49478
rect 4356 49476 4380 49478
rect 4436 49476 4460 49478
rect 4516 49476 4522 49478
rect 4214 49467 4522 49476
rect 19574 48988 19882 48997
rect 19574 48986 19580 48988
rect 19636 48986 19660 48988
rect 19716 48986 19740 48988
rect 19796 48986 19820 48988
rect 19876 48986 19882 48988
rect 19636 48934 19638 48986
rect 19818 48934 19820 48986
rect 19574 48932 19580 48934
rect 19636 48932 19660 48934
rect 19716 48932 19740 48934
rect 19796 48932 19820 48934
rect 19876 48932 19882 48934
rect 19574 48923 19882 48932
rect 4214 48444 4522 48453
rect 4214 48442 4220 48444
rect 4276 48442 4300 48444
rect 4356 48442 4380 48444
rect 4436 48442 4460 48444
rect 4516 48442 4522 48444
rect 4276 48390 4278 48442
rect 4458 48390 4460 48442
rect 4214 48388 4220 48390
rect 4276 48388 4300 48390
rect 4356 48388 4380 48390
rect 4436 48388 4460 48390
rect 4516 48388 4522 48390
rect 4214 48379 4522 48388
rect 19574 47900 19882 47909
rect 19574 47898 19580 47900
rect 19636 47898 19660 47900
rect 19716 47898 19740 47900
rect 19796 47898 19820 47900
rect 19876 47898 19882 47900
rect 19636 47846 19638 47898
rect 19818 47846 19820 47898
rect 19574 47844 19580 47846
rect 19636 47844 19660 47846
rect 19716 47844 19740 47846
rect 19796 47844 19820 47846
rect 19876 47844 19882 47846
rect 19574 47835 19882 47844
rect 4214 47356 4522 47365
rect 4214 47354 4220 47356
rect 4276 47354 4300 47356
rect 4356 47354 4380 47356
rect 4436 47354 4460 47356
rect 4516 47354 4522 47356
rect 4276 47302 4278 47354
rect 4458 47302 4460 47354
rect 4214 47300 4220 47302
rect 4276 47300 4300 47302
rect 4356 47300 4380 47302
rect 4436 47300 4460 47302
rect 4516 47300 4522 47302
rect 4214 47291 4522 47300
rect 19574 46812 19882 46821
rect 19574 46810 19580 46812
rect 19636 46810 19660 46812
rect 19716 46810 19740 46812
rect 19796 46810 19820 46812
rect 19876 46810 19882 46812
rect 19636 46758 19638 46810
rect 19818 46758 19820 46810
rect 19574 46756 19580 46758
rect 19636 46756 19660 46758
rect 19716 46756 19740 46758
rect 19796 46756 19820 46758
rect 19876 46756 19882 46758
rect 19574 46747 19882 46756
rect 4214 46268 4522 46277
rect 4214 46266 4220 46268
rect 4276 46266 4300 46268
rect 4356 46266 4380 46268
rect 4436 46266 4460 46268
rect 4516 46266 4522 46268
rect 4276 46214 4278 46266
rect 4458 46214 4460 46266
rect 4214 46212 4220 46214
rect 4276 46212 4300 46214
rect 4356 46212 4380 46214
rect 4436 46212 4460 46214
rect 4516 46212 4522 46214
rect 4214 46203 4522 46212
rect 19574 45724 19882 45733
rect 19574 45722 19580 45724
rect 19636 45722 19660 45724
rect 19716 45722 19740 45724
rect 19796 45722 19820 45724
rect 19876 45722 19882 45724
rect 19636 45670 19638 45722
rect 19818 45670 19820 45722
rect 19574 45668 19580 45670
rect 19636 45668 19660 45670
rect 19716 45668 19740 45670
rect 19796 45668 19820 45670
rect 19876 45668 19882 45670
rect 19574 45659 19882 45668
rect 4214 45180 4522 45189
rect 4214 45178 4220 45180
rect 4276 45178 4300 45180
rect 4356 45178 4380 45180
rect 4436 45178 4460 45180
rect 4516 45178 4522 45180
rect 4276 45126 4278 45178
rect 4458 45126 4460 45178
rect 4214 45124 4220 45126
rect 4276 45124 4300 45126
rect 4356 45124 4380 45126
rect 4436 45124 4460 45126
rect 4516 45124 4522 45126
rect 4214 45115 4522 45124
rect 19574 44636 19882 44645
rect 19574 44634 19580 44636
rect 19636 44634 19660 44636
rect 19716 44634 19740 44636
rect 19796 44634 19820 44636
rect 19876 44634 19882 44636
rect 19636 44582 19638 44634
rect 19818 44582 19820 44634
rect 19574 44580 19580 44582
rect 19636 44580 19660 44582
rect 19716 44580 19740 44582
rect 19796 44580 19820 44582
rect 19876 44580 19882 44582
rect 19574 44571 19882 44580
rect 4214 44092 4522 44101
rect 4214 44090 4220 44092
rect 4276 44090 4300 44092
rect 4356 44090 4380 44092
rect 4436 44090 4460 44092
rect 4516 44090 4522 44092
rect 4276 44038 4278 44090
rect 4458 44038 4460 44090
rect 4214 44036 4220 44038
rect 4276 44036 4300 44038
rect 4356 44036 4380 44038
rect 4436 44036 4460 44038
rect 4516 44036 4522 44038
rect 4214 44027 4522 44036
rect 19574 43548 19882 43557
rect 19574 43546 19580 43548
rect 19636 43546 19660 43548
rect 19716 43546 19740 43548
rect 19796 43546 19820 43548
rect 19876 43546 19882 43548
rect 19636 43494 19638 43546
rect 19818 43494 19820 43546
rect 19574 43492 19580 43494
rect 19636 43492 19660 43494
rect 19716 43492 19740 43494
rect 19796 43492 19820 43494
rect 19876 43492 19882 43494
rect 19574 43483 19882 43492
rect 4214 43004 4522 43013
rect 4214 43002 4220 43004
rect 4276 43002 4300 43004
rect 4356 43002 4380 43004
rect 4436 43002 4460 43004
rect 4516 43002 4522 43004
rect 4276 42950 4278 43002
rect 4458 42950 4460 43002
rect 4214 42948 4220 42950
rect 4276 42948 4300 42950
rect 4356 42948 4380 42950
rect 4436 42948 4460 42950
rect 4516 42948 4522 42950
rect 4214 42939 4522 42948
rect 19574 42460 19882 42469
rect 19574 42458 19580 42460
rect 19636 42458 19660 42460
rect 19716 42458 19740 42460
rect 19796 42458 19820 42460
rect 19876 42458 19882 42460
rect 19636 42406 19638 42458
rect 19818 42406 19820 42458
rect 19574 42404 19580 42406
rect 19636 42404 19660 42406
rect 19716 42404 19740 42406
rect 19796 42404 19820 42406
rect 19876 42404 19882 42406
rect 19574 42395 19882 42404
rect 4214 41916 4522 41925
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41851 4522 41860
rect 19574 41372 19882 41381
rect 19574 41370 19580 41372
rect 19636 41370 19660 41372
rect 19716 41370 19740 41372
rect 19796 41370 19820 41372
rect 19876 41370 19882 41372
rect 19636 41318 19638 41370
rect 19818 41318 19820 41370
rect 19574 41316 19580 41318
rect 19636 41316 19660 41318
rect 19716 41316 19740 41318
rect 19796 41316 19820 41318
rect 19876 41316 19882 41318
rect 19574 41307 19882 41316
rect 4214 40828 4522 40837
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40763 4522 40772
rect 19574 40284 19882 40293
rect 19574 40282 19580 40284
rect 19636 40282 19660 40284
rect 19716 40282 19740 40284
rect 19796 40282 19820 40284
rect 19876 40282 19882 40284
rect 19636 40230 19638 40282
rect 19818 40230 19820 40282
rect 19574 40228 19580 40230
rect 19636 40228 19660 40230
rect 19716 40228 19740 40230
rect 19796 40228 19820 40230
rect 19876 40228 19882 40230
rect 19574 40219 19882 40228
rect 4214 39740 4522 39749
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39675 4522 39684
rect 19574 39196 19882 39205
rect 19574 39194 19580 39196
rect 19636 39194 19660 39196
rect 19716 39194 19740 39196
rect 19796 39194 19820 39196
rect 19876 39194 19882 39196
rect 19636 39142 19638 39194
rect 19818 39142 19820 39194
rect 19574 39140 19580 39142
rect 19636 39140 19660 39142
rect 19716 39140 19740 39142
rect 19796 39140 19820 39142
rect 19876 39140 19882 39142
rect 19574 39131 19882 39140
rect 4214 38652 4522 38661
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38587 4522 38596
rect 19574 38108 19882 38117
rect 19574 38106 19580 38108
rect 19636 38106 19660 38108
rect 19716 38106 19740 38108
rect 19796 38106 19820 38108
rect 19876 38106 19882 38108
rect 19636 38054 19638 38106
rect 19818 38054 19820 38106
rect 19574 38052 19580 38054
rect 19636 38052 19660 38054
rect 19716 38052 19740 38054
rect 19796 38052 19820 38054
rect 19876 38052 19882 38054
rect 19574 38043 19882 38052
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 21652 31754 21680 56646
rect 21376 31726 21680 31754
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 7564 30252 7616 30258
rect 7564 30194 7616 30200
rect 6736 30184 6788 30190
rect 6736 30126 6788 30132
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 5080 29164 5132 29170
rect 5080 29106 5132 29112
rect 4804 28960 4856 28966
rect 4804 28902 4856 28908
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 4816 28626 4844 28902
rect 4804 28620 4856 28626
rect 4804 28562 4856 28568
rect 5092 28558 5120 29106
rect 5816 29028 5868 29034
rect 5816 28970 5868 28976
rect 5080 28552 5132 28558
rect 5080 28494 5132 28500
rect 3792 28416 3844 28422
rect 3792 28358 3844 28364
rect 3804 27674 3832 28358
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 3792 27668 3844 27674
rect 3792 27610 3844 27616
rect 1952 27532 2004 27538
rect 1952 27474 2004 27480
rect 1964 27130 1992 27474
rect 2964 27464 3016 27470
rect 2964 27406 3016 27412
rect 1952 27124 2004 27130
rect 1952 27066 2004 27072
rect 2976 26926 3004 27406
rect 5172 27396 5224 27402
rect 5172 27338 5224 27344
rect 5184 27130 5212 27338
rect 5724 27328 5776 27334
rect 5724 27270 5776 27276
rect 5736 27146 5764 27270
rect 4620 27124 4672 27130
rect 4620 27066 4672 27072
rect 5172 27124 5224 27130
rect 5172 27066 5224 27072
rect 5644 27118 5764 27146
rect 3148 26988 3200 26994
rect 3148 26930 3200 26936
rect 2964 26920 3016 26926
rect 2964 26862 3016 26868
rect 2320 25900 2372 25906
rect 2320 25842 2372 25848
rect 2504 25900 2556 25906
rect 2504 25842 2556 25848
rect 2332 24886 2360 25842
rect 2516 25498 2544 25842
rect 2504 25492 2556 25498
rect 2504 25434 2556 25440
rect 2976 25294 3004 26862
rect 3160 26042 3188 26930
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 3148 26036 3200 26042
rect 3148 25978 3200 25984
rect 3424 26036 3476 26042
rect 3476 25996 3648 26024
rect 3424 25978 3476 25984
rect 3620 25906 3648 25996
rect 3403 25900 3455 25906
rect 3608 25900 3660 25906
rect 3455 25848 3464 25888
rect 3403 25842 3464 25848
rect 3608 25842 3660 25848
rect 3436 25786 3464 25842
rect 3436 25770 3924 25786
rect 3332 25764 3384 25770
rect 3436 25764 3936 25770
rect 3436 25758 3884 25764
rect 3332 25706 3384 25712
rect 3884 25706 3936 25712
rect 3240 25696 3292 25702
rect 3240 25638 3292 25644
rect 2964 25288 3016 25294
rect 2964 25230 3016 25236
rect 2320 24880 2372 24886
rect 2320 24822 2372 24828
rect 2332 24614 2360 24822
rect 2320 24608 2372 24614
rect 2320 24550 2372 24556
rect 2976 24274 3004 25230
rect 3252 24818 3280 25638
rect 3344 25498 3372 25706
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 3332 25492 3384 25498
rect 3332 25434 3384 25440
rect 3344 24954 3372 25434
rect 4160 25220 4212 25226
rect 4160 25162 4212 25168
rect 3332 24948 3384 24954
rect 3332 24890 3384 24896
rect 3240 24812 3292 24818
rect 3240 24754 3292 24760
rect 3700 24812 3752 24818
rect 3700 24754 3752 24760
rect 2964 24268 3016 24274
rect 2964 24210 3016 24216
rect 2136 23724 2188 23730
rect 2136 23666 2188 23672
rect 2320 23724 2372 23730
rect 2320 23666 2372 23672
rect 2504 23724 2556 23730
rect 2504 23666 2556 23672
rect 2148 22982 2176 23666
rect 2332 23322 2360 23666
rect 2320 23316 2372 23322
rect 2320 23258 2372 23264
rect 2228 23044 2280 23050
rect 2228 22986 2280 22992
rect 2136 22976 2188 22982
rect 2136 22918 2188 22924
rect 2240 22710 2268 22986
rect 2228 22704 2280 22710
rect 2516 22681 2544 23666
rect 2976 23662 3004 24210
rect 3712 24070 3740 24754
rect 4172 24750 4200 25162
rect 4160 24744 4212 24750
rect 4160 24686 4212 24692
rect 4632 24682 4660 27066
rect 4712 26784 4764 26790
rect 4712 26726 4764 26732
rect 4724 26518 4752 26726
rect 4712 26512 4764 26518
rect 4712 26454 4764 26460
rect 4724 25294 4752 26454
rect 4988 25764 5040 25770
rect 4988 25706 5040 25712
rect 4712 25288 4764 25294
rect 4712 25230 4764 25236
rect 4620 24676 4672 24682
rect 4620 24618 4672 24624
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 3700 24064 3752 24070
rect 3700 24006 3752 24012
rect 3424 23860 3476 23866
rect 3424 23802 3476 23808
rect 2688 23656 2740 23662
rect 2688 23598 2740 23604
rect 2964 23656 3016 23662
rect 2964 23598 3016 23604
rect 2700 22710 2728 23598
rect 2688 22704 2740 22710
rect 2228 22646 2280 22652
rect 2502 22672 2558 22681
rect 2688 22646 2740 22652
rect 2502 22607 2558 22616
rect 2412 22024 2464 22030
rect 2516 22012 2544 22607
rect 2596 22432 2648 22438
rect 2596 22374 2648 22380
rect 2608 22166 2636 22374
rect 2700 22166 2728 22646
rect 2596 22160 2648 22166
rect 2596 22102 2648 22108
rect 2688 22160 2740 22166
rect 2688 22102 2740 22108
rect 2976 22098 3004 23598
rect 3436 23118 3464 23802
rect 3424 23112 3476 23118
rect 3424 23054 3476 23060
rect 3332 22976 3384 22982
rect 3332 22918 3384 22924
rect 2964 22092 3016 22098
rect 2964 22034 3016 22040
rect 2464 21984 2544 22012
rect 2412 21966 2464 21972
rect 2976 21554 3004 22034
rect 3240 22024 3292 22030
rect 3240 21966 3292 21972
rect 3148 21888 3200 21894
rect 3148 21830 3200 21836
rect 3160 21554 3188 21830
rect 2964 21548 3016 21554
rect 2964 21490 3016 21496
rect 3148 21548 3200 21554
rect 3148 21490 3200 21496
rect 3252 21078 3280 21966
rect 3240 21072 3292 21078
rect 3240 21014 3292 21020
rect 1492 20936 1544 20942
rect 1492 20878 1544 20884
rect 1860 20936 1912 20942
rect 1860 20878 1912 20884
rect 1400 20460 1452 20466
rect 1400 20402 1452 20408
rect 1412 17338 1440 20402
rect 1504 20398 1532 20878
rect 1492 20392 1544 20398
rect 1492 20334 1544 20340
rect 1504 19718 1532 20334
rect 1492 19712 1544 19718
rect 1492 19654 1544 19660
rect 1504 18834 1532 19654
rect 1492 18828 1544 18834
rect 1492 18770 1544 18776
rect 1768 18760 1820 18766
rect 1768 18702 1820 18708
rect 1400 17332 1452 17338
rect 1400 17274 1452 17280
rect 1412 15502 1440 17274
rect 1780 15706 1808 18702
rect 1872 17882 1900 20878
rect 3148 20256 3200 20262
rect 3148 20198 3200 20204
rect 2228 19848 2280 19854
rect 2228 19790 2280 19796
rect 2240 19514 2268 19790
rect 2228 19508 2280 19514
rect 2228 19450 2280 19456
rect 2872 19372 2924 19378
rect 2872 19314 2924 19320
rect 2780 19304 2832 19310
rect 2780 19246 2832 19252
rect 2792 18290 2820 19246
rect 2884 18426 2912 19314
rect 3160 19310 3188 20198
rect 3148 19304 3200 19310
rect 3148 19246 3200 19252
rect 2872 18420 2924 18426
rect 2872 18362 2924 18368
rect 2780 18284 2832 18290
rect 2780 18226 2832 18232
rect 2320 18080 2372 18086
rect 2320 18022 2372 18028
rect 1860 17876 1912 17882
rect 1860 17818 1912 17824
rect 1872 17610 1900 17818
rect 2332 17678 2360 18022
rect 2884 17746 2912 18362
rect 2872 17740 2924 17746
rect 2872 17682 2924 17688
rect 2320 17672 2372 17678
rect 2320 17614 2372 17620
rect 1860 17604 1912 17610
rect 1860 17546 1912 17552
rect 2332 17202 2360 17614
rect 2884 17338 2912 17682
rect 2872 17332 2924 17338
rect 2872 17274 2924 17280
rect 2320 17196 2372 17202
rect 2320 17138 2372 17144
rect 2596 17196 2648 17202
rect 2596 17138 2648 17144
rect 1952 16992 2004 16998
rect 1952 16934 2004 16940
rect 1964 16794 1992 16934
rect 1952 16788 2004 16794
rect 1952 16730 2004 16736
rect 2332 16590 2360 17138
rect 2412 17128 2464 17134
rect 2412 17070 2464 17076
rect 2320 16584 2372 16590
rect 2320 16526 2372 16532
rect 1768 15700 1820 15706
rect 1768 15642 1820 15648
rect 1400 15496 1452 15502
rect 1400 15438 1452 15444
rect 2136 15496 2188 15502
rect 2136 15438 2188 15444
rect 1492 13864 1544 13870
rect 1492 13806 1544 13812
rect 1504 10810 1532 13806
rect 2044 12844 2096 12850
rect 2044 12786 2096 12792
rect 1952 11824 2004 11830
rect 1952 11766 2004 11772
rect 1492 10804 1544 10810
rect 1492 10746 1544 10752
rect 1964 10606 1992 11766
rect 2056 11762 2084 12786
rect 2148 11898 2176 15438
rect 2320 14272 2372 14278
rect 2320 14214 2372 14220
rect 2136 11892 2188 11898
rect 2136 11834 2188 11840
rect 2044 11756 2096 11762
rect 2044 11698 2096 11704
rect 1952 10600 2004 10606
rect 1952 10542 2004 10548
rect 1964 9178 1992 10542
rect 1952 9172 2004 9178
rect 1952 9114 2004 9120
rect 2228 8900 2280 8906
rect 2228 8842 2280 8848
rect 2044 8628 2096 8634
rect 2044 8570 2096 8576
rect 1860 8492 1912 8498
rect 1860 8434 1912 8440
rect 1872 8090 1900 8434
rect 1860 8084 1912 8090
rect 1860 8026 1912 8032
rect 1768 7880 1820 7886
rect 1768 7822 1820 7828
rect 1780 6390 1808 7822
rect 2056 6798 2084 8570
rect 2136 8356 2188 8362
rect 2136 8298 2188 8304
rect 2148 7954 2176 8298
rect 2136 7948 2188 7954
rect 2136 7890 2188 7896
rect 1952 6792 2004 6798
rect 1952 6734 2004 6740
rect 2044 6792 2096 6798
rect 2044 6734 2096 6740
rect 1964 6458 1992 6734
rect 1952 6452 2004 6458
rect 1952 6394 2004 6400
rect 1768 6384 1820 6390
rect 1768 6326 1820 6332
rect 1780 4622 1808 6326
rect 1860 5636 1912 5642
rect 1860 5578 1912 5584
rect 1872 5370 1900 5578
rect 1860 5364 1912 5370
rect 1860 5306 1912 5312
rect 2056 5166 2084 6734
rect 2240 5658 2268 8842
rect 2332 7818 2360 14214
rect 2424 11898 2452 17070
rect 2608 16726 2636 17138
rect 2884 16794 2912 17274
rect 3240 17264 3292 17270
rect 3240 17206 3292 17212
rect 2964 17196 3016 17202
rect 2964 17138 3016 17144
rect 3148 17196 3200 17202
rect 3148 17138 3200 17144
rect 2976 16794 3004 17138
rect 3160 16998 3188 17138
rect 3148 16992 3200 16998
rect 3148 16934 3200 16940
rect 2872 16788 2924 16794
rect 2872 16730 2924 16736
rect 2964 16788 3016 16794
rect 2964 16730 3016 16736
rect 2596 16720 2648 16726
rect 2596 16662 2648 16668
rect 2964 16652 3016 16658
rect 2964 16594 3016 16600
rect 2780 15700 2832 15706
rect 2780 15642 2832 15648
rect 2596 15020 2648 15026
rect 2596 14962 2648 14968
rect 2504 13932 2556 13938
rect 2504 13874 2556 13880
rect 2516 13394 2544 13874
rect 2504 13388 2556 13394
rect 2504 13330 2556 13336
rect 2516 12238 2544 13330
rect 2608 13258 2636 14962
rect 2688 14068 2740 14074
rect 2688 14010 2740 14016
rect 2700 13326 2728 14010
rect 2792 13734 2820 15642
rect 2976 15570 3004 16594
rect 3160 16250 3188 16934
rect 3252 16658 3280 17206
rect 3240 16652 3292 16658
rect 3240 16594 3292 16600
rect 3148 16244 3200 16250
rect 3148 16186 3200 16192
rect 3252 16114 3280 16594
rect 3240 16108 3292 16114
rect 3068 16068 3240 16096
rect 2964 15564 3016 15570
rect 2964 15506 3016 15512
rect 2872 14612 2924 14618
rect 2872 14554 2924 14560
rect 2884 13938 2912 14554
rect 3068 14006 3096 16068
rect 3240 16050 3292 16056
rect 3148 15972 3200 15978
rect 3148 15914 3200 15920
rect 3160 15162 3188 15914
rect 3148 15156 3200 15162
rect 3148 15098 3200 15104
rect 3344 14618 3372 22918
rect 3436 22778 3464 23054
rect 3424 22772 3476 22778
rect 3424 22714 3476 22720
rect 3424 21072 3476 21078
rect 3424 21014 3476 21020
rect 3436 16114 3464 21014
rect 3424 16108 3476 16114
rect 3424 16050 3476 16056
rect 3424 15564 3476 15570
rect 3424 15506 3476 15512
rect 3332 14612 3384 14618
rect 3332 14554 3384 14560
rect 3056 14000 3108 14006
rect 3056 13942 3108 13948
rect 2872 13932 2924 13938
rect 2924 13892 3004 13920
rect 2872 13874 2924 13880
rect 2872 13796 2924 13802
rect 2872 13738 2924 13744
rect 2780 13728 2832 13734
rect 2780 13670 2832 13676
rect 2884 13530 2912 13738
rect 2976 13530 3004 13892
rect 2872 13524 2924 13530
rect 2872 13466 2924 13472
rect 2964 13524 3016 13530
rect 2964 13466 3016 13472
rect 2688 13320 2740 13326
rect 2688 13262 2740 13268
rect 3068 13258 3096 13942
rect 2596 13252 2648 13258
rect 2596 13194 2648 13200
rect 3056 13252 3108 13258
rect 3056 13194 3108 13200
rect 2608 12918 2636 13194
rect 2596 12912 2648 12918
rect 2596 12854 2648 12860
rect 2688 12640 2740 12646
rect 2688 12582 2740 12588
rect 2700 12238 2728 12582
rect 3068 12306 3096 13194
rect 3148 12844 3200 12850
rect 3148 12786 3200 12792
rect 3160 12442 3188 12786
rect 3148 12436 3200 12442
rect 3148 12378 3200 12384
rect 3056 12300 3108 12306
rect 3056 12242 3108 12248
rect 2504 12232 2556 12238
rect 2504 12174 2556 12180
rect 2688 12232 2740 12238
rect 3436 12209 3464 15506
rect 3608 15496 3660 15502
rect 3608 15438 3660 15444
rect 3620 13938 3648 15438
rect 3608 13932 3660 13938
rect 3608 13874 3660 13880
rect 3620 13734 3648 13874
rect 3608 13728 3660 13734
rect 3608 13670 3660 13676
rect 3712 12442 3740 24006
rect 4342 23896 4398 23905
rect 4342 23831 4344 23840
rect 4396 23831 4398 23840
rect 4344 23802 4396 23808
rect 4894 23760 4950 23769
rect 4894 23695 4896 23704
rect 4948 23695 4950 23704
rect 4896 23666 4948 23672
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 5000 22624 5028 25706
rect 5264 25152 5316 25158
rect 5264 25094 5316 25100
rect 5276 24682 5304 25094
rect 5264 24676 5316 24682
rect 5264 24618 5316 24624
rect 5644 24410 5672 27118
rect 5828 27062 5856 28970
rect 6748 28966 6776 30126
rect 7576 29510 7604 30194
rect 8024 29640 8076 29646
rect 8024 29582 8076 29588
rect 7932 29572 7984 29578
rect 7932 29514 7984 29520
rect 7564 29504 7616 29510
rect 7564 29446 7616 29452
rect 7012 29096 7064 29102
rect 7012 29038 7064 29044
rect 6736 28960 6788 28966
rect 6736 28902 6788 28908
rect 6920 28960 6972 28966
rect 6920 28902 6972 28908
rect 6748 28762 6776 28902
rect 6736 28756 6788 28762
rect 6736 28698 6788 28704
rect 6932 28558 6960 28902
rect 6276 28552 6328 28558
rect 6276 28494 6328 28500
rect 6920 28552 6972 28558
rect 6920 28494 6972 28500
rect 6288 28218 6316 28494
rect 6276 28212 6328 28218
rect 6276 28154 6328 28160
rect 7024 27606 7052 29038
rect 7576 28082 7604 29446
rect 7944 29238 7972 29514
rect 7932 29232 7984 29238
rect 7932 29174 7984 29180
rect 7656 28960 7708 28966
rect 7656 28902 7708 28908
rect 7668 28558 7696 28902
rect 7656 28552 7708 28558
rect 7656 28494 7708 28500
rect 7564 28076 7616 28082
rect 7564 28018 7616 28024
rect 7668 27962 7696 28494
rect 7944 28422 7972 29174
rect 8036 29034 8064 29582
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 19892 29164 19944 29170
rect 19892 29106 19944 29112
rect 8116 29096 8168 29102
rect 8116 29038 8168 29044
rect 19432 29096 19484 29102
rect 19432 29038 19484 29044
rect 8024 29028 8076 29034
rect 8024 28970 8076 28976
rect 7840 28416 7892 28422
rect 7840 28358 7892 28364
rect 7932 28416 7984 28422
rect 7932 28358 7984 28364
rect 7852 28082 7880 28358
rect 7840 28076 7892 28082
rect 7840 28018 7892 28024
rect 7576 27934 7696 27962
rect 7012 27600 7064 27606
rect 7012 27542 7064 27548
rect 7196 27328 7248 27334
rect 7196 27270 7248 27276
rect 5816 27056 5868 27062
rect 5816 26998 5868 27004
rect 7104 27056 7156 27062
rect 7104 26998 7156 27004
rect 5724 26988 5776 26994
rect 5724 26930 5776 26936
rect 5736 26314 5764 26930
rect 6276 26920 6328 26926
rect 6276 26862 6328 26868
rect 5724 26308 5776 26314
rect 5724 26250 5776 26256
rect 5632 24404 5684 24410
rect 5632 24346 5684 24352
rect 5540 24132 5592 24138
rect 5540 24074 5592 24080
rect 5264 24064 5316 24070
rect 5264 24006 5316 24012
rect 5276 23730 5304 24006
rect 5552 23866 5580 24074
rect 5540 23860 5592 23866
rect 5540 23802 5592 23808
rect 5080 23724 5132 23730
rect 5080 23666 5132 23672
rect 5264 23724 5316 23730
rect 5264 23666 5316 23672
rect 5092 23322 5120 23666
rect 5264 23588 5316 23594
rect 5264 23530 5316 23536
rect 5080 23316 5132 23322
rect 5080 23258 5132 23264
rect 5276 23254 5304 23530
rect 5644 23322 5672 24346
rect 5632 23316 5684 23322
rect 5632 23258 5684 23264
rect 5264 23248 5316 23254
rect 5264 23190 5316 23196
rect 5276 22710 5304 23190
rect 5644 23050 5672 23258
rect 5632 23044 5684 23050
rect 5632 22986 5684 22992
rect 5264 22704 5316 22710
rect 5264 22646 5316 22652
rect 5080 22636 5132 22642
rect 5000 22596 5080 22624
rect 5080 22578 5132 22584
rect 5632 22636 5684 22642
rect 5632 22578 5684 22584
rect 4620 22432 4672 22438
rect 4620 22374 4672 22380
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 4632 21350 4660 22374
rect 4620 21344 4672 21350
rect 4620 21286 4672 21292
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4632 21010 4660 21286
rect 4620 21004 4672 21010
rect 4620 20946 4672 20952
rect 4896 20392 4948 20398
rect 4896 20334 4948 20340
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4908 19854 4936 20334
rect 4620 19848 4672 19854
rect 4620 19790 4672 19796
rect 4896 19848 4948 19854
rect 4896 19790 4948 19796
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 4344 18624 4396 18630
rect 4344 18566 4396 18572
rect 4356 18222 4384 18566
rect 4632 18222 4660 19790
rect 4988 18624 5040 18630
rect 4988 18566 5040 18572
rect 5000 18358 5028 18566
rect 4988 18352 5040 18358
rect 4988 18294 5040 18300
rect 4344 18216 4396 18222
rect 4344 18158 4396 18164
rect 4620 18216 4672 18222
rect 4620 18158 4672 18164
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4632 17882 4660 18158
rect 4620 17876 4672 17882
rect 4620 17818 4672 17824
rect 4632 17270 4660 17818
rect 4620 17264 4672 17270
rect 4620 17206 4672 17212
rect 4712 17196 4764 17202
rect 4712 17138 4764 17144
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4724 16522 4752 17138
rect 4988 16992 5040 16998
rect 4988 16934 5040 16940
rect 5000 16590 5028 16934
rect 5092 16726 5120 22578
rect 5172 22432 5224 22438
rect 5172 22374 5224 22380
rect 5184 22030 5212 22374
rect 5644 22234 5672 22578
rect 5632 22228 5684 22234
rect 5632 22170 5684 22176
rect 5172 22024 5224 22030
rect 5172 21966 5224 21972
rect 5540 21480 5592 21486
rect 5460 21428 5540 21434
rect 5460 21422 5592 21428
rect 5460 21406 5580 21422
rect 5460 20398 5488 21406
rect 5736 20806 5764 26250
rect 6288 25838 6316 26862
rect 7116 26586 7144 26998
rect 7208 26586 7236 27270
rect 7104 26580 7156 26586
rect 7104 26522 7156 26528
rect 7196 26580 7248 26586
rect 7196 26522 7248 26528
rect 6644 25900 6696 25906
rect 6644 25842 6696 25848
rect 6276 25832 6328 25838
rect 6276 25774 6328 25780
rect 6000 25152 6052 25158
rect 6000 25094 6052 25100
rect 6012 24886 6040 25094
rect 6000 24880 6052 24886
rect 6000 24822 6052 24828
rect 5816 23044 5868 23050
rect 5816 22986 5868 22992
rect 5828 21690 5856 22986
rect 6012 22982 6040 24822
rect 6288 24206 6316 25774
rect 6656 25498 6684 25842
rect 6644 25492 6696 25498
rect 6644 25434 6696 25440
rect 7012 25288 7064 25294
rect 7012 25230 7064 25236
rect 6828 25152 6880 25158
rect 6828 25094 6880 25100
rect 6840 24614 6868 25094
rect 7024 24954 7052 25230
rect 7012 24948 7064 24954
rect 7012 24890 7064 24896
rect 7208 24818 7236 26522
rect 7576 26518 7604 27934
rect 7944 27470 7972 28358
rect 8036 27470 8064 28970
rect 8128 28558 8156 29038
rect 18972 29028 19024 29034
rect 18972 28970 19024 28976
rect 9404 28960 9456 28966
rect 9404 28902 9456 28908
rect 8300 28756 8352 28762
rect 8300 28698 8352 28704
rect 8116 28552 8168 28558
rect 8116 28494 8168 28500
rect 8312 27946 8340 28698
rect 9416 28558 9444 28902
rect 18984 28694 19012 28970
rect 19248 28756 19300 28762
rect 19248 28698 19300 28704
rect 9680 28688 9732 28694
rect 9680 28630 9732 28636
rect 18972 28688 19024 28694
rect 18972 28630 19024 28636
rect 9404 28552 9456 28558
rect 9404 28494 9456 28500
rect 9128 28484 9180 28490
rect 9128 28426 9180 28432
rect 9140 28218 9168 28426
rect 9128 28212 9180 28218
rect 9128 28154 9180 28160
rect 9416 28082 9444 28494
rect 9692 28218 9720 28630
rect 18604 28620 18656 28626
rect 18604 28562 18656 28568
rect 10232 28552 10284 28558
rect 10232 28494 10284 28500
rect 14004 28552 14056 28558
rect 14004 28494 14056 28500
rect 18052 28552 18104 28558
rect 18052 28494 18104 28500
rect 9680 28212 9732 28218
rect 9680 28154 9732 28160
rect 8576 28076 8628 28082
rect 8576 28018 8628 28024
rect 9404 28076 9456 28082
rect 9404 28018 9456 28024
rect 8300 27940 8352 27946
rect 8300 27882 8352 27888
rect 7748 27464 7800 27470
rect 7748 27406 7800 27412
rect 7932 27464 7984 27470
rect 7932 27406 7984 27412
rect 8024 27464 8076 27470
rect 8024 27406 8076 27412
rect 7656 26784 7708 26790
rect 7656 26726 7708 26732
rect 7564 26512 7616 26518
rect 7564 26454 7616 26460
rect 7472 25288 7524 25294
rect 7472 25230 7524 25236
rect 7484 25158 7512 25230
rect 7472 25152 7524 25158
rect 7472 25094 7524 25100
rect 7196 24812 7248 24818
rect 7196 24754 7248 24760
rect 7208 24682 7236 24754
rect 7196 24676 7248 24682
rect 7196 24618 7248 24624
rect 6828 24608 6880 24614
rect 6828 24550 6880 24556
rect 6276 24200 6328 24206
rect 6276 24142 6328 24148
rect 6288 23186 6316 24142
rect 7472 24064 7524 24070
rect 7472 24006 7524 24012
rect 7484 23798 7512 24006
rect 7472 23792 7524 23798
rect 7472 23734 7524 23740
rect 6276 23180 6328 23186
rect 6276 23122 6328 23128
rect 6000 22976 6052 22982
rect 6000 22918 6052 22924
rect 6288 22710 6316 23122
rect 6368 23112 6420 23118
rect 6368 23054 6420 23060
rect 6276 22704 6328 22710
rect 5906 22672 5962 22681
rect 6276 22646 6328 22652
rect 5906 22607 5908 22616
rect 5960 22607 5962 22616
rect 5908 22578 5960 22584
rect 6380 21962 6408 23054
rect 7380 22976 7432 22982
rect 7380 22918 7432 22924
rect 6368 21956 6420 21962
rect 6368 21898 6420 21904
rect 5816 21684 5868 21690
rect 5816 21626 5868 21632
rect 5540 20800 5592 20806
rect 5540 20742 5592 20748
rect 5724 20800 5776 20806
rect 5724 20742 5776 20748
rect 5552 20505 5580 20742
rect 5538 20496 5594 20505
rect 5538 20431 5540 20440
rect 5592 20431 5594 20440
rect 5540 20402 5592 20408
rect 5448 20392 5500 20398
rect 5448 20334 5500 20340
rect 6380 20262 6408 21898
rect 7196 21888 7248 21894
rect 7196 21830 7248 21836
rect 6644 21548 6696 21554
rect 6644 21490 6696 21496
rect 6550 21176 6606 21185
rect 6656 21146 6684 21490
rect 6550 21111 6552 21120
rect 6604 21111 6606 21120
rect 6644 21140 6696 21146
rect 6552 21082 6604 21088
rect 6644 21082 6696 21088
rect 6920 21004 6972 21010
rect 6920 20946 6972 20952
rect 6932 20398 6960 20946
rect 7208 20924 7236 21830
rect 7288 21344 7340 21350
rect 7288 21286 7340 21292
rect 7300 21078 7328 21286
rect 7288 21072 7340 21078
rect 7288 21014 7340 21020
rect 7288 20936 7340 20942
rect 7208 20896 7288 20924
rect 7288 20878 7340 20884
rect 6920 20392 6972 20398
rect 6920 20334 6972 20340
rect 6368 20256 6420 20262
rect 6368 20198 6420 20204
rect 6380 19446 6408 20198
rect 7288 20052 7340 20058
rect 7288 19994 7340 20000
rect 7104 19848 7156 19854
rect 7104 19790 7156 19796
rect 6920 19712 6972 19718
rect 6920 19654 6972 19660
rect 6368 19440 6420 19446
rect 6368 19382 6420 19388
rect 6932 19378 6960 19654
rect 6920 19372 6972 19378
rect 6920 19314 6972 19320
rect 7116 19156 7144 19790
rect 7300 19310 7328 19994
rect 7288 19304 7340 19310
rect 7288 19246 7340 19252
rect 7288 19168 7340 19174
rect 7116 19128 7288 19156
rect 7288 19110 7340 19116
rect 7300 18970 7328 19110
rect 7288 18964 7340 18970
rect 7288 18906 7340 18912
rect 5816 18760 5868 18766
rect 5816 18702 5868 18708
rect 5264 17536 5316 17542
rect 5264 17478 5316 17484
rect 5276 17270 5304 17478
rect 5264 17264 5316 17270
rect 5264 17206 5316 17212
rect 5080 16720 5132 16726
rect 5080 16662 5132 16668
rect 4988 16584 5040 16590
rect 4988 16526 5040 16532
rect 4712 16516 4764 16522
rect 4712 16458 4764 16464
rect 4724 15910 4752 16458
rect 3884 15904 3936 15910
rect 3884 15846 3936 15852
rect 4712 15904 4764 15910
rect 4712 15846 4764 15852
rect 3896 15502 3924 15846
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 3884 15496 3936 15502
rect 3884 15438 3936 15444
rect 4724 15094 4752 15846
rect 5276 15450 5304 17206
rect 5448 16584 5500 16590
rect 5448 16526 5500 16532
rect 5356 16448 5408 16454
rect 5356 16390 5408 16396
rect 5184 15422 5304 15450
rect 4896 15360 4948 15366
rect 4896 15302 4948 15308
rect 4908 15162 4936 15302
rect 4896 15156 4948 15162
rect 4896 15098 4948 15104
rect 4712 15088 4764 15094
rect 4712 15030 4764 15036
rect 5184 15026 5212 15422
rect 5264 15360 5316 15366
rect 5264 15302 5316 15308
rect 5172 15020 5224 15026
rect 5172 14962 5224 14968
rect 5276 14958 5304 15302
rect 5368 15026 5396 16390
rect 5356 15020 5408 15026
rect 5356 14962 5408 14968
rect 5264 14952 5316 14958
rect 5460 14929 5488 16526
rect 5264 14894 5316 14900
rect 5446 14920 5502 14929
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 5276 14346 5304 14894
rect 5446 14855 5502 14864
rect 5460 14822 5488 14855
rect 5448 14816 5500 14822
rect 5448 14758 5500 14764
rect 5264 14340 5316 14346
rect 5264 14282 5316 14288
rect 5632 14272 5684 14278
rect 5632 14214 5684 14220
rect 3792 13728 3844 13734
rect 3792 13670 3844 13676
rect 3804 12918 3832 13670
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 5644 13326 5672 14214
rect 5632 13320 5684 13326
rect 5632 13262 5684 13268
rect 4620 12980 4672 12986
rect 4620 12922 4672 12928
rect 3792 12912 3844 12918
rect 3792 12854 3844 12860
rect 3700 12436 3752 12442
rect 3700 12378 3752 12384
rect 3712 12238 3740 12378
rect 3804 12238 3832 12854
rect 4632 12753 4660 12922
rect 4618 12744 4674 12753
rect 4618 12679 4620 12688
rect 4672 12679 4674 12688
rect 4620 12650 4672 12656
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 3700 12232 3752 12238
rect 2688 12174 2740 12180
rect 3422 12200 3478 12209
rect 3700 12174 3752 12180
rect 3792 12232 3844 12238
rect 3792 12174 3844 12180
rect 3422 12135 3478 12144
rect 3148 12096 3200 12102
rect 3148 12038 3200 12044
rect 2412 11892 2464 11898
rect 2412 11834 2464 11840
rect 2504 11688 2556 11694
rect 2504 11630 2556 11636
rect 2516 11558 2544 11630
rect 2504 11552 2556 11558
rect 2504 11494 2556 11500
rect 2516 11014 2544 11494
rect 3160 11150 3188 12038
rect 3240 11620 3292 11626
rect 3240 11562 3292 11568
rect 3148 11144 3200 11150
rect 3148 11086 3200 11092
rect 2504 11008 2556 11014
rect 2504 10950 2556 10956
rect 2516 10674 2544 10950
rect 2504 10668 2556 10674
rect 2504 10610 2556 10616
rect 2516 10470 2544 10610
rect 2504 10464 2556 10470
rect 2504 10406 2556 10412
rect 2412 8900 2464 8906
rect 2412 8842 2464 8848
rect 2424 8498 2452 8842
rect 2412 8492 2464 8498
rect 2412 8434 2464 8440
rect 2320 7812 2372 7818
rect 2320 7754 2372 7760
rect 2332 7206 2360 7754
rect 2424 7546 2452 8434
rect 2516 8090 2544 10406
rect 2780 8968 2832 8974
rect 2780 8910 2832 8916
rect 2792 8838 2820 8910
rect 2780 8832 2832 8838
rect 2780 8774 2832 8780
rect 3056 8832 3108 8838
rect 3056 8774 3108 8780
rect 2504 8084 2556 8090
rect 2504 8026 2556 8032
rect 2412 7540 2464 7546
rect 2412 7482 2464 7488
rect 2320 7200 2372 7206
rect 2320 7142 2372 7148
rect 2424 6610 2452 7482
rect 3068 6798 3096 8774
rect 3056 6792 3108 6798
rect 3056 6734 3108 6740
rect 2964 6724 3016 6730
rect 2964 6666 3016 6672
rect 2504 6656 2556 6662
rect 2424 6604 2504 6610
rect 2424 6598 2556 6604
rect 2424 6582 2544 6598
rect 2780 6384 2832 6390
rect 2780 6326 2832 6332
rect 2792 5914 2820 6326
rect 2976 6322 3004 6666
rect 2964 6316 3016 6322
rect 2964 6258 3016 6264
rect 3056 6112 3108 6118
rect 3056 6054 3108 6060
rect 2780 5908 2832 5914
rect 2780 5850 2832 5856
rect 2148 5630 2268 5658
rect 2044 5160 2096 5166
rect 2044 5102 2096 5108
rect 1768 4616 1820 4622
rect 1768 4558 1820 4564
rect 2148 4146 2176 5630
rect 2320 5228 2372 5234
rect 2320 5170 2372 5176
rect 2504 5228 2556 5234
rect 2504 5170 2556 5176
rect 2332 4826 2360 5170
rect 2412 5160 2464 5166
rect 2412 5102 2464 5108
rect 2320 4820 2372 4826
rect 2320 4762 2372 4768
rect 2228 4684 2280 4690
rect 2228 4626 2280 4632
rect 2136 4140 2188 4146
rect 2136 4082 2188 4088
rect 2148 3942 2176 4082
rect 2136 3936 2188 3942
rect 2136 3878 2188 3884
rect 2240 3738 2268 4626
rect 2320 4480 2372 4486
rect 2320 4422 2372 4428
rect 2332 4146 2360 4422
rect 2424 4214 2452 5102
rect 2412 4208 2464 4214
rect 2412 4150 2464 4156
rect 2516 4146 2544 5170
rect 3068 5030 3096 6054
rect 3056 5024 3108 5030
rect 3056 4966 3108 4972
rect 3160 4554 3188 11086
rect 3252 5914 3280 11562
rect 3804 11150 3832 12174
rect 4632 11898 4660 12650
rect 5828 12434 5856 18702
rect 7300 18358 7328 18906
rect 7288 18352 7340 18358
rect 7288 18294 7340 18300
rect 6920 18284 6972 18290
rect 6920 18226 6972 18232
rect 7104 18284 7156 18290
rect 7104 18226 7156 18232
rect 6460 18080 6512 18086
rect 6460 18022 6512 18028
rect 6472 17610 6500 18022
rect 6460 17604 6512 17610
rect 6460 17546 6512 17552
rect 6932 17338 6960 18226
rect 7012 17536 7064 17542
rect 7012 17478 7064 17484
rect 6920 17332 6972 17338
rect 6920 17274 6972 17280
rect 7024 17218 7052 17478
rect 6932 17190 7052 17218
rect 6932 16114 6960 17190
rect 7116 17066 7144 18226
rect 7104 17060 7156 17066
rect 7104 17002 7156 17008
rect 7012 16448 7064 16454
rect 7012 16390 7064 16396
rect 6920 16108 6972 16114
rect 6920 16050 6972 16056
rect 7024 15978 7052 16390
rect 7196 16040 7248 16046
rect 7196 15982 7248 15988
rect 7012 15972 7064 15978
rect 7012 15914 7064 15920
rect 6552 15904 6604 15910
rect 6552 15846 6604 15852
rect 6460 15700 6512 15706
rect 6460 15642 6512 15648
rect 6472 15502 6500 15642
rect 6564 15502 6592 15846
rect 6460 15496 6512 15502
rect 6460 15438 6512 15444
rect 6552 15496 6604 15502
rect 6552 15438 6604 15444
rect 7024 15434 7052 15914
rect 7208 15570 7236 15982
rect 7196 15564 7248 15570
rect 7196 15506 7248 15512
rect 7012 15428 7064 15434
rect 7012 15370 7064 15376
rect 6644 15360 6696 15366
rect 6644 15302 6696 15308
rect 6184 14816 6236 14822
rect 6184 14758 6236 14764
rect 6092 13932 6144 13938
rect 6092 13874 6144 13880
rect 6104 13530 6132 13874
rect 6092 13524 6144 13530
rect 6092 13466 6144 13472
rect 5828 12406 5948 12434
rect 5816 12368 5868 12374
rect 5816 12310 5868 12316
rect 5724 12096 5776 12102
rect 5724 12038 5776 12044
rect 4620 11892 4672 11898
rect 4620 11834 4672 11840
rect 5736 11830 5764 12038
rect 5724 11824 5776 11830
rect 5724 11766 5776 11772
rect 5828 11762 5856 12310
rect 5816 11756 5868 11762
rect 5816 11698 5868 11704
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 3792 11144 3844 11150
rect 3792 11086 3844 11092
rect 3804 10130 3832 11086
rect 5080 11076 5132 11082
rect 5080 11018 5132 11024
rect 5092 10810 5120 11018
rect 5632 11008 5684 11014
rect 5632 10950 5684 10956
rect 5080 10804 5132 10810
rect 5080 10746 5132 10752
rect 5644 10674 5672 10950
rect 4712 10668 4764 10674
rect 4712 10610 4764 10616
rect 5540 10668 5592 10674
rect 5540 10610 5592 10616
rect 5632 10668 5684 10674
rect 5632 10610 5684 10616
rect 4724 10577 4752 10610
rect 4710 10568 4766 10577
rect 4710 10503 4766 10512
rect 5448 10464 5500 10470
rect 5448 10406 5500 10412
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 3792 10124 3844 10130
rect 3792 10066 3844 10072
rect 5172 9716 5224 9722
rect 5172 9658 5224 9664
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 5184 9178 5212 9658
rect 5460 9586 5488 10406
rect 5552 10130 5580 10610
rect 5540 10124 5592 10130
rect 5540 10066 5592 10072
rect 5448 9580 5500 9586
rect 5448 9522 5500 9528
rect 5724 9580 5776 9586
rect 5724 9522 5776 9528
rect 5172 9172 5224 9178
rect 5172 9114 5224 9120
rect 3516 8968 3568 8974
rect 3516 8910 3568 8916
rect 3528 8566 3556 8910
rect 5080 8900 5132 8906
rect 5080 8842 5132 8848
rect 5092 8634 5120 8842
rect 5080 8628 5132 8634
rect 5080 8570 5132 8576
rect 3516 8560 3568 8566
rect 3516 8502 3568 8508
rect 3528 7410 3556 8502
rect 5184 8498 5212 9114
rect 5264 8968 5316 8974
rect 5264 8910 5316 8916
rect 5276 8566 5304 8910
rect 5264 8560 5316 8566
rect 5264 8502 5316 8508
rect 5172 8492 5224 8498
rect 5172 8434 5224 8440
rect 3792 8356 3844 8362
rect 3792 8298 3844 8304
rect 3804 8090 3832 8298
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 3792 8084 3844 8090
rect 3792 8026 3844 8032
rect 5460 7886 5488 9522
rect 5632 9376 5684 9382
rect 5632 9318 5684 9324
rect 5644 8634 5672 9318
rect 5632 8628 5684 8634
rect 5632 8570 5684 8576
rect 5736 8378 5764 9522
rect 5644 8350 5764 8378
rect 5448 7880 5500 7886
rect 5448 7822 5500 7828
rect 3516 7404 3568 7410
rect 3516 7346 3568 7352
rect 5540 7404 5592 7410
rect 5540 7346 5592 7352
rect 3528 6984 3556 7346
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 3436 6956 3556 6984
rect 3436 6390 3464 6956
rect 4068 6928 4120 6934
rect 4068 6870 4120 6876
rect 4080 6798 4108 6870
rect 5552 6866 5580 7346
rect 5540 6860 5592 6866
rect 5540 6802 5592 6808
rect 4068 6792 4120 6798
rect 4068 6734 4120 6740
rect 3516 6656 3568 6662
rect 3516 6598 3568 6604
rect 3424 6384 3476 6390
rect 3424 6326 3476 6332
rect 3240 5908 3292 5914
rect 3240 5850 3292 5856
rect 3252 5302 3280 5850
rect 3240 5296 3292 5302
rect 3240 5238 3292 5244
rect 3436 5166 3464 6326
rect 3528 5370 3556 6598
rect 4080 6458 4108 6734
rect 4068 6452 4120 6458
rect 4068 6394 4120 6400
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 5644 5817 5672 8350
rect 5722 7848 5778 7857
rect 5722 7783 5724 7792
rect 5776 7783 5778 7792
rect 5724 7754 5776 7760
rect 5736 7546 5764 7754
rect 5724 7540 5776 7546
rect 5724 7482 5776 7488
rect 5724 6792 5776 6798
rect 5724 6734 5776 6740
rect 5736 6202 5764 6734
rect 5828 6322 5856 11698
rect 5920 10826 5948 12406
rect 6000 11756 6052 11762
rect 6000 11698 6052 11704
rect 6012 11558 6040 11698
rect 6000 11552 6052 11558
rect 6000 11494 6052 11500
rect 6012 11082 6040 11494
rect 6092 11212 6144 11218
rect 6092 11154 6144 11160
rect 6000 11076 6052 11082
rect 6000 11018 6052 11024
rect 5920 10798 6040 10826
rect 5908 10668 5960 10674
rect 5908 10610 5960 10616
rect 5920 8430 5948 10610
rect 5908 8424 5960 8430
rect 5908 8366 5960 8372
rect 6012 8022 6040 10798
rect 6104 10062 6132 11154
rect 6092 10056 6144 10062
rect 6092 9998 6144 10004
rect 6104 9926 6132 9957
rect 6092 9920 6144 9926
rect 6090 9888 6092 9897
rect 6144 9888 6146 9897
rect 6090 9823 6146 9832
rect 6104 9654 6132 9823
rect 6092 9648 6144 9654
rect 6092 9590 6144 9596
rect 6000 8016 6052 8022
rect 6000 7958 6052 7964
rect 6000 7744 6052 7750
rect 6000 7686 6052 7692
rect 5906 7032 5962 7041
rect 5906 6967 5962 6976
rect 5816 6316 5868 6322
rect 5816 6258 5868 6264
rect 5736 6174 5856 6202
rect 5828 6118 5856 6174
rect 5816 6112 5868 6118
rect 5816 6054 5868 6060
rect 5828 5846 5856 6054
rect 5816 5840 5868 5846
rect 5630 5808 5686 5817
rect 5630 5743 5686 5752
rect 5736 5800 5816 5828
rect 5644 5710 5672 5743
rect 5632 5704 5684 5710
rect 5632 5646 5684 5652
rect 5356 5568 5408 5574
rect 5356 5510 5408 5516
rect 3516 5364 3568 5370
rect 3516 5306 3568 5312
rect 5368 5302 5396 5510
rect 5356 5296 5408 5302
rect 5356 5238 5408 5244
rect 3424 5160 3476 5166
rect 3424 5102 3476 5108
rect 3974 5128 4030 5137
rect 3148 4548 3200 4554
rect 3148 4490 3200 4496
rect 3436 4214 3464 5102
rect 3974 5063 4030 5072
rect 3988 4826 4016 5063
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 3976 4820 4028 4826
rect 3976 4762 4028 4768
rect 5632 4820 5684 4826
rect 5632 4762 5684 4768
rect 3988 4554 4016 4762
rect 3976 4548 4028 4554
rect 3976 4490 4028 4496
rect 5540 4480 5592 4486
rect 5540 4422 5592 4428
rect 3424 4208 3476 4214
rect 3424 4150 3476 4156
rect 4986 4176 5042 4185
rect 2320 4140 2372 4146
rect 2320 4082 2372 4088
rect 2504 4140 2556 4146
rect 2504 4082 2556 4088
rect 2516 3738 2544 4082
rect 2228 3732 2280 3738
rect 2228 3674 2280 3680
rect 2504 3732 2556 3738
rect 2504 3674 2556 3680
rect 3436 3466 3464 4150
rect 4986 4111 4988 4120
rect 5040 4111 5042 4120
rect 4988 4082 5040 4088
rect 5552 4010 5580 4422
rect 5644 4214 5672 4762
rect 5736 4690 5764 5800
rect 5816 5782 5868 5788
rect 5816 5704 5868 5710
rect 5816 5646 5868 5652
rect 5828 5370 5856 5646
rect 5816 5364 5868 5370
rect 5816 5306 5868 5312
rect 5724 4684 5776 4690
rect 5724 4626 5776 4632
rect 5632 4208 5684 4214
rect 5632 4150 5684 4156
rect 5540 4004 5592 4010
rect 5540 3946 5592 3952
rect 4620 3936 4672 3942
rect 4620 3878 4672 3884
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4632 3777 4660 3878
rect 4618 3768 4674 3777
rect 4618 3703 4674 3712
rect 3424 3460 3476 3466
rect 3424 3402 3476 3408
rect 5644 3398 5672 4150
rect 4160 3392 4212 3398
rect 4160 3334 4212 3340
rect 5632 3392 5684 3398
rect 5632 3334 5684 3340
rect 4172 3058 4200 3334
rect 4160 3052 4212 3058
rect 4160 2994 4212 3000
rect 4896 2984 4948 2990
rect 4896 2926 4948 2932
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 4908 2446 4936 2926
rect 5920 2922 5948 6967
rect 6012 6798 6040 7686
rect 6196 6934 6224 14758
rect 6368 13864 6420 13870
rect 6368 13806 6420 13812
rect 6380 12442 6408 13806
rect 6552 13320 6604 13326
rect 6552 13262 6604 13268
rect 6564 12714 6592 13262
rect 6552 12708 6604 12714
rect 6552 12650 6604 12656
rect 6368 12436 6420 12442
rect 6368 12378 6420 12384
rect 6380 12238 6408 12378
rect 6368 12232 6420 12238
rect 6368 12174 6420 12180
rect 6656 11082 6684 15302
rect 7024 14822 7052 15370
rect 7012 14816 7064 14822
rect 7012 14758 7064 14764
rect 7104 14816 7156 14822
rect 7104 14758 7156 14764
rect 7116 14074 7144 14758
rect 7208 14414 7236 15506
rect 7196 14408 7248 14414
rect 7196 14350 7248 14356
rect 7104 14068 7156 14074
rect 7104 14010 7156 14016
rect 7392 13258 7420 22918
rect 7472 22636 7524 22642
rect 7472 22578 7524 22584
rect 7484 19854 7512 22578
rect 7576 20602 7604 26454
rect 7668 26382 7696 26726
rect 7656 26376 7708 26382
rect 7656 26318 7708 26324
rect 7668 26042 7696 26318
rect 7656 26036 7708 26042
rect 7656 25978 7708 25984
rect 7656 25696 7708 25702
rect 7656 25638 7708 25644
rect 7668 25294 7696 25638
rect 7656 25288 7708 25294
rect 7656 25230 7708 25236
rect 7656 23520 7708 23526
rect 7656 23462 7708 23468
rect 7668 23118 7696 23462
rect 7656 23112 7708 23118
rect 7656 23054 7708 23060
rect 7760 21146 7788 27406
rect 7944 26858 7972 27406
rect 8588 27334 8616 28018
rect 9588 28008 9640 28014
rect 9588 27950 9640 27956
rect 9496 27940 9548 27946
rect 9496 27882 9548 27888
rect 9220 27872 9272 27878
rect 9220 27814 9272 27820
rect 9312 27872 9364 27878
rect 9312 27814 9364 27820
rect 8024 27328 8076 27334
rect 8024 27270 8076 27276
rect 8576 27328 8628 27334
rect 8576 27270 8628 27276
rect 7932 26852 7984 26858
rect 7932 26794 7984 26800
rect 7932 25288 7984 25294
rect 7932 25230 7984 25236
rect 7944 24954 7972 25230
rect 7932 24948 7984 24954
rect 7932 24890 7984 24896
rect 8036 24410 8064 27270
rect 8116 25288 8168 25294
rect 8116 25230 8168 25236
rect 8128 24886 8156 25230
rect 8300 25152 8352 25158
rect 8300 25094 8352 25100
rect 8116 24880 8168 24886
rect 8168 24840 8248 24868
rect 8116 24822 8168 24828
rect 8024 24404 8076 24410
rect 8024 24346 8076 24352
rect 8036 24290 8064 24346
rect 7944 24262 8064 24290
rect 7944 24206 7972 24262
rect 7932 24200 7984 24206
rect 7932 24142 7984 24148
rect 8116 24200 8168 24206
rect 8116 24142 8168 24148
rect 7840 23724 7892 23730
rect 7840 23666 7892 23672
rect 7852 23050 7880 23666
rect 7840 23044 7892 23050
rect 7840 22986 7892 22992
rect 8128 22982 8156 24142
rect 8220 23118 8248 24840
rect 8312 23730 8340 25094
rect 8588 23905 8616 27270
rect 8760 25900 8812 25906
rect 8760 25842 8812 25848
rect 8772 25498 8800 25842
rect 8760 25492 8812 25498
rect 8760 25434 8812 25440
rect 8668 24608 8720 24614
rect 8668 24550 8720 24556
rect 8574 23896 8630 23905
rect 8574 23831 8630 23840
rect 8482 23760 8538 23769
rect 8300 23724 8352 23730
rect 8482 23695 8484 23704
rect 8300 23666 8352 23672
rect 8536 23695 8538 23704
rect 8484 23666 8536 23672
rect 8208 23112 8260 23118
rect 8208 23054 8260 23060
rect 8116 22976 8168 22982
rect 8116 22918 8168 22924
rect 8312 22234 8340 23666
rect 8300 22228 8352 22234
rect 8300 22170 8352 22176
rect 7932 22092 7984 22098
rect 7932 22034 7984 22040
rect 7840 21480 7892 21486
rect 7840 21422 7892 21428
rect 7748 21140 7800 21146
rect 7748 21082 7800 21088
rect 7852 20874 7880 21422
rect 7840 20868 7892 20874
rect 7840 20810 7892 20816
rect 7748 20800 7800 20806
rect 7748 20742 7800 20748
rect 7564 20596 7616 20602
rect 7564 20538 7616 20544
rect 7472 19848 7524 19854
rect 7472 19790 7524 19796
rect 7656 18216 7708 18222
rect 7656 18158 7708 18164
rect 7668 17882 7696 18158
rect 7656 17876 7708 17882
rect 7656 17818 7708 17824
rect 7760 17678 7788 20742
rect 7852 19990 7880 20810
rect 7944 20754 7972 22034
rect 8300 22024 8352 22030
rect 8352 21984 8432 22012
rect 8300 21966 8352 21972
rect 8116 21956 8168 21962
rect 8116 21898 8168 21904
rect 8128 21536 8156 21898
rect 8208 21548 8260 21554
rect 8128 21508 8208 21536
rect 8208 21490 8260 21496
rect 8300 21548 8352 21554
rect 8300 21490 8352 21496
rect 8114 21040 8170 21049
rect 8114 20975 8170 20984
rect 8128 20942 8156 20975
rect 8116 20936 8168 20942
rect 8116 20878 8168 20884
rect 7944 20726 8064 20754
rect 7932 20392 7984 20398
rect 7932 20334 7984 20340
rect 7840 19984 7892 19990
rect 7840 19926 7892 19932
rect 7852 19718 7880 19926
rect 7944 19786 7972 20334
rect 8036 19922 8064 20726
rect 8128 20602 8156 20878
rect 8116 20596 8168 20602
rect 8116 20538 8168 20544
rect 8220 20466 8248 21490
rect 8312 20942 8340 21490
rect 8404 21350 8432 21984
rect 8484 21888 8536 21894
rect 8484 21830 8536 21836
rect 8392 21344 8444 21350
rect 8392 21286 8444 21292
rect 8300 20936 8352 20942
rect 8300 20878 8352 20884
rect 8404 20874 8432 21286
rect 8496 21078 8524 21830
rect 8484 21072 8536 21078
rect 8484 21014 8536 21020
rect 8392 20868 8444 20874
rect 8392 20810 8444 20816
rect 8208 20460 8260 20466
rect 8208 20402 8260 20408
rect 8116 20052 8168 20058
rect 8116 19994 8168 20000
rect 8024 19916 8076 19922
rect 8024 19858 8076 19864
rect 7932 19780 7984 19786
rect 7932 19722 7984 19728
rect 7840 19712 7892 19718
rect 7840 19654 7892 19660
rect 7840 19440 7892 19446
rect 7840 19382 7892 19388
rect 7748 17672 7800 17678
rect 7748 17614 7800 17620
rect 7472 17128 7524 17134
rect 7472 17070 7524 17076
rect 7484 16590 7512 17070
rect 7760 16726 7788 17614
rect 7748 16720 7800 16726
rect 7748 16662 7800 16668
rect 7472 16584 7524 16590
rect 7472 16526 7524 16532
rect 7656 16584 7708 16590
rect 7656 16526 7708 16532
rect 7484 15094 7512 16526
rect 7668 16250 7696 16526
rect 7656 16244 7708 16250
rect 7656 16186 7708 16192
rect 7668 15502 7696 16186
rect 7656 15496 7708 15502
rect 7656 15438 7708 15444
rect 7852 15162 7880 19382
rect 7944 19174 7972 19722
rect 8036 19514 8064 19858
rect 8024 19508 8076 19514
rect 8024 19450 8076 19456
rect 8128 19378 8156 19994
rect 8220 19446 8248 20402
rect 8484 20324 8536 20330
rect 8484 20266 8536 20272
rect 8496 19922 8524 20266
rect 8484 19916 8536 19922
rect 8484 19858 8536 19864
rect 8208 19440 8260 19446
rect 8208 19382 8260 19388
rect 8116 19372 8168 19378
rect 8116 19314 8168 19320
rect 7932 19168 7984 19174
rect 7932 19110 7984 19116
rect 7944 17762 7972 19110
rect 8024 18284 8076 18290
rect 8024 18226 8076 18232
rect 8036 17882 8064 18226
rect 8024 17876 8076 17882
rect 8024 17818 8076 17824
rect 7944 17734 8064 17762
rect 7932 15564 7984 15570
rect 7932 15506 7984 15512
rect 7840 15156 7892 15162
rect 7840 15098 7892 15104
rect 7472 15088 7524 15094
rect 7472 15030 7524 15036
rect 7484 14482 7512 15030
rect 7564 15020 7616 15026
rect 7564 14962 7616 14968
rect 7472 14476 7524 14482
rect 7472 14418 7524 14424
rect 7380 13252 7432 13258
rect 7380 13194 7432 13200
rect 6828 13184 6880 13190
rect 6828 13126 6880 13132
rect 6840 12374 6868 13126
rect 7472 12640 7524 12646
rect 7472 12582 7524 12588
rect 7104 12436 7156 12442
rect 7104 12378 7156 12384
rect 6828 12368 6880 12374
rect 6828 12310 6880 12316
rect 6920 12300 6972 12306
rect 6920 12242 6972 12248
rect 6736 12232 6788 12238
rect 6736 12174 6788 12180
rect 6828 12232 6880 12238
rect 6828 12174 6880 12180
rect 6748 11898 6776 12174
rect 6736 11892 6788 11898
rect 6736 11834 6788 11840
rect 6644 11076 6696 11082
rect 6644 11018 6696 11024
rect 6656 10266 6684 11018
rect 6840 10810 6868 12174
rect 6828 10804 6880 10810
rect 6828 10746 6880 10752
rect 6828 10668 6880 10674
rect 6828 10610 6880 10616
rect 6644 10260 6696 10266
rect 6644 10202 6696 10208
rect 6840 10062 6868 10610
rect 6932 10198 6960 12242
rect 7116 11694 7144 12378
rect 7484 12238 7512 12582
rect 7472 12232 7524 12238
rect 7472 12174 7524 12180
rect 7196 12096 7248 12102
rect 7196 12038 7248 12044
rect 7208 11898 7236 12038
rect 7196 11892 7248 11898
rect 7196 11834 7248 11840
rect 7104 11688 7156 11694
rect 7104 11630 7156 11636
rect 7116 11218 7144 11630
rect 7104 11212 7156 11218
rect 7104 11154 7156 11160
rect 7116 10674 7144 11154
rect 7104 10668 7156 10674
rect 7104 10610 7156 10616
rect 7380 10668 7432 10674
rect 7380 10610 7432 10616
rect 7288 10464 7340 10470
rect 7288 10406 7340 10412
rect 6920 10192 6972 10198
rect 6920 10134 6972 10140
rect 6276 10056 6328 10062
rect 6276 9998 6328 10004
rect 6828 10056 6880 10062
rect 6828 9998 6880 10004
rect 6288 9761 6316 9998
rect 6932 9994 6960 10134
rect 6920 9988 6972 9994
rect 6920 9930 6972 9936
rect 6274 9752 6330 9761
rect 6274 9687 6330 9696
rect 6288 7954 6316 9687
rect 6932 9586 6960 9930
rect 7104 9920 7156 9926
rect 7104 9862 7156 9868
rect 6920 9580 6972 9586
rect 6920 9522 6972 9528
rect 6552 9512 6604 9518
rect 6552 9454 6604 9460
rect 6276 7948 6328 7954
rect 6276 7890 6328 7896
rect 6184 6928 6236 6934
rect 6184 6870 6236 6876
rect 6288 6798 6316 7890
rect 6460 7812 6512 7818
rect 6460 7754 6512 7760
rect 6472 7410 6500 7754
rect 6460 7404 6512 7410
rect 6460 7346 6512 7352
rect 6000 6792 6052 6798
rect 6000 6734 6052 6740
rect 6276 6792 6328 6798
rect 6276 6734 6328 6740
rect 6288 5710 6316 6734
rect 6472 6458 6500 7346
rect 6460 6452 6512 6458
rect 6460 6394 6512 6400
rect 6276 5704 6328 5710
rect 6276 5646 6328 5652
rect 6472 5302 6500 6394
rect 6564 5710 6592 9454
rect 7116 9450 7144 9862
rect 7300 9518 7328 10406
rect 7392 10266 7420 10610
rect 7576 10266 7604 14962
rect 7748 14408 7800 14414
rect 7748 14350 7800 14356
rect 7760 14074 7788 14350
rect 7748 14068 7800 14074
rect 7748 14010 7800 14016
rect 7760 13977 7788 14010
rect 7746 13968 7802 13977
rect 7746 13903 7802 13912
rect 7748 12844 7800 12850
rect 7748 12786 7800 12792
rect 7656 12368 7708 12374
rect 7656 12310 7708 12316
rect 7668 12238 7696 12310
rect 7656 12232 7708 12238
rect 7656 12174 7708 12180
rect 7380 10260 7432 10266
rect 7380 10202 7432 10208
rect 7564 10260 7616 10266
rect 7564 10202 7616 10208
rect 7288 9512 7340 9518
rect 7288 9454 7340 9460
rect 7104 9444 7156 9450
rect 7104 9386 7156 9392
rect 6920 8968 6972 8974
rect 6920 8910 6972 8916
rect 6932 8498 6960 8910
rect 7012 8832 7064 8838
rect 7012 8774 7064 8780
rect 7024 8566 7052 8774
rect 7012 8560 7064 8566
rect 7012 8502 7064 8508
rect 7116 8498 7144 9386
rect 7288 8832 7340 8838
rect 7286 8800 7288 8809
rect 7340 8800 7342 8809
rect 7286 8735 7342 8744
rect 6920 8492 6972 8498
rect 6920 8434 6972 8440
rect 7104 8492 7156 8498
rect 7668 8480 7696 12174
rect 7760 11014 7788 12786
rect 7748 11008 7800 11014
rect 7748 10950 7800 10956
rect 7728 10056 7780 10062
rect 7780 10004 7788 10044
rect 7728 9998 7788 10004
rect 7760 9466 7788 9998
rect 7944 9500 7972 15506
rect 8036 13841 8064 17734
rect 8128 15434 8156 19314
rect 8484 18420 8536 18426
rect 8484 18362 8536 18368
rect 8496 17202 8524 18362
rect 8208 17196 8260 17202
rect 8208 17138 8260 17144
rect 8484 17196 8536 17202
rect 8484 17138 8536 17144
rect 8220 16794 8248 17138
rect 8208 16788 8260 16794
rect 8208 16730 8260 16736
rect 8392 15496 8444 15502
rect 8392 15438 8444 15444
rect 8484 15496 8536 15502
rect 8484 15438 8536 15444
rect 8116 15428 8168 15434
rect 8116 15370 8168 15376
rect 8404 15026 8432 15438
rect 8392 15020 8444 15026
rect 8392 14962 8444 14968
rect 8392 14884 8444 14890
rect 8392 14826 8444 14832
rect 8300 13932 8352 13938
rect 8300 13874 8352 13880
rect 8022 13832 8078 13841
rect 8022 13767 8078 13776
rect 8312 12186 8340 13874
rect 8404 13326 8432 14826
rect 8392 13320 8444 13326
rect 8392 13262 8444 13268
rect 8392 12640 8444 12646
rect 8392 12582 8444 12588
rect 8404 12374 8432 12582
rect 8392 12368 8444 12374
rect 8392 12310 8444 12316
rect 8312 12158 8432 12186
rect 8024 12096 8076 12102
rect 8024 12038 8076 12044
rect 8300 12096 8352 12102
rect 8300 12038 8352 12044
rect 8036 11762 8064 12038
rect 8024 11756 8076 11762
rect 8024 11698 8076 11704
rect 8312 11082 8340 12038
rect 8300 11076 8352 11082
rect 8300 11018 8352 11024
rect 8116 10056 8168 10062
rect 8116 9998 8168 10004
rect 8128 9761 8156 9998
rect 8114 9752 8170 9761
rect 8114 9687 8170 9696
rect 8312 9654 8340 11018
rect 8300 9648 8352 9654
rect 8300 9590 8352 9596
rect 7944 9472 8156 9500
rect 7760 9438 7880 9466
rect 7748 9376 7800 9382
rect 7748 9318 7800 9324
rect 7760 8974 7788 9318
rect 7748 8968 7800 8974
rect 7748 8910 7800 8916
rect 7852 8809 7880 9438
rect 8128 8974 8156 9472
rect 7932 8968 7984 8974
rect 7932 8910 7984 8916
rect 8116 8968 8168 8974
rect 8404 8922 8432 12158
rect 8496 11830 8524 15438
rect 8588 14618 8616 23831
rect 8680 23662 8708 24550
rect 9128 24200 9180 24206
rect 9128 24142 9180 24148
rect 8852 24064 8904 24070
rect 8852 24006 8904 24012
rect 8864 23730 8892 24006
rect 8852 23724 8904 23730
rect 8852 23666 8904 23672
rect 9039 23724 9091 23730
rect 9039 23666 9091 23672
rect 8668 23656 8720 23662
rect 8668 23598 8720 23604
rect 8760 23520 8812 23526
rect 8760 23462 8812 23468
rect 8668 22976 8720 22982
rect 8668 22918 8720 22924
rect 8680 21026 8708 22918
rect 8772 22030 8800 23462
rect 9048 23322 9076 23666
rect 9036 23316 9088 23322
rect 9036 23258 9088 23264
rect 9140 23186 9168 24142
rect 8944 23180 8996 23186
rect 8944 23122 8996 23128
rect 9128 23180 9180 23186
rect 9128 23122 9180 23128
rect 8956 22098 8984 23122
rect 9036 22228 9088 22234
rect 9036 22170 9088 22176
rect 8944 22092 8996 22098
rect 8944 22034 8996 22040
rect 8760 22024 8812 22030
rect 8760 21966 8812 21972
rect 8772 21486 8800 21966
rect 8956 21894 8984 22034
rect 8944 21888 8996 21894
rect 8944 21830 8996 21836
rect 8760 21480 8812 21486
rect 8760 21422 8812 21428
rect 8758 21176 8814 21185
rect 8758 21111 8760 21120
rect 8812 21111 8814 21120
rect 8760 21082 8812 21088
rect 8680 20998 8800 21026
rect 8668 20936 8720 20942
rect 8668 20878 8720 20884
rect 8680 20398 8708 20878
rect 8668 20392 8720 20398
rect 8668 20334 8720 20340
rect 8680 18834 8708 20334
rect 8668 18828 8720 18834
rect 8668 18770 8720 18776
rect 8680 18358 8708 18770
rect 8772 18426 8800 20998
rect 8852 20868 8904 20874
rect 8852 20810 8904 20816
rect 8760 18420 8812 18426
rect 8760 18362 8812 18368
rect 8668 18352 8720 18358
rect 8668 18294 8720 18300
rect 8680 16658 8708 18294
rect 8760 18216 8812 18222
rect 8760 18158 8812 18164
rect 8772 18086 8800 18158
rect 8760 18080 8812 18086
rect 8760 18022 8812 18028
rect 8772 17746 8800 18022
rect 8760 17740 8812 17746
rect 8760 17682 8812 17688
rect 8772 17270 8800 17682
rect 8760 17264 8812 17270
rect 8760 17206 8812 17212
rect 8760 16992 8812 16998
rect 8760 16934 8812 16940
rect 8668 16652 8720 16658
rect 8668 16594 8720 16600
rect 8772 16590 8800 16934
rect 8760 16584 8812 16590
rect 8760 16526 8812 16532
rect 8864 15434 8892 20810
rect 8852 15428 8904 15434
rect 8852 15370 8904 15376
rect 8956 15162 8984 21830
rect 9048 21554 9076 22170
rect 9036 21548 9088 21554
rect 9036 21490 9088 21496
rect 9048 21010 9076 21490
rect 9036 21004 9088 21010
rect 9036 20946 9088 20952
rect 9232 20058 9260 27814
rect 9324 27674 9352 27814
rect 9312 27668 9364 27674
rect 9312 27610 9364 27616
rect 9404 27464 9456 27470
rect 9404 27406 9456 27412
rect 9416 27130 9444 27406
rect 9404 27124 9456 27130
rect 9404 27066 9456 27072
rect 9404 24132 9456 24138
rect 9404 24074 9456 24080
rect 9416 23866 9444 24074
rect 9404 23860 9456 23866
rect 9404 23802 9456 23808
rect 9404 22636 9456 22642
rect 9404 22578 9456 22584
rect 9312 22432 9364 22438
rect 9312 22374 9364 22380
rect 9324 21078 9352 22374
rect 9312 21072 9364 21078
rect 9312 21014 9364 21020
rect 9220 20052 9272 20058
rect 9220 19994 9272 20000
rect 9107 19845 9159 19851
rect 9159 19793 9168 19836
rect 9107 19787 9168 19793
rect 9140 19514 9168 19787
rect 9128 19508 9180 19514
rect 9128 19450 9180 19456
rect 9324 19334 9352 21014
rect 9416 20806 9444 22578
rect 9508 22522 9536 27882
rect 9600 27606 9628 27950
rect 10244 27674 10272 28494
rect 11612 28076 11664 28082
rect 11612 28018 11664 28024
rect 12164 28076 12216 28082
rect 12164 28018 12216 28024
rect 10876 27872 10928 27878
rect 10876 27814 10928 27820
rect 10232 27668 10284 27674
rect 10232 27610 10284 27616
rect 9588 27600 9640 27606
rect 9588 27542 9640 27548
rect 9600 26518 9628 27542
rect 9784 27526 9996 27554
rect 10888 27538 10916 27814
rect 9784 27470 9812 27526
rect 9772 27464 9824 27470
rect 9772 27406 9824 27412
rect 9968 27334 9996 27526
rect 10876 27532 10928 27538
rect 10876 27474 10928 27480
rect 10692 27396 10744 27402
rect 10692 27338 10744 27344
rect 9956 27328 10008 27334
rect 9956 27270 10008 27276
rect 10704 27130 10732 27338
rect 9680 27124 9732 27130
rect 9680 27066 9732 27072
rect 10692 27124 10744 27130
rect 10692 27066 10744 27072
rect 9588 26512 9640 26518
rect 9588 26454 9640 26460
rect 9588 24200 9640 24206
rect 9588 24142 9640 24148
rect 9600 22710 9628 24142
rect 9692 24070 9720 27066
rect 10048 26988 10100 26994
rect 10048 26930 10100 26936
rect 10060 26246 10088 26930
rect 10888 26790 10916 27474
rect 11520 27464 11572 27470
rect 11520 27406 11572 27412
rect 10876 26784 10928 26790
rect 10876 26726 10928 26732
rect 10888 26586 10916 26726
rect 10876 26580 10928 26586
rect 10876 26522 10928 26528
rect 11244 26444 11296 26450
rect 11244 26386 11296 26392
rect 10784 26376 10836 26382
rect 10784 26318 10836 26324
rect 10048 26240 10100 26246
rect 10048 26182 10100 26188
rect 10060 25702 10088 26182
rect 10692 26036 10744 26042
rect 10692 25978 10744 25984
rect 10048 25696 10100 25702
rect 10048 25638 10100 25644
rect 10060 24614 10088 25638
rect 10704 25294 10732 25978
rect 10796 25430 10824 26318
rect 11060 26240 11112 26246
rect 11060 26182 11112 26188
rect 10784 25424 10836 25430
rect 10784 25366 10836 25372
rect 10140 25288 10192 25294
rect 10140 25230 10192 25236
rect 10692 25288 10744 25294
rect 10692 25230 10744 25236
rect 10048 24608 10100 24614
rect 10048 24550 10100 24556
rect 9772 24336 9824 24342
rect 9772 24278 9824 24284
rect 9680 24064 9732 24070
rect 9680 24006 9732 24012
rect 9692 23866 9720 24006
rect 9680 23860 9732 23866
rect 9680 23802 9732 23808
rect 9784 23662 9812 24278
rect 9864 23792 9916 23798
rect 9864 23734 9916 23740
rect 9772 23656 9824 23662
rect 9772 23598 9824 23604
rect 9588 22704 9640 22710
rect 9588 22646 9640 22652
rect 9508 22494 9628 22522
rect 9600 21418 9628 22494
rect 9680 21480 9732 21486
rect 9678 21448 9680 21457
rect 9732 21448 9734 21457
rect 9588 21412 9640 21418
rect 9678 21383 9734 21392
rect 9588 21354 9640 21360
rect 9680 21344 9732 21350
rect 9680 21286 9732 21292
rect 9692 20942 9720 21286
rect 9680 20936 9732 20942
rect 9680 20878 9732 20884
rect 9404 20800 9456 20806
rect 9404 20742 9456 20748
rect 9416 20534 9444 20742
rect 9404 20528 9456 20534
rect 9404 20470 9456 20476
rect 9416 19854 9444 20470
rect 9772 19916 9824 19922
rect 9772 19858 9824 19864
rect 9404 19848 9456 19854
rect 9404 19790 9456 19796
rect 9324 19306 9444 19334
rect 9784 19310 9812 19858
rect 9128 18080 9180 18086
rect 9128 18022 9180 18028
rect 9140 17610 9168 18022
rect 9220 17672 9272 17678
rect 9220 17614 9272 17620
rect 9128 17604 9180 17610
rect 9128 17546 9180 17552
rect 9232 16182 9260 17614
rect 9220 16176 9272 16182
rect 9220 16118 9272 16124
rect 9312 16108 9364 16114
rect 9312 16050 9364 16056
rect 9324 15706 9352 16050
rect 9312 15700 9364 15706
rect 9312 15642 9364 15648
rect 8944 15156 8996 15162
rect 8944 15098 8996 15104
rect 8852 15020 8904 15026
rect 8852 14962 8904 14968
rect 8576 14612 8628 14618
rect 8576 14554 8628 14560
rect 8760 14612 8812 14618
rect 8760 14554 8812 14560
rect 8772 14006 8800 14554
rect 8760 14000 8812 14006
rect 8760 13942 8812 13948
rect 8864 13938 8892 14962
rect 9036 14612 9088 14618
rect 9036 14554 9088 14560
rect 9048 14074 9076 14554
rect 9416 14346 9444 19306
rect 9772 19304 9824 19310
rect 9772 19246 9824 19252
rect 9876 18442 9904 23734
rect 10152 20466 10180 25230
rect 10796 25226 10824 25366
rect 10784 25220 10836 25226
rect 10784 25162 10836 25168
rect 11072 24682 11100 26182
rect 11256 25362 11284 26386
rect 11428 26240 11480 26246
rect 11428 26182 11480 26188
rect 11440 25974 11468 26182
rect 11428 25968 11480 25974
rect 11428 25910 11480 25916
rect 11532 25906 11560 27406
rect 11624 27130 11652 28018
rect 11612 27124 11664 27130
rect 11612 27066 11664 27072
rect 12176 26858 12204 28018
rect 14016 28014 14044 28494
rect 15384 28484 15436 28490
rect 15384 28426 15436 28432
rect 16764 28484 16816 28490
rect 16764 28426 16816 28432
rect 17776 28484 17828 28490
rect 17776 28426 17828 28432
rect 14004 28008 14056 28014
rect 14004 27950 14056 27956
rect 13912 27872 13964 27878
rect 13912 27814 13964 27820
rect 13820 27532 13872 27538
rect 13820 27474 13872 27480
rect 13452 27396 13504 27402
rect 13452 27338 13504 27344
rect 13084 27328 13136 27334
rect 13084 27270 13136 27276
rect 13096 26926 13124 27270
rect 13464 27130 13492 27338
rect 13452 27124 13504 27130
rect 13452 27066 13504 27072
rect 13832 26994 13860 27474
rect 13924 26994 13952 27814
rect 14016 27334 14044 27950
rect 15396 27946 15424 28426
rect 15384 27940 15436 27946
rect 15384 27882 15436 27888
rect 14556 27872 14608 27878
rect 14556 27814 14608 27820
rect 14568 27470 14596 27814
rect 14556 27464 14608 27470
rect 14556 27406 14608 27412
rect 14740 27464 14792 27470
rect 14740 27406 14792 27412
rect 16580 27464 16632 27470
rect 16580 27406 16632 27412
rect 14004 27328 14056 27334
rect 14004 27270 14056 27276
rect 14096 27328 14148 27334
rect 14096 27270 14148 27276
rect 13820 26988 13872 26994
rect 13820 26930 13872 26936
rect 13912 26988 13964 26994
rect 13912 26930 13964 26936
rect 12992 26920 13044 26926
rect 12992 26862 13044 26868
rect 13084 26920 13136 26926
rect 13084 26862 13136 26868
rect 12164 26852 12216 26858
rect 12164 26794 12216 26800
rect 12176 26314 12204 26794
rect 12900 26376 12952 26382
rect 12900 26318 12952 26324
rect 12164 26308 12216 26314
rect 12164 26250 12216 26256
rect 11520 25900 11572 25906
rect 11520 25842 11572 25848
rect 11244 25356 11296 25362
rect 11244 25298 11296 25304
rect 11060 24676 11112 24682
rect 11060 24618 11112 24624
rect 10968 24608 11020 24614
rect 10968 24550 11020 24556
rect 10876 22636 10928 22642
rect 10876 22578 10928 22584
rect 10888 22234 10916 22578
rect 10876 22228 10928 22234
rect 10876 22170 10928 22176
rect 10600 22024 10652 22030
rect 10600 21966 10652 21972
rect 10612 21690 10640 21966
rect 10508 21684 10560 21690
rect 10508 21626 10560 21632
rect 10600 21684 10652 21690
rect 10600 21626 10652 21632
rect 10232 21548 10284 21554
rect 10232 21490 10284 21496
rect 10244 21350 10272 21490
rect 10232 21344 10284 21350
rect 10232 21286 10284 21292
rect 10140 20460 10192 20466
rect 10140 20402 10192 20408
rect 10140 19712 10192 19718
rect 10140 19654 10192 19660
rect 10048 19440 10100 19446
rect 10048 19382 10100 19388
rect 9876 18426 9996 18442
rect 9864 18420 9996 18426
rect 9916 18414 9996 18420
rect 9864 18362 9916 18368
rect 9864 18284 9916 18290
rect 9864 18226 9916 18232
rect 9876 17882 9904 18226
rect 9864 17876 9916 17882
rect 9864 17818 9916 17824
rect 9968 17814 9996 18414
rect 9956 17808 10008 17814
rect 9956 17750 10008 17756
rect 9968 17270 9996 17750
rect 9956 17264 10008 17270
rect 9956 17206 10008 17212
rect 9588 17196 9640 17202
rect 9588 17138 9640 17144
rect 9600 17105 9628 17138
rect 9586 17096 9642 17105
rect 9586 17031 9642 17040
rect 9496 16448 9548 16454
rect 9496 16390 9548 16396
rect 9508 16114 9536 16390
rect 9496 16108 9548 16114
rect 9496 16050 9548 16056
rect 9588 15564 9640 15570
rect 9588 15506 9640 15512
rect 9600 15434 9628 15506
rect 9772 15496 9824 15502
rect 9772 15438 9824 15444
rect 9588 15428 9640 15434
rect 9588 15370 9640 15376
rect 9404 14340 9456 14346
rect 9404 14282 9456 14288
rect 9128 14272 9180 14278
rect 9128 14214 9180 14220
rect 9140 14074 9168 14214
rect 9036 14068 9088 14074
rect 9036 14010 9088 14016
rect 9128 14068 9180 14074
rect 9128 14010 9180 14016
rect 9600 14006 9628 15370
rect 9588 14000 9640 14006
rect 9588 13942 9640 13948
rect 8668 13932 8720 13938
rect 8668 13874 8720 13880
rect 8852 13932 8904 13938
rect 8852 13874 8904 13880
rect 9404 13932 9456 13938
rect 9404 13874 9456 13880
rect 8680 13394 8708 13874
rect 8668 13388 8720 13394
rect 8668 13330 8720 13336
rect 9416 13326 9444 13874
rect 9600 13394 9628 13942
rect 9588 13388 9640 13394
rect 9588 13330 9640 13336
rect 8944 13320 8996 13326
rect 8944 13262 8996 13268
rect 9404 13320 9456 13326
rect 9404 13262 9456 13268
rect 8852 13184 8904 13190
rect 8852 13126 8904 13132
rect 8484 11824 8536 11830
rect 8484 11766 8536 11772
rect 8864 10674 8892 13126
rect 8956 12918 8984 13262
rect 8944 12912 8996 12918
rect 8944 12854 8996 12860
rect 8956 11898 8984 12854
rect 9680 12844 9732 12850
rect 9680 12786 9732 12792
rect 8944 11892 8996 11898
rect 8944 11834 8996 11840
rect 8944 11008 8996 11014
rect 8944 10950 8996 10956
rect 8484 10668 8536 10674
rect 8484 10610 8536 10616
rect 8852 10668 8904 10674
rect 8852 10610 8904 10616
rect 8116 8910 8168 8916
rect 7838 8800 7894 8809
rect 7838 8735 7894 8744
rect 7944 8634 7972 8910
rect 7932 8628 7984 8634
rect 7932 8570 7984 8576
rect 7932 8492 7984 8498
rect 7668 8452 7932 8480
rect 7104 8434 7156 8440
rect 7932 8434 7984 8440
rect 7012 8424 7064 8430
rect 7012 8366 7064 8372
rect 7472 8424 7524 8430
rect 7944 8401 7972 8434
rect 7472 8366 7524 8372
rect 7930 8392 7986 8401
rect 6736 6724 6788 6730
rect 6736 6666 6788 6672
rect 6644 6316 6696 6322
rect 6644 6258 6696 6264
rect 6552 5704 6604 5710
rect 6552 5646 6604 5652
rect 6656 5522 6684 6258
rect 6748 6254 6776 6666
rect 6736 6248 6788 6254
rect 6736 6190 6788 6196
rect 6748 5778 6776 6190
rect 6736 5772 6788 5778
rect 6736 5714 6788 5720
rect 6828 5704 6880 5710
rect 6828 5646 6880 5652
rect 6564 5494 6684 5522
rect 6460 5296 6512 5302
rect 6460 5238 6512 5244
rect 6460 5024 6512 5030
rect 6460 4966 6512 4972
rect 6368 3936 6420 3942
rect 6368 3878 6420 3884
rect 6380 3466 6408 3878
rect 6368 3460 6420 3466
rect 6368 3402 6420 3408
rect 6472 3233 6500 4966
rect 6564 4214 6592 5494
rect 6644 4548 6696 4554
rect 6644 4490 6696 4496
rect 6552 4208 6604 4214
rect 6552 4150 6604 4156
rect 6564 3942 6592 4150
rect 6656 4146 6684 4490
rect 6840 4282 6868 5646
rect 6920 4616 6972 4622
rect 6920 4558 6972 4564
rect 6828 4276 6880 4282
rect 6828 4218 6880 4224
rect 6644 4140 6696 4146
rect 6644 4082 6696 4088
rect 6552 3936 6604 3942
rect 6552 3878 6604 3884
rect 6458 3224 6514 3233
rect 6458 3159 6514 3168
rect 6472 2922 6500 3159
rect 5632 2916 5684 2922
rect 5632 2858 5684 2864
rect 5908 2916 5960 2922
rect 5908 2858 5960 2864
rect 6460 2916 6512 2922
rect 6460 2858 6512 2864
rect 4896 2440 4948 2446
rect 4896 2382 4948 2388
rect 4436 2304 4488 2310
rect 4436 2246 4488 2252
rect 4448 2106 4476 2246
rect 4436 2100 4488 2106
rect 4436 2042 4488 2048
rect 4908 1766 4936 2382
rect 5080 2304 5132 2310
rect 5080 2246 5132 2252
rect 5092 2038 5120 2246
rect 5080 2032 5132 2038
rect 5080 1974 5132 1980
rect 5644 1970 5672 2858
rect 6656 2774 6684 4082
rect 6736 3460 6788 3466
rect 6736 3402 6788 3408
rect 6748 3058 6776 3402
rect 6736 3052 6788 3058
rect 6736 2994 6788 3000
rect 6748 2922 6776 2994
rect 6736 2916 6788 2922
rect 6736 2858 6788 2864
rect 6840 2802 6868 4218
rect 6932 3534 6960 4558
rect 7024 4146 7052 8366
rect 7484 7886 7512 8366
rect 8128 8362 8156 8910
rect 8312 8894 8432 8922
rect 7930 8327 7986 8336
rect 8116 8356 8168 8362
rect 8116 8298 8168 8304
rect 7472 7880 7524 7886
rect 7472 7822 7524 7828
rect 7104 7200 7156 7206
rect 7104 7142 7156 7148
rect 7116 6798 7144 7142
rect 7484 6798 7512 7822
rect 7932 7812 7984 7818
rect 7932 7754 7984 7760
rect 7564 7404 7616 7410
rect 7564 7346 7616 7352
rect 7576 7002 7604 7346
rect 7944 7206 7972 7754
rect 8312 7324 8340 8894
rect 8392 8832 8444 8838
rect 8392 8774 8444 8780
rect 8404 8566 8432 8774
rect 8392 8560 8444 8566
rect 8392 8502 8444 8508
rect 8390 8392 8446 8401
rect 8390 8327 8446 8336
rect 8404 7750 8432 8327
rect 8392 7744 8444 7750
rect 8392 7686 8444 7692
rect 8312 7296 8432 7324
rect 7932 7200 7984 7206
rect 7932 7142 7984 7148
rect 7564 6996 7616 7002
rect 7564 6938 7616 6944
rect 7104 6792 7156 6798
rect 7104 6734 7156 6740
rect 7288 6792 7340 6798
rect 7288 6734 7340 6740
rect 7472 6792 7524 6798
rect 7472 6734 7524 6740
rect 7300 6118 7328 6734
rect 7288 6112 7340 6118
rect 7288 6054 7340 6060
rect 7300 5137 7328 6054
rect 7944 5710 7972 7142
rect 8300 6656 8352 6662
rect 8300 6598 8352 6604
rect 8312 6186 8340 6598
rect 8300 6180 8352 6186
rect 8300 6122 8352 6128
rect 8116 5840 8168 5846
rect 8116 5782 8168 5788
rect 7932 5704 7984 5710
rect 7932 5646 7984 5652
rect 7748 5568 7800 5574
rect 7748 5510 7800 5516
rect 7286 5128 7342 5137
rect 7286 5063 7342 5072
rect 7760 4622 7788 5510
rect 7840 5228 7892 5234
rect 7840 5170 7892 5176
rect 7748 4616 7800 4622
rect 7748 4558 7800 4564
rect 7012 4140 7064 4146
rect 7012 4082 7064 4088
rect 6920 3528 6972 3534
rect 6920 3470 6972 3476
rect 6932 3058 6960 3470
rect 6920 3052 6972 3058
rect 6920 2994 6972 3000
rect 6472 2746 6684 2774
rect 6748 2774 6868 2802
rect 5724 2304 5776 2310
rect 5724 2246 5776 2252
rect 5632 1964 5684 1970
rect 5632 1906 5684 1912
rect 4896 1760 4948 1766
rect 4896 1702 4948 1708
rect 5736 1630 5764 2246
rect 6472 2145 6500 2746
rect 6748 2514 6776 2774
rect 6736 2508 6788 2514
rect 6736 2450 6788 2456
rect 7024 2446 7052 4082
rect 7654 4040 7710 4049
rect 7654 3975 7656 3984
rect 7708 3975 7710 3984
rect 7748 4004 7800 4010
rect 7656 3946 7708 3952
rect 7748 3946 7800 3952
rect 7564 3936 7616 3942
rect 7564 3878 7616 3884
rect 7576 3602 7604 3878
rect 7564 3596 7616 3602
rect 7564 3538 7616 3544
rect 7760 3534 7788 3946
rect 7852 3534 7880 5170
rect 7748 3528 7800 3534
rect 7748 3470 7800 3476
rect 7840 3528 7892 3534
rect 7840 3470 7892 3476
rect 7380 3392 7432 3398
rect 7380 3334 7432 3340
rect 7748 3392 7800 3398
rect 7748 3334 7800 3340
rect 7392 2446 7420 3334
rect 7760 3194 7788 3334
rect 7852 3194 7880 3470
rect 7748 3188 7800 3194
rect 7748 3130 7800 3136
rect 7840 3188 7892 3194
rect 7840 3130 7892 3136
rect 7840 3052 7892 3058
rect 7840 2994 7892 3000
rect 7852 2650 7880 2994
rect 7944 2689 7972 5646
rect 8128 4729 8156 5782
rect 8208 5704 8260 5710
rect 8208 5646 8260 5652
rect 8220 5370 8248 5646
rect 8208 5364 8260 5370
rect 8208 5306 8260 5312
rect 8404 5166 8432 7296
rect 8496 5234 8524 10610
rect 8956 10062 8984 10950
rect 9692 10826 9720 12786
rect 9784 11150 9812 15438
rect 10060 12986 10088 19382
rect 10152 19378 10180 19654
rect 10140 19372 10192 19378
rect 10140 19314 10192 19320
rect 10048 12980 10100 12986
rect 10048 12922 10100 12928
rect 10048 12708 10100 12714
rect 10048 12650 10100 12656
rect 10060 12238 10088 12650
rect 9864 12232 9916 12238
rect 9864 12174 9916 12180
rect 10048 12232 10100 12238
rect 10048 12174 10100 12180
rect 9772 11144 9824 11150
rect 9772 11086 9824 11092
rect 9600 10798 9720 10826
rect 9876 10810 9904 12174
rect 10152 12170 10180 19314
rect 10244 18358 10272 21286
rect 10520 20874 10548 21626
rect 10508 20868 10560 20874
rect 10508 20810 10560 20816
rect 10416 20800 10468 20806
rect 10416 20742 10468 20748
rect 10324 18692 10376 18698
rect 10324 18634 10376 18640
rect 10336 18426 10364 18634
rect 10324 18420 10376 18426
rect 10324 18362 10376 18368
rect 10232 18352 10284 18358
rect 10232 18294 10284 18300
rect 10324 15496 10376 15502
rect 10428 15484 10456 20742
rect 10980 20074 11008 24550
rect 11532 24274 11560 25842
rect 11520 24268 11572 24274
rect 11520 24210 11572 24216
rect 11796 24132 11848 24138
rect 11796 24074 11848 24080
rect 11152 24064 11204 24070
rect 11152 24006 11204 24012
rect 11164 23730 11192 24006
rect 11152 23724 11204 23730
rect 11152 23666 11204 23672
rect 11060 22432 11112 22438
rect 11060 22374 11112 22380
rect 11072 22234 11100 22374
rect 11060 22228 11112 22234
rect 11060 22170 11112 22176
rect 10980 20058 11100 20074
rect 10980 20052 11112 20058
rect 10980 20046 11060 20052
rect 11060 19994 11112 20000
rect 11060 18216 11112 18222
rect 11060 18158 11112 18164
rect 11072 17270 11100 18158
rect 10692 17264 10744 17270
rect 10692 17206 10744 17212
rect 11060 17264 11112 17270
rect 11060 17206 11112 17212
rect 10704 16658 10732 17206
rect 10692 16652 10744 16658
rect 10692 16594 10744 16600
rect 10980 16522 11100 16538
rect 10968 16516 11100 16522
rect 11020 16510 11100 16516
rect 10968 16458 11020 16464
rect 10376 15456 10456 15484
rect 10692 15496 10744 15502
rect 10598 15464 10654 15473
rect 10324 15438 10376 15444
rect 10692 15438 10744 15444
rect 10598 15399 10654 15408
rect 10612 15366 10640 15399
rect 10600 15360 10652 15366
rect 10600 15302 10652 15308
rect 10232 15020 10284 15026
rect 10232 14962 10284 14968
rect 10140 12164 10192 12170
rect 10140 12106 10192 12112
rect 9956 12096 10008 12102
rect 10244 12084 10272 14962
rect 10704 14498 10732 15438
rect 11072 15162 11100 16510
rect 11060 15156 11112 15162
rect 11060 15098 11112 15104
rect 10428 14470 10732 14498
rect 10428 14414 10456 14470
rect 10416 14408 10468 14414
rect 10416 14350 10468 14356
rect 10508 14408 10560 14414
rect 10508 14350 10560 14356
rect 10416 14272 10468 14278
rect 10416 14214 10468 14220
rect 10428 14113 10456 14214
rect 10414 14104 10470 14113
rect 10414 14039 10470 14048
rect 10324 13864 10376 13870
rect 10324 13806 10376 13812
rect 10336 12238 10364 13806
rect 10520 12434 10548 14350
rect 10704 13734 10732 14470
rect 10968 14476 11020 14482
rect 10968 14418 11020 14424
rect 10692 13728 10744 13734
rect 10692 13670 10744 13676
rect 10704 12850 10732 13670
rect 10876 13184 10928 13190
rect 10876 13126 10928 13132
rect 10888 12986 10916 13126
rect 10876 12980 10928 12986
rect 10876 12922 10928 12928
rect 10692 12844 10744 12850
rect 10692 12786 10744 12792
rect 10428 12406 10548 12434
rect 10324 12232 10376 12238
rect 10324 12174 10376 12180
rect 10244 12056 10364 12084
rect 9956 12038 10008 12044
rect 9968 11354 9996 12038
rect 10048 11824 10100 11830
rect 10048 11766 10100 11772
rect 9956 11348 10008 11354
rect 9956 11290 10008 11296
rect 9864 10804 9916 10810
rect 9494 10704 9550 10713
rect 9494 10639 9496 10648
rect 9548 10639 9550 10648
rect 9496 10610 9548 10616
rect 9126 10568 9182 10577
rect 9126 10503 9182 10512
rect 9140 10470 9168 10503
rect 9128 10464 9180 10470
rect 9128 10406 9180 10412
rect 8944 10056 8996 10062
rect 8944 9998 8996 10004
rect 8760 9512 8812 9518
rect 8760 9454 8812 9460
rect 9600 9466 9628 10798
rect 9864 10746 9916 10752
rect 9680 10668 9732 10674
rect 9680 10610 9732 10616
rect 9692 9586 9720 10610
rect 9876 10062 9904 10746
rect 9968 10674 9996 11290
rect 9956 10668 10008 10674
rect 9956 10610 10008 10616
rect 9956 10532 10008 10538
rect 9956 10474 10008 10480
rect 9864 10056 9916 10062
rect 9864 9998 9916 10004
rect 9864 9920 9916 9926
rect 9968 9874 9996 10474
rect 10060 9897 10088 11766
rect 10232 11076 10284 11082
rect 10232 11018 10284 11024
rect 10244 10810 10272 11018
rect 10232 10804 10284 10810
rect 10232 10746 10284 10752
rect 10336 10130 10364 12056
rect 10324 10124 10376 10130
rect 10324 10066 10376 10072
rect 10140 10056 10192 10062
rect 10140 9998 10192 10004
rect 9916 9868 9996 9874
rect 9864 9862 9996 9868
rect 9876 9846 9996 9862
rect 10046 9888 10102 9897
rect 9680 9580 9732 9586
rect 9680 9522 9732 9528
rect 9772 9580 9824 9586
rect 9772 9522 9824 9528
rect 8772 8430 8800 9454
rect 9600 9438 9720 9466
rect 8760 8424 8812 8430
rect 8760 8366 8812 8372
rect 8668 8084 8720 8090
rect 8668 8026 8720 8032
rect 8576 8016 8628 8022
rect 8576 7958 8628 7964
rect 8484 5228 8536 5234
rect 8484 5170 8536 5176
rect 8392 5160 8444 5166
rect 8392 5102 8444 5108
rect 8404 4826 8432 5102
rect 8392 4820 8444 4826
rect 8392 4762 8444 4768
rect 8114 4720 8170 4729
rect 8114 4655 8170 4664
rect 8588 4146 8616 7958
rect 8680 7546 8708 8026
rect 8668 7540 8720 7546
rect 8668 7482 8720 7488
rect 8772 7478 8800 8366
rect 9312 7744 9364 7750
rect 9312 7686 9364 7692
rect 8760 7472 8812 7478
rect 8760 7414 8812 7420
rect 8772 6866 8800 7414
rect 9036 7268 9088 7274
rect 9036 7210 9088 7216
rect 8668 6860 8720 6866
rect 8668 6802 8720 6808
rect 8760 6860 8812 6866
rect 8760 6802 8812 6808
rect 8680 6322 8708 6802
rect 8668 6316 8720 6322
rect 9048 6304 9076 7210
rect 9220 6724 9272 6730
rect 9220 6666 9272 6672
rect 9232 6458 9260 6666
rect 9220 6452 9272 6458
rect 9220 6394 9272 6400
rect 8720 6276 9076 6304
rect 8668 6258 8720 6264
rect 8668 6180 8720 6186
rect 8668 6122 8720 6128
rect 8576 4140 8628 4146
rect 8576 4082 8628 4088
rect 8208 3936 8260 3942
rect 8208 3878 8260 3884
rect 8220 3738 8248 3878
rect 8208 3732 8260 3738
rect 8208 3674 8260 3680
rect 8576 3460 8628 3466
rect 8576 3402 8628 3408
rect 8588 3194 8616 3402
rect 8680 3233 8708 6122
rect 9048 5914 9076 6276
rect 9128 6316 9180 6322
rect 9128 6258 9180 6264
rect 9036 5908 9088 5914
rect 9036 5850 9088 5856
rect 9140 5234 9168 6258
rect 9220 6248 9272 6254
rect 9218 6216 9220 6225
rect 9272 6216 9274 6225
rect 9218 6151 9274 6160
rect 9128 5228 9180 5234
rect 9128 5170 9180 5176
rect 9128 5024 9180 5030
rect 9128 4966 9180 4972
rect 8944 4208 8996 4214
rect 8942 4176 8944 4185
rect 8996 4176 8998 4185
rect 8942 4111 8998 4120
rect 9036 3528 9088 3534
rect 9036 3470 9088 3476
rect 8666 3224 8722 3233
rect 8576 3188 8628 3194
rect 8666 3159 8722 3168
rect 8576 3130 8628 3136
rect 7930 2680 7986 2689
rect 7840 2644 7892 2650
rect 7930 2615 7986 2624
rect 7840 2586 7892 2592
rect 7012 2440 7064 2446
rect 7012 2382 7064 2388
rect 7380 2440 7432 2446
rect 7380 2382 7432 2388
rect 7564 2440 7616 2446
rect 7564 2382 7616 2388
rect 6736 2372 6788 2378
rect 6736 2314 6788 2320
rect 6458 2136 6514 2145
rect 6458 2071 6514 2080
rect 6748 2009 6776 2314
rect 6734 2000 6790 2009
rect 6734 1935 6790 1944
rect 7576 1698 7604 2382
rect 9048 1873 9076 3470
rect 9140 3058 9168 4966
rect 9324 3505 9352 7686
rect 9692 5370 9720 9438
rect 9784 8294 9812 9522
rect 9876 9042 9904 9846
rect 10046 9823 10102 9832
rect 9864 9036 9916 9042
rect 9864 8978 9916 8984
rect 9772 8288 9824 8294
rect 9772 8230 9824 8236
rect 9772 7948 9824 7954
rect 9772 7890 9824 7896
rect 9784 7546 9812 7890
rect 9772 7540 9824 7546
rect 9772 7482 9824 7488
rect 9784 6458 9812 7482
rect 9772 6452 9824 6458
rect 9824 6412 9904 6440
rect 9772 6394 9824 6400
rect 9680 5364 9732 5370
rect 9680 5306 9732 5312
rect 9772 5364 9824 5370
rect 9772 5306 9824 5312
rect 9588 5160 9640 5166
rect 9588 5102 9640 5108
rect 9600 3534 9628 5102
rect 9784 4826 9812 5306
rect 9876 5030 9904 6412
rect 9956 6112 10008 6118
rect 9956 6054 10008 6060
rect 9864 5024 9916 5030
rect 9864 4966 9916 4972
rect 9772 4820 9824 4826
rect 9772 4762 9824 4768
rect 9968 4593 9996 6054
rect 9770 4584 9826 4593
rect 9770 4519 9826 4528
rect 9954 4584 10010 4593
rect 9954 4519 10010 4528
rect 9784 4486 9812 4519
rect 9772 4480 9824 4486
rect 9772 4422 9824 4428
rect 9680 4276 9732 4282
rect 9680 4218 9732 4224
rect 9692 4146 9720 4218
rect 9864 4208 9916 4214
rect 9864 4150 9916 4156
rect 9680 4140 9732 4146
rect 9680 4082 9732 4088
rect 9876 3534 9904 4150
rect 9588 3528 9640 3534
rect 9310 3496 9366 3505
rect 9588 3470 9640 3476
rect 9864 3528 9916 3534
rect 9864 3470 9916 3476
rect 9310 3431 9366 3440
rect 9600 3126 9628 3470
rect 9588 3120 9640 3126
rect 9588 3062 9640 3068
rect 9128 3052 9180 3058
rect 9128 2994 9180 3000
rect 9586 2816 9642 2825
rect 9586 2751 9642 2760
rect 9496 2644 9548 2650
rect 9496 2586 9548 2592
rect 9508 2446 9536 2586
rect 9600 2446 9628 2751
rect 9496 2440 9548 2446
rect 9496 2382 9548 2388
rect 9588 2440 9640 2446
rect 10060 2417 10088 9823
rect 10152 8974 10180 9998
rect 10324 9988 10376 9994
rect 10324 9930 10376 9936
rect 10336 9586 10364 9930
rect 10324 9580 10376 9586
rect 10324 9522 10376 9528
rect 10336 9178 10364 9522
rect 10324 9172 10376 9178
rect 10324 9114 10376 9120
rect 10140 8968 10192 8974
rect 10140 8910 10192 8916
rect 10232 7200 10284 7206
rect 10232 7142 10284 7148
rect 10140 4548 10192 4554
rect 10140 4490 10192 4496
rect 9588 2382 9640 2388
rect 10046 2408 10102 2417
rect 10046 2343 10102 2352
rect 10060 2310 10088 2343
rect 9588 2304 9640 2310
rect 9588 2246 9640 2252
rect 10048 2304 10100 2310
rect 10048 2246 10100 2252
rect 9034 1864 9090 1873
rect 9034 1799 9090 1808
rect 7564 1692 7616 1698
rect 7564 1634 7616 1640
rect 5724 1624 5776 1630
rect 5724 1566 5776 1572
rect 9600 1222 9628 2246
rect 10152 2038 10180 4490
rect 10244 4282 10272 7142
rect 10428 6662 10456 12406
rect 10876 11552 10928 11558
rect 10876 11494 10928 11500
rect 10508 11076 10560 11082
rect 10508 11018 10560 11024
rect 10520 9586 10548 11018
rect 10782 10704 10838 10713
rect 10782 10639 10784 10648
rect 10836 10639 10838 10648
rect 10784 10610 10836 10616
rect 10888 10470 10916 11494
rect 10876 10464 10928 10470
rect 10876 10406 10928 10412
rect 10692 10124 10744 10130
rect 10692 10066 10744 10072
rect 10508 9580 10560 9586
rect 10508 9522 10560 9528
rect 10704 8974 10732 10066
rect 10784 9580 10836 9586
rect 10784 9522 10836 9528
rect 10692 8968 10744 8974
rect 10692 8910 10744 8916
rect 10796 8838 10824 9522
rect 10784 8832 10836 8838
rect 10784 8774 10836 8780
rect 10692 8288 10744 8294
rect 10692 8230 10744 8236
rect 10416 6656 10468 6662
rect 10416 6598 10468 6604
rect 10428 6390 10456 6598
rect 10600 6452 10652 6458
rect 10600 6394 10652 6400
rect 10416 6384 10468 6390
rect 10416 6326 10468 6332
rect 10416 5704 10468 5710
rect 10416 5646 10468 5652
rect 10324 4616 10376 4622
rect 10324 4558 10376 4564
rect 10232 4276 10284 4282
rect 10232 4218 10284 4224
rect 10232 4140 10284 4146
rect 10232 4082 10284 4088
rect 10244 3346 10272 4082
rect 10336 4049 10364 4558
rect 10322 4040 10378 4049
rect 10322 3975 10378 3984
rect 10244 3318 10364 3346
rect 10232 2440 10284 2446
rect 10232 2382 10284 2388
rect 10140 2032 10192 2038
rect 10140 1974 10192 1980
rect 10244 1970 10272 2382
rect 10232 1964 10284 1970
rect 10232 1906 10284 1912
rect 10336 1426 10364 3318
rect 10428 3194 10456 5646
rect 10508 5024 10560 5030
rect 10508 4966 10560 4972
rect 10520 4146 10548 4966
rect 10612 4826 10640 6394
rect 10600 4820 10652 4826
rect 10600 4762 10652 4768
rect 10508 4140 10560 4146
rect 10508 4082 10560 4088
rect 10598 4040 10654 4049
rect 10598 3975 10654 3984
rect 10506 3904 10562 3913
rect 10506 3839 10562 3848
rect 10416 3188 10468 3194
rect 10416 3130 10468 3136
rect 10416 2984 10468 2990
rect 10416 2926 10468 2932
rect 10428 2446 10456 2926
rect 10416 2440 10468 2446
rect 10416 2382 10468 2388
rect 10520 2378 10548 3839
rect 10508 2372 10560 2378
rect 10508 2314 10560 2320
rect 10324 1420 10376 1426
rect 10324 1362 10376 1368
rect 9588 1216 9640 1222
rect 9588 1158 9640 1164
rect 10612 800 10640 3975
rect 10704 3534 10732 8230
rect 10876 6384 10928 6390
rect 10876 6326 10928 6332
rect 10888 6089 10916 6326
rect 10874 6080 10930 6089
rect 10874 6015 10930 6024
rect 10784 5568 10836 5574
rect 10784 5510 10836 5516
rect 10692 3528 10744 3534
rect 10692 3470 10744 3476
rect 10692 3392 10744 3398
rect 10692 3334 10744 3340
rect 10704 800 10732 3334
rect 10796 800 10824 5510
rect 10980 5370 11008 14418
rect 11164 14414 11192 23666
rect 11808 23322 11836 24074
rect 12072 23520 12124 23526
rect 12072 23462 12124 23468
rect 11796 23316 11848 23322
rect 11796 23258 11848 23264
rect 11336 23112 11388 23118
rect 11336 23054 11388 23060
rect 11348 22506 11376 23054
rect 11336 22500 11388 22506
rect 11336 22442 11388 22448
rect 12084 21962 12112 23462
rect 12348 23180 12400 23186
rect 12348 23122 12400 23128
rect 12624 23180 12676 23186
rect 12808 23180 12860 23186
rect 12676 23140 12808 23168
rect 12624 23122 12676 23128
rect 12808 23122 12860 23128
rect 12256 23112 12308 23118
rect 12256 23054 12308 23060
rect 12268 22778 12296 23054
rect 12256 22772 12308 22778
rect 12256 22714 12308 22720
rect 12360 22658 12388 23122
rect 12440 23112 12492 23118
rect 12440 23054 12492 23060
rect 12268 22630 12388 22658
rect 12072 21956 12124 21962
rect 12072 21898 12124 21904
rect 12268 21622 12296 22630
rect 12452 22030 12480 23054
rect 12716 22772 12768 22778
rect 12716 22714 12768 22720
rect 12532 22636 12584 22642
rect 12532 22578 12584 22584
rect 12440 22024 12492 22030
rect 12440 21966 12492 21972
rect 12348 21956 12400 21962
rect 12348 21898 12400 21904
rect 12256 21616 12308 21622
rect 12256 21558 12308 21564
rect 11704 21548 11756 21554
rect 11704 21490 11756 21496
rect 11716 21457 11744 21490
rect 12256 21480 12308 21486
rect 11702 21448 11758 21457
rect 12256 21422 12308 21428
rect 11702 21383 11758 21392
rect 11704 21344 11756 21350
rect 11704 21286 11756 21292
rect 11716 20942 11744 21286
rect 11612 20936 11664 20942
rect 11612 20878 11664 20884
rect 11704 20936 11756 20942
rect 11704 20878 11756 20884
rect 11624 19854 11652 20878
rect 12268 20602 12296 21422
rect 12256 20596 12308 20602
rect 12256 20538 12308 20544
rect 11612 19848 11664 19854
rect 11612 19790 11664 19796
rect 12164 19848 12216 19854
rect 12164 19790 12216 19796
rect 12176 19378 12204 19790
rect 12164 19372 12216 19378
rect 12164 19314 12216 19320
rect 11980 19304 12032 19310
rect 11980 19246 12032 19252
rect 11704 18624 11756 18630
rect 11704 18566 11756 18572
rect 11716 17678 11744 18566
rect 11992 18193 12020 19246
rect 11978 18184 12034 18193
rect 11978 18119 12034 18128
rect 11704 17672 11756 17678
rect 11704 17614 11756 17620
rect 11612 17604 11664 17610
rect 11612 17546 11664 17552
rect 11244 17536 11296 17542
rect 11296 17484 11376 17490
rect 11244 17478 11376 17484
rect 11256 17462 11376 17478
rect 11244 16584 11296 16590
rect 11244 16526 11296 16532
rect 11256 16250 11284 16526
rect 11244 16244 11296 16250
rect 11244 16186 11296 16192
rect 11348 15502 11376 17462
rect 11520 17196 11572 17202
rect 11520 17138 11572 17144
rect 11428 17128 11480 17134
rect 11428 17070 11480 17076
rect 11440 16998 11468 17070
rect 11428 16992 11480 16998
rect 11428 16934 11480 16940
rect 11428 16584 11480 16590
rect 11426 16552 11428 16561
rect 11480 16552 11482 16561
rect 11426 16487 11482 16496
rect 11532 16114 11560 17138
rect 11520 16108 11572 16114
rect 11520 16050 11572 16056
rect 11336 15496 11388 15502
rect 11336 15438 11388 15444
rect 11348 15366 11376 15438
rect 11336 15360 11388 15366
rect 11336 15302 11388 15308
rect 11532 14634 11560 16050
rect 11624 15502 11652 17546
rect 11716 16810 11744 17614
rect 11796 17536 11848 17542
rect 11796 17478 11848 17484
rect 11808 17202 11836 17478
rect 11992 17202 12020 18119
rect 12176 17746 12204 19314
rect 12164 17740 12216 17746
rect 12164 17682 12216 17688
rect 11796 17196 11848 17202
rect 11796 17138 11848 17144
rect 11980 17196 12032 17202
rect 11980 17138 12032 17144
rect 12072 17128 12124 17134
rect 12072 17070 12124 17076
rect 11716 16782 11928 16810
rect 11796 16448 11848 16454
rect 11796 16390 11848 16396
rect 11808 16182 11836 16390
rect 11796 16176 11848 16182
rect 11796 16118 11848 16124
rect 11704 16108 11756 16114
rect 11704 16050 11756 16056
rect 11612 15496 11664 15502
rect 11612 15438 11664 15444
rect 11716 15434 11744 16050
rect 11808 15570 11836 16118
rect 11900 15706 11928 16782
rect 12084 16046 12112 17070
rect 12176 16658 12204 17682
rect 12256 17604 12308 17610
rect 12256 17546 12308 17552
rect 12268 17338 12296 17546
rect 12256 17332 12308 17338
rect 12256 17274 12308 17280
rect 12360 17218 12388 21898
rect 12452 21554 12480 21966
rect 12440 21548 12492 21554
rect 12440 21490 12492 21496
rect 12544 20534 12572 22578
rect 12624 21684 12676 21690
rect 12624 21626 12676 21632
rect 12532 20528 12584 20534
rect 12532 20470 12584 20476
rect 12268 17190 12388 17218
rect 12164 16652 12216 16658
rect 12164 16594 12216 16600
rect 12072 16040 12124 16046
rect 12072 15982 12124 15988
rect 11980 15972 12032 15978
rect 11980 15914 12032 15920
rect 11992 15706 12020 15914
rect 11888 15700 11940 15706
rect 11888 15642 11940 15648
rect 11980 15700 12032 15706
rect 11980 15642 12032 15648
rect 11900 15609 11928 15642
rect 11886 15600 11942 15609
rect 11796 15564 11848 15570
rect 11886 15535 11942 15544
rect 11796 15506 11848 15512
rect 11704 15428 11756 15434
rect 11704 15370 11756 15376
rect 11704 15088 11756 15094
rect 11704 15030 11756 15036
rect 11716 14958 11744 15030
rect 11796 15020 11848 15026
rect 11796 14962 11848 14968
rect 11980 15020 12032 15026
rect 11980 14962 12032 14968
rect 11704 14952 11756 14958
rect 11704 14894 11756 14900
rect 11532 14606 11652 14634
rect 11152 14408 11204 14414
rect 11152 14350 11204 14356
rect 11244 14408 11296 14414
rect 11244 14350 11296 14356
rect 11256 13870 11284 14350
rect 11428 14340 11480 14346
rect 11428 14282 11480 14288
rect 11244 13864 11296 13870
rect 11244 13806 11296 13812
rect 11256 13297 11284 13806
rect 11336 13456 11388 13462
rect 11336 13398 11388 13404
rect 11242 13288 11298 13297
rect 11242 13223 11298 13232
rect 11348 12986 11376 13398
rect 11440 13326 11468 14282
rect 11520 13864 11572 13870
rect 11520 13806 11572 13812
rect 11532 13394 11560 13806
rect 11520 13388 11572 13394
rect 11520 13330 11572 13336
rect 11428 13320 11480 13326
rect 11428 13262 11480 13268
rect 11336 12980 11388 12986
rect 11336 12922 11388 12928
rect 11440 12850 11468 13262
rect 11624 12918 11652 14606
rect 11808 14278 11836 14962
rect 11992 14822 12020 14962
rect 11980 14816 12032 14822
rect 11980 14758 12032 14764
rect 11796 14272 11848 14278
rect 11796 14214 11848 14220
rect 11704 12980 11756 12986
rect 11704 12922 11756 12928
rect 12072 12980 12124 12986
rect 12072 12922 12124 12928
rect 11612 12912 11664 12918
rect 11612 12854 11664 12860
rect 11428 12844 11480 12850
rect 11428 12786 11480 12792
rect 11336 12232 11388 12238
rect 11336 12174 11388 12180
rect 11060 12164 11112 12170
rect 11060 12106 11112 12112
rect 11072 11558 11100 12106
rect 11348 11762 11376 12174
rect 11336 11756 11388 11762
rect 11336 11698 11388 11704
rect 11060 11552 11112 11558
rect 11058 11520 11060 11529
rect 11112 11520 11114 11529
rect 11058 11455 11114 11464
rect 11348 11082 11376 11698
rect 11520 11620 11572 11626
rect 11520 11562 11572 11568
rect 11428 11280 11480 11286
rect 11428 11222 11480 11228
rect 11336 11076 11388 11082
rect 11336 11018 11388 11024
rect 11152 10668 11204 10674
rect 11152 10610 11204 10616
rect 11164 10062 11192 10610
rect 11440 10130 11468 11222
rect 11532 11082 11560 11562
rect 11624 11286 11652 12854
rect 11716 12238 11744 12922
rect 12084 12238 12112 12922
rect 12268 12646 12296 17190
rect 12636 16561 12664 21626
rect 12622 16552 12678 16561
rect 12622 16487 12678 16496
rect 12624 15496 12676 15502
rect 12624 15438 12676 15444
rect 12636 15162 12664 15438
rect 12624 15156 12676 15162
rect 12624 15098 12676 15104
rect 12532 15020 12584 15026
rect 12532 14962 12584 14968
rect 12544 14618 12572 14962
rect 12532 14612 12584 14618
rect 12532 14554 12584 14560
rect 12348 14408 12400 14414
rect 12636 14396 12664 15098
rect 12728 15026 12756 22714
rect 12808 22432 12860 22438
rect 12808 22374 12860 22380
rect 12820 22166 12848 22374
rect 12808 22160 12860 22166
rect 12808 22102 12860 22108
rect 12912 21622 12940 26318
rect 13004 23662 13032 26862
rect 13268 26376 13320 26382
rect 13268 26318 13320 26324
rect 13280 25702 13308 26318
rect 13268 25696 13320 25702
rect 13268 25638 13320 25644
rect 13280 24750 13308 25638
rect 13820 25152 13872 25158
rect 13820 25094 13872 25100
rect 13268 24744 13320 24750
rect 13268 24686 13320 24692
rect 13082 24440 13138 24449
rect 13082 24375 13084 24384
rect 13136 24375 13138 24384
rect 13084 24346 13136 24352
rect 12992 23656 13044 23662
rect 12992 23598 13044 23604
rect 13096 23202 13124 24346
rect 13004 23174 13124 23202
rect 13004 22778 13032 23174
rect 13084 23112 13136 23118
rect 13084 23054 13136 23060
rect 13096 22778 13124 23054
rect 12992 22772 13044 22778
rect 12992 22714 13044 22720
rect 13084 22772 13136 22778
rect 13084 22714 13136 22720
rect 13176 22092 13228 22098
rect 13176 22034 13228 22040
rect 12900 21616 12952 21622
rect 12900 21558 12952 21564
rect 12912 21457 12940 21558
rect 13188 21554 13216 22034
rect 13176 21548 13228 21554
rect 13176 21490 13228 21496
rect 12898 21448 12954 21457
rect 12898 21383 12954 21392
rect 12808 15428 12860 15434
rect 12808 15370 12860 15376
rect 12716 15020 12768 15026
rect 12716 14962 12768 14968
rect 12716 14408 12768 14414
rect 12400 14368 12480 14396
rect 12636 14368 12716 14396
rect 12348 14350 12400 14356
rect 12452 13394 12480 14368
rect 12716 14350 12768 14356
rect 12728 13410 12756 14350
rect 12820 13870 12848 15370
rect 12808 13864 12860 13870
rect 12808 13806 12860 13812
rect 12912 13705 12940 21383
rect 12992 20800 13044 20806
rect 12992 20742 13044 20748
rect 13004 20602 13032 20742
rect 12992 20596 13044 20602
rect 12992 20538 13044 20544
rect 13004 20398 13032 20538
rect 12992 20392 13044 20398
rect 12992 20334 13044 20340
rect 13188 19310 13216 21490
rect 13280 19922 13308 24686
rect 13544 24132 13596 24138
rect 13544 24074 13596 24080
rect 13360 23656 13412 23662
rect 13360 23598 13412 23604
rect 13372 23118 13400 23598
rect 13556 23322 13584 24074
rect 13832 23866 13860 25094
rect 13820 23860 13872 23866
rect 13820 23802 13872 23808
rect 13544 23316 13596 23322
rect 13544 23258 13596 23264
rect 13360 23112 13412 23118
rect 13360 23054 13412 23060
rect 13452 22228 13504 22234
rect 13452 22170 13504 22176
rect 13268 19916 13320 19922
rect 13268 19858 13320 19864
rect 13176 19304 13228 19310
rect 13176 19246 13228 19252
rect 13464 18766 13492 22170
rect 14016 20942 14044 27270
rect 14108 26994 14136 27270
rect 14372 27124 14424 27130
rect 14372 27066 14424 27072
rect 14096 26988 14148 26994
rect 14096 26930 14148 26936
rect 14108 26450 14136 26930
rect 14384 26790 14412 27066
rect 14752 27062 14780 27406
rect 14740 27056 14792 27062
rect 14740 26998 14792 27004
rect 14556 26920 14608 26926
rect 14556 26862 14608 26868
rect 14372 26784 14424 26790
rect 14372 26726 14424 26732
rect 14280 26580 14332 26586
rect 14280 26522 14332 26528
rect 14096 26444 14148 26450
rect 14096 26386 14148 26392
rect 14188 26376 14240 26382
rect 14188 26318 14240 26324
rect 14200 26042 14228 26318
rect 14188 26036 14240 26042
rect 14188 25978 14240 25984
rect 14292 25702 14320 26522
rect 14280 25696 14332 25702
rect 14280 25638 14332 25644
rect 14292 23662 14320 25638
rect 14568 24818 14596 26862
rect 14556 24812 14608 24818
rect 14556 24754 14608 24760
rect 14648 24200 14700 24206
rect 14648 24142 14700 24148
rect 14280 23656 14332 23662
rect 14280 23598 14332 23604
rect 14292 22778 14320 23598
rect 14372 23520 14424 23526
rect 14372 23462 14424 23468
rect 14384 23118 14412 23462
rect 14660 23118 14688 24142
rect 14372 23112 14424 23118
rect 14372 23054 14424 23060
rect 14648 23112 14700 23118
rect 14648 23054 14700 23060
rect 14280 22772 14332 22778
rect 14280 22714 14332 22720
rect 14384 22094 14412 23054
rect 14752 22234 14780 26998
rect 16304 26852 16356 26858
rect 16304 26794 16356 26800
rect 15568 26376 15620 26382
rect 15568 26318 15620 26324
rect 15384 25900 15436 25906
rect 15384 25842 15436 25848
rect 15396 25498 15424 25842
rect 15384 25492 15436 25498
rect 15384 25434 15436 25440
rect 14924 25288 14976 25294
rect 14924 25230 14976 25236
rect 14740 22228 14792 22234
rect 14740 22170 14792 22176
rect 14384 22066 14504 22094
rect 14004 20936 14056 20942
rect 14004 20878 14056 20884
rect 14476 19786 14504 22066
rect 14936 21962 14964 25230
rect 15292 25220 15344 25226
rect 15292 25162 15344 25168
rect 15304 24886 15332 25162
rect 15476 24948 15528 24954
rect 15476 24890 15528 24896
rect 15292 24880 15344 24886
rect 15292 24822 15344 24828
rect 15016 24812 15068 24818
rect 15016 24754 15068 24760
rect 15200 24812 15252 24818
rect 15200 24754 15252 24760
rect 15028 22234 15056 24754
rect 15212 23662 15240 24754
rect 15292 24404 15344 24410
rect 15292 24346 15344 24352
rect 15200 23656 15252 23662
rect 15200 23598 15252 23604
rect 15108 23112 15160 23118
rect 15108 23054 15160 23060
rect 15016 22228 15068 22234
rect 15016 22170 15068 22176
rect 15120 22030 15148 23054
rect 15200 22636 15252 22642
rect 15200 22578 15252 22584
rect 15108 22024 15160 22030
rect 15108 21966 15160 21972
rect 14924 21956 14976 21962
rect 14924 21898 14976 21904
rect 15212 21894 15240 22578
rect 15304 22574 15332 24346
rect 15292 22568 15344 22574
rect 15292 22510 15344 22516
rect 15200 21888 15252 21894
rect 15200 21830 15252 21836
rect 14832 21344 14884 21350
rect 14832 21286 14884 21292
rect 14648 20936 14700 20942
rect 14648 20878 14700 20884
rect 14556 20256 14608 20262
rect 14556 20198 14608 20204
rect 14464 19780 14516 19786
rect 14464 19722 14516 19728
rect 14372 19712 14424 19718
rect 14372 19654 14424 19660
rect 14384 19446 14412 19654
rect 14372 19440 14424 19446
rect 14372 19382 14424 19388
rect 14096 19372 14148 19378
rect 14096 19314 14148 19320
rect 13912 19168 13964 19174
rect 13912 19110 13964 19116
rect 13924 18970 13952 19110
rect 14108 18970 14136 19314
rect 14464 19304 14516 19310
rect 14464 19246 14516 19252
rect 13912 18964 13964 18970
rect 13912 18906 13964 18912
rect 14096 18964 14148 18970
rect 14096 18906 14148 18912
rect 14476 18766 14504 19246
rect 14568 18766 14596 20198
rect 13452 18760 13504 18766
rect 13452 18702 13504 18708
rect 14188 18760 14240 18766
rect 14188 18702 14240 18708
rect 14464 18760 14516 18766
rect 14464 18702 14516 18708
rect 14556 18760 14608 18766
rect 14556 18702 14608 18708
rect 14096 18216 14148 18222
rect 14096 18158 14148 18164
rect 14004 18080 14056 18086
rect 14004 18022 14056 18028
rect 13636 17060 13688 17066
rect 13636 17002 13688 17008
rect 13084 16516 13136 16522
rect 13084 16458 13136 16464
rect 12992 15632 13044 15638
rect 12992 15574 13044 15580
rect 13004 15026 13032 15574
rect 13096 15502 13124 16458
rect 13648 16182 13676 17002
rect 13636 16176 13688 16182
rect 13636 16118 13688 16124
rect 13084 15496 13136 15502
rect 13084 15438 13136 15444
rect 13176 15428 13228 15434
rect 13176 15370 13228 15376
rect 13188 15094 13216 15370
rect 13544 15360 13596 15366
rect 13544 15302 13596 15308
rect 13176 15088 13228 15094
rect 13176 15030 13228 15036
rect 12992 15020 13044 15026
rect 12992 14962 13044 14968
rect 13004 14822 13032 14962
rect 12992 14816 13044 14822
rect 12992 14758 13044 14764
rect 13004 13938 13032 14758
rect 13452 14272 13504 14278
rect 13452 14214 13504 14220
rect 13464 13938 13492 14214
rect 12992 13932 13044 13938
rect 12992 13874 13044 13880
rect 13452 13932 13504 13938
rect 13452 13874 13504 13880
rect 13268 13796 13320 13802
rect 13268 13738 13320 13744
rect 12898 13696 12954 13705
rect 12898 13631 12954 13640
rect 12898 13424 12954 13433
rect 12440 13388 12492 13394
rect 12728 13382 12898 13410
rect 12898 13359 12954 13368
rect 12440 13330 12492 13336
rect 12912 13326 12940 13359
rect 12900 13320 12952 13326
rect 12900 13262 12952 13268
rect 13280 12986 13308 13738
rect 13452 13388 13504 13394
rect 13452 13330 13504 13336
rect 13268 12980 13320 12986
rect 13268 12922 13320 12928
rect 12530 12880 12586 12889
rect 12530 12815 12532 12824
rect 12584 12815 12586 12824
rect 12532 12786 12584 12792
rect 12256 12640 12308 12646
rect 12256 12582 12308 12588
rect 12544 12434 12572 12786
rect 13280 12442 13308 12922
rect 13360 12844 13412 12850
rect 13360 12786 13412 12792
rect 13268 12436 13320 12442
rect 12544 12406 12664 12434
rect 11704 12232 11756 12238
rect 11704 12174 11756 12180
rect 12072 12232 12124 12238
rect 12072 12174 12124 12180
rect 11612 11280 11664 11286
rect 11612 11222 11664 11228
rect 11612 11144 11664 11150
rect 11612 11086 11664 11092
rect 11520 11076 11572 11082
rect 11520 11018 11572 11024
rect 11624 10606 11652 11086
rect 11716 10742 11744 12174
rect 12256 12164 12308 12170
rect 12256 12106 12308 12112
rect 12072 11552 12124 11558
rect 12072 11494 12124 11500
rect 11888 11144 11940 11150
rect 11888 11086 11940 11092
rect 11704 10736 11756 10742
rect 11704 10678 11756 10684
rect 11796 10736 11848 10742
rect 11796 10678 11848 10684
rect 11612 10600 11664 10606
rect 11612 10542 11664 10548
rect 11428 10124 11480 10130
rect 11428 10066 11480 10072
rect 11152 10056 11204 10062
rect 11152 9998 11204 10004
rect 11164 9586 11192 9998
rect 11428 9648 11480 9654
rect 11428 9590 11480 9596
rect 11152 9580 11204 9586
rect 11152 9522 11204 9528
rect 11440 9382 11468 9590
rect 11428 9376 11480 9382
rect 11428 9318 11480 9324
rect 11624 9042 11652 10542
rect 11808 9450 11836 10678
rect 11900 10674 11928 11086
rect 12084 10674 12112 11494
rect 12268 11132 12296 12106
rect 12636 11558 12664 12406
rect 13268 12378 13320 12384
rect 12806 12200 12862 12209
rect 12806 12135 12862 12144
rect 12820 12102 12848 12135
rect 12808 12096 12860 12102
rect 12808 12038 12860 12044
rect 13176 11824 13228 11830
rect 13176 11766 13228 11772
rect 12624 11552 12676 11558
rect 12624 11494 12676 11500
rect 12440 11144 12492 11150
rect 12268 11104 12440 11132
rect 12360 10742 12388 11104
rect 12440 11086 12492 11092
rect 12348 10736 12400 10742
rect 12348 10678 12400 10684
rect 11888 10668 11940 10674
rect 11888 10610 11940 10616
rect 12072 10668 12124 10674
rect 12072 10610 12124 10616
rect 12256 10668 12308 10674
rect 12256 10610 12308 10616
rect 12268 10266 12296 10610
rect 12256 10260 12308 10266
rect 12256 10202 12308 10208
rect 11888 10056 11940 10062
rect 11888 9998 11940 10004
rect 12256 10056 12308 10062
rect 12256 9998 12308 10004
rect 11900 9674 11928 9998
rect 12268 9722 12296 9998
rect 12256 9716 12308 9722
rect 11900 9646 12020 9674
rect 12256 9658 12308 9664
rect 11992 9586 12020 9646
rect 11980 9580 12032 9586
rect 11980 9522 12032 9528
rect 11796 9444 11848 9450
rect 11796 9386 11848 9392
rect 12532 9444 12584 9450
rect 12532 9386 12584 9392
rect 11808 9110 11836 9386
rect 12164 9376 12216 9382
rect 12164 9318 12216 9324
rect 11796 9104 11848 9110
rect 11796 9046 11848 9052
rect 11612 9036 11664 9042
rect 11612 8978 11664 8984
rect 12176 8974 12204 9318
rect 12164 8968 12216 8974
rect 11058 8936 11114 8945
rect 12164 8910 12216 8916
rect 11058 8871 11114 8880
rect 11072 7041 11100 8871
rect 11152 8832 11204 8838
rect 11150 8800 11152 8809
rect 11204 8800 11206 8809
rect 11150 8735 11206 8744
rect 11152 8016 11204 8022
rect 11152 7958 11204 7964
rect 11164 7478 11192 7958
rect 12256 7812 12308 7818
rect 12256 7754 12308 7760
rect 12268 7546 12296 7754
rect 12256 7540 12308 7546
rect 12256 7482 12308 7488
rect 11152 7472 11204 7478
rect 11152 7414 11204 7420
rect 11702 7440 11758 7449
rect 11520 7404 11572 7410
rect 11702 7375 11704 7384
rect 11520 7346 11572 7352
rect 11756 7375 11758 7384
rect 11704 7346 11756 7352
rect 11336 7200 11388 7206
rect 11336 7142 11388 7148
rect 11058 7032 11114 7041
rect 11348 7002 11376 7142
rect 11058 6967 11114 6976
rect 11336 6996 11388 7002
rect 11336 6938 11388 6944
rect 11348 6798 11376 6938
rect 11532 6934 11560 7346
rect 12544 7342 12572 9386
rect 11612 7336 11664 7342
rect 11612 7278 11664 7284
rect 12532 7336 12584 7342
rect 12532 7278 12584 7284
rect 11624 7002 11652 7278
rect 12544 7154 12572 7278
rect 12452 7126 12572 7154
rect 12452 7018 12480 7126
rect 12360 7002 12480 7018
rect 11612 6996 11664 7002
rect 11612 6938 11664 6944
rect 12348 6996 12480 7002
rect 12400 6990 12480 6996
rect 12532 6996 12584 7002
rect 12348 6938 12400 6944
rect 12532 6938 12584 6944
rect 11520 6928 11572 6934
rect 11426 6896 11482 6905
rect 12256 6928 12308 6934
rect 11520 6870 11572 6876
rect 11978 6896 12034 6905
rect 11426 6831 11482 6840
rect 12256 6870 12308 6876
rect 11978 6831 12034 6840
rect 11440 6798 11468 6831
rect 11060 6792 11112 6798
rect 11060 6734 11112 6740
rect 11336 6792 11388 6798
rect 11336 6734 11388 6740
rect 11428 6792 11480 6798
rect 11428 6734 11480 6740
rect 11072 6322 11100 6734
rect 11992 6322 12020 6831
rect 11060 6316 11112 6322
rect 11980 6316 12032 6322
rect 11060 6258 11112 6264
rect 11808 6276 11980 6304
rect 11072 5953 11100 6258
rect 11244 6248 11296 6254
rect 11244 6190 11296 6196
rect 11058 5944 11114 5953
rect 11058 5879 11114 5888
rect 10968 5364 11020 5370
rect 10968 5306 11020 5312
rect 11256 4826 11284 6190
rect 11428 6180 11480 6186
rect 11428 6122 11480 6128
rect 11244 4820 11296 4826
rect 11244 4762 11296 4768
rect 11152 4684 11204 4690
rect 11152 4626 11204 4632
rect 10876 4548 10928 4554
rect 10876 4490 10928 4496
rect 10888 3641 10916 4490
rect 11060 4140 11112 4146
rect 11060 4082 11112 4088
rect 10966 4040 11022 4049
rect 10966 3975 10968 3984
rect 11020 3975 11022 3984
rect 10968 3946 11020 3952
rect 10874 3632 10930 3641
rect 11072 3602 11100 4082
rect 10874 3567 10930 3576
rect 11060 3596 11112 3602
rect 11060 3538 11112 3544
rect 10876 3528 10928 3534
rect 10876 3470 10928 3476
rect 10888 2145 10916 3470
rect 11060 3392 11112 3398
rect 11060 3334 11112 3340
rect 10874 2136 10930 2145
rect 10874 2071 10930 2080
rect 10876 1760 10928 1766
rect 10876 1702 10928 1708
rect 10888 800 10916 1702
rect 10968 1420 11020 1426
rect 10968 1362 11020 1368
rect 10980 800 11008 1362
rect 11072 800 11100 3334
rect 11164 1358 11192 4626
rect 11256 4622 11284 4762
rect 11334 4720 11390 4729
rect 11334 4655 11390 4664
rect 11244 4616 11296 4622
rect 11244 4558 11296 4564
rect 11348 4486 11376 4655
rect 11336 4480 11388 4486
rect 11336 4422 11388 4428
rect 11440 4264 11468 6122
rect 11612 6112 11664 6118
rect 11612 6054 11664 6060
rect 11520 5568 11572 5574
rect 11520 5510 11572 5516
rect 11348 4236 11468 4264
rect 11244 3936 11296 3942
rect 11348 3913 11376 4236
rect 11426 4176 11482 4185
rect 11426 4111 11482 4120
rect 11244 3878 11296 3884
rect 11334 3904 11390 3913
rect 11256 3398 11284 3878
rect 11334 3839 11390 3848
rect 11336 3732 11388 3738
rect 11336 3674 11388 3680
rect 11244 3392 11296 3398
rect 11244 3334 11296 3340
rect 11244 3120 11296 3126
rect 11244 3062 11296 3068
rect 11152 1352 11204 1358
rect 11152 1294 11204 1300
rect 11152 1216 11204 1222
rect 11152 1158 11204 1164
rect 11164 800 11192 1158
rect 11256 800 11284 3062
rect 11348 800 11376 3674
rect 11440 1442 11468 4111
rect 11532 3618 11560 5510
rect 11624 5370 11652 6054
rect 11808 5710 11836 6276
rect 11980 6258 12032 6264
rect 12164 6316 12216 6322
rect 12164 6258 12216 6264
rect 12072 6112 12124 6118
rect 12072 6054 12124 6060
rect 11796 5704 11848 5710
rect 11796 5646 11848 5652
rect 11980 5568 12032 5574
rect 11980 5510 12032 5516
rect 11612 5364 11664 5370
rect 11612 5306 11664 5312
rect 11992 5234 12020 5510
rect 11704 5228 11756 5234
rect 11704 5170 11756 5176
rect 11980 5228 12032 5234
rect 11980 5170 12032 5176
rect 11716 5137 11744 5170
rect 11702 5128 11758 5137
rect 11702 5063 11704 5072
rect 11756 5063 11758 5072
rect 11704 5034 11756 5040
rect 11716 5003 11744 5034
rect 11978 4992 12034 5001
rect 11978 4927 12034 4936
rect 11612 4752 11664 4758
rect 11612 4694 11664 4700
rect 11624 3738 11652 4694
rect 11992 4622 12020 4927
rect 12084 4690 12112 6054
rect 12176 5953 12204 6258
rect 12162 5944 12218 5953
rect 12162 5879 12218 5888
rect 12176 5710 12204 5879
rect 12164 5704 12216 5710
rect 12164 5646 12216 5652
rect 12162 5400 12218 5409
rect 12162 5335 12218 5344
rect 12176 5234 12204 5335
rect 12268 5234 12296 6870
rect 12440 6724 12492 6730
rect 12440 6666 12492 6672
rect 12348 6656 12400 6662
rect 12348 6598 12400 6604
rect 12360 6186 12388 6598
rect 12452 6390 12480 6666
rect 12440 6384 12492 6390
rect 12440 6326 12492 6332
rect 12348 6180 12400 6186
rect 12348 6122 12400 6128
rect 12452 5778 12480 6326
rect 12440 5772 12492 5778
rect 12440 5714 12492 5720
rect 12348 5636 12400 5642
rect 12348 5578 12400 5584
rect 12164 5228 12216 5234
rect 12164 5170 12216 5176
rect 12256 5228 12308 5234
rect 12256 5170 12308 5176
rect 12164 4820 12216 4826
rect 12164 4762 12216 4768
rect 12072 4684 12124 4690
rect 12072 4626 12124 4632
rect 11980 4616 12032 4622
rect 11980 4558 12032 4564
rect 11888 4548 11940 4554
rect 11888 4490 11940 4496
rect 11796 4276 11848 4282
rect 11796 4218 11848 4224
rect 11612 3732 11664 3738
rect 11612 3674 11664 3680
rect 11532 3590 11744 3618
rect 11612 3528 11664 3534
rect 11612 3470 11664 3476
rect 11518 2952 11574 2961
rect 11518 2887 11574 2896
rect 11532 2514 11560 2887
rect 11520 2508 11572 2514
rect 11520 2450 11572 2456
rect 11440 1414 11560 1442
rect 11428 1352 11480 1358
rect 11428 1294 11480 1300
rect 11440 800 11468 1294
rect 11532 800 11560 1414
rect 11624 800 11652 3470
rect 11716 800 11744 3590
rect 11808 1426 11836 4218
rect 11900 3534 11928 4490
rect 11980 4480 12032 4486
rect 11980 4422 12032 4428
rect 11888 3528 11940 3534
rect 11888 3470 11940 3476
rect 11886 2816 11942 2825
rect 11886 2751 11942 2760
rect 11796 1420 11848 1426
rect 11796 1362 11848 1368
rect 11900 800 11928 2751
rect 11992 2650 12020 4422
rect 12176 4162 12204 4762
rect 12268 4758 12296 5170
rect 12256 4752 12308 4758
rect 12256 4694 12308 4700
rect 12360 4622 12388 5578
rect 12544 5574 12572 6938
rect 12636 6225 12664 11494
rect 13188 10674 13216 11766
rect 13372 11354 13400 12786
rect 13360 11348 13412 11354
rect 13360 11290 13412 11296
rect 13176 10668 13228 10674
rect 13176 10610 13228 10616
rect 13268 10260 13320 10266
rect 13268 10202 13320 10208
rect 12716 9512 12768 9518
rect 12716 9454 12768 9460
rect 12728 7886 12756 9454
rect 13280 9178 13308 10202
rect 13268 9172 13320 9178
rect 13268 9114 13320 9120
rect 13360 8832 13412 8838
rect 13360 8774 13412 8780
rect 12716 7880 12768 7886
rect 12716 7822 12768 7828
rect 12728 7342 12756 7822
rect 13084 7540 13136 7546
rect 13084 7482 13136 7488
rect 12716 7336 12768 7342
rect 12716 7278 12768 7284
rect 12808 6656 12860 6662
rect 12808 6598 12860 6604
rect 12622 6216 12678 6225
rect 12622 6151 12678 6160
rect 12624 5908 12676 5914
rect 12624 5850 12676 5856
rect 12532 5568 12584 5574
rect 12532 5510 12584 5516
rect 12544 5166 12572 5510
rect 12532 5160 12584 5166
rect 12532 5102 12584 5108
rect 12544 4690 12572 5102
rect 12532 4684 12584 4690
rect 12452 4644 12532 4672
rect 12348 4616 12400 4622
rect 12348 4558 12400 4564
rect 12360 4282 12388 4558
rect 12348 4276 12400 4282
rect 12348 4218 12400 4224
rect 12452 4214 12480 4644
rect 12532 4626 12584 4632
rect 12532 4480 12584 4486
rect 12532 4422 12584 4428
rect 12544 4214 12572 4422
rect 12440 4208 12492 4214
rect 12176 4134 12388 4162
rect 12440 4150 12492 4156
rect 12532 4208 12584 4214
rect 12532 4150 12584 4156
rect 12162 3632 12218 3641
rect 12162 3567 12218 3576
rect 12072 2848 12124 2854
rect 12070 2816 12072 2825
rect 12124 2816 12126 2825
rect 12070 2751 12126 2760
rect 11980 2644 12032 2650
rect 11980 2586 12032 2592
rect 12072 2644 12124 2650
rect 12072 2586 12124 2592
rect 12084 2038 12112 2586
rect 12176 2378 12204 3567
rect 12256 3392 12308 3398
rect 12256 3334 12308 3340
rect 12268 3058 12296 3334
rect 12256 3052 12308 3058
rect 12256 2994 12308 3000
rect 12268 2650 12296 2994
rect 12256 2644 12308 2650
rect 12256 2586 12308 2592
rect 12164 2372 12216 2378
rect 12164 2314 12216 2320
rect 12072 2032 12124 2038
rect 12072 1974 12124 1980
rect 12176 1902 12204 2314
rect 12256 2304 12308 2310
rect 12256 2246 12308 2252
rect 12164 1896 12216 1902
rect 12164 1838 12216 1844
rect 11980 1760 12032 1766
rect 11980 1702 12032 1708
rect 11992 800 12020 1702
rect 12268 1562 12296 2246
rect 12256 1556 12308 1562
rect 12256 1498 12308 1504
rect 12072 1488 12124 1494
rect 12072 1430 12124 1436
rect 12084 800 12112 1430
rect 12256 1420 12308 1426
rect 12256 1362 12308 1368
rect 12268 800 12296 1362
rect 12360 800 12388 4134
rect 12440 4072 12492 4078
rect 12440 4014 12492 4020
rect 12452 3738 12480 4014
rect 12440 3732 12492 3738
rect 12440 3674 12492 3680
rect 12636 3466 12664 5850
rect 12716 5160 12768 5166
rect 12716 5102 12768 5108
rect 12624 3460 12676 3466
rect 12624 3402 12676 3408
rect 12440 3188 12492 3194
rect 12440 3130 12492 3136
rect 12452 800 12480 3130
rect 12728 2990 12756 5102
rect 12716 2984 12768 2990
rect 12716 2926 12768 2932
rect 12532 2848 12584 2854
rect 12532 2790 12584 2796
rect 12544 1970 12572 2790
rect 12716 2576 12768 2582
rect 12716 2518 12768 2524
rect 12624 2440 12676 2446
rect 12624 2382 12676 2388
rect 12636 2106 12664 2382
rect 12624 2100 12676 2106
rect 12624 2042 12676 2048
rect 12532 1964 12584 1970
rect 12532 1906 12584 1912
rect 12544 1426 12572 1906
rect 12532 1420 12584 1426
rect 12532 1362 12584 1368
rect 12636 800 12664 2042
rect 12728 1442 12756 2518
rect 12820 1698 12848 6598
rect 13096 5166 13124 7482
rect 13268 5364 13320 5370
rect 13268 5306 13320 5312
rect 13084 5160 13136 5166
rect 13084 5102 13136 5108
rect 13280 4486 13308 5306
rect 13268 4480 13320 4486
rect 13188 4440 13268 4468
rect 12900 4140 12952 4146
rect 12900 4082 12952 4088
rect 12808 1692 12860 1698
rect 12808 1634 12860 1640
rect 12728 1414 12848 1442
rect 12714 1320 12770 1329
rect 12714 1255 12770 1264
rect 12728 800 12756 1255
rect 12820 800 12848 1414
rect 12912 1329 12940 4082
rect 13084 3936 13136 3942
rect 13084 3878 13136 3884
rect 12992 3528 13044 3534
rect 12992 3470 13044 3476
rect 13004 2582 13032 3470
rect 12992 2576 13044 2582
rect 12992 2518 13044 2524
rect 12992 2032 13044 2038
rect 12992 1974 13044 1980
rect 12898 1320 12954 1329
rect 12898 1255 12954 1264
rect 12900 1216 12952 1222
rect 12900 1158 12952 1164
rect 12912 800 12940 1158
rect 13004 800 13032 1974
rect 13096 800 13124 3878
rect 13188 800 13216 4440
rect 13268 4422 13320 4428
rect 13372 3534 13400 8774
rect 13464 6202 13492 13330
rect 13556 11354 13584 15302
rect 13728 15020 13780 15026
rect 13728 14962 13780 14968
rect 13636 14272 13688 14278
rect 13636 14214 13688 14220
rect 13648 13870 13676 14214
rect 13636 13864 13688 13870
rect 13636 13806 13688 13812
rect 13740 13530 13768 14962
rect 14016 14618 14044 18022
rect 14108 17882 14136 18158
rect 14096 17876 14148 17882
rect 14096 17818 14148 17824
rect 14096 16584 14148 16590
rect 14096 16526 14148 16532
rect 14108 15076 14136 16526
rect 14200 15201 14228 18702
rect 14660 18306 14688 20878
rect 14844 18426 14872 21286
rect 15292 20936 15344 20942
rect 15292 20878 15344 20884
rect 15016 20800 15068 20806
rect 15016 20742 15068 20748
rect 14924 18760 14976 18766
rect 14924 18702 14976 18708
rect 14832 18420 14884 18426
rect 14832 18362 14884 18368
rect 14568 18278 14688 18306
rect 14280 15496 14332 15502
rect 14280 15438 14332 15444
rect 14186 15192 14242 15201
rect 14186 15127 14242 15136
rect 14188 15088 14240 15094
rect 14108 15048 14188 15076
rect 14188 15030 14240 15036
rect 14292 15026 14320 15438
rect 14372 15360 14424 15366
rect 14372 15302 14424 15308
rect 14280 15020 14332 15026
rect 14280 14962 14332 14968
rect 14004 14612 14056 14618
rect 14004 14554 14056 14560
rect 14384 13734 14412 15302
rect 13820 13728 13872 13734
rect 13820 13670 13872 13676
rect 14372 13728 14424 13734
rect 14372 13670 14424 13676
rect 13832 13530 13860 13670
rect 13728 13524 13780 13530
rect 13728 13466 13780 13472
rect 13820 13524 13872 13530
rect 13820 13466 13872 13472
rect 14384 13002 14412 13670
rect 14568 13530 14596 18278
rect 14648 18216 14700 18222
rect 14648 18158 14700 18164
rect 14660 16114 14688 18158
rect 14844 17882 14872 18362
rect 14936 18086 14964 18702
rect 14924 18080 14976 18086
rect 14924 18022 14976 18028
rect 14832 17876 14884 17882
rect 14832 17818 14884 17824
rect 14936 17610 14964 18022
rect 14924 17604 14976 17610
rect 14924 17546 14976 17552
rect 14924 16652 14976 16658
rect 14924 16594 14976 16600
rect 14648 16108 14700 16114
rect 14648 16050 14700 16056
rect 14832 16108 14884 16114
rect 14832 16050 14884 16056
rect 14844 15502 14872 16050
rect 14936 15706 14964 16594
rect 15028 16504 15056 20742
rect 15200 20528 15252 20534
rect 15200 20470 15252 20476
rect 15108 19780 15160 19786
rect 15108 19722 15160 19728
rect 15120 16574 15148 19722
rect 15212 19514 15240 20470
rect 15304 19786 15332 20878
rect 15488 20584 15516 24890
rect 15580 23662 15608 26318
rect 15844 26308 15896 26314
rect 15844 26250 15896 26256
rect 15660 25356 15712 25362
rect 15660 25298 15712 25304
rect 15672 24886 15700 25298
rect 15660 24880 15712 24886
rect 15660 24822 15712 24828
rect 15672 24342 15700 24822
rect 15856 24750 15884 26250
rect 15936 25696 15988 25702
rect 15936 25638 15988 25644
rect 15948 25294 15976 25638
rect 15936 25288 15988 25294
rect 15936 25230 15988 25236
rect 15948 24954 15976 25230
rect 15936 24948 15988 24954
rect 15936 24890 15988 24896
rect 16028 24812 16080 24818
rect 16028 24754 16080 24760
rect 15844 24744 15896 24750
rect 15844 24686 15896 24692
rect 15936 24744 15988 24750
rect 15936 24686 15988 24692
rect 15948 24410 15976 24686
rect 16040 24410 16068 24754
rect 16212 24676 16264 24682
rect 16212 24618 16264 24624
rect 15936 24404 15988 24410
rect 15936 24346 15988 24352
rect 16028 24404 16080 24410
rect 16028 24346 16080 24352
rect 15660 24336 15712 24342
rect 15660 24278 15712 24284
rect 16224 24206 16252 24618
rect 16212 24200 16264 24206
rect 16212 24142 16264 24148
rect 16224 23730 16252 24142
rect 16212 23724 16264 23730
rect 16212 23666 16264 23672
rect 15568 23656 15620 23662
rect 15568 23598 15620 23604
rect 15936 23520 15988 23526
rect 15936 23462 15988 23468
rect 15568 22636 15620 22642
rect 15568 22578 15620 22584
rect 15844 22636 15896 22642
rect 15844 22578 15896 22584
rect 15580 21554 15608 22578
rect 15856 22094 15884 22578
rect 15764 22066 15884 22094
rect 15764 21894 15792 22066
rect 15948 21978 15976 23462
rect 16224 23050 16252 23666
rect 16212 23044 16264 23050
rect 16212 22986 16264 22992
rect 15856 21950 15976 21978
rect 16212 22024 16264 22030
rect 16212 21966 16264 21972
rect 15752 21888 15804 21894
rect 15752 21830 15804 21836
rect 15764 21554 15792 21830
rect 15568 21548 15620 21554
rect 15568 21490 15620 21496
rect 15752 21548 15804 21554
rect 15752 21490 15804 21496
rect 15856 21350 15884 21950
rect 15936 21888 15988 21894
rect 15936 21830 15988 21836
rect 15844 21344 15896 21350
rect 15844 21286 15896 21292
rect 15948 20942 15976 21830
rect 16224 21690 16252 21966
rect 16212 21684 16264 21690
rect 16212 21626 16264 21632
rect 16028 21548 16080 21554
rect 16028 21490 16080 21496
rect 15936 20936 15988 20942
rect 15936 20878 15988 20884
rect 15488 20556 15884 20584
rect 15384 20528 15436 20534
rect 15384 20470 15436 20476
rect 15396 20262 15424 20470
rect 15476 20460 15528 20466
rect 15476 20402 15528 20408
rect 15752 20460 15804 20466
rect 15752 20402 15804 20408
rect 15384 20256 15436 20262
rect 15384 20198 15436 20204
rect 15292 19780 15344 19786
rect 15292 19722 15344 19728
rect 15396 19666 15424 20198
rect 15304 19638 15424 19666
rect 15200 19508 15252 19514
rect 15200 19450 15252 19456
rect 15304 19446 15332 19638
rect 15292 19440 15344 19446
rect 15292 19382 15344 19388
rect 15198 18456 15254 18465
rect 15198 18391 15254 18400
rect 15212 18358 15240 18391
rect 15200 18352 15252 18358
rect 15200 18294 15252 18300
rect 15120 16546 15240 16574
rect 15028 16476 15148 16504
rect 15016 16108 15068 16114
rect 15016 16050 15068 16056
rect 14924 15700 14976 15706
rect 14924 15642 14976 15648
rect 15028 15570 15056 16050
rect 15016 15564 15068 15570
rect 15016 15506 15068 15512
rect 14832 15496 14884 15502
rect 14832 15438 14884 15444
rect 14924 15496 14976 15502
rect 14924 15438 14976 15444
rect 14936 15366 14964 15438
rect 14924 15360 14976 15366
rect 14924 15302 14976 15308
rect 14648 15088 14700 15094
rect 14648 15030 14700 15036
rect 14660 14929 14688 15030
rect 15028 15026 15056 15506
rect 15016 15020 15068 15026
rect 15016 14962 15068 14968
rect 14646 14920 14702 14929
rect 14646 14855 14702 14864
rect 14648 14612 14700 14618
rect 14648 14554 14700 14560
rect 14660 14346 14688 14554
rect 14648 14340 14700 14346
rect 14648 14282 14700 14288
rect 14740 14340 14792 14346
rect 14740 14282 14792 14288
rect 14752 13977 14780 14282
rect 14738 13968 14794 13977
rect 14738 13903 14794 13912
rect 14556 13524 14608 13530
rect 14556 13466 14608 13472
rect 14646 13288 14702 13297
rect 14646 13223 14648 13232
rect 14700 13223 14702 13232
rect 14648 13194 14700 13200
rect 14384 12974 14596 13002
rect 14464 12640 14516 12646
rect 14464 12582 14516 12588
rect 14476 12238 14504 12582
rect 13820 12232 13872 12238
rect 13820 12174 13872 12180
rect 14464 12232 14516 12238
rect 14464 12174 14516 12180
rect 13636 12164 13688 12170
rect 13636 12106 13688 12112
rect 13544 11348 13596 11354
rect 13544 11290 13596 11296
rect 13544 11076 13596 11082
rect 13544 11018 13596 11024
rect 13556 6780 13584 11018
rect 13648 10198 13676 12106
rect 13832 11150 13860 12174
rect 14568 12170 14596 12974
rect 14924 12640 14976 12646
rect 14924 12582 14976 12588
rect 14936 12238 14964 12582
rect 15120 12238 15148 16476
rect 15212 15570 15240 16546
rect 15200 15564 15252 15570
rect 15200 15506 15252 15512
rect 14740 12232 14792 12238
rect 14924 12232 14976 12238
rect 14740 12174 14792 12180
rect 14922 12200 14924 12209
rect 15108 12232 15160 12238
rect 14976 12200 14978 12209
rect 14556 12164 14608 12170
rect 14556 12106 14608 12112
rect 14752 11286 14780 12174
rect 15108 12174 15160 12180
rect 14922 12135 14978 12144
rect 14832 12096 14884 12102
rect 14832 12038 14884 12044
rect 14844 11286 14872 12038
rect 15106 11928 15162 11937
rect 15106 11863 15162 11872
rect 15120 11354 15148 11863
rect 15212 11762 15240 15506
rect 15304 15026 15332 19382
rect 15384 18896 15436 18902
rect 15384 18838 15436 18844
rect 15396 18766 15424 18838
rect 15384 18760 15436 18766
rect 15384 18702 15436 18708
rect 15384 18624 15436 18630
rect 15384 18566 15436 18572
rect 15396 18290 15424 18566
rect 15384 18284 15436 18290
rect 15384 18226 15436 18232
rect 15488 18222 15516 20402
rect 15660 20392 15712 20398
rect 15764 20369 15792 20402
rect 15660 20334 15712 20340
rect 15750 20360 15806 20369
rect 15672 19854 15700 20334
rect 15750 20295 15806 20304
rect 15660 19848 15712 19854
rect 15660 19790 15712 19796
rect 15568 19780 15620 19786
rect 15568 19722 15620 19728
rect 15752 19780 15804 19786
rect 15752 19722 15804 19728
rect 15476 18216 15528 18222
rect 15476 18158 15528 18164
rect 15384 18080 15436 18086
rect 15384 18022 15436 18028
rect 15396 17678 15424 18022
rect 15384 17672 15436 17678
rect 15476 17672 15528 17678
rect 15384 17614 15436 17620
rect 15474 17640 15476 17649
rect 15580 17660 15608 19722
rect 15660 19372 15712 19378
rect 15660 19314 15712 19320
rect 15672 18970 15700 19314
rect 15660 18964 15712 18970
rect 15660 18906 15712 18912
rect 15672 18766 15700 18906
rect 15764 18902 15792 19722
rect 15856 19174 15884 20556
rect 15844 19168 15896 19174
rect 15844 19110 15896 19116
rect 15752 18896 15804 18902
rect 15752 18838 15804 18844
rect 15660 18760 15712 18766
rect 15660 18702 15712 18708
rect 15660 18284 15712 18290
rect 15660 18226 15712 18232
rect 15672 17814 15700 18226
rect 15764 17864 15792 18838
rect 15936 18624 15988 18630
rect 15936 18566 15988 18572
rect 15764 17836 15884 17864
rect 15660 17808 15712 17814
rect 15660 17750 15712 17756
rect 15528 17640 15608 17660
rect 15530 17632 15608 17640
rect 15474 17575 15530 17584
rect 15660 17196 15712 17202
rect 15660 17138 15712 17144
rect 15672 16794 15700 17138
rect 15660 16788 15712 16794
rect 15660 16730 15712 16736
rect 15568 15904 15620 15910
rect 15568 15846 15620 15852
rect 15292 15020 15344 15026
rect 15292 14962 15344 14968
rect 15292 14816 15344 14822
rect 15292 14758 15344 14764
rect 15200 11756 15252 11762
rect 15200 11698 15252 11704
rect 15108 11348 15160 11354
rect 15108 11290 15160 11296
rect 14740 11280 14792 11286
rect 14740 11222 14792 11228
rect 14832 11280 14884 11286
rect 14832 11222 14884 11228
rect 13820 11144 13872 11150
rect 13820 11086 13872 11092
rect 14648 11076 14700 11082
rect 14648 11018 14700 11024
rect 13636 10192 13688 10198
rect 13636 10134 13688 10140
rect 13648 8362 13676 10134
rect 14096 10056 14148 10062
rect 14096 9998 14148 10004
rect 14188 10056 14240 10062
rect 14188 9998 14240 10004
rect 13636 8356 13688 8362
rect 13636 8298 13688 8304
rect 13820 7744 13872 7750
rect 13820 7686 13872 7692
rect 13728 7200 13780 7206
rect 13728 7142 13780 7148
rect 13556 6752 13676 6780
rect 13464 6174 13584 6202
rect 13450 6080 13506 6089
rect 13450 6015 13506 6024
rect 13464 5234 13492 6015
rect 13452 5228 13504 5234
rect 13452 5170 13504 5176
rect 13556 4298 13584 6174
rect 13464 4270 13584 4298
rect 13464 3670 13492 4270
rect 13544 4140 13596 4146
rect 13544 4082 13596 4088
rect 13452 3664 13504 3670
rect 13452 3606 13504 3612
rect 13360 3528 13412 3534
rect 13360 3470 13412 3476
rect 13452 3460 13504 3466
rect 13452 3402 13504 3408
rect 13268 3120 13320 3126
rect 13268 3062 13320 3068
rect 13280 800 13308 3062
rect 13360 1556 13412 1562
rect 13360 1498 13412 1504
rect 13372 800 13400 1498
rect 13464 800 13492 3402
rect 13556 3058 13584 4082
rect 13648 3942 13676 6752
rect 13740 4622 13768 7142
rect 13728 4616 13780 4622
rect 13728 4558 13780 4564
rect 13740 4146 13768 4558
rect 13832 4146 13860 7686
rect 14004 6792 14056 6798
rect 14004 6734 14056 6740
rect 14016 6118 14044 6734
rect 14108 6254 14136 9998
rect 14200 9178 14228 9998
rect 14556 9988 14608 9994
rect 14556 9930 14608 9936
rect 14568 9722 14596 9930
rect 14556 9716 14608 9722
rect 14556 9658 14608 9664
rect 14188 9172 14240 9178
rect 14188 9114 14240 9120
rect 14096 6248 14148 6254
rect 14096 6190 14148 6196
rect 13912 6112 13964 6118
rect 13912 6054 13964 6060
rect 14004 6112 14056 6118
rect 14004 6054 14056 6060
rect 13728 4140 13780 4146
rect 13728 4082 13780 4088
rect 13820 4140 13872 4146
rect 13820 4082 13872 4088
rect 13636 3936 13688 3942
rect 13636 3878 13688 3884
rect 13636 3392 13688 3398
rect 13636 3334 13688 3340
rect 13544 3052 13596 3058
rect 13544 2994 13596 3000
rect 13544 1828 13596 1834
rect 13544 1770 13596 1776
rect 13556 800 13584 1770
rect 13648 800 13676 3334
rect 13832 800 13860 4082
rect 13924 3126 13952 6054
rect 14200 5710 14228 9114
rect 14372 8628 14424 8634
rect 14372 8570 14424 8576
rect 14384 8430 14412 8570
rect 14464 8492 14516 8498
rect 14464 8434 14516 8440
rect 14372 8424 14424 8430
rect 14372 8366 14424 8372
rect 14280 7744 14332 7750
rect 14280 7686 14332 7692
rect 14292 7478 14320 7686
rect 14280 7472 14332 7478
rect 14280 7414 14332 7420
rect 14476 7206 14504 8434
rect 14660 8022 14688 11018
rect 14752 9586 14780 11222
rect 15212 10470 15240 11698
rect 15304 11694 15332 14758
rect 15476 13932 15528 13938
rect 15476 13874 15528 13880
rect 15488 13530 15516 13874
rect 15476 13524 15528 13530
rect 15476 13466 15528 13472
rect 15476 12232 15528 12238
rect 15476 12174 15528 12180
rect 15488 11801 15516 12174
rect 15474 11792 15530 11801
rect 15474 11727 15530 11736
rect 15292 11688 15344 11694
rect 15292 11630 15344 11636
rect 15580 11354 15608 15846
rect 15752 15496 15804 15502
rect 15752 15438 15804 15444
rect 15764 15026 15792 15438
rect 15856 15416 15884 17836
rect 15948 16522 15976 18566
rect 15936 16516 15988 16522
rect 15936 16458 15988 16464
rect 15936 15428 15988 15434
rect 15856 15388 15936 15416
rect 15752 15020 15804 15026
rect 15752 14962 15804 14968
rect 15764 14890 15792 14962
rect 15752 14884 15804 14890
rect 15752 14826 15804 14832
rect 15856 14618 15884 15388
rect 15936 15370 15988 15376
rect 15936 14816 15988 14822
rect 15936 14758 15988 14764
rect 15844 14612 15896 14618
rect 15844 14554 15896 14560
rect 15856 14414 15884 14554
rect 15844 14408 15896 14414
rect 15844 14350 15896 14356
rect 15856 14006 15884 14350
rect 15844 14000 15896 14006
rect 15844 13942 15896 13948
rect 15844 13524 15896 13530
rect 15844 13466 15896 13472
rect 15660 13388 15712 13394
rect 15712 13348 15792 13376
rect 15660 13330 15712 13336
rect 15764 12238 15792 13348
rect 15856 13326 15884 13466
rect 15844 13320 15896 13326
rect 15844 13262 15896 13268
rect 15844 13184 15896 13190
rect 15844 13126 15896 13132
rect 15660 12232 15712 12238
rect 15660 12174 15712 12180
rect 15752 12232 15804 12238
rect 15752 12174 15804 12180
rect 15568 11348 15620 11354
rect 15568 11290 15620 11296
rect 15476 11144 15528 11150
rect 15476 11086 15528 11092
rect 15200 10464 15252 10470
rect 15200 10406 15252 10412
rect 15212 9926 15240 10406
rect 15488 10062 15516 11086
rect 15476 10056 15528 10062
rect 15476 9998 15528 10004
rect 14832 9920 14884 9926
rect 14832 9862 14884 9868
rect 15200 9920 15252 9926
rect 15200 9862 15252 9868
rect 14740 9580 14792 9586
rect 14740 9522 14792 9528
rect 14844 9518 14872 9862
rect 15212 9654 15240 9862
rect 15200 9648 15252 9654
rect 15672 9602 15700 12174
rect 15752 12096 15804 12102
rect 15752 12038 15804 12044
rect 15764 11762 15792 12038
rect 15752 11756 15804 11762
rect 15752 11698 15804 11704
rect 15200 9590 15252 9596
rect 15476 9580 15528 9586
rect 15476 9522 15528 9528
rect 15580 9574 15700 9602
rect 14832 9512 14884 9518
rect 14832 9454 14884 9460
rect 15384 9444 15436 9450
rect 15384 9386 15436 9392
rect 15016 8560 15068 8566
rect 15016 8502 15068 8508
rect 14740 8288 14792 8294
rect 14740 8230 14792 8236
rect 14832 8288 14884 8294
rect 14832 8230 14884 8236
rect 14648 8016 14700 8022
rect 14648 7958 14700 7964
rect 14752 7886 14780 8230
rect 14740 7880 14792 7886
rect 14740 7822 14792 7828
rect 14464 7200 14516 7206
rect 14464 7142 14516 7148
rect 14740 7200 14792 7206
rect 14740 7142 14792 7148
rect 14280 6792 14332 6798
rect 14280 6734 14332 6740
rect 14292 6186 14320 6734
rect 14372 6316 14424 6322
rect 14372 6258 14424 6264
rect 14280 6180 14332 6186
rect 14280 6122 14332 6128
rect 14188 5704 14240 5710
rect 14188 5646 14240 5652
rect 14280 5704 14332 5710
rect 14280 5646 14332 5652
rect 14292 5302 14320 5646
rect 14384 5370 14412 6258
rect 14372 5364 14424 5370
rect 14372 5306 14424 5312
rect 14280 5296 14332 5302
rect 14280 5238 14332 5244
rect 14372 5228 14424 5234
rect 14372 5170 14424 5176
rect 14096 5160 14148 5166
rect 14096 5102 14148 5108
rect 14108 4826 14136 5102
rect 14280 5024 14332 5030
rect 14280 4966 14332 4972
rect 14096 4820 14148 4826
rect 14096 4762 14148 4768
rect 14096 3936 14148 3942
rect 14096 3878 14148 3884
rect 14108 3777 14136 3878
rect 14094 3768 14150 3777
rect 14094 3703 14150 3712
rect 14188 3392 14240 3398
rect 14188 3334 14240 3340
rect 13912 3120 13964 3126
rect 13912 3062 13964 3068
rect 14094 2952 14150 2961
rect 14094 2887 14150 2896
rect 13912 2848 13964 2854
rect 13912 2790 13964 2796
rect 13924 800 13952 2790
rect 14108 800 14136 2887
rect 14200 800 14228 3334
rect 14292 1630 14320 4966
rect 14384 3058 14412 5170
rect 14372 3052 14424 3058
rect 14372 2994 14424 3000
rect 14372 2576 14424 2582
rect 14372 2518 14424 2524
rect 14280 1624 14332 1630
rect 14280 1566 14332 1572
rect 14384 800 14412 2518
rect 14476 2514 14504 7142
rect 14648 6112 14700 6118
rect 14648 6054 14700 6060
rect 14464 2508 14516 2514
rect 14464 2450 14516 2456
rect 14556 2440 14608 2446
rect 14556 2382 14608 2388
rect 14464 2304 14516 2310
rect 14464 2246 14516 2252
rect 14476 800 14504 2246
rect 14568 2106 14596 2382
rect 14556 2100 14608 2106
rect 14556 2042 14608 2048
rect 14660 800 14688 6054
rect 14752 5642 14780 7142
rect 14740 5636 14792 5642
rect 14740 5578 14792 5584
rect 14752 5370 14780 5578
rect 14740 5364 14792 5370
rect 14740 5306 14792 5312
rect 14844 2774 14872 8230
rect 15028 7750 15056 8502
rect 15108 8492 15160 8498
rect 15108 8434 15160 8440
rect 14924 7744 14976 7750
rect 14924 7686 14976 7692
rect 15016 7744 15068 7750
rect 15016 7686 15068 7692
rect 14936 6730 14964 7686
rect 15028 7342 15056 7686
rect 15016 7336 15068 7342
rect 15016 7278 15068 7284
rect 15016 6860 15068 6866
rect 15016 6802 15068 6808
rect 14924 6724 14976 6730
rect 14924 6666 14976 6672
rect 14936 6458 14964 6666
rect 14924 6452 14976 6458
rect 14924 6394 14976 6400
rect 14936 6322 14964 6394
rect 14924 6316 14976 6322
rect 14924 6258 14976 6264
rect 14922 5536 14978 5545
rect 14922 5471 14978 5480
rect 14936 4146 14964 5471
rect 14924 4140 14976 4146
rect 14924 4082 14976 4088
rect 14924 3188 14976 3194
rect 14924 3130 14976 3136
rect 14936 3058 14964 3130
rect 14924 3052 14976 3058
rect 14924 2994 14976 3000
rect 14752 2746 14872 2774
rect 14752 2582 14780 2746
rect 14740 2576 14792 2582
rect 14740 2518 14792 2524
rect 14752 2428 14780 2518
rect 14924 2440 14976 2446
rect 14752 2400 14924 2428
rect 14924 2382 14976 2388
rect 14740 2304 14792 2310
rect 14740 2246 14792 2252
rect 14752 800 14780 2246
rect 15028 800 15056 6802
rect 15120 5778 15148 8434
rect 15292 8356 15344 8362
rect 15292 8298 15344 8304
rect 15200 6112 15252 6118
rect 15200 6054 15252 6060
rect 15108 5772 15160 5778
rect 15108 5714 15160 5720
rect 15120 5234 15148 5714
rect 15108 5228 15160 5234
rect 15108 5170 15160 5176
rect 15212 4554 15240 6054
rect 15200 4548 15252 4554
rect 15200 4490 15252 4496
rect 15108 3664 15160 3670
rect 15106 3632 15108 3641
rect 15160 3632 15162 3641
rect 15106 3567 15162 3576
rect 15200 3052 15252 3058
rect 15200 2994 15252 3000
rect 15212 2961 15240 2994
rect 15198 2952 15254 2961
rect 15198 2887 15254 2896
rect 15200 2372 15252 2378
rect 15200 2314 15252 2320
rect 15212 1970 15240 2314
rect 15200 1964 15252 1970
rect 15200 1906 15252 1912
rect 15304 800 15332 8298
rect 15396 6322 15424 9386
rect 15488 8838 15516 9522
rect 15476 8832 15528 8838
rect 15476 8774 15528 8780
rect 15580 8090 15608 9574
rect 15660 9376 15712 9382
rect 15660 9318 15712 9324
rect 15672 8974 15700 9318
rect 15660 8968 15712 8974
rect 15660 8910 15712 8916
rect 15568 8084 15620 8090
rect 15568 8026 15620 8032
rect 15752 7948 15804 7954
rect 15752 7890 15804 7896
rect 15568 7880 15620 7886
rect 15568 7822 15620 7828
rect 15384 6316 15436 6322
rect 15384 6258 15436 6264
rect 15476 6316 15528 6322
rect 15476 6258 15528 6264
rect 15382 5808 15438 5817
rect 15382 5743 15438 5752
rect 15396 4010 15424 5743
rect 15488 5370 15516 6258
rect 15476 5364 15528 5370
rect 15476 5306 15528 5312
rect 15384 4004 15436 4010
rect 15384 3946 15436 3952
rect 15384 3528 15436 3534
rect 15384 3470 15436 3476
rect 15396 1834 15424 3470
rect 15384 1828 15436 1834
rect 15384 1770 15436 1776
rect 15580 800 15608 7822
rect 15660 6792 15712 6798
rect 15660 6734 15712 6740
rect 15672 6322 15700 6734
rect 15660 6316 15712 6322
rect 15660 6258 15712 6264
rect 15764 3466 15792 7890
rect 15856 7857 15884 13126
rect 15948 12646 15976 14758
rect 16040 14550 16068 21490
rect 16316 20398 16344 26794
rect 16592 26382 16620 27406
rect 16580 26376 16632 26382
rect 16580 26318 16632 26324
rect 16592 25906 16620 26318
rect 16580 25900 16632 25906
rect 16580 25842 16632 25848
rect 16672 25900 16724 25906
rect 16672 25842 16724 25848
rect 16684 24614 16712 25842
rect 16672 24608 16724 24614
rect 16672 24550 16724 24556
rect 16488 24336 16540 24342
rect 16488 24278 16540 24284
rect 16500 23798 16528 24278
rect 16580 24064 16632 24070
rect 16580 24006 16632 24012
rect 16684 24018 16712 24550
rect 16776 24449 16804 28426
rect 17224 27940 17276 27946
rect 17224 27882 17276 27888
rect 17236 27334 17264 27882
rect 17408 27872 17460 27878
rect 17408 27814 17460 27820
rect 17420 27470 17448 27814
rect 17408 27464 17460 27470
rect 17408 27406 17460 27412
rect 17224 27328 17276 27334
rect 17224 27270 17276 27276
rect 17132 26920 17184 26926
rect 17132 26862 17184 26868
rect 17144 26518 17172 26862
rect 17132 26512 17184 26518
rect 17132 26454 17184 26460
rect 17040 26308 17092 26314
rect 17040 26250 17092 26256
rect 16856 25696 16908 25702
rect 16856 25638 16908 25644
rect 16868 24886 16896 25638
rect 16856 24880 16908 24886
rect 16856 24822 16908 24828
rect 16762 24440 16818 24449
rect 16762 24375 16818 24384
rect 16764 24200 16816 24206
rect 16868 24188 16896 24822
rect 17052 24818 17080 26250
rect 17132 25288 17184 25294
rect 17132 25230 17184 25236
rect 17040 24812 17092 24818
rect 17040 24754 17092 24760
rect 17040 24676 17092 24682
rect 17040 24618 17092 24624
rect 16816 24160 16896 24188
rect 16764 24142 16816 24148
rect 16488 23792 16540 23798
rect 16488 23734 16540 23740
rect 16592 23730 16620 24006
rect 16684 23990 16804 24018
rect 16580 23724 16632 23730
rect 16580 23666 16632 23672
rect 16592 23594 16620 23666
rect 16580 23588 16632 23594
rect 16580 23530 16632 23536
rect 16672 23588 16724 23594
rect 16672 23530 16724 23536
rect 16592 22030 16620 23530
rect 16396 22024 16448 22030
rect 16396 21966 16448 21972
rect 16580 22024 16632 22030
rect 16580 21966 16632 21972
rect 16408 21690 16436 21966
rect 16396 21684 16448 21690
rect 16396 21626 16448 21632
rect 16580 21480 16632 21486
rect 16580 21422 16632 21428
rect 16592 21350 16620 21422
rect 16580 21344 16632 21350
rect 16580 21286 16632 21292
rect 16684 20534 16712 23530
rect 16776 21554 16804 23990
rect 16856 23724 16908 23730
rect 16856 23666 16908 23672
rect 16868 23322 16896 23666
rect 16948 23588 17000 23594
rect 16948 23530 17000 23536
rect 16856 23316 16908 23322
rect 16856 23258 16908 23264
rect 16960 22094 16988 23530
rect 16868 22066 16988 22094
rect 16868 21570 16896 22066
rect 16764 21548 16816 21554
rect 16868 21542 16988 21570
rect 16764 21490 16816 21496
rect 16672 20528 16724 20534
rect 16672 20470 16724 20476
rect 16304 20392 16356 20398
rect 16304 20334 16356 20340
rect 16316 19786 16344 20334
rect 16672 19916 16724 19922
rect 16672 19858 16724 19864
rect 16304 19780 16356 19786
rect 16304 19722 16356 19728
rect 16488 19712 16540 19718
rect 16488 19654 16540 19660
rect 16120 18692 16172 18698
rect 16120 18634 16172 18640
rect 16132 18329 16160 18634
rect 16210 18456 16266 18465
rect 16210 18391 16266 18400
rect 16224 18358 16252 18391
rect 16212 18352 16264 18358
rect 16118 18320 16174 18329
rect 16212 18294 16264 18300
rect 16118 18255 16120 18264
rect 16172 18255 16174 18264
rect 16120 18226 16172 18232
rect 16132 17338 16160 18226
rect 16212 18216 16264 18222
rect 16212 18158 16264 18164
rect 16224 17746 16252 18158
rect 16212 17740 16264 17746
rect 16212 17682 16264 17688
rect 16224 17338 16252 17682
rect 16304 17672 16356 17678
rect 16304 17614 16356 17620
rect 16394 17640 16450 17649
rect 16120 17332 16172 17338
rect 16120 17274 16172 17280
rect 16212 17332 16264 17338
rect 16212 17274 16264 17280
rect 16212 17196 16264 17202
rect 16212 17138 16264 17144
rect 16224 16726 16252 17138
rect 16212 16720 16264 16726
rect 16212 16662 16264 16668
rect 16316 16658 16344 17614
rect 16394 17575 16450 17584
rect 16408 17270 16436 17575
rect 16396 17264 16448 17270
rect 16396 17206 16448 17212
rect 16304 16652 16356 16658
rect 16304 16594 16356 16600
rect 16304 14884 16356 14890
rect 16304 14826 16356 14832
rect 16028 14544 16080 14550
rect 16028 14486 16080 14492
rect 16316 14482 16344 14826
rect 16304 14476 16356 14482
rect 16304 14418 16356 14424
rect 16396 13864 16448 13870
rect 16396 13806 16448 13812
rect 16026 13424 16082 13433
rect 16026 13359 16082 13368
rect 16040 13326 16068 13359
rect 16028 13320 16080 13326
rect 16028 13262 16080 13268
rect 16304 13184 16356 13190
rect 16304 13126 16356 13132
rect 16120 12844 16172 12850
rect 16120 12786 16172 12792
rect 16212 12844 16264 12850
rect 16212 12786 16264 12792
rect 15936 12640 15988 12646
rect 15936 12582 15988 12588
rect 16132 12345 16160 12786
rect 16118 12336 16174 12345
rect 16118 12271 16174 12280
rect 16224 11830 16252 12786
rect 16212 11824 16264 11830
rect 16212 11766 16264 11772
rect 15936 11552 15988 11558
rect 15936 11494 15988 11500
rect 15842 7848 15898 7857
rect 15842 7783 15898 7792
rect 15844 7200 15896 7206
rect 15844 7142 15896 7148
rect 15856 3534 15884 7142
rect 15948 5001 15976 11494
rect 16028 9920 16080 9926
rect 16028 9862 16080 9868
rect 16040 6390 16068 9862
rect 16224 9042 16252 11766
rect 16316 11762 16344 13126
rect 16304 11756 16356 11762
rect 16304 11698 16356 11704
rect 16304 11076 16356 11082
rect 16304 11018 16356 11024
rect 16212 9036 16264 9042
rect 16212 8978 16264 8984
rect 16316 7886 16344 11018
rect 16304 7880 16356 7886
rect 16304 7822 16356 7828
rect 16120 7812 16172 7818
rect 16120 7754 16172 7760
rect 16132 6798 16160 7754
rect 16408 7732 16436 13806
rect 16500 13530 16528 19654
rect 16684 19378 16712 19858
rect 16776 19514 16804 21490
rect 16854 21176 16910 21185
rect 16854 21111 16856 21120
rect 16908 21111 16910 21120
rect 16856 21082 16908 21088
rect 16960 19530 16988 21542
rect 17052 19854 17080 24618
rect 17144 24188 17172 25230
rect 17236 24834 17264 27270
rect 17420 26586 17448 27406
rect 17500 27328 17552 27334
rect 17500 27270 17552 27276
rect 17684 27328 17736 27334
rect 17684 27270 17736 27276
rect 17512 27062 17540 27270
rect 17500 27056 17552 27062
rect 17500 26998 17552 27004
rect 17696 26994 17724 27270
rect 17684 26988 17736 26994
rect 17684 26930 17736 26936
rect 17408 26580 17460 26586
rect 17408 26522 17460 26528
rect 17696 26382 17724 26930
rect 17684 26376 17736 26382
rect 17684 26318 17736 26324
rect 17696 25906 17724 26318
rect 17684 25900 17736 25906
rect 17684 25842 17736 25848
rect 17316 25288 17368 25294
rect 17316 25230 17368 25236
rect 17328 24954 17356 25230
rect 17316 24948 17368 24954
rect 17316 24890 17368 24896
rect 17696 24886 17724 25842
rect 17684 24880 17736 24886
rect 17236 24806 17356 24834
rect 17684 24822 17736 24828
rect 17224 24200 17276 24206
rect 17144 24160 17224 24188
rect 17224 24142 17276 24148
rect 17236 24070 17264 24142
rect 17224 24064 17276 24070
rect 17224 24006 17276 24012
rect 17132 22636 17184 22642
rect 17132 22578 17184 22584
rect 17224 22636 17276 22642
rect 17224 22578 17276 22584
rect 17144 21146 17172 22578
rect 17236 21622 17264 22578
rect 17224 21616 17276 21622
rect 17224 21558 17276 21564
rect 17224 21480 17276 21486
rect 17224 21422 17276 21428
rect 17236 21185 17264 21422
rect 17328 21350 17356 24806
rect 17684 24744 17736 24750
rect 17684 24686 17736 24692
rect 17408 24404 17460 24410
rect 17408 24346 17460 24352
rect 17316 21344 17368 21350
rect 17316 21286 17368 21292
rect 17222 21176 17278 21185
rect 17132 21140 17184 21146
rect 17222 21111 17278 21120
rect 17132 21082 17184 21088
rect 17132 20800 17184 20806
rect 17132 20742 17184 20748
rect 17144 20466 17172 20742
rect 17132 20460 17184 20466
rect 17132 20402 17184 20408
rect 17224 20460 17276 20466
rect 17224 20402 17276 20408
rect 17040 19848 17092 19854
rect 17040 19790 17092 19796
rect 16764 19508 16816 19514
rect 16764 19450 16816 19456
rect 16868 19502 16988 19530
rect 16672 19372 16724 19378
rect 16672 19314 16724 19320
rect 16764 19304 16816 19310
rect 16764 19246 16816 19252
rect 16672 19168 16724 19174
rect 16672 19110 16724 19116
rect 16684 17814 16712 19110
rect 16776 18630 16804 19246
rect 16764 18624 16816 18630
rect 16764 18566 16816 18572
rect 16672 17808 16724 17814
rect 16672 17750 16724 17756
rect 16580 17536 16632 17542
rect 16580 17478 16632 17484
rect 16592 15094 16620 17478
rect 16670 17096 16726 17105
rect 16670 17031 16726 17040
rect 16580 15088 16632 15094
rect 16580 15030 16632 15036
rect 16580 14544 16632 14550
rect 16580 14486 16632 14492
rect 16592 14414 16620 14486
rect 16580 14408 16632 14414
rect 16580 14350 16632 14356
rect 16578 13696 16634 13705
rect 16578 13631 16634 13640
rect 16488 13524 16540 13530
rect 16488 13466 16540 13472
rect 16486 13424 16542 13433
rect 16592 13394 16620 13631
rect 16486 13359 16488 13368
rect 16540 13359 16542 13368
rect 16580 13388 16632 13394
rect 16488 13330 16540 13336
rect 16580 13330 16632 13336
rect 16684 12442 16712 17031
rect 16776 13258 16804 18566
rect 16868 16726 16896 19502
rect 16948 19440 17000 19446
rect 16948 19382 17000 19388
rect 16960 17678 16988 19382
rect 17144 19310 17172 20402
rect 17132 19304 17184 19310
rect 17132 19246 17184 19252
rect 17132 19168 17184 19174
rect 17132 19110 17184 19116
rect 17040 18624 17092 18630
rect 17040 18566 17092 18572
rect 16948 17672 17000 17678
rect 16948 17614 17000 17620
rect 17052 17490 17080 18566
rect 17144 18426 17172 19110
rect 17236 18630 17264 20402
rect 17328 18766 17356 21286
rect 17316 18760 17368 18766
rect 17316 18702 17368 18708
rect 17224 18624 17276 18630
rect 17420 18612 17448 24346
rect 17696 24342 17724 24686
rect 17684 24336 17736 24342
rect 17684 24278 17736 24284
rect 17684 24200 17736 24206
rect 17684 24142 17736 24148
rect 17696 24070 17724 24142
rect 17684 24064 17736 24070
rect 17684 24006 17736 24012
rect 17696 23594 17724 24006
rect 17684 23588 17736 23594
rect 17684 23530 17736 23536
rect 17592 23520 17644 23526
rect 17592 23462 17644 23468
rect 17604 23050 17632 23462
rect 17592 23044 17644 23050
rect 17592 22986 17644 22992
rect 17788 22778 17816 28426
rect 18064 28150 18092 28494
rect 18052 28144 18104 28150
rect 18052 28086 18104 28092
rect 18236 28076 18288 28082
rect 18236 28018 18288 28024
rect 18248 27962 18276 28018
rect 18248 27946 18368 27962
rect 18248 27940 18380 27946
rect 18248 27934 18328 27940
rect 18328 27882 18380 27888
rect 17960 27872 18012 27878
rect 17960 27814 18012 27820
rect 17972 27470 18000 27814
rect 17960 27464 18012 27470
rect 17960 27406 18012 27412
rect 18236 27124 18288 27130
rect 18236 27066 18288 27072
rect 17960 25900 18012 25906
rect 17960 25842 18012 25848
rect 17972 25498 18000 25842
rect 17960 25492 18012 25498
rect 17960 25434 18012 25440
rect 17868 24200 17920 24206
rect 17868 24142 17920 24148
rect 17880 23526 17908 24142
rect 17868 23520 17920 23526
rect 17868 23462 17920 23468
rect 17776 22772 17828 22778
rect 17776 22714 17828 22720
rect 17880 22642 17908 23462
rect 17960 22976 18012 22982
rect 17960 22918 18012 22924
rect 17500 22636 17552 22642
rect 17500 22578 17552 22584
rect 17868 22636 17920 22642
rect 17868 22578 17920 22584
rect 17512 20466 17540 22578
rect 17972 22098 18000 22918
rect 17960 22092 18012 22098
rect 18248 22094 18276 27066
rect 18340 26790 18368 27882
rect 18328 26784 18380 26790
rect 18328 26726 18380 26732
rect 18328 24812 18380 24818
rect 18328 24754 18380 24760
rect 18420 24812 18472 24818
rect 18420 24754 18472 24760
rect 18340 23186 18368 24754
rect 18432 24410 18460 24754
rect 18420 24404 18472 24410
rect 18420 24346 18472 24352
rect 18328 23180 18380 23186
rect 18328 23122 18380 23128
rect 18248 22066 18368 22094
rect 17960 22034 18012 22040
rect 17592 22024 17644 22030
rect 18142 21992 18198 22001
rect 17644 21972 17724 21978
rect 17592 21966 17724 21972
rect 17604 21950 17724 21966
rect 17592 21888 17644 21894
rect 17592 21830 17644 21836
rect 17604 21418 17632 21830
rect 17696 21690 17724 21950
rect 18142 21927 18198 21936
rect 17684 21684 17736 21690
rect 17684 21626 17736 21632
rect 17868 21548 17920 21554
rect 17868 21490 17920 21496
rect 17592 21412 17644 21418
rect 17592 21354 17644 21360
rect 17500 20460 17552 20466
rect 17500 20402 17552 20408
rect 17500 19712 17552 19718
rect 17500 19654 17552 19660
rect 17684 19712 17736 19718
rect 17684 19654 17736 19660
rect 17224 18566 17276 18572
rect 17328 18584 17448 18612
rect 17328 18442 17356 18584
rect 17132 18420 17184 18426
rect 17132 18362 17184 18368
rect 17236 18414 17356 18442
rect 17236 17542 17264 18414
rect 17420 18290 17448 18584
rect 17408 18284 17460 18290
rect 17408 18226 17460 18232
rect 16960 17462 17080 17490
rect 17224 17536 17276 17542
rect 17224 17478 17276 17484
rect 16856 16720 16908 16726
rect 16856 16662 16908 16668
rect 16856 15496 16908 15502
rect 16854 15464 16856 15473
rect 16908 15464 16910 15473
rect 16854 15399 16910 15408
rect 16960 15162 16988 17462
rect 17236 17105 17264 17478
rect 17222 17096 17278 17105
rect 17222 17031 17278 17040
rect 17132 16448 17184 16454
rect 17132 16390 17184 16396
rect 17040 15904 17092 15910
rect 17040 15846 17092 15852
rect 17052 15502 17080 15846
rect 17040 15496 17092 15502
rect 17040 15438 17092 15444
rect 16948 15156 17000 15162
rect 16948 15098 17000 15104
rect 17038 14104 17094 14113
rect 17038 14039 17094 14048
rect 17052 13938 17080 14039
rect 17040 13932 17092 13938
rect 17040 13874 17092 13880
rect 17144 13818 17172 16390
rect 17222 15600 17278 15609
rect 17222 15535 17278 15544
rect 17236 15502 17264 15535
rect 17224 15496 17276 15502
rect 17224 15438 17276 15444
rect 17316 15496 17368 15502
rect 17316 15438 17368 15444
rect 17224 15156 17276 15162
rect 17224 15098 17276 15104
rect 17236 13938 17264 15098
rect 17328 14414 17356 15438
rect 17512 15076 17540 19654
rect 17592 18692 17644 18698
rect 17592 18634 17644 18640
rect 17604 18426 17632 18634
rect 17592 18420 17644 18426
rect 17592 18362 17644 18368
rect 17696 16153 17724 19654
rect 17776 17672 17828 17678
rect 17776 17614 17828 17620
rect 17788 16182 17816 17614
rect 17776 16176 17828 16182
rect 17682 16144 17738 16153
rect 17776 16118 17828 16124
rect 17682 16079 17738 16088
rect 17684 15088 17736 15094
rect 17512 15048 17684 15076
rect 17684 15030 17736 15036
rect 17408 14952 17460 14958
rect 17408 14894 17460 14900
rect 17420 14521 17448 14894
rect 17696 14890 17724 15030
rect 17788 15026 17816 16118
rect 17880 15638 17908 21490
rect 18156 20942 18184 21927
rect 17960 20936 18012 20942
rect 17960 20878 18012 20884
rect 18144 20936 18196 20942
rect 18144 20878 18196 20884
rect 18236 20936 18288 20942
rect 18236 20878 18288 20884
rect 17972 20602 18000 20878
rect 17960 20596 18012 20602
rect 17960 20538 18012 20544
rect 17972 19378 18000 20538
rect 18052 20256 18104 20262
rect 18052 20198 18104 20204
rect 18064 20058 18092 20198
rect 18052 20052 18104 20058
rect 18052 19994 18104 20000
rect 17960 19372 18012 19378
rect 17960 19314 18012 19320
rect 17960 16992 18012 16998
rect 17960 16934 18012 16940
rect 17972 16590 18000 16934
rect 17960 16584 18012 16590
rect 17960 16526 18012 16532
rect 17972 16114 18000 16526
rect 18248 16250 18276 20878
rect 18340 19922 18368 22066
rect 18512 21888 18564 21894
rect 18512 21830 18564 21836
rect 18420 20800 18472 20806
rect 18420 20742 18472 20748
rect 18328 19916 18380 19922
rect 18328 19858 18380 19864
rect 18340 19514 18368 19858
rect 18328 19508 18380 19514
rect 18328 19450 18380 19456
rect 18326 16552 18382 16561
rect 18326 16487 18382 16496
rect 18236 16244 18288 16250
rect 18236 16186 18288 16192
rect 17960 16108 18012 16114
rect 17960 16050 18012 16056
rect 18052 16108 18104 16114
rect 18052 16050 18104 16056
rect 17868 15632 17920 15638
rect 17868 15574 17920 15580
rect 18064 15502 18092 16050
rect 18144 15972 18196 15978
rect 18144 15914 18196 15920
rect 18052 15496 18104 15502
rect 18052 15438 18104 15444
rect 18064 15162 18092 15438
rect 18052 15156 18104 15162
rect 18052 15098 18104 15104
rect 17776 15020 17828 15026
rect 17776 14962 17828 14968
rect 17684 14884 17736 14890
rect 17684 14826 17736 14832
rect 17406 14512 17462 14521
rect 17406 14447 17462 14456
rect 17316 14408 17368 14414
rect 17368 14368 17540 14396
rect 17316 14350 17368 14356
rect 17512 13938 17540 14368
rect 17592 14340 17644 14346
rect 17592 14282 17644 14288
rect 17604 14074 17632 14282
rect 17592 14068 17644 14074
rect 17592 14010 17644 14016
rect 17696 13938 17724 14826
rect 17776 14816 17828 14822
rect 17776 14758 17828 14764
rect 17960 14816 18012 14822
rect 17960 14758 18012 14764
rect 17224 13932 17276 13938
rect 17224 13874 17276 13880
rect 17408 13932 17460 13938
rect 17408 13874 17460 13880
rect 17500 13932 17552 13938
rect 17500 13874 17552 13880
rect 17684 13932 17736 13938
rect 17684 13874 17736 13880
rect 17420 13818 17448 13874
rect 17144 13790 17448 13818
rect 16764 13252 16816 13258
rect 16764 13194 16816 13200
rect 17500 13252 17552 13258
rect 17500 13194 17552 13200
rect 17224 12980 17276 12986
rect 17224 12922 17276 12928
rect 17132 12844 17184 12850
rect 17132 12786 17184 12792
rect 16672 12436 16724 12442
rect 16672 12378 16724 12384
rect 17144 12306 17172 12786
rect 17132 12300 17184 12306
rect 17132 12242 17184 12248
rect 16764 12232 16816 12238
rect 16764 12174 16816 12180
rect 16672 12096 16724 12102
rect 16776 12073 16804 12174
rect 16672 12038 16724 12044
rect 16762 12064 16818 12073
rect 16580 11552 16632 11558
rect 16580 11494 16632 11500
rect 16486 11248 16542 11257
rect 16486 11183 16488 11192
rect 16540 11183 16542 11192
rect 16488 11154 16540 11160
rect 16224 7704 16436 7732
rect 16120 6792 16172 6798
rect 16120 6734 16172 6740
rect 16120 6452 16172 6458
rect 16120 6394 16172 6400
rect 16028 6384 16080 6390
rect 16028 6326 16080 6332
rect 15934 4992 15990 5001
rect 15934 4927 15990 4936
rect 15844 3528 15896 3534
rect 15844 3470 15896 3476
rect 15752 3460 15804 3466
rect 15752 3402 15804 3408
rect 15660 3188 15712 3194
rect 15660 3130 15712 3136
rect 15672 3097 15700 3130
rect 15658 3088 15714 3097
rect 15658 3023 15714 3032
rect 15660 2304 15712 2310
rect 15660 2246 15712 2252
rect 15672 2145 15700 2246
rect 15658 2136 15714 2145
rect 15658 2071 15714 2080
rect 15842 1864 15898 1873
rect 15842 1799 15898 1808
rect 15856 800 15884 1799
rect 16132 800 16160 6394
rect 16224 5409 16252 7704
rect 16488 7268 16540 7274
rect 16488 7210 16540 7216
rect 16304 6792 16356 6798
rect 16304 6734 16356 6740
rect 16316 5914 16344 6734
rect 16396 6112 16448 6118
rect 16396 6054 16448 6060
rect 16304 5908 16356 5914
rect 16304 5850 16356 5856
rect 16408 5710 16436 6054
rect 16396 5704 16448 5710
rect 16396 5646 16448 5652
rect 16210 5400 16266 5409
rect 16210 5335 16266 5344
rect 16302 3904 16358 3913
rect 16302 3839 16358 3848
rect 16316 3534 16344 3839
rect 16304 3528 16356 3534
rect 16304 3470 16356 3476
rect 16408 3126 16436 5646
rect 16396 3120 16448 3126
rect 16396 3062 16448 3068
rect 16500 2774 16528 7210
rect 16592 6866 16620 11494
rect 16684 10062 16712 12038
rect 16762 11999 16818 12008
rect 17132 11892 17184 11898
rect 17132 11834 17184 11840
rect 17144 11762 17172 11834
rect 17132 11756 17184 11762
rect 17132 11698 17184 11704
rect 17040 11620 17092 11626
rect 17040 11562 17092 11568
rect 17052 11150 17080 11562
rect 16764 11144 16816 11150
rect 16762 11112 16764 11121
rect 17040 11144 17092 11150
rect 16816 11112 16818 11121
rect 17040 11086 17092 11092
rect 16762 11047 16818 11056
rect 16948 11008 17000 11014
rect 17144 10962 17172 11698
rect 16948 10950 17000 10956
rect 16960 10810 16988 10950
rect 17052 10934 17172 10962
rect 16948 10804 17000 10810
rect 16948 10746 17000 10752
rect 16672 10056 16724 10062
rect 16672 9998 16724 10004
rect 16856 9920 16908 9926
rect 16856 9862 16908 9868
rect 16868 9586 16896 9862
rect 16856 9580 16908 9586
rect 16856 9522 16908 9528
rect 16764 8492 16816 8498
rect 16764 8434 16816 8440
rect 16672 8424 16724 8430
rect 16672 8366 16724 8372
rect 16580 6860 16632 6866
rect 16580 6802 16632 6808
rect 16684 6390 16712 8366
rect 16776 8090 16804 8434
rect 16764 8084 16816 8090
rect 16764 8026 16816 8032
rect 16764 7880 16816 7886
rect 16764 7822 16816 7828
rect 16776 7342 16804 7822
rect 16764 7336 16816 7342
rect 16764 7278 16816 7284
rect 16776 6934 16804 7278
rect 16764 6928 16816 6934
rect 16868 6905 16896 9522
rect 17052 8634 17080 10934
rect 17130 9616 17186 9625
rect 17236 9586 17264 12922
rect 17406 12608 17462 12617
rect 17406 12543 17462 12552
rect 17420 11626 17448 12543
rect 17408 11620 17460 11626
rect 17408 11562 17460 11568
rect 17314 11384 17370 11393
rect 17314 11319 17370 11328
rect 17328 11218 17356 11319
rect 17316 11212 17368 11218
rect 17316 11154 17368 11160
rect 17328 10810 17356 11154
rect 17316 10804 17368 10810
rect 17316 10746 17368 10752
rect 17316 10464 17368 10470
rect 17316 10406 17368 10412
rect 17328 10266 17356 10406
rect 17316 10260 17368 10266
rect 17316 10202 17368 10208
rect 17130 9551 17132 9560
rect 17184 9551 17186 9560
rect 17224 9580 17276 9586
rect 17132 9522 17184 9528
rect 17224 9522 17276 9528
rect 17144 9178 17172 9522
rect 17512 9178 17540 13194
rect 17788 12442 17816 14758
rect 17868 14612 17920 14618
rect 17868 14554 17920 14560
rect 17776 12436 17828 12442
rect 17776 12378 17828 12384
rect 17684 12232 17736 12238
rect 17880 12209 17908 14554
rect 17972 14482 18000 14758
rect 17960 14476 18012 14482
rect 17960 14418 18012 14424
rect 18052 13796 18104 13802
rect 18052 13738 18104 13744
rect 18064 12986 18092 13738
rect 18156 13190 18184 15914
rect 18340 15706 18368 16487
rect 18328 15700 18380 15706
rect 18328 15642 18380 15648
rect 18432 15586 18460 20742
rect 18340 15558 18460 15586
rect 18236 15360 18288 15366
rect 18236 15302 18288 15308
rect 18144 13184 18196 13190
rect 18144 13126 18196 13132
rect 18052 12980 18104 12986
rect 18052 12922 18104 12928
rect 17684 12174 17736 12180
rect 17866 12200 17922 12209
rect 17696 11286 17724 12174
rect 17866 12135 17922 12144
rect 17868 12096 17920 12102
rect 17866 12064 17868 12073
rect 17920 12064 17922 12073
rect 17866 11999 17922 12008
rect 18248 11694 18276 15302
rect 18340 14906 18368 15558
rect 18420 15428 18472 15434
rect 18420 15370 18472 15376
rect 18432 15094 18460 15370
rect 18420 15088 18472 15094
rect 18418 15056 18420 15065
rect 18472 15056 18474 15065
rect 18418 14991 18474 15000
rect 18340 14878 18460 14906
rect 18328 14068 18380 14074
rect 18328 14010 18380 14016
rect 18236 11688 18288 11694
rect 18236 11630 18288 11636
rect 17684 11280 17736 11286
rect 17684 11222 17736 11228
rect 18340 11218 18368 14010
rect 18432 11354 18460 14878
rect 18524 11937 18552 21830
rect 18616 20534 18644 28562
rect 19260 27946 19288 28698
rect 19340 28552 19392 28558
rect 19340 28494 19392 28500
rect 19352 28234 19380 28494
rect 19444 28422 19472 29038
rect 19904 28558 19932 29106
rect 19892 28552 19944 28558
rect 19892 28494 19944 28500
rect 20076 28552 20128 28558
rect 20128 28500 20208 28506
rect 20076 28494 20208 28500
rect 20088 28478 20208 28494
rect 19432 28416 19484 28422
rect 19432 28358 19484 28364
rect 20076 28416 20128 28422
rect 20076 28358 20128 28364
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 19352 28206 19472 28234
rect 19340 28076 19392 28082
rect 19444 28064 19472 28206
rect 20088 28082 20116 28358
rect 19524 28076 19576 28082
rect 19444 28036 19524 28064
rect 19340 28018 19392 28024
rect 19524 28018 19576 28024
rect 20076 28076 20128 28082
rect 20076 28018 20128 28024
rect 19248 27940 19300 27946
rect 19248 27882 19300 27888
rect 19352 27674 19380 28018
rect 19536 27878 19564 28018
rect 19984 28008 20036 28014
rect 19984 27950 20036 27956
rect 19524 27872 19576 27878
rect 19524 27814 19576 27820
rect 19340 27668 19392 27674
rect 19340 27610 19392 27616
rect 19800 27532 19852 27538
rect 19800 27474 19852 27480
rect 19812 27402 19840 27474
rect 19996 27470 20024 27950
rect 19892 27464 19944 27470
rect 19892 27406 19944 27412
rect 19984 27464 20036 27470
rect 19984 27406 20036 27412
rect 19800 27396 19852 27402
rect 19800 27338 19852 27344
rect 19904 27316 19932 27406
rect 19904 27288 20024 27316
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 19996 27130 20024 27288
rect 20180 27146 20208 28478
rect 21272 27668 21324 27674
rect 21272 27610 21324 27616
rect 20352 27600 20404 27606
rect 20352 27542 20404 27548
rect 20260 27464 20312 27470
rect 20260 27406 20312 27412
rect 20272 27334 20300 27406
rect 20364 27402 20392 27542
rect 20352 27396 20404 27402
rect 20352 27338 20404 27344
rect 20260 27328 20312 27334
rect 20260 27270 20312 27276
rect 19984 27124 20036 27130
rect 19984 27066 20036 27072
rect 20088 27118 20208 27146
rect 18972 26784 19024 26790
rect 18972 26726 19024 26732
rect 18788 23724 18840 23730
rect 18788 23666 18840 23672
rect 18800 21010 18828 23666
rect 18880 22024 18932 22030
rect 18880 21966 18932 21972
rect 18892 21185 18920 21966
rect 18878 21176 18934 21185
rect 18878 21111 18934 21120
rect 18892 21010 18920 21111
rect 18788 21004 18840 21010
rect 18788 20946 18840 20952
rect 18880 21004 18932 21010
rect 18880 20946 18932 20952
rect 18604 20528 18656 20534
rect 18604 20470 18656 20476
rect 18880 19848 18932 19854
rect 18880 19790 18932 19796
rect 18788 19372 18840 19378
rect 18788 19314 18840 19320
rect 18696 18420 18748 18426
rect 18696 18362 18748 18368
rect 18708 18193 18736 18362
rect 18800 18329 18828 19314
rect 18892 19310 18920 19790
rect 18880 19304 18932 19310
rect 18880 19246 18932 19252
rect 18892 18902 18920 19246
rect 18880 18896 18932 18902
rect 18880 18838 18932 18844
rect 18786 18320 18842 18329
rect 18786 18255 18788 18264
rect 18840 18255 18842 18264
rect 18788 18226 18840 18232
rect 18800 18195 18828 18226
rect 18694 18184 18750 18193
rect 18694 18119 18750 18128
rect 18708 17338 18736 18119
rect 18788 17876 18840 17882
rect 18788 17818 18840 17824
rect 18696 17332 18748 17338
rect 18696 17274 18748 17280
rect 18800 17066 18828 17818
rect 18788 17060 18840 17066
rect 18788 17002 18840 17008
rect 18984 16980 19012 26726
rect 19248 26308 19300 26314
rect 19248 26250 19300 26256
rect 19260 26042 19288 26250
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 19248 26036 19300 26042
rect 19248 25978 19300 25984
rect 19260 25770 19288 25978
rect 19984 25832 20036 25838
rect 19984 25774 20036 25780
rect 19248 25764 19300 25770
rect 19248 25706 19300 25712
rect 19996 25362 20024 25774
rect 19984 25356 20036 25362
rect 19984 25298 20036 25304
rect 19340 25152 19392 25158
rect 19340 25094 19392 25100
rect 19352 24682 19380 25094
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 19340 24676 19392 24682
rect 19260 24636 19340 24664
rect 19064 21548 19116 21554
rect 19064 21490 19116 21496
rect 19076 20602 19104 21490
rect 19156 21480 19208 21486
rect 19156 21422 19208 21428
rect 19168 20874 19196 21422
rect 19156 20868 19208 20874
rect 19156 20810 19208 20816
rect 19064 20596 19116 20602
rect 19064 20538 19116 20544
rect 19076 19310 19104 20538
rect 19064 19304 19116 19310
rect 19064 19246 19116 19252
rect 19260 18426 19288 24636
rect 19340 24618 19392 24624
rect 19432 24608 19484 24614
rect 19432 24550 19484 24556
rect 19444 24138 19472 24550
rect 19996 24206 20024 25298
rect 20088 24274 20116 27118
rect 20168 26988 20220 26994
rect 20168 26930 20220 26936
rect 20180 26314 20208 26930
rect 20168 26308 20220 26314
rect 20168 26250 20220 26256
rect 20168 24812 20220 24818
rect 20168 24754 20220 24760
rect 20180 24614 20208 24754
rect 20168 24608 20220 24614
rect 20168 24550 20220 24556
rect 20076 24268 20128 24274
rect 20076 24210 20128 24216
rect 19984 24200 20036 24206
rect 19984 24142 20036 24148
rect 20168 24200 20220 24206
rect 20168 24142 20220 24148
rect 19432 24132 19484 24138
rect 19432 24074 19484 24080
rect 19340 23724 19392 23730
rect 19340 23666 19392 23672
rect 19352 23322 19380 23666
rect 19340 23316 19392 23322
rect 19340 23258 19392 23264
rect 19352 22642 19380 23258
rect 19340 22636 19392 22642
rect 19340 22578 19392 22584
rect 19444 22234 19472 24074
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 20180 23662 20208 24142
rect 20168 23656 20220 23662
rect 20168 23598 20220 23604
rect 20076 23520 20128 23526
rect 20076 23462 20128 23468
rect 20088 23118 20116 23462
rect 20076 23112 20128 23118
rect 20076 23054 20128 23060
rect 19984 23044 20036 23050
rect 19984 22986 20036 22992
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 19996 22642 20024 22986
rect 19984 22636 20036 22642
rect 19984 22578 20036 22584
rect 19432 22228 19484 22234
rect 19432 22170 19484 22176
rect 20076 22228 20128 22234
rect 20076 22170 20128 22176
rect 19432 22024 19484 22030
rect 19432 21966 19484 21972
rect 19984 22024 20036 22030
rect 19984 21966 20036 21972
rect 19340 21956 19392 21962
rect 19340 21898 19392 21904
rect 19352 21418 19380 21898
rect 19444 21554 19472 21966
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 19800 21616 19852 21622
rect 19800 21558 19852 21564
rect 19432 21548 19484 21554
rect 19432 21490 19484 21496
rect 19340 21412 19392 21418
rect 19340 21354 19392 21360
rect 19444 20942 19472 21490
rect 19432 20936 19484 20942
rect 19432 20878 19484 20884
rect 19340 20868 19392 20874
rect 19340 20810 19392 20816
rect 19352 20534 19380 20810
rect 19340 20528 19392 20534
rect 19340 20470 19392 20476
rect 19352 19990 19380 20470
rect 19444 20466 19472 20878
rect 19812 20806 19840 21558
rect 19800 20800 19852 20806
rect 19800 20742 19852 20748
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 19432 20460 19484 20466
rect 19432 20402 19484 20408
rect 19340 19984 19392 19990
rect 19340 19926 19392 19932
rect 19444 19922 19472 20402
rect 19432 19916 19484 19922
rect 19432 19858 19484 19864
rect 19996 19802 20024 21966
rect 20088 21622 20116 22170
rect 20180 21690 20208 23598
rect 20272 22506 20300 27270
rect 20364 26926 20392 27338
rect 21284 26994 21312 27610
rect 21272 26988 21324 26994
rect 21272 26930 21324 26936
rect 20352 26920 20404 26926
rect 20352 26862 20404 26868
rect 20364 25906 20392 26862
rect 21284 26586 21312 26930
rect 21272 26580 21324 26586
rect 21272 26522 21324 26528
rect 20536 26308 20588 26314
rect 20536 26250 20588 26256
rect 20352 25900 20404 25906
rect 20352 25842 20404 25848
rect 20444 24948 20496 24954
rect 20444 24890 20496 24896
rect 20352 24812 20404 24818
rect 20352 24754 20404 24760
rect 20364 24410 20392 24754
rect 20456 24410 20484 24890
rect 20352 24404 20404 24410
rect 20352 24346 20404 24352
rect 20444 24404 20496 24410
rect 20444 24346 20496 24352
rect 20444 23044 20496 23050
rect 20444 22986 20496 22992
rect 20260 22500 20312 22506
rect 20260 22442 20312 22448
rect 20260 21888 20312 21894
rect 20260 21830 20312 21836
rect 20168 21684 20220 21690
rect 20168 21626 20220 21632
rect 20076 21616 20128 21622
rect 20076 21558 20128 21564
rect 20272 21554 20300 21830
rect 20456 21706 20484 22986
rect 20548 22030 20576 26250
rect 20720 25288 20772 25294
rect 20720 25230 20772 25236
rect 20732 24886 20760 25230
rect 21272 25152 21324 25158
rect 21272 25094 21324 25100
rect 20720 24880 20772 24886
rect 20720 24822 20772 24828
rect 20732 24750 20760 24822
rect 20720 24744 20772 24750
rect 20720 24686 20772 24692
rect 20628 24268 20680 24274
rect 20628 24210 20680 24216
rect 20640 23866 20668 24210
rect 21284 24206 21312 25094
rect 21272 24200 21324 24206
rect 21272 24142 21324 24148
rect 20628 23860 20680 23866
rect 20628 23802 20680 23808
rect 20628 23724 20680 23730
rect 20628 23666 20680 23672
rect 20536 22024 20588 22030
rect 20536 21966 20588 21972
rect 20456 21678 20576 21706
rect 20260 21548 20312 21554
rect 20444 21548 20496 21554
rect 20312 21508 20392 21536
rect 20260 21490 20312 21496
rect 20260 21412 20312 21418
rect 20260 21354 20312 21360
rect 20076 21344 20128 21350
rect 20076 21286 20128 21292
rect 19352 19774 20024 19802
rect 19248 18420 19300 18426
rect 19248 18362 19300 18368
rect 19260 18290 19288 18362
rect 19064 18284 19116 18290
rect 19064 18226 19116 18232
rect 19248 18284 19300 18290
rect 19248 18226 19300 18232
rect 19076 17746 19104 18226
rect 19064 17740 19116 17746
rect 19064 17682 19116 17688
rect 19076 17134 19104 17682
rect 19156 17604 19208 17610
rect 19156 17546 19208 17552
rect 19064 17128 19116 17134
rect 19064 17070 19116 17076
rect 18984 16952 19104 16980
rect 18972 16516 19024 16522
rect 18972 16458 19024 16464
rect 18984 16182 19012 16458
rect 18972 16176 19024 16182
rect 18972 16118 19024 16124
rect 18984 15434 19012 16118
rect 18972 15428 19024 15434
rect 18972 15370 19024 15376
rect 19076 15162 19104 16952
rect 19168 16522 19196 17546
rect 19248 17196 19300 17202
rect 19248 17138 19300 17144
rect 19260 16794 19288 17138
rect 19248 16788 19300 16794
rect 19248 16730 19300 16736
rect 19156 16516 19208 16522
rect 19156 16458 19208 16464
rect 19248 16448 19300 16454
rect 19248 16390 19300 16396
rect 19064 15156 19116 15162
rect 19064 15098 19116 15104
rect 19260 15094 19288 16390
rect 19352 15201 19380 19774
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 19984 18828 20036 18834
rect 19984 18770 20036 18776
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 19996 18290 20024 18770
rect 19984 18284 20036 18290
rect 19984 18226 20036 18232
rect 19616 18148 19668 18154
rect 19616 18090 19668 18096
rect 19628 17882 19656 18090
rect 19616 17876 19668 17882
rect 19616 17818 19668 17824
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 19996 17270 20024 18226
rect 19984 17264 20036 17270
rect 19984 17206 20036 17212
rect 19432 17196 19484 17202
rect 19432 17138 19484 17144
rect 19708 17196 19760 17202
rect 19708 17138 19760 17144
rect 19444 16250 19472 17138
rect 19614 16552 19670 16561
rect 19720 16538 19748 17138
rect 19996 16658 20024 17206
rect 19984 16652 20036 16658
rect 19984 16594 20036 16600
rect 19670 16510 19748 16538
rect 19984 16516 20036 16522
rect 19614 16487 19670 16496
rect 19628 16454 19656 16487
rect 19984 16458 20036 16464
rect 19616 16448 19668 16454
rect 19616 16390 19668 16396
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 19432 16244 19484 16250
rect 19432 16186 19484 16192
rect 19996 15706 20024 16458
rect 19984 15700 20036 15706
rect 19984 15642 20036 15648
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19338 15192 19394 15201
rect 19574 15195 19882 15204
rect 19338 15127 19394 15136
rect 19248 15088 19300 15094
rect 19248 15030 19300 15036
rect 18880 14952 18932 14958
rect 18880 14894 18932 14900
rect 18788 12980 18840 12986
rect 18788 12922 18840 12928
rect 18510 11928 18566 11937
rect 18800 11898 18828 12922
rect 18892 12918 18920 14894
rect 19352 14550 19380 15127
rect 19984 14884 20036 14890
rect 19984 14826 20036 14832
rect 19156 14544 19208 14550
rect 19156 14486 19208 14492
rect 19340 14544 19392 14550
rect 19340 14486 19392 14492
rect 19168 14006 19196 14486
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 19892 14068 19944 14074
rect 19892 14010 19944 14016
rect 19156 14000 19208 14006
rect 19156 13942 19208 13948
rect 19708 13932 19760 13938
rect 19708 13874 19760 13880
rect 19432 13864 19484 13870
rect 19432 13806 19484 13812
rect 18972 13796 19024 13802
rect 18972 13738 19024 13744
rect 18984 13394 19012 13738
rect 18972 13388 19024 13394
rect 18972 13330 19024 13336
rect 19064 13388 19116 13394
rect 19064 13330 19116 13336
rect 18984 12986 19012 13330
rect 19076 13297 19104 13330
rect 19444 13326 19472 13806
rect 19616 13728 19668 13734
rect 19616 13670 19668 13676
rect 19340 13320 19392 13326
rect 19062 13288 19118 13297
rect 19340 13262 19392 13268
rect 19432 13320 19484 13326
rect 19432 13262 19484 13268
rect 19062 13223 19118 13232
rect 18972 12980 19024 12986
rect 18972 12922 19024 12928
rect 18880 12912 18932 12918
rect 18880 12854 18932 12860
rect 19352 12850 19380 13262
rect 19340 12844 19392 12850
rect 19340 12786 19392 12792
rect 19154 12200 19210 12209
rect 19154 12135 19210 12144
rect 18510 11863 18566 11872
rect 18788 11892 18840 11898
rect 18788 11834 18840 11840
rect 18512 11756 18564 11762
rect 18512 11698 18564 11704
rect 18420 11348 18472 11354
rect 18420 11290 18472 11296
rect 18328 11212 18380 11218
rect 18328 11154 18380 11160
rect 18236 11144 18288 11150
rect 18236 11086 18288 11092
rect 18248 10033 18276 11086
rect 18328 11076 18380 11082
rect 18328 11018 18380 11024
rect 18340 10606 18368 11018
rect 18524 10674 18552 11698
rect 18972 11552 19024 11558
rect 18972 11494 19024 11500
rect 18604 11076 18656 11082
rect 18604 11018 18656 11024
rect 18512 10668 18564 10674
rect 18512 10610 18564 10616
rect 18328 10600 18380 10606
rect 18380 10560 18460 10588
rect 18328 10542 18380 10548
rect 18432 10062 18460 10560
rect 18420 10056 18472 10062
rect 18234 10024 18290 10033
rect 18420 9998 18472 10004
rect 18234 9959 18290 9968
rect 18432 9654 18460 9998
rect 18420 9648 18472 9654
rect 18420 9590 18472 9596
rect 18236 9444 18288 9450
rect 18236 9386 18288 9392
rect 18512 9444 18564 9450
rect 18512 9386 18564 9392
rect 17132 9172 17184 9178
rect 17132 9114 17184 9120
rect 17500 9172 17552 9178
rect 17500 9114 17552 9120
rect 17040 8628 17092 8634
rect 17040 8570 17092 8576
rect 17408 8288 17460 8294
rect 17408 8230 17460 8236
rect 17420 7886 17448 8230
rect 18248 7886 18276 9386
rect 18524 9178 18552 9386
rect 18512 9172 18564 9178
rect 18512 9114 18564 9120
rect 17132 7880 17184 7886
rect 17132 7822 17184 7828
rect 17408 7880 17460 7886
rect 17408 7822 17460 7828
rect 18236 7880 18288 7886
rect 18236 7822 18288 7828
rect 18512 7880 18564 7886
rect 18512 7822 18564 7828
rect 16948 7200 17000 7206
rect 16948 7142 17000 7148
rect 16764 6870 16816 6876
rect 16854 6896 16910 6905
rect 16854 6831 16910 6840
rect 16856 6656 16908 6662
rect 16856 6598 16908 6604
rect 16672 6384 16724 6390
rect 16672 6326 16724 6332
rect 16580 5092 16632 5098
rect 16580 5034 16632 5040
rect 16592 4554 16620 5034
rect 16684 4690 16712 6326
rect 16868 6322 16896 6598
rect 16856 6316 16908 6322
rect 16856 6258 16908 6264
rect 16764 5296 16816 5302
rect 16764 5238 16816 5244
rect 16672 4684 16724 4690
rect 16672 4626 16724 4632
rect 16580 4548 16632 4554
rect 16580 4490 16632 4496
rect 16592 4078 16620 4490
rect 16776 4486 16804 5238
rect 16764 4480 16816 4486
rect 16764 4422 16816 4428
rect 16580 4072 16632 4078
rect 16580 4014 16632 4020
rect 16592 3602 16620 4014
rect 16672 3936 16724 3942
rect 16672 3878 16724 3884
rect 16580 3596 16632 3602
rect 16580 3538 16632 3544
rect 16408 2746 16528 2774
rect 16408 800 16436 2746
rect 16684 800 16712 3878
rect 16776 3466 16804 4422
rect 16856 4140 16908 4146
rect 16856 4082 16908 4088
rect 16868 3534 16896 4082
rect 16856 3528 16908 3534
rect 16856 3470 16908 3476
rect 16764 3460 16816 3466
rect 16764 3402 16816 3408
rect 16764 2916 16816 2922
rect 16764 2858 16816 2864
rect 16776 2802 16804 2858
rect 16776 2774 16896 2802
rect 16868 2650 16896 2774
rect 16856 2644 16908 2650
rect 16856 2586 16908 2592
rect 16960 800 16988 7142
rect 17144 5710 17172 7822
rect 17224 6792 17276 6798
rect 17224 6734 17276 6740
rect 17132 5704 17184 5710
rect 17132 5646 17184 5652
rect 17040 4480 17092 4486
rect 17040 4422 17092 4428
rect 17052 4146 17080 4422
rect 17040 4140 17092 4146
rect 17040 4082 17092 4088
rect 17040 3528 17092 3534
rect 17092 3488 17172 3516
rect 17040 3470 17092 3476
rect 17040 2848 17092 2854
rect 17040 2790 17092 2796
rect 17052 1494 17080 2790
rect 17144 2582 17172 3488
rect 17132 2576 17184 2582
rect 17132 2518 17184 2524
rect 17040 1488 17092 1494
rect 17040 1430 17092 1436
rect 17236 800 17264 6734
rect 17420 5545 17448 7822
rect 18524 7750 18552 7822
rect 18328 7744 18380 7750
rect 18328 7686 18380 7692
rect 18512 7744 18564 7750
rect 18512 7686 18564 7692
rect 18340 7546 18368 7686
rect 18328 7540 18380 7546
rect 18328 7482 18380 7488
rect 17960 6792 18012 6798
rect 17960 6734 18012 6740
rect 17500 5704 17552 5710
rect 17500 5646 17552 5652
rect 17776 5704 17828 5710
rect 17776 5646 17828 5652
rect 17406 5536 17462 5545
rect 17406 5471 17462 5480
rect 17408 5160 17460 5166
rect 17314 5128 17370 5137
rect 17408 5102 17460 5108
rect 17314 5063 17370 5072
rect 17328 3058 17356 5063
rect 17420 4690 17448 5102
rect 17408 4684 17460 4690
rect 17408 4626 17460 4632
rect 17420 4214 17448 4626
rect 17408 4208 17460 4214
rect 17408 4150 17460 4156
rect 17316 3052 17368 3058
rect 17316 2994 17368 3000
rect 17512 800 17540 5646
rect 17592 5228 17644 5234
rect 17592 5170 17644 5176
rect 17604 4554 17632 5170
rect 17592 4548 17644 4554
rect 17592 4490 17644 4496
rect 17604 4010 17632 4490
rect 17592 4004 17644 4010
rect 17592 3946 17644 3952
rect 17604 3534 17632 3946
rect 17592 3528 17644 3534
rect 17592 3470 17644 3476
rect 17604 2650 17632 3470
rect 17592 2644 17644 2650
rect 17592 2586 17644 2592
rect 17788 800 17816 5646
rect 17868 4616 17920 4622
rect 17868 4558 17920 4564
rect 17880 4146 17908 4558
rect 17868 4140 17920 4146
rect 17868 4082 17920 4088
rect 17972 3942 18000 6734
rect 18512 6656 18564 6662
rect 18512 6598 18564 6604
rect 18328 5704 18380 5710
rect 18328 5646 18380 5652
rect 18144 5092 18196 5098
rect 18144 5034 18196 5040
rect 18052 4752 18104 4758
rect 18052 4694 18104 4700
rect 17960 3936 18012 3942
rect 17960 3878 18012 3884
rect 18064 800 18092 4694
rect 18156 3670 18184 5034
rect 18236 4140 18288 4146
rect 18236 4082 18288 4088
rect 18248 3738 18276 4082
rect 18236 3732 18288 3738
rect 18236 3674 18288 3680
rect 18144 3664 18196 3670
rect 18144 3606 18196 3612
rect 18234 2680 18290 2689
rect 18234 2615 18236 2624
rect 18288 2615 18290 2624
rect 18236 2586 18288 2592
rect 18248 2514 18276 2586
rect 18236 2508 18288 2514
rect 18236 2450 18288 2456
rect 18340 800 18368 5646
rect 18524 5302 18552 6598
rect 18616 6390 18644 11018
rect 18984 10577 19012 11494
rect 18970 10568 19026 10577
rect 18970 10503 19026 10512
rect 18788 9580 18840 9586
rect 18788 9522 18840 9528
rect 18800 8906 18828 9522
rect 18788 8900 18840 8906
rect 18788 8842 18840 8848
rect 19168 8838 19196 12135
rect 19248 11620 19300 11626
rect 19248 11562 19300 11568
rect 19156 8832 19208 8838
rect 19156 8774 19208 8780
rect 19260 8634 19288 11562
rect 19352 9994 19380 12786
rect 19444 12646 19472 13262
rect 19628 13190 19656 13670
rect 19720 13569 19748 13874
rect 19904 13841 19932 14010
rect 19890 13832 19946 13841
rect 19890 13767 19946 13776
rect 19706 13560 19762 13569
rect 19996 13530 20024 14826
rect 19706 13495 19762 13504
rect 19984 13524 20036 13530
rect 19984 13466 20036 13472
rect 19984 13320 20036 13326
rect 19984 13262 20036 13268
rect 19616 13184 19668 13190
rect 19616 13126 19668 13132
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 19432 12640 19484 12646
rect 19432 12582 19484 12588
rect 19996 12306 20024 13262
rect 19432 12300 19484 12306
rect 19432 12242 19484 12248
rect 19984 12300 20036 12306
rect 19984 12242 20036 12248
rect 19444 11540 19472 12242
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 20088 11762 20116 21286
rect 20168 21004 20220 21010
rect 20168 20946 20220 20952
rect 20180 20346 20208 20946
rect 20272 20466 20300 21354
rect 20364 20534 20392 21508
rect 20444 21490 20496 21496
rect 20456 21146 20484 21490
rect 20444 21140 20496 21146
rect 20444 21082 20496 21088
rect 20548 20754 20576 21678
rect 20640 21010 20668 23666
rect 20996 21956 21048 21962
rect 20996 21898 21048 21904
rect 21008 21690 21036 21898
rect 20996 21684 21048 21690
rect 20996 21626 21048 21632
rect 20904 21548 20956 21554
rect 20904 21490 20956 21496
rect 20628 21004 20680 21010
rect 20628 20946 20680 20952
rect 20916 20913 20944 21490
rect 21376 21078 21404 31726
rect 27172 29850 27200 56986
rect 30116 30258 30144 57190
rect 34934 57148 35242 57157
rect 34934 57146 34940 57148
rect 34996 57146 35020 57148
rect 35076 57146 35100 57148
rect 35156 57146 35180 57148
rect 35236 57146 35242 57148
rect 34996 57094 34998 57146
rect 35178 57094 35180 57146
rect 34934 57092 34940 57094
rect 34996 57092 35020 57094
rect 35076 57092 35100 57094
rect 35156 57092 35180 57094
rect 35236 57092 35242 57094
rect 34934 57083 35242 57092
rect 34934 56060 35242 56069
rect 34934 56058 34940 56060
rect 34996 56058 35020 56060
rect 35076 56058 35100 56060
rect 35156 56058 35180 56060
rect 35236 56058 35242 56060
rect 34996 56006 34998 56058
rect 35178 56006 35180 56058
rect 34934 56004 34940 56006
rect 34996 56004 35020 56006
rect 35076 56004 35100 56006
rect 35156 56004 35180 56006
rect 35236 56004 35242 56006
rect 34934 55995 35242 56004
rect 34934 54972 35242 54981
rect 34934 54970 34940 54972
rect 34996 54970 35020 54972
rect 35076 54970 35100 54972
rect 35156 54970 35180 54972
rect 35236 54970 35242 54972
rect 34996 54918 34998 54970
rect 35178 54918 35180 54970
rect 34934 54916 34940 54918
rect 34996 54916 35020 54918
rect 35076 54916 35100 54918
rect 35156 54916 35180 54918
rect 35236 54916 35242 54918
rect 34934 54907 35242 54916
rect 34934 53884 35242 53893
rect 34934 53882 34940 53884
rect 34996 53882 35020 53884
rect 35076 53882 35100 53884
rect 35156 53882 35180 53884
rect 35236 53882 35242 53884
rect 34996 53830 34998 53882
rect 35178 53830 35180 53882
rect 34934 53828 34940 53830
rect 34996 53828 35020 53830
rect 35076 53828 35100 53830
rect 35156 53828 35180 53830
rect 35236 53828 35242 53830
rect 34934 53819 35242 53828
rect 34934 52796 35242 52805
rect 34934 52794 34940 52796
rect 34996 52794 35020 52796
rect 35076 52794 35100 52796
rect 35156 52794 35180 52796
rect 35236 52794 35242 52796
rect 34996 52742 34998 52794
rect 35178 52742 35180 52794
rect 34934 52740 34940 52742
rect 34996 52740 35020 52742
rect 35076 52740 35100 52742
rect 35156 52740 35180 52742
rect 35236 52740 35242 52742
rect 34934 52731 35242 52740
rect 34934 51708 35242 51717
rect 34934 51706 34940 51708
rect 34996 51706 35020 51708
rect 35076 51706 35100 51708
rect 35156 51706 35180 51708
rect 35236 51706 35242 51708
rect 34996 51654 34998 51706
rect 35178 51654 35180 51706
rect 34934 51652 34940 51654
rect 34996 51652 35020 51654
rect 35076 51652 35100 51654
rect 35156 51652 35180 51654
rect 35236 51652 35242 51654
rect 34934 51643 35242 51652
rect 34934 50620 35242 50629
rect 34934 50618 34940 50620
rect 34996 50618 35020 50620
rect 35076 50618 35100 50620
rect 35156 50618 35180 50620
rect 35236 50618 35242 50620
rect 34996 50566 34998 50618
rect 35178 50566 35180 50618
rect 34934 50564 34940 50566
rect 34996 50564 35020 50566
rect 35076 50564 35100 50566
rect 35156 50564 35180 50566
rect 35236 50564 35242 50566
rect 34934 50555 35242 50564
rect 34934 49532 35242 49541
rect 34934 49530 34940 49532
rect 34996 49530 35020 49532
rect 35076 49530 35100 49532
rect 35156 49530 35180 49532
rect 35236 49530 35242 49532
rect 34996 49478 34998 49530
rect 35178 49478 35180 49530
rect 34934 49476 34940 49478
rect 34996 49476 35020 49478
rect 35076 49476 35100 49478
rect 35156 49476 35180 49478
rect 35236 49476 35242 49478
rect 34934 49467 35242 49476
rect 34934 48444 35242 48453
rect 34934 48442 34940 48444
rect 34996 48442 35020 48444
rect 35076 48442 35100 48444
rect 35156 48442 35180 48444
rect 35236 48442 35242 48444
rect 34996 48390 34998 48442
rect 35178 48390 35180 48442
rect 34934 48388 34940 48390
rect 34996 48388 35020 48390
rect 35076 48388 35100 48390
rect 35156 48388 35180 48390
rect 35236 48388 35242 48390
rect 34934 48379 35242 48388
rect 34934 47356 35242 47365
rect 34934 47354 34940 47356
rect 34996 47354 35020 47356
rect 35076 47354 35100 47356
rect 35156 47354 35180 47356
rect 35236 47354 35242 47356
rect 34996 47302 34998 47354
rect 35178 47302 35180 47354
rect 34934 47300 34940 47302
rect 34996 47300 35020 47302
rect 35076 47300 35100 47302
rect 35156 47300 35180 47302
rect 35236 47300 35242 47302
rect 34934 47291 35242 47300
rect 34934 46268 35242 46277
rect 34934 46266 34940 46268
rect 34996 46266 35020 46268
rect 35076 46266 35100 46268
rect 35156 46266 35180 46268
rect 35236 46266 35242 46268
rect 34996 46214 34998 46266
rect 35178 46214 35180 46266
rect 34934 46212 34940 46214
rect 34996 46212 35020 46214
rect 35076 46212 35100 46214
rect 35156 46212 35180 46214
rect 35236 46212 35242 46214
rect 34934 46203 35242 46212
rect 34934 45180 35242 45189
rect 34934 45178 34940 45180
rect 34996 45178 35020 45180
rect 35076 45178 35100 45180
rect 35156 45178 35180 45180
rect 35236 45178 35242 45180
rect 34996 45126 34998 45178
rect 35178 45126 35180 45178
rect 34934 45124 34940 45126
rect 34996 45124 35020 45126
rect 35076 45124 35100 45126
rect 35156 45124 35180 45126
rect 35236 45124 35242 45126
rect 34934 45115 35242 45124
rect 34934 44092 35242 44101
rect 34934 44090 34940 44092
rect 34996 44090 35020 44092
rect 35076 44090 35100 44092
rect 35156 44090 35180 44092
rect 35236 44090 35242 44092
rect 34996 44038 34998 44090
rect 35178 44038 35180 44090
rect 34934 44036 34940 44038
rect 34996 44036 35020 44038
rect 35076 44036 35100 44038
rect 35156 44036 35180 44038
rect 35236 44036 35242 44038
rect 34934 44027 35242 44036
rect 34934 43004 35242 43013
rect 34934 43002 34940 43004
rect 34996 43002 35020 43004
rect 35076 43002 35100 43004
rect 35156 43002 35180 43004
rect 35236 43002 35242 43004
rect 34996 42950 34998 43002
rect 35178 42950 35180 43002
rect 34934 42948 34940 42950
rect 34996 42948 35020 42950
rect 35076 42948 35100 42950
rect 35156 42948 35180 42950
rect 35236 42948 35242 42950
rect 34934 42939 35242 42948
rect 34934 41916 35242 41925
rect 34934 41914 34940 41916
rect 34996 41914 35020 41916
rect 35076 41914 35100 41916
rect 35156 41914 35180 41916
rect 35236 41914 35242 41916
rect 34996 41862 34998 41914
rect 35178 41862 35180 41914
rect 34934 41860 34940 41862
rect 34996 41860 35020 41862
rect 35076 41860 35100 41862
rect 35156 41860 35180 41862
rect 35236 41860 35242 41862
rect 34934 41851 35242 41860
rect 34934 40828 35242 40837
rect 34934 40826 34940 40828
rect 34996 40826 35020 40828
rect 35076 40826 35100 40828
rect 35156 40826 35180 40828
rect 35236 40826 35242 40828
rect 34996 40774 34998 40826
rect 35178 40774 35180 40826
rect 34934 40772 34940 40774
rect 34996 40772 35020 40774
rect 35076 40772 35100 40774
rect 35156 40772 35180 40774
rect 35236 40772 35242 40774
rect 34934 40763 35242 40772
rect 34934 39740 35242 39749
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39675 35242 39684
rect 34934 38652 35242 38661
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38587 35242 38596
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 30104 30252 30156 30258
rect 30104 30194 30156 30200
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 27160 29844 27212 29850
rect 27160 29786 27212 29792
rect 25780 29640 25832 29646
rect 25780 29582 25832 29588
rect 26424 29640 26476 29646
rect 26424 29582 26476 29588
rect 25044 29164 25096 29170
rect 25044 29106 25096 29112
rect 24400 28960 24452 28966
rect 24400 28902 24452 28908
rect 24412 28558 24440 28902
rect 25056 28558 25084 29106
rect 25792 28948 25820 29582
rect 25700 28920 25820 28948
rect 25700 28626 25728 28920
rect 26056 28756 26108 28762
rect 26056 28698 26108 28704
rect 25688 28620 25740 28626
rect 25688 28562 25740 28568
rect 22008 28552 22060 28558
rect 22008 28494 22060 28500
rect 23204 28552 23256 28558
rect 23204 28494 23256 28500
rect 23296 28552 23348 28558
rect 23296 28494 23348 28500
rect 24400 28552 24452 28558
rect 24400 28494 24452 28500
rect 25044 28552 25096 28558
rect 25044 28494 25096 28500
rect 25136 28552 25188 28558
rect 25136 28494 25188 28500
rect 22020 28422 22048 28494
rect 22008 28416 22060 28422
rect 22008 28358 22060 28364
rect 23216 28218 23244 28494
rect 23308 28218 23336 28494
rect 23572 28416 23624 28422
rect 23572 28358 23624 28364
rect 23204 28212 23256 28218
rect 23204 28154 23256 28160
rect 23296 28212 23348 28218
rect 23296 28154 23348 28160
rect 22376 28144 22428 28150
rect 22376 28086 22428 28092
rect 21456 26376 21508 26382
rect 21456 26318 21508 26324
rect 21468 25294 21496 26318
rect 21916 25696 21968 25702
rect 21916 25638 21968 25644
rect 22284 25696 22336 25702
rect 22284 25638 22336 25644
rect 21456 25288 21508 25294
rect 21456 25230 21508 25236
rect 21364 21072 21416 21078
rect 21364 21014 21416 21020
rect 20902 20904 20958 20913
rect 20628 20868 20680 20874
rect 20902 20839 20958 20848
rect 20628 20810 20680 20816
rect 20456 20726 20576 20754
rect 20352 20528 20404 20534
rect 20352 20470 20404 20476
rect 20260 20460 20312 20466
rect 20260 20402 20312 20408
rect 20180 20318 20300 20346
rect 20168 18760 20220 18766
rect 20168 18702 20220 18708
rect 20076 11756 20128 11762
rect 20076 11698 20128 11704
rect 19524 11552 19576 11558
rect 19444 11512 19524 11540
rect 19524 11494 19576 11500
rect 20076 11552 20128 11558
rect 20076 11494 20128 11500
rect 19432 11212 19484 11218
rect 19432 11154 19484 11160
rect 19340 9988 19392 9994
rect 19340 9930 19392 9936
rect 19340 9512 19392 9518
rect 19340 9454 19392 9460
rect 19352 8974 19380 9454
rect 19340 8968 19392 8974
rect 19340 8910 19392 8916
rect 19444 8786 19472 11154
rect 20088 11150 20116 11494
rect 20180 11354 20208 18702
rect 20272 17202 20300 20318
rect 20364 19854 20392 20470
rect 20352 19848 20404 19854
rect 20352 19790 20404 19796
rect 20352 19712 20404 19718
rect 20352 19654 20404 19660
rect 20260 17196 20312 17202
rect 20260 17138 20312 17144
rect 20260 16992 20312 16998
rect 20260 16934 20312 16940
rect 20272 16590 20300 16934
rect 20260 16584 20312 16590
rect 20260 16526 20312 16532
rect 20260 15496 20312 15502
rect 20260 15438 20312 15444
rect 20272 15162 20300 15438
rect 20260 15156 20312 15162
rect 20260 15098 20312 15104
rect 20258 13968 20314 13977
rect 20258 13903 20260 13912
rect 20312 13903 20314 13912
rect 20260 13874 20312 13880
rect 20364 13818 20392 19654
rect 20456 19242 20484 20726
rect 20534 20632 20590 20641
rect 20534 20567 20590 20576
rect 20548 20466 20576 20567
rect 20536 20460 20588 20466
rect 20536 20402 20588 20408
rect 20640 19990 20668 20810
rect 20916 20806 20944 20839
rect 20904 20800 20956 20806
rect 20904 20742 20956 20748
rect 20628 19984 20680 19990
rect 20628 19926 20680 19932
rect 20996 19304 21048 19310
rect 20996 19246 21048 19252
rect 20444 19236 20496 19242
rect 20444 19178 20496 19184
rect 20456 18834 20484 19178
rect 20536 19168 20588 19174
rect 20536 19110 20588 19116
rect 20444 18828 20496 18834
rect 20444 18770 20496 18776
rect 20548 18714 20576 19110
rect 20628 18760 20680 18766
rect 20456 18708 20628 18714
rect 20456 18702 20680 18708
rect 20456 18686 20668 18702
rect 20456 16998 20484 18686
rect 20628 18624 20680 18630
rect 20628 18566 20680 18572
rect 20444 16992 20496 16998
rect 20444 16934 20496 16940
rect 20456 14618 20484 16934
rect 20444 14612 20496 14618
rect 20640 14600 20668 18566
rect 20904 17808 20956 17814
rect 20904 17750 20956 17756
rect 20916 17270 20944 17750
rect 20904 17264 20956 17270
rect 20904 17206 20956 17212
rect 20916 17066 20944 17206
rect 20904 17060 20956 17066
rect 20904 17002 20956 17008
rect 20904 15020 20956 15026
rect 21008 15008 21036 19246
rect 21272 18080 21324 18086
rect 21272 18022 21324 18028
rect 21284 17678 21312 18022
rect 21468 17882 21496 25230
rect 21824 24812 21876 24818
rect 21824 24754 21876 24760
rect 21836 24614 21864 24754
rect 21824 24608 21876 24614
rect 21824 24550 21876 24556
rect 21732 24064 21784 24070
rect 21732 24006 21784 24012
rect 21640 23792 21692 23798
rect 21640 23734 21692 23740
rect 21548 21888 21600 21894
rect 21548 21830 21600 21836
rect 21560 20942 21588 21830
rect 21548 20936 21600 20942
rect 21548 20878 21600 20884
rect 21652 20534 21680 23734
rect 21744 23526 21772 24006
rect 21732 23520 21784 23526
rect 21732 23462 21784 23468
rect 21744 20942 21772 23462
rect 21836 23186 21864 24550
rect 21928 23798 21956 25638
rect 22008 24812 22060 24818
rect 22008 24754 22060 24760
rect 22192 24812 22244 24818
rect 22192 24754 22244 24760
rect 22020 24410 22048 24754
rect 22008 24404 22060 24410
rect 22008 24346 22060 24352
rect 22204 24342 22232 24754
rect 22192 24336 22244 24342
rect 22192 24278 22244 24284
rect 21916 23792 21968 23798
rect 21916 23734 21968 23740
rect 22192 23724 22244 23730
rect 22192 23666 22244 23672
rect 22204 23322 22232 23666
rect 21916 23316 21968 23322
rect 21916 23258 21968 23264
rect 22192 23316 22244 23322
rect 22192 23258 22244 23264
rect 21824 23180 21876 23186
rect 21824 23122 21876 23128
rect 21928 22030 21956 23258
rect 22296 22710 22324 25638
rect 22388 23866 22416 28086
rect 23480 28076 23532 28082
rect 23480 28018 23532 28024
rect 22468 27872 22520 27878
rect 22468 27814 22520 27820
rect 22480 27334 22508 27814
rect 23492 27713 23520 28018
rect 23478 27704 23534 27713
rect 23478 27639 23534 27648
rect 22468 27328 22520 27334
rect 22468 27270 22520 27276
rect 23204 27328 23256 27334
rect 23204 27270 23256 27276
rect 22468 25900 22520 25906
rect 22468 25842 22520 25848
rect 22480 24750 22508 25842
rect 22560 25152 22612 25158
rect 22560 25094 22612 25100
rect 22572 24818 22600 25094
rect 22560 24812 22612 24818
rect 22560 24754 22612 24760
rect 22468 24744 22520 24750
rect 22468 24686 22520 24692
rect 22468 24608 22520 24614
rect 22468 24550 22520 24556
rect 22744 24608 22796 24614
rect 22744 24550 22796 24556
rect 22480 24206 22508 24550
rect 22468 24200 22520 24206
rect 22468 24142 22520 24148
rect 22376 23860 22428 23866
rect 22376 23802 22428 23808
rect 22284 22704 22336 22710
rect 22284 22646 22336 22652
rect 22652 22636 22704 22642
rect 22652 22578 22704 22584
rect 22664 22234 22692 22578
rect 22652 22228 22704 22234
rect 22652 22170 22704 22176
rect 21824 22024 21876 22030
rect 21824 21966 21876 21972
rect 21916 22024 21968 22030
rect 21916 21966 21968 21972
rect 22192 22024 22244 22030
rect 22192 21966 22244 21972
rect 21836 21010 21864 21966
rect 22006 21448 22062 21457
rect 22204 21418 22232 21966
rect 22468 21956 22520 21962
rect 22468 21898 22520 21904
rect 22376 21548 22428 21554
rect 22376 21490 22428 21496
rect 22006 21383 22062 21392
rect 22192 21412 22244 21418
rect 21916 21344 21968 21350
rect 21916 21286 21968 21292
rect 21928 21078 21956 21286
rect 21916 21072 21968 21078
rect 21916 21014 21968 21020
rect 21824 21004 21876 21010
rect 21824 20946 21876 20952
rect 21732 20936 21784 20942
rect 21732 20878 21784 20884
rect 21732 20800 21784 20806
rect 21732 20742 21784 20748
rect 21640 20528 21692 20534
rect 21640 20470 21692 20476
rect 21744 19310 21772 20742
rect 21824 20596 21876 20602
rect 21824 20538 21876 20544
rect 21836 20262 21864 20538
rect 21928 20466 21956 21014
rect 22020 20942 22048 21383
rect 22192 21354 22244 21360
rect 22008 20936 22060 20942
rect 22008 20878 22060 20884
rect 22284 20596 22336 20602
rect 22284 20538 22336 20544
rect 21916 20460 21968 20466
rect 21916 20402 21968 20408
rect 22100 20460 22152 20466
rect 22100 20402 22152 20408
rect 22112 20330 22140 20402
rect 22100 20324 22152 20330
rect 22100 20266 22152 20272
rect 21824 20256 21876 20262
rect 21824 20198 21876 20204
rect 21824 19780 21876 19786
rect 21824 19722 21876 19728
rect 21732 19304 21784 19310
rect 21732 19246 21784 19252
rect 21836 19122 21864 19722
rect 21744 19094 21864 19122
rect 21744 18290 21772 19094
rect 21916 18760 21968 18766
rect 21916 18702 21968 18708
rect 21928 18426 21956 18702
rect 22112 18698 22140 20266
rect 22192 20052 22244 20058
rect 22192 19994 22244 20000
rect 22100 18692 22152 18698
rect 22100 18634 22152 18640
rect 21916 18420 21968 18426
rect 21916 18362 21968 18368
rect 21732 18284 21784 18290
rect 21732 18226 21784 18232
rect 21456 17876 21508 17882
rect 21456 17818 21508 17824
rect 21744 17678 21772 18226
rect 21928 17814 21956 18362
rect 22008 18284 22060 18290
rect 22008 18226 22060 18232
rect 22020 18193 22048 18226
rect 22006 18184 22062 18193
rect 22006 18119 22008 18128
rect 22060 18119 22062 18128
rect 22008 18090 22060 18096
rect 22020 18059 22048 18090
rect 21916 17808 21968 17814
rect 21916 17750 21968 17756
rect 21272 17672 21324 17678
rect 21272 17614 21324 17620
rect 21732 17672 21784 17678
rect 21732 17614 21784 17620
rect 21744 17542 21772 17614
rect 21732 17536 21784 17542
rect 21732 17478 21784 17484
rect 22112 17320 22140 18634
rect 22020 17292 22140 17320
rect 21272 17196 21324 17202
rect 21272 17138 21324 17144
rect 21284 15434 21312 17138
rect 22020 16590 22048 17292
rect 22204 17218 22232 19994
rect 22112 17190 22232 17218
rect 22112 16998 22140 17190
rect 22192 17128 22244 17134
rect 22192 17070 22244 17076
rect 22100 16992 22152 16998
rect 22100 16934 22152 16940
rect 22204 16726 22232 17070
rect 22192 16720 22244 16726
rect 22192 16662 22244 16668
rect 22008 16584 22060 16590
rect 22008 16526 22060 16532
rect 22100 16584 22152 16590
rect 22100 16526 22152 16532
rect 21732 16448 21784 16454
rect 21732 16390 21784 16396
rect 21744 16182 21772 16390
rect 21732 16176 21784 16182
rect 21732 16118 21784 16124
rect 22112 16046 22140 16526
rect 22100 16040 22152 16046
rect 22100 15982 22152 15988
rect 21272 15428 21324 15434
rect 21272 15370 21324 15376
rect 21824 15428 21876 15434
rect 21824 15370 21876 15376
rect 22008 15428 22060 15434
rect 22008 15370 22060 15376
rect 20956 14980 21036 15008
rect 20904 14962 20956 14968
rect 20812 14952 20864 14958
rect 20812 14894 20864 14900
rect 20444 14554 20496 14560
rect 20548 14572 20668 14600
rect 20442 14512 20498 14521
rect 20442 14447 20498 14456
rect 20456 14414 20484 14447
rect 20444 14408 20496 14414
rect 20444 14350 20496 14356
rect 20548 13870 20576 14572
rect 20628 14476 20680 14482
rect 20628 14418 20680 14424
rect 20272 13790 20392 13818
rect 20536 13864 20588 13870
rect 20536 13806 20588 13812
rect 20272 13734 20300 13790
rect 20260 13728 20312 13734
rect 20260 13670 20312 13676
rect 20352 13388 20404 13394
rect 20352 13330 20404 13336
rect 20260 12232 20312 12238
rect 20260 12174 20312 12180
rect 20272 11694 20300 12174
rect 20260 11688 20312 11694
rect 20260 11630 20312 11636
rect 20168 11348 20220 11354
rect 20168 11290 20220 11296
rect 20076 11144 20128 11150
rect 20076 11086 20128 11092
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 20088 10266 20116 11086
rect 20076 10260 20128 10266
rect 20076 10202 20128 10208
rect 20076 10124 20128 10130
rect 20076 10066 20128 10072
rect 19984 9920 20036 9926
rect 19984 9862 20036 9868
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 19996 9586 20024 9862
rect 19984 9580 20036 9586
rect 19984 9522 20036 9528
rect 20088 9178 20116 10066
rect 20180 10062 20208 11290
rect 20272 11082 20300 11630
rect 20260 11076 20312 11082
rect 20260 11018 20312 11024
rect 20168 10056 20220 10062
rect 20168 9998 20220 10004
rect 20168 9920 20220 9926
rect 20168 9862 20220 9868
rect 20076 9172 20128 9178
rect 20076 9114 20128 9120
rect 20180 8974 20208 9862
rect 20168 8968 20220 8974
rect 20168 8910 20220 8916
rect 19352 8758 19472 8786
rect 20076 8832 20128 8838
rect 20076 8774 20128 8780
rect 19248 8628 19300 8634
rect 19248 8570 19300 8576
rect 18696 8492 18748 8498
rect 18696 8434 18748 8440
rect 18972 8492 19024 8498
rect 18972 8434 19024 8440
rect 19156 8492 19208 8498
rect 19156 8434 19208 8440
rect 18708 7002 18736 8434
rect 18984 8090 19012 8434
rect 18972 8084 19024 8090
rect 18972 8026 19024 8032
rect 19168 7410 19196 8434
rect 19248 7812 19300 7818
rect 19248 7754 19300 7760
rect 19156 7404 19208 7410
rect 19156 7346 19208 7352
rect 18696 6996 18748 7002
rect 18696 6938 18748 6944
rect 18604 6384 18656 6390
rect 18604 6326 18656 6332
rect 18708 6322 18736 6938
rect 19168 6866 19196 7346
rect 19156 6860 19208 6866
rect 19156 6802 19208 6808
rect 19168 6322 19196 6802
rect 19260 6798 19288 7754
rect 19248 6792 19300 6798
rect 19248 6734 19300 6740
rect 18696 6316 18748 6322
rect 18696 6258 18748 6264
rect 18880 6316 18932 6322
rect 18880 6258 18932 6264
rect 19156 6316 19208 6322
rect 19156 6258 19208 6264
rect 18892 5914 18920 6258
rect 18880 5908 18932 5914
rect 18880 5850 18932 5856
rect 19260 5710 19288 6734
rect 19248 5704 19300 5710
rect 19248 5646 19300 5652
rect 19352 5370 19380 8758
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 20088 8566 20116 8774
rect 20076 8560 20128 8566
rect 20076 8502 20128 8508
rect 19432 8288 19484 8294
rect 19432 8230 19484 8236
rect 19444 7818 19472 8230
rect 19892 7880 19944 7886
rect 19892 7822 19944 7828
rect 19432 7812 19484 7818
rect 19432 7754 19484 7760
rect 19904 7732 19932 7822
rect 19904 7704 20024 7732
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 19432 7540 19484 7546
rect 19432 7482 19484 7488
rect 19444 6798 19472 7482
rect 19996 6866 20024 7704
rect 20088 7546 20116 8502
rect 20076 7540 20128 7546
rect 20076 7482 20128 7488
rect 19984 6860 20036 6866
rect 19984 6802 20036 6808
rect 19432 6792 19484 6798
rect 19432 6734 19484 6740
rect 19444 5710 19472 6734
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 19996 6254 20024 6802
rect 20076 6724 20128 6730
rect 20076 6666 20128 6672
rect 20088 6458 20116 6666
rect 20076 6452 20128 6458
rect 20076 6394 20128 6400
rect 19984 6248 20036 6254
rect 19984 6190 20036 6196
rect 19432 5704 19484 5710
rect 19432 5646 19484 5652
rect 19984 5704 20036 5710
rect 19984 5646 20036 5652
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 19340 5364 19392 5370
rect 19340 5306 19392 5312
rect 18512 5296 18564 5302
rect 18512 5238 18564 5244
rect 19708 5296 19760 5302
rect 19708 5238 19760 5244
rect 19432 5160 19484 5166
rect 19432 5102 19484 5108
rect 19340 5092 19392 5098
rect 19340 5034 19392 5040
rect 18880 5024 18932 5030
rect 18880 4966 18932 4972
rect 18604 4752 18656 4758
rect 18604 4694 18656 4700
rect 18512 3936 18564 3942
rect 18512 3878 18564 3884
rect 18420 3732 18472 3738
rect 18420 3674 18472 3680
rect 18432 2774 18460 3674
rect 18524 3670 18552 3878
rect 18512 3664 18564 3670
rect 18512 3606 18564 3612
rect 18432 2746 18552 2774
rect 18420 2440 18472 2446
rect 18420 2382 18472 2388
rect 18432 1766 18460 2382
rect 18420 1760 18472 1766
rect 18420 1702 18472 1708
rect 18524 1426 18552 2746
rect 18512 1420 18564 1426
rect 18512 1362 18564 1368
rect 18616 800 18644 4694
rect 18696 4072 18748 4078
rect 18696 4014 18748 4020
rect 18708 3738 18736 4014
rect 18696 3732 18748 3738
rect 18696 3674 18748 3680
rect 18892 800 18920 4966
rect 19156 4684 19208 4690
rect 19156 4626 19208 4632
rect 19064 4616 19116 4622
rect 19064 4558 19116 4564
rect 19076 2009 19104 4558
rect 19062 2000 19118 2009
rect 19062 1935 19118 1944
rect 19168 800 19196 4626
rect 19352 4622 19380 5034
rect 19444 4622 19472 5102
rect 19720 4622 19748 5238
rect 19996 5234 20024 5646
rect 19984 5228 20036 5234
rect 19984 5170 20036 5176
rect 19996 5030 20024 5170
rect 19984 5024 20036 5030
rect 19984 4966 20036 4972
rect 19996 4622 20024 4966
rect 19340 4616 19392 4622
rect 19340 4558 19392 4564
rect 19432 4616 19484 4622
rect 19432 4558 19484 4564
rect 19708 4616 19760 4622
rect 19708 4558 19760 4564
rect 19984 4616 20036 4622
rect 19984 4558 20036 4564
rect 19340 4140 19392 4146
rect 19340 4082 19392 4088
rect 19248 3392 19300 3398
rect 19248 3334 19300 3340
rect 19260 1902 19288 3334
rect 19352 2310 19380 4082
rect 19444 4049 19472 4558
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 19996 4146 20024 4558
rect 20180 4486 20208 8910
rect 20272 5370 20300 11018
rect 20364 10266 20392 13330
rect 20444 13252 20496 13258
rect 20444 13194 20496 13200
rect 20456 12434 20484 13194
rect 20456 12406 20576 12434
rect 20444 12096 20496 12102
rect 20444 12038 20496 12044
rect 20352 10260 20404 10266
rect 20352 10202 20404 10208
rect 20352 10124 20404 10130
rect 20352 10066 20404 10072
rect 20364 9994 20392 10066
rect 20352 9988 20404 9994
rect 20352 9930 20404 9936
rect 20364 8974 20392 9930
rect 20352 8968 20404 8974
rect 20456 8956 20484 12038
rect 20548 11762 20576 12406
rect 20536 11756 20588 11762
rect 20536 11698 20588 11704
rect 20548 11218 20576 11698
rect 20536 11212 20588 11218
rect 20536 11154 20588 11160
rect 20536 10600 20588 10606
rect 20536 10542 20588 10548
rect 20548 10062 20576 10542
rect 20640 10305 20668 14418
rect 20824 14346 20852 14894
rect 20812 14340 20864 14346
rect 20812 14282 20864 14288
rect 20904 14000 20956 14006
rect 20904 13942 20956 13948
rect 20720 13932 20772 13938
rect 20720 13874 20772 13880
rect 20732 13326 20760 13874
rect 20720 13320 20772 13326
rect 20720 13262 20772 13268
rect 20812 13252 20864 13258
rect 20812 13194 20864 13200
rect 20824 13025 20852 13194
rect 20810 13016 20866 13025
rect 20810 12951 20866 12960
rect 20720 12640 20772 12646
rect 20720 12582 20772 12588
rect 20732 12102 20760 12582
rect 20824 12442 20852 12951
rect 20916 12850 20944 13942
rect 21008 12986 21036 14980
rect 21272 14816 21324 14822
rect 21272 14758 21324 14764
rect 21088 14272 21140 14278
rect 21088 14214 21140 14220
rect 20996 12980 21048 12986
rect 20996 12922 21048 12928
rect 20904 12844 20956 12850
rect 20904 12786 20956 12792
rect 20812 12436 20864 12442
rect 20812 12378 20864 12384
rect 20720 12096 20772 12102
rect 20720 12038 20772 12044
rect 20720 11552 20772 11558
rect 20720 11494 20772 11500
rect 20732 11234 20760 11494
rect 20732 11218 20852 11234
rect 20732 11212 20864 11218
rect 20732 11206 20812 11212
rect 20626 10296 20682 10305
rect 20626 10231 20682 10240
rect 20732 10130 20760 11206
rect 20812 11154 20864 11160
rect 20916 11098 20944 12786
rect 20996 12436 21048 12442
rect 20996 12378 21048 12384
rect 21008 12170 21036 12378
rect 20996 12164 21048 12170
rect 20996 12106 21048 12112
rect 20996 11688 21048 11694
rect 20996 11630 21048 11636
rect 20824 11082 20944 11098
rect 20812 11076 20944 11082
rect 20864 11070 20944 11076
rect 20812 11018 20864 11024
rect 20720 10124 20772 10130
rect 20720 10066 20772 10072
rect 20536 10056 20588 10062
rect 20536 9998 20588 10004
rect 20548 9722 20576 9998
rect 20536 9716 20588 9722
rect 20536 9658 20588 9664
rect 20628 8968 20680 8974
rect 20456 8928 20628 8956
rect 20352 8910 20404 8916
rect 20628 8910 20680 8916
rect 20364 8786 20392 8910
rect 20364 8758 20576 8786
rect 20352 6656 20404 6662
rect 20352 6598 20404 6604
rect 20364 5778 20392 6598
rect 20444 6112 20496 6118
rect 20444 6054 20496 6060
rect 20352 5772 20404 5778
rect 20352 5714 20404 5720
rect 20260 5364 20312 5370
rect 20260 5306 20312 5312
rect 20168 4480 20220 4486
rect 20168 4422 20220 4428
rect 19984 4140 20036 4146
rect 19984 4082 20036 4088
rect 19430 4040 19486 4049
rect 19430 3975 19486 3984
rect 19432 3936 19484 3942
rect 19432 3878 19484 3884
rect 19984 3936 20036 3942
rect 19984 3878 20036 3884
rect 19444 3602 19472 3878
rect 19432 3596 19484 3602
rect 19432 3538 19484 3544
rect 19996 3466 20024 3878
rect 20076 3664 20128 3670
rect 20076 3606 20128 3612
rect 19432 3460 19484 3466
rect 19432 3402 19484 3408
rect 19984 3460 20036 3466
rect 19984 3402 20036 3408
rect 19340 2304 19392 2310
rect 19340 2246 19392 2252
rect 19248 1896 19300 1902
rect 19248 1838 19300 1844
rect 19352 1766 19380 2246
rect 19340 1760 19392 1766
rect 19340 1702 19392 1708
rect 19248 1420 19300 1426
rect 19248 1362 19300 1368
rect 19260 800 19288 1362
rect 19444 800 19472 3402
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 20088 3194 20116 3606
rect 20168 3528 20220 3534
rect 20168 3470 20220 3476
rect 20076 3188 20128 3194
rect 20076 3130 20128 3136
rect 20180 3074 20208 3470
rect 20088 3046 20208 3074
rect 19984 2984 20036 2990
rect 19984 2926 20036 2932
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 19800 1760 19852 1766
rect 19800 1702 19852 1708
rect 19708 1556 19760 1562
rect 19708 1498 19760 1504
rect 19524 1420 19576 1426
rect 19524 1362 19576 1368
rect 19536 800 19564 1362
rect 19720 800 19748 1498
rect 19812 800 19840 1702
rect 19996 800 20024 2926
rect 20088 1562 20116 3046
rect 20168 2984 20220 2990
rect 20168 2926 20220 2932
rect 20076 1556 20128 1562
rect 20076 1498 20128 1504
rect 20180 1442 20208 2926
rect 20260 2848 20312 2854
rect 20260 2790 20312 2796
rect 20088 1414 20208 1442
rect 20088 800 20116 1414
rect 20272 800 20300 2790
rect 20364 2106 20392 5714
rect 20456 5710 20484 6054
rect 20444 5704 20496 5710
rect 20444 5646 20496 5652
rect 20456 5574 20484 5646
rect 20444 5568 20496 5574
rect 20444 5510 20496 5516
rect 20456 5302 20484 5510
rect 20444 5296 20496 5302
rect 20444 5238 20496 5244
rect 20548 5114 20576 8758
rect 20456 5086 20576 5114
rect 20456 3913 20484 5086
rect 20536 4548 20588 4554
rect 20536 4490 20588 4496
rect 20548 4146 20576 4490
rect 20536 4140 20588 4146
rect 20536 4082 20588 4088
rect 20442 3904 20498 3913
rect 20442 3839 20498 3848
rect 20444 3528 20496 3534
rect 20444 3470 20496 3476
rect 20352 2100 20404 2106
rect 20352 2042 20404 2048
rect 20456 800 20484 3470
rect 20548 3194 20576 4082
rect 20640 4078 20668 8910
rect 20732 5778 20760 10066
rect 20824 10062 20852 11018
rect 20812 10056 20864 10062
rect 20812 9998 20864 10004
rect 20904 10056 20956 10062
rect 20904 9998 20956 10004
rect 20824 9722 20852 9998
rect 20812 9716 20864 9722
rect 20812 9658 20864 9664
rect 20812 9580 20864 9586
rect 20916 9568 20944 9998
rect 20864 9540 20944 9568
rect 20812 9522 20864 9528
rect 20824 9042 20852 9522
rect 21008 9518 21036 11630
rect 20996 9512 21048 9518
rect 20996 9454 21048 9460
rect 21100 9382 21128 14214
rect 21284 13394 21312 14758
rect 21272 13388 21324 13394
rect 21272 13330 21324 13336
rect 21640 13320 21692 13326
rect 21640 13262 21692 13268
rect 21652 12986 21680 13262
rect 21640 12980 21692 12986
rect 21640 12922 21692 12928
rect 21836 11665 21864 15370
rect 22020 14482 22048 15370
rect 22296 15178 22324 20538
rect 22388 20466 22416 21490
rect 22480 21486 22508 21898
rect 22468 21480 22520 21486
rect 22468 21422 22520 21428
rect 22480 20874 22508 21422
rect 22468 20868 22520 20874
rect 22468 20810 22520 20816
rect 22376 20460 22428 20466
rect 22376 20402 22428 20408
rect 22388 19378 22416 20402
rect 22376 19372 22428 19378
rect 22376 19314 22428 19320
rect 22388 18834 22416 19314
rect 22376 18828 22428 18834
rect 22376 18770 22428 18776
rect 22388 17610 22416 18770
rect 22376 17604 22428 17610
rect 22376 17546 22428 17552
rect 22376 16516 22428 16522
rect 22376 16458 22428 16464
rect 22388 16250 22416 16458
rect 22376 16244 22428 16250
rect 22376 16186 22428 16192
rect 22376 16108 22428 16114
rect 22376 16050 22428 16056
rect 22388 15994 22416 16050
rect 22480 15994 22508 20810
rect 22756 20369 22784 24550
rect 23112 23588 23164 23594
rect 23112 23530 23164 23536
rect 23124 23322 23152 23530
rect 23112 23316 23164 23322
rect 23112 23258 23164 23264
rect 22836 22772 22888 22778
rect 22836 22714 22888 22720
rect 22848 22642 22876 22714
rect 22836 22636 22888 22642
rect 22836 22578 22888 22584
rect 22836 22432 22888 22438
rect 22836 22374 22888 22380
rect 22742 20360 22798 20369
rect 22742 20295 22798 20304
rect 22560 19168 22612 19174
rect 22560 19110 22612 19116
rect 22572 18766 22600 19110
rect 22560 18760 22612 18766
rect 22560 18702 22612 18708
rect 22572 17882 22600 18702
rect 22560 17876 22612 17882
rect 22560 17818 22612 17824
rect 22848 17320 22876 22374
rect 22928 22024 22980 22030
rect 22928 21966 22980 21972
rect 23020 22024 23072 22030
rect 23020 21966 23072 21972
rect 22940 21865 22968 21966
rect 22926 21856 22982 21865
rect 22926 21791 22982 21800
rect 23032 21554 23060 21966
rect 23216 21894 23244 27270
rect 23584 27062 23612 28358
rect 24412 28082 24440 28494
rect 24400 28076 24452 28082
rect 24400 28018 24452 28024
rect 24308 27872 24360 27878
rect 24308 27814 24360 27820
rect 23572 27056 23624 27062
rect 23572 26998 23624 27004
rect 23572 26920 23624 26926
rect 23572 26862 23624 26868
rect 23480 25900 23532 25906
rect 23480 25842 23532 25848
rect 23492 25226 23520 25842
rect 23584 25838 23612 26862
rect 23756 26784 23808 26790
rect 23756 26726 23808 26732
rect 23572 25832 23624 25838
rect 23572 25774 23624 25780
rect 23480 25220 23532 25226
rect 23480 25162 23532 25168
rect 23664 25220 23716 25226
rect 23664 25162 23716 25168
rect 23386 24712 23442 24721
rect 23386 24647 23442 24656
rect 23400 24614 23428 24647
rect 23388 24608 23440 24614
rect 23388 24550 23440 24556
rect 23492 23798 23520 25162
rect 23676 24614 23704 25162
rect 23768 24818 23796 26726
rect 23848 25900 23900 25906
rect 23848 25842 23900 25848
rect 23860 25498 23888 25842
rect 23848 25492 23900 25498
rect 23848 25434 23900 25440
rect 23860 25378 23888 25434
rect 23860 25350 23980 25378
rect 23848 25220 23900 25226
rect 23848 25162 23900 25168
rect 23756 24812 23808 24818
rect 23756 24754 23808 24760
rect 23664 24608 23716 24614
rect 23664 24550 23716 24556
rect 23768 24426 23796 24754
rect 23676 24398 23796 24426
rect 23480 23792 23532 23798
rect 23480 23734 23532 23740
rect 23296 23724 23348 23730
rect 23296 23666 23348 23672
rect 23308 23050 23336 23666
rect 23492 23050 23520 23734
rect 23296 23044 23348 23050
rect 23296 22986 23348 22992
rect 23480 23044 23532 23050
rect 23480 22986 23532 22992
rect 23388 22976 23440 22982
rect 23388 22918 23440 22924
rect 23400 22438 23428 22918
rect 23480 22636 23532 22642
rect 23480 22578 23532 22584
rect 23388 22432 23440 22438
rect 23388 22374 23440 22380
rect 23492 22234 23520 22578
rect 23572 22432 23624 22438
rect 23572 22374 23624 22380
rect 23584 22273 23612 22374
rect 23570 22264 23626 22273
rect 23480 22228 23532 22234
rect 23570 22199 23626 22208
rect 23480 22170 23532 22176
rect 23492 22114 23520 22170
rect 23492 22086 23612 22114
rect 23204 21888 23256 21894
rect 23204 21830 23256 21836
rect 23388 21616 23440 21622
rect 23388 21558 23440 21564
rect 23480 21616 23532 21622
rect 23480 21558 23532 21564
rect 23020 21548 23072 21554
rect 23020 21490 23072 21496
rect 23032 20806 23060 21490
rect 23400 21185 23428 21558
rect 23386 21176 23442 21185
rect 23386 21111 23442 21120
rect 23020 20800 23072 20806
rect 23020 20742 23072 20748
rect 22928 20460 22980 20466
rect 22928 20402 22980 20408
rect 23388 20460 23440 20466
rect 23492 20448 23520 21558
rect 23584 21554 23612 22086
rect 23676 22094 23704 24398
rect 23676 22066 23796 22094
rect 23664 21888 23716 21894
rect 23664 21830 23716 21836
rect 23572 21548 23624 21554
rect 23572 21490 23624 21496
rect 23584 20602 23612 21490
rect 23572 20596 23624 20602
rect 23572 20538 23624 20544
rect 23676 20466 23704 21830
rect 23768 20874 23796 22066
rect 23756 20868 23808 20874
rect 23756 20810 23808 20816
rect 23440 20420 23520 20448
rect 23388 20402 23440 20408
rect 22940 20262 22968 20402
rect 22928 20256 22980 20262
rect 22928 20198 22980 20204
rect 23296 20256 23348 20262
rect 23296 20198 23348 20204
rect 23112 17876 23164 17882
rect 23112 17818 23164 17824
rect 22664 17292 22876 17320
rect 22558 16144 22614 16153
rect 22558 16079 22560 16088
rect 22612 16079 22614 16088
rect 22560 16050 22612 16056
rect 22388 15966 22508 15994
rect 22204 15150 22324 15178
rect 22008 14476 22060 14482
rect 22008 14418 22060 14424
rect 21916 14408 21968 14414
rect 21916 14350 21968 14356
rect 21928 12209 21956 14350
rect 22204 14346 22232 15150
rect 22284 15020 22336 15026
rect 22284 14962 22336 14968
rect 22296 14906 22324 14962
rect 22296 14878 22416 14906
rect 22192 14340 22244 14346
rect 22192 14282 22244 14288
rect 22388 14278 22416 14878
rect 22376 14272 22428 14278
rect 22376 14214 22428 14220
rect 22192 14068 22244 14074
rect 22192 14010 22244 14016
rect 22008 13320 22060 13326
rect 22008 13262 22060 13268
rect 22020 12646 22048 13262
rect 22204 12918 22232 14010
rect 22284 12980 22336 12986
rect 22284 12922 22336 12928
rect 22192 12912 22244 12918
rect 22192 12854 22244 12860
rect 22008 12640 22060 12646
rect 22008 12582 22060 12588
rect 22296 12434 22324 12922
rect 22388 12753 22416 14214
rect 22480 13530 22508 15966
rect 22560 14816 22612 14822
rect 22560 14758 22612 14764
rect 22572 14074 22600 14758
rect 22560 14068 22612 14074
rect 22560 14010 22612 14016
rect 22468 13524 22520 13530
rect 22468 13466 22520 13472
rect 22560 13320 22612 13326
rect 22560 13262 22612 13268
rect 22572 12986 22600 13262
rect 22560 12980 22612 12986
rect 22560 12922 22612 12928
rect 22374 12744 22430 12753
rect 22374 12679 22430 12688
rect 22204 12406 22324 12434
rect 22204 12238 22232 12406
rect 22192 12232 22244 12238
rect 21914 12200 21970 12209
rect 22192 12174 22244 12180
rect 21914 12135 21970 12144
rect 22100 12164 22152 12170
rect 22100 12106 22152 12112
rect 21822 11656 21878 11665
rect 21822 11591 21878 11600
rect 22112 11354 22140 12106
rect 22204 11642 22232 12174
rect 22376 11756 22428 11762
rect 22376 11698 22428 11704
rect 22204 11626 22324 11642
rect 22204 11620 22336 11626
rect 22204 11614 22284 11620
rect 22100 11348 22152 11354
rect 22100 11290 22152 11296
rect 22204 11150 22232 11614
rect 22284 11562 22336 11568
rect 22388 11354 22416 11698
rect 22376 11348 22428 11354
rect 22376 11290 22428 11296
rect 22192 11144 22244 11150
rect 22192 11086 22244 11092
rect 22204 10810 22232 11086
rect 22560 11076 22612 11082
rect 22560 11018 22612 11024
rect 22192 10804 22244 10810
rect 22192 10746 22244 10752
rect 22284 10668 22336 10674
rect 22284 10610 22336 10616
rect 22296 9994 22324 10610
rect 22284 9988 22336 9994
rect 22284 9930 22336 9936
rect 21272 9648 21324 9654
rect 21272 9590 21324 9596
rect 21088 9376 21140 9382
rect 21088 9318 21140 9324
rect 20812 9036 20864 9042
rect 20812 8978 20864 8984
rect 20720 5772 20772 5778
rect 20720 5714 20772 5720
rect 20720 5636 20772 5642
rect 20720 5578 20772 5584
rect 20732 5080 20760 5578
rect 20824 5370 20852 8978
rect 21178 8936 21234 8945
rect 21178 8871 21180 8880
rect 21232 8871 21234 8880
rect 21180 8842 21232 8848
rect 21088 7880 21140 7886
rect 21088 7822 21140 7828
rect 21100 7410 21128 7822
rect 21088 7404 21140 7410
rect 21088 7346 21140 7352
rect 21100 6798 21128 7346
rect 21088 6792 21140 6798
rect 21088 6734 21140 6740
rect 21100 6322 21128 6734
rect 21088 6316 21140 6322
rect 21088 6258 21140 6264
rect 20904 6112 20956 6118
rect 20904 6054 20956 6060
rect 20812 5364 20864 5370
rect 20812 5306 20864 5312
rect 20812 5092 20864 5098
rect 20732 5052 20812 5080
rect 20812 5034 20864 5040
rect 20824 4146 20852 5034
rect 20812 4140 20864 4146
rect 20812 4082 20864 4088
rect 20628 4072 20680 4078
rect 20824 4049 20852 4082
rect 20628 4014 20680 4020
rect 20810 4040 20866 4049
rect 20916 4010 20944 6054
rect 21088 5160 21140 5166
rect 21088 5102 21140 5108
rect 21100 4146 21128 5102
rect 21284 4826 21312 9590
rect 22296 9586 22324 9930
rect 22572 9654 22600 11018
rect 22664 10470 22692 17292
rect 22836 17196 22888 17202
rect 22836 17138 22888 17144
rect 22744 15904 22796 15910
rect 22744 15846 22796 15852
rect 22756 15162 22784 15846
rect 22848 15366 22876 17138
rect 22836 15360 22888 15366
rect 22836 15302 22888 15308
rect 22744 15156 22796 15162
rect 22744 15098 22796 15104
rect 22928 15088 22980 15094
rect 22928 15030 22980 15036
rect 22836 13864 22888 13870
rect 22836 13806 22888 13812
rect 22652 10464 22704 10470
rect 22652 10406 22704 10412
rect 22560 9648 22612 9654
rect 22560 9590 22612 9596
rect 22284 9580 22336 9586
rect 22284 9522 22336 9528
rect 21640 8900 21692 8906
rect 21640 8842 21692 8848
rect 21652 7954 21680 8842
rect 22100 8832 22152 8838
rect 22100 8774 22152 8780
rect 22112 8498 22140 8774
rect 22100 8492 22152 8498
rect 22100 8434 22152 8440
rect 21640 7948 21692 7954
rect 21640 7890 21692 7896
rect 22112 6866 22140 8434
rect 22192 7812 22244 7818
rect 22192 7754 22244 7760
rect 22204 7478 22232 7754
rect 22192 7472 22244 7478
rect 22192 7414 22244 7420
rect 22192 7200 22244 7206
rect 22192 7142 22244 7148
rect 22100 6860 22152 6866
rect 22100 6802 22152 6808
rect 22112 5234 22140 6802
rect 22204 6798 22232 7142
rect 22192 6792 22244 6798
rect 22192 6734 22244 6740
rect 22192 6316 22244 6322
rect 22192 6258 22244 6264
rect 22100 5228 22152 5234
rect 22100 5170 22152 5176
rect 22204 4826 22232 6258
rect 21272 4820 21324 4826
rect 21272 4762 21324 4768
rect 22192 4820 22244 4826
rect 22192 4762 22244 4768
rect 22204 4622 22232 4762
rect 22192 4616 22244 4622
rect 22192 4558 22244 4564
rect 22192 4480 22244 4486
rect 22192 4422 22244 4428
rect 22204 4282 22232 4422
rect 22192 4276 22244 4282
rect 22192 4218 22244 4224
rect 22296 4214 22324 9522
rect 22560 7472 22612 7478
rect 22560 7414 22612 7420
rect 22468 7404 22520 7410
rect 22468 7346 22520 7352
rect 22376 7268 22428 7274
rect 22376 7210 22428 7216
rect 22284 4208 22336 4214
rect 22284 4150 22336 4156
rect 21088 4140 21140 4146
rect 21088 4082 21140 4088
rect 20810 3975 20866 3984
rect 20904 4004 20956 4010
rect 20904 3946 20956 3952
rect 20628 3936 20680 3942
rect 20628 3878 20680 3884
rect 20536 3188 20588 3194
rect 20536 3130 20588 3136
rect 20640 1426 20668 3878
rect 22388 3738 22416 7210
rect 22480 6458 22508 7346
rect 22468 6452 22520 6458
rect 22468 6394 22520 6400
rect 22572 4758 22600 7414
rect 22652 7404 22704 7410
rect 22652 7346 22704 7352
rect 22664 6322 22692 7346
rect 22652 6316 22704 6322
rect 22652 6258 22704 6264
rect 22652 5772 22704 5778
rect 22652 5714 22704 5720
rect 22664 5234 22692 5714
rect 22848 5370 22876 13806
rect 22940 12306 22968 15030
rect 23020 14544 23072 14550
rect 23020 14486 23072 14492
rect 22928 12300 22980 12306
rect 22928 12242 22980 12248
rect 22940 12102 22968 12133
rect 22928 12096 22980 12102
rect 22926 12064 22928 12073
rect 22980 12064 22982 12073
rect 22926 11999 22982 12008
rect 22940 11762 22968 11999
rect 22928 11756 22980 11762
rect 22928 11698 22980 11704
rect 23032 10470 23060 14486
rect 23020 10464 23072 10470
rect 23020 10406 23072 10412
rect 23124 8974 23152 17818
rect 23204 16176 23256 16182
rect 23204 16118 23256 16124
rect 23216 14618 23244 16118
rect 23204 14612 23256 14618
rect 23204 14554 23256 14560
rect 23308 12434 23336 20198
rect 23388 19916 23440 19922
rect 23388 19858 23440 19864
rect 23400 13326 23428 19858
rect 23492 19854 23520 20420
rect 23664 20460 23716 20466
rect 23664 20402 23716 20408
rect 23480 19848 23532 19854
rect 23480 19790 23532 19796
rect 23480 19372 23532 19378
rect 23480 19314 23532 19320
rect 23492 16794 23520 19314
rect 23572 19304 23624 19310
rect 23572 19246 23624 19252
rect 23584 18358 23612 19246
rect 23572 18352 23624 18358
rect 23572 18294 23624 18300
rect 23584 17882 23612 18294
rect 23664 18080 23716 18086
rect 23664 18022 23716 18028
rect 23572 17876 23624 17882
rect 23572 17818 23624 17824
rect 23480 16788 23532 16794
rect 23480 16730 23532 16736
rect 23584 16726 23612 17818
rect 23572 16720 23624 16726
rect 23572 16662 23624 16668
rect 23480 15904 23532 15910
rect 23480 15846 23532 15852
rect 23492 15026 23520 15846
rect 23570 15056 23626 15065
rect 23480 15020 23532 15026
rect 23570 14991 23626 15000
rect 23480 14962 23532 14968
rect 23388 13320 23440 13326
rect 23388 13262 23440 13268
rect 23216 12406 23336 12434
rect 23216 11830 23244 12406
rect 23296 11892 23348 11898
rect 23296 11834 23348 11840
rect 23204 11824 23256 11830
rect 23308 11801 23336 11834
rect 23204 11766 23256 11772
rect 23294 11792 23350 11801
rect 23294 11727 23350 11736
rect 23400 11642 23428 13262
rect 23478 13016 23534 13025
rect 23478 12951 23534 12960
rect 23492 12918 23520 12951
rect 23480 12912 23532 12918
rect 23480 12854 23532 12860
rect 23478 12744 23534 12753
rect 23478 12679 23534 12688
rect 23492 12306 23520 12679
rect 23480 12300 23532 12306
rect 23480 12242 23532 12248
rect 23480 11756 23532 11762
rect 23480 11698 23532 11704
rect 23492 11642 23520 11698
rect 23400 11614 23520 11642
rect 23400 10606 23428 11614
rect 23388 10600 23440 10606
rect 23388 10542 23440 10548
rect 23296 10464 23348 10470
rect 23296 10406 23348 10412
rect 23308 10062 23336 10406
rect 23296 10056 23348 10062
rect 23296 9998 23348 10004
rect 23112 8968 23164 8974
rect 23112 8910 23164 8916
rect 23112 7744 23164 7750
rect 23112 7686 23164 7692
rect 22836 5364 22888 5370
rect 22836 5306 22888 5312
rect 22652 5228 22704 5234
rect 22652 5170 22704 5176
rect 22560 4752 22612 4758
rect 22560 4694 22612 4700
rect 22664 4146 22692 5170
rect 22848 4729 22876 5306
rect 22928 5228 22980 5234
rect 22928 5170 22980 5176
rect 22940 4826 22968 5170
rect 22928 4820 22980 4826
rect 22928 4762 22980 4768
rect 22834 4720 22890 4729
rect 22834 4655 22890 4664
rect 22848 4622 22876 4655
rect 22836 4616 22888 4622
rect 22836 4558 22888 4564
rect 22652 4140 22704 4146
rect 22652 4082 22704 4088
rect 22376 3732 22428 3738
rect 22376 3674 22428 3680
rect 21548 3528 21600 3534
rect 21548 3470 21600 3476
rect 22376 3528 22428 3534
rect 22376 3470 22428 3476
rect 20996 2848 21048 2854
rect 20996 2790 21048 2796
rect 20720 2440 20772 2446
rect 20720 2382 20772 2388
rect 20628 1420 20680 1426
rect 20628 1362 20680 1368
rect 20732 800 20760 2382
rect 21008 800 21036 2790
rect 21272 2576 21324 2582
rect 21272 2518 21324 2524
rect 21284 800 21312 2518
rect 21560 800 21588 3470
rect 21732 3052 21784 3058
rect 21732 2994 21784 3000
rect 21744 2650 21772 2994
rect 21824 2984 21876 2990
rect 21824 2926 21876 2932
rect 21732 2644 21784 2650
rect 21732 2586 21784 2592
rect 21836 800 21864 2926
rect 22100 2440 22152 2446
rect 22100 2382 22152 2388
rect 22112 800 22140 2382
rect 22388 800 22416 3470
rect 22652 2848 22704 2854
rect 22652 2790 22704 2796
rect 22928 2848 22980 2854
rect 22928 2790 22980 2796
rect 22664 800 22692 2790
rect 22940 800 22968 2790
rect 23124 2650 23152 7686
rect 23308 7342 23336 9998
rect 23388 9580 23440 9586
rect 23388 9522 23440 9528
rect 23400 9178 23428 9522
rect 23388 9172 23440 9178
rect 23388 9114 23440 9120
rect 23584 8498 23612 14991
rect 23676 13258 23704 18022
rect 23860 17338 23888 25162
rect 23952 24750 23980 25350
rect 24216 25288 24268 25294
rect 24216 25230 24268 25236
rect 24228 24818 24256 25230
rect 24216 24812 24268 24818
rect 24216 24754 24268 24760
rect 23940 24744 23992 24750
rect 23940 24686 23992 24692
rect 23952 22794 23980 24686
rect 24124 24132 24176 24138
rect 24124 24074 24176 24080
rect 23952 22778 24072 22794
rect 23952 22772 24084 22778
rect 23952 22766 24032 22772
rect 24032 22714 24084 22720
rect 23940 22704 23992 22710
rect 23940 22646 23992 22652
rect 23952 21622 23980 22646
rect 23940 21616 23992 21622
rect 23940 21558 23992 21564
rect 24032 21344 24084 21350
rect 24032 21286 24084 21292
rect 24044 20777 24072 21286
rect 24030 20768 24086 20777
rect 24030 20703 24086 20712
rect 23940 18216 23992 18222
rect 23940 18158 23992 18164
rect 23952 17814 23980 18158
rect 23940 17808 23992 17814
rect 23940 17750 23992 17756
rect 23848 17332 23900 17338
rect 23848 17274 23900 17280
rect 23952 17202 23980 17750
rect 23940 17196 23992 17202
rect 23940 17138 23992 17144
rect 23756 16652 23808 16658
rect 23756 16594 23808 16600
rect 23768 16114 23796 16594
rect 24136 16250 24164 24074
rect 24228 23730 24256 24754
rect 24216 23724 24268 23730
rect 24216 23666 24268 23672
rect 24228 23186 24256 23666
rect 24216 23180 24268 23186
rect 24216 23122 24268 23128
rect 24320 22094 24348 27814
rect 25056 27674 25084 28494
rect 25148 28422 25176 28494
rect 25700 28490 25728 28562
rect 26068 28558 26096 28698
rect 26056 28552 26108 28558
rect 26056 28494 26108 28500
rect 25688 28484 25740 28490
rect 25688 28426 25740 28432
rect 25136 28416 25188 28422
rect 25136 28358 25188 28364
rect 25596 28416 25648 28422
rect 25596 28358 25648 28364
rect 25148 28082 25176 28358
rect 25608 28082 25636 28358
rect 25700 28218 25728 28426
rect 25688 28212 25740 28218
rect 25688 28154 25740 28160
rect 25136 28076 25188 28082
rect 25136 28018 25188 28024
rect 25596 28076 25648 28082
rect 25596 28018 25648 28024
rect 25044 27668 25096 27674
rect 25044 27610 25096 27616
rect 25148 27130 25176 28018
rect 26436 27878 26464 29582
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 26792 28416 26844 28422
rect 26792 28358 26844 28364
rect 26424 27872 26476 27878
rect 26424 27814 26476 27820
rect 26804 27674 26832 28358
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 26792 27668 26844 27674
rect 26792 27610 26844 27616
rect 27896 27464 27948 27470
rect 27896 27406 27948 27412
rect 26976 27396 27028 27402
rect 26976 27338 27028 27344
rect 26988 27130 27016 27338
rect 25136 27124 25188 27130
rect 25136 27066 25188 27072
rect 26976 27124 27028 27130
rect 26976 27066 27028 27072
rect 25320 27056 25372 27062
rect 25320 26998 25372 27004
rect 25332 26586 25360 26998
rect 25780 26988 25832 26994
rect 25780 26930 25832 26936
rect 25320 26580 25372 26586
rect 25320 26522 25372 26528
rect 25792 26382 25820 26930
rect 25320 26376 25372 26382
rect 25320 26318 25372 26324
rect 25780 26376 25832 26382
rect 25780 26318 25832 26324
rect 25136 25900 25188 25906
rect 25136 25842 25188 25848
rect 24768 25832 24820 25838
rect 24768 25774 24820 25780
rect 24400 25696 24452 25702
rect 24400 25638 24452 25644
rect 24584 25696 24636 25702
rect 24584 25638 24636 25644
rect 24412 24818 24440 25638
rect 24596 25226 24624 25638
rect 24676 25424 24728 25430
rect 24676 25366 24728 25372
rect 24584 25220 24636 25226
rect 24584 25162 24636 25168
rect 24688 24954 24716 25366
rect 24492 24948 24544 24954
rect 24492 24890 24544 24896
rect 24676 24948 24728 24954
rect 24676 24890 24728 24896
rect 24400 24812 24452 24818
rect 24400 24754 24452 24760
rect 24504 23730 24532 24890
rect 24676 24676 24728 24682
rect 24676 24618 24728 24624
rect 24688 24410 24716 24618
rect 24676 24404 24728 24410
rect 24676 24346 24728 24352
rect 24780 24206 24808 25774
rect 25148 25498 25176 25842
rect 25136 25492 25188 25498
rect 25136 25434 25188 25440
rect 24768 24200 24820 24206
rect 24768 24142 24820 24148
rect 24676 24132 24728 24138
rect 24676 24074 24728 24080
rect 24860 24132 24912 24138
rect 24860 24074 24912 24080
rect 24688 23730 24716 24074
rect 24872 23866 24900 24074
rect 24860 23860 24912 23866
rect 24860 23802 24912 23808
rect 24492 23724 24544 23730
rect 24492 23666 24544 23672
rect 24676 23724 24728 23730
rect 24676 23666 24728 23672
rect 25042 23080 25098 23089
rect 25042 23015 25044 23024
rect 25096 23015 25098 23024
rect 25044 22986 25096 22992
rect 24860 22704 24912 22710
rect 24860 22646 24912 22652
rect 24768 22636 24820 22642
rect 24768 22578 24820 22584
rect 24320 22066 24440 22094
rect 24412 22001 24440 22066
rect 24780 22030 24808 22578
rect 24768 22024 24820 22030
rect 24398 21992 24454 22001
rect 24768 21966 24820 21972
rect 24398 21927 24454 21936
rect 24492 21888 24544 21894
rect 24490 21856 24492 21865
rect 24544 21856 24546 21865
rect 24490 21791 24546 21800
rect 24308 21548 24360 21554
rect 24308 21490 24360 21496
rect 24320 21049 24348 21490
rect 24306 21040 24362 21049
rect 24306 20975 24362 20984
rect 24400 20460 24452 20466
rect 24400 20402 24452 20408
rect 24412 20058 24440 20402
rect 24400 20052 24452 20058
rect 24400 19994 24452 20000
rect 24504 19553 24532 21791
rect 24676 21548 24728 21554
rect 24676 21490 24728 21496
rect 24688 21078 24716 21490
rect 24676 21072 24728 21078
rect 24676 21014 24728 21020
rect 24780 21010 24808 21966
rect 24872 21554 24900 22646
rect 24860 21548 24912 21554
rect 24860 21490 24912 21496
rect 24768 21004 24820 21010
rect 24768 20946 24820 20952
rect 24674 20496 24730 20505
rect 24674 20431 24730 20440
rect 24688 20058 24716 20431
rect 24676 20052 24728 20058
rect 24676 19994 24728 20000
rect 25056 19854 25084 22986
rect 25136 22636 25188 22642
rect 25136 22578 25188 22584
rect 25148 21962 25176 22578
rect 25136 21956 25188 21962
rect 25136 21898 25188 21904
rect 25148 20874 25176 21898
rect 25136 20868 25188 20874
rect 25136 20810 25188 20816
rect 25332 20505 25360 26318
rect 26056 25696 26108 25702
rect 26056 25638 26108 25644
rect 26068 24614 26096 25638
rect 27908 25294 27936 27406
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 36832 26586 36860 57462
rect 67652 57458 67680 57559
rect 56324 57452 56376 57458
rect 56324 57394 56376 57400
rect 67640 57452 67692 57458
rect 67640 57394 67692 57400
rect 39304 57384 39356 57390
rect 39304 57326 39356 57332
rect 39212 57248 39264 57254
rect 39212 57190 39264 57196
rect 39224 57050 39252 57190
rect 39212 57044 39264 57050
rect 39212 56986 39264 56992
rect 39316 45554 39344 57326
rect 56336 57254 56364 57394
rect 56324 57248 56376 57254
rect 56324 57190 56376 57196
rect 50294 56604 50602 56613
rect 50294 56602 50300 56604
rect 50356 56602 50380 56604
rect 50436 56602 50460 56604
rect 50516 56602 50540 56604
rect 50596 56602 50602 56604
rect 50356 56550 50358 56602
rect 50538 56550 50540 56602
rect 50294 56548 50300 56550
rect 50356 56548 50380 56550
rect 50436 56548 50460 56550
rect 50516 56548 50540 56550
rect 50596 56548 50602 56550
rect 50294 56539 50602 56548
rect 50294 55516 50602 55525
rect 50294 55514 50300 55516
rect 50356 55514 50380 55516
rect 50436 55514 50460 55516
rect 50516 55514 50540 55516
rect 50596 55514 50602 55516
rect 50356 55462 50358 55514
rect 50538 55462 50540 55514
rect 50294 55460 50300 55462
rect 50356 55460 50380 55462
rect 50436 55460 50460 55462
rect 50516 55460 50540 55462
rect 50596 55460 50602 55462
rect 50294 55451 50602 55460
rect 50294 54428 50602 54437
rect 50294 54426 50300 54428
rect 50356 54426 50380 54428
rect 50436 54426 50460 54428
rect 50516 54426 50540 54428
rect 50596 54426 50602 54428
rect 50356 54374 50358 54426
rect 50538 54374 50540 54426
rect 50294 54372 50300 54374
rect 50356 54372 50380 54374
rect 50436 54372 50460 54374
rect 50516 54372 50540 54374
rect 50596 54372 50602 54374
rect 50294 54363 50602 54372
rect 50294 53340 50602 53349
rect 50294 53338 50300 53340
rect 50356 53338 50380 53340
rect 50436 53338 50460 53340
rect 50516 53338 50540 53340
rect 50596 53338 50602 53340
rect 50356 53286 50358 53338
rect 50538 53286 50540 53338
rect 50294 53284 50300 53286
rect 50356 53284 50380 53286
rect 50436 53284 50460 53286
rect 50516 53284 50540 53286
rect 50596 53284 50602 53286
rect 50294 53275 50602 53284
rect 50294 52252 50602 52261
rect 50294 52250 50300 52252
rect 50356 52250 50380 52252
rect 50436 52250 50460 52252
rect 50516 52250 50540 52252
rect 50596 52250 50602 52252
rect 50356 52198 50358 52250
rect 50538 52198 50540 52250
rect 50294 52196 50300 52198
rect 50356 52196 50380 52198
rect 50436 52196 50460 52198
rect 50516 52196 50540 52198
rect 50596 52196 50602 52198
rect 50294 52187 50602 52196
rect 50294 51164 50602 51173
rect 50294 51162 50300 51164
rect 50356 51162 50380 51164
rect 50436 51162 50460 51164
rect 50516 51162 50540 51164
rect 50596 51162 50602 51164
rect 50356 51110 50358 51162
rect 50538 51110 50540 51162
rect 50294 51108 50300 51110
rect 50356 51108 50380 51110
rect 50436 51108 50460 51110
rect 50516 51108 50540 51110
rect 50596 51108 50602 51110
rect 50294 51099 50602 51108
rect 50294 50076 50602 50085
rect 50294 50074 50300 50076
rect 50356 50074 50380 50076
rect 50436 50074 50460 50076
rect 50516 50074 50540 50076
rect 50596 50074 50602 50076
rect 50356 50022 50358 50074
rect 50538 50022 50540 50074
rect 50294 50020 50300 50022
rect 50356 50020 50380 50022
rect 50436 50020 50460 50022
rect 50516 50020 50540 50022
rect 50596 50020 50602 50022
rect 50294 50011 50602 50020
rect 50294 48988 50602 48997
rect 50294 48986 50300 48988
rect 50356 48986 50380 48988
rect 50436 48986 50460 48988
rect 50516 48986 50540 48988
rect 50596 48986 50602 48988
rect 50356 48934 50358 48986
rect 50538 48934 50540 48986
rect 50294 48932 50300 48934
rect 50356 48932 50380 48934
rect 50436 48932 50460 48934
rect 50516 48932 50540 48934
rect 50596 48932 50602 48934
rect 50294 48923 50602 48932
rect 50294 47900 50602 47909
rect 50294 47898 50300 47900
rect 50356 47898 50380 47900
rect 50436 47898 50460 47900
rect 50516 47898 50540 47900
rect 50596 47898 50602 47900
rect 50356 47846 50358 47898
rect 50538 47846 50540 47898
rect 50294 47844 50300 47846
rect 50356 47844 50380 47846
rect 50436 47844 50460 47846
rect 50516 47844 50540 47846
rect 50596 47844 50602 47846
rect 50294 47835 50602 47844
rect 50294 46812 50602 46821
rect 50294 46810 50300 46812
rect 50356 46810 50380 46812
rect 50436 46810 50460 46812
rect 50516 46810 50540 46812
rect 50596 46810 50602 46812
rect 50356 46758 50358 46810
rect 50538 46758 50540 46810
rect 50294 46756 50300 46758
rect 50356 46756 50380 46758
rect 50436 46756 50460 46758
rect 50516 46756 50540 46758
rect 50596 46756 50602 46758
rect 50294 46747 50602 46756
rect 50294 45724 50602 45733
rect 50294 45722 50300 45724
rect 50356 45722 50380 45724
rect 50436 45722 50460 45724
rect 50516 45722 50540 45724
rect 50596 45722 50602 45724
rect 50356 45670 50358 45722
rect 50538 45670 50540 45722
rect 50294 45668 50300 45670
rect 50356 45668 50380 45670
rect 50436 45668 50460 45670
rect 50516 45668 50540 45670
rect 50596 45668 50602 45670
rect 50294 45659 50602 45668
rect 39224 45526 39344 45554
rect 39224 35894 39252 45526
rect 50294 44636 50602 44645
rect 50294 44634 50300 44636
rect 50356 44634 50380 44636
rect 50436 44634 50460 44636
rect 50516 44634 50540 44636
rect 50596 44634 50602 44636
rect 50356 44582 50358 44634
rect 50538 44582 50540 44634
rect 50294 44580 50300 44582
rect 50356 44580 50380 44582
rect 50436 44580 50460 44582
rect 50516 44580 50540 44582
rect 50596 44580 50602 44582
rect 50294 44571 50602 44580
rect 50294 43548 50602 43557
rect 50294 43546 50300 43548
rect 50356 43546 50380 43548
rect 50436 43546 50460 43548
rect 50516 43546 50540 43548
rect 50596 43546 50602 43548
rect 50356 43494 50358 43546
rect 50538 43494 50540 43546
rect 50294 43492 50300 43494
rect 50356 43492 50380 43494
rect 50436 43492 50460 43494
rect 50516 43492 50540 43494
rect 50596 43492 50602 43494
rect 50294 43483 50602 43492
rect 50294 42460 50602 42469
rect 50294 42458 50300 42460
rect 50356 42458 50380 42460
rect 50436 42458 50460 42460
rect 50516 42458 50540 42460
rect 50596 42458 50602 42460
rect 50356 42406 50358 42458
rect 50538 42406 50540 42458
rect 50294 42404 50300 42406
rect 50356 42404 50380 42406
rect 50436 42404 50460 42406
rect 50516 42404 50540 42406
rect 50596 42404 50602 42406
rect 50294 42395 50602 42404
rect 50294 41372 50602 41381
rect 50294 41370 50300 41372
rect 50356 41370 50380 41372
rect 50436 41370 50460 41372
rect 50516 41370 50540 41372
rect 50596 41370 50602 41372
rect 50356 41318 50358 41370
rect 50538 41318 50540 41370
rect 50294 41316 50300 41318
rect 50356 41316 50380 41318
rect 50436 41316 50460 41318
rect 50516 41316 50540 41318
rect 50596 41316 50602 41318
rect 50294 41307 50602 41316
rect 50294 40284 50602 40293
rect 50294 40282 50300 40284
rect 50356 40282 50380 40284
rect 50436 40282 50460 40284
rect 50516 40282 50540 40284
rect 50596 40282 50602 40284
rect 50356 40230 50358 40282
rect 50538 40230 50540 40282
rect 50294 40228 50300 40230
rect 50356 40228 50380 40230
rect 50436 40228 50460 40230
rect 50516 40228 50540 40230
rect 50596 40228 50602 40230
rect 50294 40219 50602 40228
rect 50294 39196 50602 39205
rect 50294 39194 50300 39196
rect 50356 39194 50380 39196
rect 50436 39194 50460 39196
rect 50516 39194 50540 39196
rect 50596 39194 50602 39196
rect 50356 39142 50358 39194
rect 50538 39142 50540 39194
rect 50294 39140 50300 39142
rect 50356 39140 50380 39142
rect 50436 39140 50460 39142
rect 50516 39140 50540 39142
rect 50596 39140 50602 39142
rect 50294 39131 50602 39140
rect 50294 38108 50602 38117
rect 50294 38106 50300 38108
rect 50356 38106 50380 38108
rect 50436 38106 50460 38108
rect 50516 38106 50540 38108
rect 50596 38106 50602 38108
rect 50356 38054 50358 38106
rect 50538 38054 50540 38106
rect 50294 38052 50300 38054
rect 50356 38052 50380 38054
rect 50436 38052 50460 38054
rect 50516 38052 50540 38054
rect 50596 38052 50602 38054
rect 50294 38043 50602 38052
rect 50294 37020 50602 37029
rect 50294 37018 50300 37020
rect 50356 37018 50380 37020
rect 50436 37018 50460 37020
rect 50516 37018 50540 37020
rect 50596 37018 50602 37020
rect 50356 36966 50358 37018
rect 50538 36966 50540 37018
rect 50294 36964 50300 36966
rect 50356 36964 50380 36966
rect 50436 36964 50460 36966
rect 50516 36964 50540 36966
rect 50596 36964 50602 36966
rect 50294 36955 50602 36964
rect 50294 35932 50602 35941
rect 50294 35930 50300 35932
rect 50356 35930 50380 35932
rect 50436 35930 50460 35932
rect 50516 35930 50540 35932
rect 50596 35930 50602 35932
rect 39224 35866 39344 35894
rect 50356 35878 50358 35930
rect 50538 35878 50540 35930
rect 50294 35876 50300 35878
rect 50356 35876 50380 35878
rect 50436 35876 50460 35878
rect 50516 35876 50540 35878
rect 50596 35876 50602 35878
rect 50294 35867 50602 35876
rect 39316 31754 39344 35866
rect 50294 34844 50602 34853
rect 50294 34842 50300 34844
rect 50356 34842 50380 34844
rect 50436 34842 50460 34844
rect 50516 34842 50540 34844
rect 50596 34842 50602 34844
rect 50356 34790 50358 34842
rect 50538 34790 50540 34842
rect 50294 34788 50300 34790
rect 50356 34788 50380 34790
rect 50436 34788 50460 34790
rect 50516 34788 50540 34790
rect 50596 34788 50602 34790
rect 50294 34779 50602 34788
rect 50294 33756 50602 33765
rect 50294 33754 50300 33756
rect 50356 33754 50380 33756
rect 50436 33754 50460 33756
rect 50516 33754 50540 33756
rect 50596 33754 50602 33756
rect 50356 33702 50358 33754
rect 50538 33702 50540 33754
rect 50294 33700 50300 33702
rect 50356 33700 50380 33702
rect 50436 33700 50460 33702
rect 50516 33700 50540 33702
rect 50596 33700 50602 33702
rect 50294 33691 50602 33700
rect 50294 32668 50602 32677
rect 50294 32666 50300 32668
rect 50356 32666 50380 32668
rect 50436 32666 50460 32668
rect 50516 32666 50540 32668
rect 50596 32666 50602 32668
rect 50356 32614 50358 32666
rect 50538 32614 50540 32666
rect 50294 32612 50300 32614
rect 50356 32612 50380 32614
rect 50436 32612 50460 32614
rect 50516 32612 50540 32614
rect 50596 32612 50602 32614
rect 50294 32603 50602 32612
rect 39316 31726 39436 31754
rect 36820 26580 36872 26586
rect 36820 26522 36872 26528
rect 32220 26376 32272 26382
rect 32220 26318 32272 26324
rect 32404 26376 32456 26382
rect 32404 26318 32456 26324
rect 35164 26376 35216 26382
rect 35164 26318 35216 26324
rect 35808 26376 35860 26382
rect 35808 26318 35860 26324
rect 36084 26376 36136 26382
rect 36084 26318 36136 26324
rect 32232 25702 32260 26318
rect 32220 25696 32272 25702
rect 32220 25638 32272 25644
rect 32232 25362 32260 25638
rect 32220 25356 32272 25362
rect 32220 25298 32272 25304
rect 27896 25288 27948 25294
rect 27896 25230 27948 25236
rect 28356 25288 28408 25294
rect 28356 25230 28408 25236
rect 30656 25288 30708 25294
rect 30656 25230 30708 25236
rect 26240 25220 26292 25226
rect 26240 25162 26292 25168
rect 26252 24750 26280 25162
rect 28368 24750 28396 25230
rect 28448 24812 28500 24818
rect 28448 24754 28500 24760
rect 26240 24744 26292 24750
rect 26240 24686 26292 24692
rect 28356 24744 28408 24750
rect 28356 24686 28408 24692
rect 26056 24608 26108 24614
rect 26056 24550 26108 24556
rect 25964 24064 26016 24070
rect 25964 24006 26016 24012
rect 25976 23662 26004 24006
rect 25964 23656 26016 23662
rect 25964 23598 26016 23604
rect 25778 22808 25834 22817
rect 25778 22743 25834 22752
rect 25792 22642 25820 22743
rect 25780 22636 25832 22642
rect 25780 22578 25832 22584
rect 25872 22636 25924 22642
rect 25872 22578 25924 22584
rect 25884 22030 25912 22578
rect 25976 22030 26004 23598
rect 26068 22710 26096 24550
rect 28368 24206 28396 24686
rect 28356 24200 28408 24206
rect 28356 24142 28408 24148
rect 27068 24132 27120 24138
rect 27068 24074 27120 24080
rect 27080 23322 27108 24074
rect 27804 24064 27856 24070
rect 27804 24006 27856 24012
rect 27068 23316 27120 23322
rect 27068 23258 27120 23264
rect 26332 23248 26384 23254
rect 26332 23190 26384 23196
rect 26056 22704 26108 22710
rect 26056 22646 26108 22652
rect 26344 22642 26372 23190
rect 27252 23112 27304 23118
rect 27252 23054 27304 23060
rect 27436 23112 27488 23118
rect 27620 23112 27672 23118
rect 27436 23054 27488 23060
rect 27618 23080 27620 23089
rect 27672 23080 27674 23089
rect 27160 22976 27212 22982
rect 27160 22918 27212 22924
rect 27172 22710 27200 22918
rect 27160 22704 27212 22710
rect 27160 22646 27212 22652
rect 26148 22636 26200 22642
rect 26148 22578 26200 22584
rect 26332 22636 26384 22642
rect 26332 22578 26384 22584
rect 26976 22636 27028 22642
rect 26976 22578 27028 22584
rect 25872 22024 25924 22030
rect 25872 21966 25924 21972
rect 25964 22024 26016 22030
rect 25964 21966 26016 21972
rect 26160 21962 26188 22578
rect 26988 22166 27016 22578
rect 26976 22160 27028 22166
rect 26976 22102 27028 22108
rect 26148 21956 26200 21962
rect 26148 21898 26200 21904
rect 25596 21616 25648 21622
rect 25596 21558 25648 21564
rect 25608 20874 25636 21558
rect 26240 20936 26292 20942
rect 26240 20878 26292 20884
rect 25412 20868 25464 20874
rect 25412 20810 25464 20816
rect 25596 20868 25648 20874
rect 25596 20810 25648 20816
rect 26148 20868 26200 20874
rect 26148 20810 26200 20816
rect 25424 20602 25452 20810
rect 25688 20800 25740 20806
rect 25688 20742 25740 20748
rect 25412 20596 25464 20602
rect 25412 20538 25464 20544
rect 25318 20496 25374 20505
rect 25318 20431 25374 20440
rect 25136 20392 25188 20398
rect 25136 20334 25188 20340
rect 25320 20392 25372 20398
rect 25320 20334 25372 20340
rect 24584 19848 24636 19854
rect 24584 19790 24636 19796
rect 25044 19848 25096 19854
rect 25044 19790 25096 19796
rect 24490 19544 24546 19553
rect 24490 19479 24546 19488
rect 24596 19378 24624 19790
rect 24952 19780 25004 19786
rect 24952 19722 25004 19728
rect 24584 19372 24636 19378
rect 24584 19314 24636 19320
rect 24964 18902 24992 19722
rect 24952 18896 25004 18902
rect 24952 18838 25004 18844
rect 25056 18290 25084 19790
rect 25148 18698 25176 20334
rect 25228 20256 25280 20262
rect 25228 20198 25280 20204
rect 25240 19310 25268 20198
rect 25332 19922 25360 20334
rect 25320 19916 25372 19922
rect 25320 19858 25372 19864
rect 25332 19514 25360 19858
rect 25320 19508 25372 19514
rect 25320 19450 25372 19456
rect 25228 19304 25280 19310
rect 25228 19246 25280 19252
rect 25136 18692 25188 18698
rect 25136 18634 25188 18640
rect 25136 18352 25188 18358
rect 25136 18294 25188 18300
rect 24860 18284 24912 18290
rect 24860 18226 24912 18232
rect 25044 18284 25096 18290
rect 25044 18226 25096 18232
rect 24584 18148 24636 18154
rect 24584 18090 24636 18096
rect 24596 17610 24624 18090
rect 24872 17882 24900 18226
rect 24860 17876 24912 17882
rect 24860 17818 24912 17824
rect 24860 17672 24912 17678
rect 24860 17614 24912 17620
rect 24584 17604 24636 17610
rect 24584 17546 24636 17552
rect 24872 16590 24900 17614
rect 25044 16992 25096 16998
rect 25044 16934 25096 16940
rect 25056 16590 25084 16934
rect 24860 16584 24912 16590
rect 25044 16584 25096 16590
rect 24860 16526 24912 16532
rect 25042 16552 25044 16561
rect 25096 16552 25098 16561
rect 25042 16487 25098 16496
rect 24124 16244 24176 16250
rect 24124 16186 24176 16192
rect 23756 16108 23808 16114
rect 23756 16050 23808 16056
rect 24584 16108 24636 16114
rect 24584 16050 24636 16056
rect 24400 15496 24452 15502
rect 24400 15438 24452 15444
rect 24412 15065 24440 15438
rect 24398 15056 24454 15065
rect 24398 14991 24454 15000
rect 24216 14952 24268 14958
rect 24214 14920 24216 14929
rect 24268 14920 24270 14929
rect 24214 14855 24270 14864
rect 24412 14618 24440 14991
rect 24400 14612 24452 14618
rect 24400 14554 24452 14560
rect 24032 13524 24084 13530
rect 24032 13466 24084 13472
rect 23756 13320 23808 13326
rect 23754 13288 23756 13297
rect 23808 13288 23810 13297
rect 23664 13252 23716 13258
rect 23754 13223 23810 13232
rect 23664 13194 23716 13200
rect 24044 12850 24072 13466
rect 24308 13456 24360 13462
rect 24308 13398 24360 13404
rect 23756 12844 23808 12850
rect 23756 12786 23808 12792
rect 24032 12844 24084 12850
rect 24032 12786 24084 12792
rect 23768 12434 23796 12786
rect 23940 12708 23992 12714
rect 23940 12650 23992 12656
rect 23952 12434 23980 12650
rect 23676 12406 23796 12434
rect 23860 12406 23980 12434
rect 23572 8492 23624 8498
rect 23572 8434 23624 8440
rect 23584 7750 23612 8434
rect 23572 7744 23624 7750
rect 23572 7686 23624 7692
rect 23296 7336 23348 7342
rect 23296 7278 23348 7284
rect 23676 6662 23704 12406
rect 23756 11620 23808 11626
rect 23756 11562 23808 11568
rect 23768 11354 23796 11562
rect 23756 11348 23808 11354
rect 23756 11290 23808 11296
rect 23860 11150 23888 12406
rect 23940 11824 23992 11830
rect 23940 11766 23992 11772
rect 23952 11626 23980 11766
rect 23940 11620 23992 11626
rect 23940 11562 23992 11568
rect 23952 11218 23980 11562
rect 23940 11212 23992 11218
rect 23940 11154 23992 11160
rect 23848 11144 23900 11150
rect 23848 11086 23900 11092
rect 23860 10198 23888 11086
rect 23848 10192 23900 10198
rect 23848 10134 23900 10140
rect 24044 9586 24072 12786
rect 24124 12776 24176 12782
rect 24124 12718 24176 12724
rect 24136 11830 24164 12718
rect 24124 11824 24176 11830
rect 24124 11766 24176 11772
rect 24122 11656 24178 11665
rect 24122 11591 24178 11600
rect 24032 9580 24084 9586
rect 24032 9522 24084 9528
rect 23848 8832 23900 8838
rect 23848 8774 23900 8780
rect 23860 8430 23888 8774
rect 23848 8424 23900 8430
rect 23848 8366 23900 8372
rect 23860 7818 23888 8366
rect 23848 7812 23900 7818
rect 23848 7754 23900 7760
rect 24136 7750 24164 11591
rect 24216 10464 24268 10470
rect 24216 10406 24268 10412
rect 24228 9518 24256 10406
rect 24216 9512 24268 9518
rect 24216 9454 24268 9460
rect 24228 9042 24256 9454
rect 24216 9036 24268 9042
rect 24216 8978 24268 8984
rect 24320 8922 24348 13398
rect 24492 12640 24544 12646
rect 24492 12582 24544 12588
rect 24400 12096 24452 12102
rect 24400 12038 24452 12044
rect 24228 8894 24348 8922
rect 24124 7744 24176 7750
rect 24124 7686 24176 7692
rect 23756 7200 23808 7206
rect 23756 7142 23808 7148
rect 23664 6656 23716 6662
rect 23664 6598 23716 6604
rect 23480 6452 23532 6458
rect 23480 6394 23532 6400
rect 23492 6322 23520 6394
rect 23676 6390 23704 6598
rect 23664 6384 23716 6390
rect 23664 6326 23716 6332
rect 23480 6316 23532 6322
rect 23480 6258 23532 6264
rect 23492 4214 23520 6258
rect 23480 4208 23532 4214
rect 23480 4150 23532 4156
rect 23480 3528 23532 3534
rect 23480 3470 23532 3476
rect 23112 2644 23164 2650
rect 23112 2586 23164 2592
rect 23204 2576 23256 2582
rect 23204 2518 23256 2524
rect 23216 800 23244 2518
rect 23492 800 23520 3470
rect 23768 3097 23796 7142
rect 24228 6390 24256 8894
rect 24308 8832 24360 8838
rect 24308 8774 24360 8780
rect 24320 8498 24348 8774
rect 24412 8566 24440 12038
rect 24504 9654 24532 12582
rect 24596 12374 24624 16050
rect 24676 15972 24728 15978
rect 24676 15914 24728 15920
rect 24688 15337 24716 15914
rect 24674 15328 24730 15337
rect 24674 15263 24730 15272
rect 24768 15088 24820 15094
rect 24768 15030 24820 15036
rect 24780 13297 24808 15030
rect 24952 15020 25004 15026
rect 24952 14962 25004 14968
rect 25044 15020 25096 15026
rect 25044 14962 25096 14968
rect 24860 14884 24912 14890
rect 24860 14826 24912 14832
rect 24766 13288 24822 13297
rect 24766 13223 24822 13232
rect 24676 13184 24728 13190
rect 24676 13126 24728 13132
rect 24688 12889 24716 13126
rect 24674 12880 24730 12889
rect 24674 12815 24730 12824
rect 24676 12436 24728 12442
rect 24676 12378 24728 12384
rect 24584 12368 24636 12374
rect 24584 12310 24636 12316
rect 24584 12232 24636 12238
rect 24584 12174 24636 12180
rect 24596 11762 24624 12174
rect 24584 11756 24636 11762
rect 24584 11698 24636 11704
rect 24688 11354 24716 12378
rect 24768 12368 24820 12374
rect 24768 12310 24820 12316
rect 24780 11937 24808 12310
rect 24766 11928 24822 11937
rect 24766 11863 24822 11872
rect 24768 11824 24820 11830
rect 24768 11766 24820 11772
rect 24676 11348 24728 11354
rect 24676 11290 24728 11296
rect 24780 11150 24808 11766
rect 24768 11144 24820 11150
rect 24768 11086 24820 11092
rect 24492 9648 24544 9654
rect 24492 9590 24544 9596
rect 24584 9376 24636 9382
rect 24584 9318 24636 9324
rect 24596 8888 24624 9318
rect 24676 8900 24728 8906
rect 24596 8860 24676 8888
rect 24492 8832 24544 8838
rect 24492 8774 24544 8780
rect 24504 8634 24532 8774
rect 24492 8628 24544 8634
rect 24492 8570 24544 8576
rect 24400 8560 24452 8566
rect 24400 8502 24452 8508
rect 24308 8492 24360 8498
rect 24308 8434 24360 8440
rect 24308 7472 24360 7478
rect 24308 7414 24360 7420
rect 24320 6798 24348 7414
rect 24412 7410 24440 8502
rect 24492 7744 24544 7750
rect 24492 7686 24544 7692
rect 24400 7404 24452 7410
rect 24400 7346 24452 7352
rect 24412 6866 24440 7346
rect 24400 6860 24452 6866
rect 24400 6802 24452 6808
rect 24308 6792 24360 6798
rect 24308 6734 24360 6740
rect 24216 6384 24268 6390
rect 24216 6326 24268 6332
rect 24228 5370 24256 6326
rect 24216 5364 24268 5370
rect 24216 5306 24268 5312
rect 23848 4820 23900 4826
rect 23848 4762 23900 4768
rect 23754 3088 23810 3097
rect 23754 3023 23810 3032
rect 23860 2825 23888 4762
rect 24228 4282 24256 5306
rect 24400 4480 24452 4486
rect 24400 4422 24452 4428
rect 24216 4276 24268 4282
rect 24216 4218 24268 4224
rect 24412 4214 24440 4422
rect 24400 4208 24452 4214
rect 24400 4150 24452 4156
rect 24504 3777 24532 7686
rect 24596 6390 24624 8860
rect 24676 8842 24728 8848
rect 24676 7812 24728 7818
rect 24676 7754 24728 7760
rect 24688 7342 24716 7754
rect 24676 7336 24728 7342
rect 24676 7278 24728 7284
rect 24584 6384 24636 6390
rect 24584 6326 24636 6332
rect 24596 5710 24624 6326
rect 24584 5704 24636 5710
rect 24584 5646 24636 5652
rect 24584 4820 24636 4826
rect 24584 4762 24636 4768
rect 24596 4622 24624 4762
rect 24584 4616 24636 4622
rect 24584 4558 24636 4564
rect 24688 4486 24716 7278
rect 24872 7206 24900 14826
rect 24964 14074 24992 14962
rect 24952 14068 25004 14074
rect 24952 14010 25004 14016
rect 25056 13258 25084 14962
rect 25148 14385 25176 18294
rect 25240 18222 25268 19246
rect 25424 18834 25452 20538
rect 25700 19854 25728 20742
rect 25872 20256 25924 20262
rect 25872 20198 25924 20204
rect 25688 19848 25740 19854
rect 25688 19790 25740 19796
rect 25884 19718 25912 20198
rect 26160 20058 26188 20810
rect 26252 20602 26280 20878
rect 26240 20596 26292 20602
rect 26240 20538 26292 20544
rect 26988 20534 27016 22102
rect 26976 20528 27028 20534
rect 26976 20470 27028 20476
rect 26608 20460 26660 20466
rect 26608 20402 26660 20408
rect 26148 20052 26200 20058
rect 26148 19994 26200 20000
rect 26620 19854 26648 20402
rect 26988 20058 27016 20470
rect 26976 20052 27028 20058
rect 26976 19994 27028 20000
rect 25964 19848 26016 19854
rect 25964 19790 26016 19796
rect 26608 19848 26660 19854
rect 26608 19790 26660 19796
rect 25872 19712 25924 19718
rect 25872 19654 25924 19660
rect 25596 19440 25648 19446
rect 25596 19382 25648 19388
rect 25504 18964 25556 18970
rect 25504 18906 25556 18912
rect 25516 18834 25544 18906
rect 25412 18828 25464 18834
rect 25412 18770 25464 18776
rect 25504 18828 25556 18834
rect 25504 18770 25556 18776
rect 25424 18358 25452 18770
rect 25608 18442 25636 19382
rect 25688 19372 25740 19378
rect 25688 19314 25740 19320
rect 25700 18970 25728 19314
rect 25688 18964 25740 18970
rect 25688 18906 25740 18912
rect 25976 18834 26004 19790
rect 26424 19168 26476 19174
rect 26424 19110 26476 19116
rect 26056 18896 26108 18902
rect 26056 18838 26108 18844
rect 25964 18828 26016 18834
rect 25964 18770 26016 18776
rect 25516 18414 25636 18442
rect 25412 18352 25464 18358
rect 25412 18294 25464 18300
rect 25228 18216 25280 18222
rect 25228 18158 25280 18164
rect 25240 17746 25268 18158
rect 25228 17740 25280 17746
rect 25228 17682 25280 17688
rect 25240 17338 25268 17682
rect 25320 17672 25372 17678
rect 25424 17660 25452 18294
rect 25516 17678 25544 18414
rect 26068 18290 26096 18838
rect 26436 18766 26464 19110
rect 26424 18760 26476 18766
rect 26424 18702 26476 18708
rect 25688 18284 25740 18290
rect 25608 18244 25688 18272
rect 25372 17632 25452 17660
rect 25504 17672 25556 17678
rect 25320 17614 25372 17620
rect 25504 17614 25556 17620
rect 25516 17338 25544 17614
rect 25228 17332 25280 17338
rect 25228 17274 25280 17280
rect 25320 17332 25372 17338
rect 25320 17274 25372 17280
rect 25504 17332 25556 17338
rect 25504 17274 25556 17280
rect 25332 16794 25360 17274
rect 25608 17082 25636 18244
rect 25688 18226 25740 18232
rect 26056 18284 26108 18290
rect 26056 18226 26108 18232
rect 26056 18080 26108 18086
rect 26056 18022 26108 18028
rect 25688 17808 25740 17814
rect 25688 17750 25740 17756
rect 25516 17054 25636 17082
rect 25320 16788 25372 16794
rect 25320 16730 25372 16736
rect 25320 16584 25372 16590
rect 25320 16526 25372 16532
rect 25228 16516 25280 16522
rect 25228 16458 25280 16464
rect 25240 15502 25268 16458
rect 25228 15496 25280 15502
rect 25228 15438 25280 15444
rect 25240 14890 25268 15438
rect 25332 15434 25360 16526
rect 25320 15428 25372 15434
rect 25320 15370 25372 15376
rect 25228 14884 25280 14890
rect 25228 14826 25280 14832
rect 25332 14770 25360 15370
rect 25240 14742 25360 14770
rect 25412 14816 25464 14822
rect 25412 14758 25464 14764
rect 25134 14376 25190 14385
rect 25134 14311 25190 14320
rect 25148 13938 25176 14311
rect 25136 13932 25188 13938
rect 25136 13874 25188 13880
rect 25136 13388 25188 13394
rect 25136 13330 25188 13336
rect 25044 13252 25096 13258
rect 25044 13194 25096 13200
rect 25056 11150 25084 13194
rect 25148 12442 25176 13330
rect 25136 12436 25188 12442
rect 25136 12378 25188 12384
rect 25136 12232 25188 12238
rect 25136 12174 25188 12180
rect 25148 12073 25176 12174
rect 25134 12064 25190 12073
rect 25134 11999 25190 12008
rect 25136 11824 25188 11830
rect 25134 11792 25136 11801
rect 25188 11792 25190 11801
rect 25134 11727 25190 11736
rect 24952 11144 25004 11150
rect 24952 11086 25004 11092
rect 25044 11144 25096 11150
rect 25044 11086 25096 11092
rect 24860 7200 24912 7206
rect 24860 7142 24912 7148
rect 24964 6322 24992 11086
rect 25136 11076 25188 11082
rect 25136 11018 25188 11024
rect 25148 9926 25176 11018
rect 25136 9920 25188 9926
rect 25136 9862 25188 9868
rect 25240 8650 25268 14742
rect 25320 14408 25372 14414
rect 25320 14350 25372 14356
rect 25332 14074 25360 14350
rect 25320 14068 25372 14074
rect 25320 14010 25372 14016
rect 25424 13938 25452 14758
rect 25412 13932 25464 13938
rect 25412 13874 25464 13880
rect 25410 13016 25466 13025
rect 25410 12951 25412 12960
rect 25464 12951 25466 12960
rect 25412 12922 25464 12928
rect 25318 12472 25374 12481
rect 25318 12407 25374 12416
rect 25332 10674 25360 12407
rect 25412 12368 25464 12374
rect 25410 12336 25412 12345
rect 25464 12336 25466 12345
rect 25410 12271 25466 12280
rect 25412 12164 25464 12170
rect 25412 12106 25464 12112
rect 25424 11830 25452 12106
rect 25516 11898 25544 17054
rect 25700 16114 25728 17750
rect 26068 17610 26096 18022
rect 26332 17740 26384 17746
rect 26332 17682 26384 17688
rect 26056 17604 26108 17610
rect 26056 17546 26108 17552
rect 26240 17536 26292 17542
rect 26240 17478 26292 17484
rect 25872 16448 25924 16454
rect 25872 16390 25924 16396
rect 25884 16153 25912 16390
rect 25870 16144 25926 16153
rect 25688 16108 25740 16114
rect 25870 16079 25926 16088
rect 25688 16050 25740 16056
rect 25962 16008 26018 16017
rect 25962 15943 26018 15952
rect 25976 15638 26004 15943
rect 25964 15632 26016 15638
rect 25964 15574 26016 15580
rect 25688 15360 25740 15366
rect 25688 15302 25740 15308
rect 25700 15026 25728 15302
rect 25688 15020 25740 15026
rect 25688 14962 25740 14968
rect 25596 14272 25648 14278
rect 25596 14214 25648 14220
rect 25608 13938 25636 14214
rect 25596 13932 25648 13938
rect 25596 13874 25648 13880
rect 25596 13320 25648 13326
rect 25596 13262 25648 13268
rect 25504 11892 25556 11898
rect 25504 11834 25556 11840
rect 25412 11824 25464 11830
rect 25412 11766 25464 11772
rect 25424 11626 25452 11766
rect 25412 11620 25464 11626
rect 25412 11562 25464 11568
rect 25608 10962 25636 13262
rect 25700 12238 25728 14962
rect 25780 14476 25832 14482
rect 25780 14418 25832 14424
rect 25792 14006 25820 14418
rect 25780 14000 25832 14006
rect 25780 13942 25832 13948
rect 25792 13870 25820 13942
rect 25780 13864 25832 13870
rect 25780 13806 25832 13812
rect 25976 13818 26004 15574
rect 26252 15094 26280 17478
rect 26344 16998 26372 17682
rect 26516 17128 26568 17134
rect 26516 17070 26568 17076
rect 26332 16992 26384 16998
rect 26332 16934 26384 16940
rect 26528 16794 26556 17070
rect 26516 16788 26568 16794
rect 26516 16730 26568 16736
rect 26240 15088 26292 15094
rect 26240 15030 26292 15036
rect 26238 14920 26294 14929
rect 26238 14855 26294 14864
rect 26252 14414 26280 14855
rect 26056 14408 26108 14414
rect 26056 14350 26108 14356
rect 26240 14408 26292 14414
rect 26240 14350 26292 14356
rect 26068 14006 26096 14350
rect 26056 14000 26108 14006
rect 26056 13942 26108 13948
rect 26148 13932 26200 13938
rect 26148 13874 26200 13880
rect 25792 12986 25820 13806
rect 25976 13790 26096 13818
rect 25964 13184 26016 13190
rect 25964 13126 26016 13132
rect 25780 12980 25832 12986
rect 25780 12922 25832 12928
rect 25976 12918 26004 13126
rect 25964 12912 26016 12918
rect 25964 12854 26016 12860
rect 25964 12640 26016 12646
rect 25964 12582 26016 12588
rect 25872 12436 25924 12442
rect 25872 12378 25924 12384
rect 25688 12232 25740 12238
rect 25688 12174 25740 12180
rect 25884 12170 25912 12378
rect 25976 12220 26004 12582
rect 26068 12434 26096 13790
rect 26160 13258 26188 13874
rect 26252 13802 26280 14350
rect 26332 14272 26384 14278
rect 26332 14214 26384 14220
rect 26240 13796 26292 13802
rect 26240 13738 26292 13744
rect 26344 13410 26372 14214
rect 26528 13462 26556 16730
rect 27158 16416 27214 16425
rect 27158 16351 27214 16360
rect 27172 15910 27200 16351
rect 27264 16153 27292 23054
rect 27448 22778 27476 23054
rect 27618 23015 27674 23024
rect 27436 22772 27488 22778
rect 27436 22714 27488 22720
rect 27816 22710 27844 24006
rect 28264 23520 28316 23526
rect 28264 23462 28316 23468
rect 28276 23050 28304 23462
rect 28264 23044 28316 23050
rect 28264 22986 28316 22992
rect 27988 22976 28040 22982
rect 27988 22918 28040 22924
rect 28000 22710 28028 22918
rect 27804 22704 27856 22710
rect 27804 22646 27856 22652
rect 27988 22704 28040 22710
rect 27988 22646 28040 22652
rect 27620 21956 27672 21962
rect 27620 21898 27672 21904
rect 27632 21486 27660 21898
rect 27712 21548 27764 21554
rect 27712 21490 27764 21496
rect 27620 21480 27672 21486
rect 27620 21422 27672 21428
rect 27342 21176 27398 21185
rect 27724 21146 27752 21490
rect 27816 21350 27844 22646
rect 28000 22030 28028 22646
rect 28172 22092 28224 22098
rect 28172 22034 28224 22040
rect 27988 22024 28040 22030
rect 27988 21966 28040 21972
rect 27896 21616 27948 21622
rect 27894 21584 27896 21593
rect 27948 21584 27950 21593
rect 27894 21519 27950 21528
rect 27804 21344 27856 21350
rect 27804 21286 27856 21292
rect 27342 21111 27398 21120
rect 27712 21140 27764 21146
rect 27356 21010 27384 21111
rect 27712 21082 27764 21088
rect 27344 21004 27396 21010
rect 27344 20946 27396 20952
rect 28184 20942 28212 22034
rect 28172 20936 28224 20942
rect 28172 20878 28224 20884
rect 27436 20460 27488 20466
rect 27436 20402 27488 20408
rect 27448 19990 27476 20402
rect 28080 20392 28132 20398
rect 28080 20334 28132 20340
rect 27896 20256 27948 20262
rect 27896 20198 27948 20204
rect 27436 19984 27488 19990
rect 27436 19926 27488 19932
rect 27712 19984 27764 19990
rect 27712 19926 27764 19932
rect 27724 19854 27752 19926
rect 27908 19854 27936 20198
rect 28092 19854 28120 20334
rect 28184 19922 28212 20878
rect 28276 20466 28304 22986
rect 28460 22778 28488 24754
rect 29736 24608 29788 24614
rect 29736 24550 29788 24556
rect 29368 24200 29420 24206
rect 29368 24142 29420 24148
rect 28632 23112 28684 23118
rect 28632 23054 28684 23060
rect 29092 23112 29144 23118
rect 29092 23054 29144 23060
rect 28448 22772 28500 22778
rect 28448 22714 28500 22720
rect 28644 22658 28672 23054
rect 28906 22808 28962 22817
rect 28906 22743 28908 22752
rect 28960 22743 28962 22752
rect 28908 22714 28960 22720
rect 28644 22642 29040 22658
rect 28644 22636 29052 22642
rect 28644 22630 29000 22636
rect 28644 21554 28672 22630
rect 29000 22578 29052 22584
rect 29104 21690 29132 23054
rect 29380 23050 29408 24142
rect 29644 23724 29696 23730
rect 29644 23666 29696 23672
rect 29460 23520 29512 23526
rect 29460 23462 29512 23468
rect 29368 23044 29420 23050
rect 29368 22986 29420 22992
rect 29184 22704 29236 22710
rect 29184 22646 29236 22652
rect 29092 21684 29144 21690
rect 29092 21626 29144 21632
rect 28998 21584 29054 21593
rect 28632 21548 28684 21554
rect 28632 21490 28684 21496
rect 28724 21548 28776 21554
rect 28998 21519 29000 21528
rect 28724 21490 28776 21496
rect 29052 21519 29054 21528
rect 29000 21490 29052 21496
rect 28736 21146 28764 21490
rect 29196 21486 29224 22646
rect 29380 21554 29408 22986
rect 29368 21548 29420 21554
rect 29368 21490 29420 21496
rect 29184 21480 29236 21486
rect 29184 21422 29236 21428
rect 28724 21140 28776 21146
rect 28724 21082 28776 21088
rect 28908 21140 28960 21146
rect 28908 21082 28960 21088
rect 28920 20942 28948 21082
rect 28908 20936 28960 20942
rect 28908 20878 28960 20884
rect 29092 20936 29144 20942
rect 29092 20878 29144 20884
rect 28448 20868 28500 20874
rect 28448 20810 28500 20816
rect 28264 20460 28316 20466
rect 28264 20402 28316 20408
rect 28172 19916 28224 19922
rect 28172 19858 28224 19864
rect 27712 19848 27764 19854
rect 27712 19790 27764 19796
rect 27896 19848 27948 19854
rect 27896 19790 27948 19796
rect 28080 19848 28132 19854
rect 28080 19790 28132 19796
rect 27620 19780 27672 19786
rect 27540 19740 27620 19768
rect 27344 19168 27396 19174
rect 27344 19110 27396 19116
rect 27356 18902 27384 19110
rect 27344 18896 27396 18902
rect 27344 18838 27396 18844
rect 27250 16144 27306 16153
rect 27250 16079 27306 16088
rect 27160 15904 27212 15910
rect 27160 15846 27212 15852
rect 27540 15570 27568 19740
rect 27620 19722 27672 19728
rect 27804 19168 27856 19174
rect 28092 19156 28120 19790
rect 28276 19786 28304 20402
rect 28460 20398 28488 20810
rect 29104 20641 29132 20878
rect 29090 20632 29146 20641
rect 29090 20567 29146 20576
rect 28448 20392 28500 20398
rect 28448 20334 28500 20340
rect 28356 19984 28408 19990
rect 28356 19926 28408 19932
rect 28264 19780 28316 19786
rect 28264 19722 28316 19728
rect 27856 19128 28120 19156
rect 27804 19110 27856 19116
rect 27620 18692 27672 18698
rect 27620 18634 27672 18640
rect 27632 18358 27660 18634
rect 27712 18624 27764 18630
rect 27712 18566 27764 18572
rect 27620 18352 27672 18358
rect 27620 18294 27672 18300
rect 27620 18216 27672 18222
rect 27620 18158 27672 18164
rect 27632 17882 27660 18158
rect 27724 18086 27752 18566
rect 27712 18080 27764 18086
rect 27712 18022 27764 18028
rect 27620 17876 27672 17882
rect 27620 17818 27672 17824
rect 27712 16108 27764 16114
rect 27712 16050 27764 16056
rect 27528 15564 27580 15570
rect 27528 15506 27580 15512
rect 26884 15496 26936 15502
rect 26884 15438 26936 15444
rect 27620 15496 27672 15502
rect 27620 15438 27672 15444
rect 26792 13864 26844 13870
rect 26792 13806 26844 13812
rect 26252 13382 26372 13410
rect 26516 13456 26568 13462
rect 26516 13398 26568 13404
rect 26148 13252 26200 13258
rect 26148 13194 26200 13200
rect 26146 13016 26202 13025
rect 26146 12951 26148 12960
rect 26200 12951 26202 12960
rect 26148 12922 26200 12928
rect 26252 12850 26280 13382
rect 26332 13252 26384 13258
rect 26332 13194 26384 13200
rect 26344 12889 26372 13194
rect 26330 12880 26386 12889
rect 26240 12844 26292 12850
rect 26330 12815 26386 12824
rect 26424 12844 26476 12850
rect 26240 12786 26292 12792
rect 26068 12406 26188 12434
rect 26056 12232 26108 12238
rect 25976 12192 26056 12220
rect 25872 12164 25924 12170
rect 25872 12106 25924 12112
rect 25976 11082 26004 12192
rect 26056 12174 26108 12180
rect 26056 11144 26108 11150
rect 26056 11086 26108 11092
rect 25964 11076 26016 11082
rect 25964 11018 26016 11024
rect 25608 10934 25728 10962
rect 25320 10668 25372 10674
rect 25320 10610 25372 10616
rect 25596 10668 25648 10674
rect 25596 10610 25648 10616
rect 25608 10266 25636 10610
rect 25596 10260 25648 10266
rect 25596 10202 25648 10208
rect 25320 9920 25372 9926
rect 25320 9862 25372 9868
rect 25056 8622 25268 8650
rect 25332 8634 25360 9862
rect 25700 9722 25728 10934
rect 25976 10810 26004 11018
rect 26068 10810 26096 11086
rect 25964 10804 26016 10810
rect 25964 10746 26016 10752
rect 26056 10804 26108 10810
rect 26056 10746 26108 10752
rect 26068 10266 26096 10746
rect 26056 10260 26108 10266
rect 26056 10202 26108 10208
rect 25688 9716 25740 9722
rect 25688 9658 25740 9664
rect 25320 8628 25372 8634
rect 24768 6316 24820 6322
rect 24768 6258 24820 6264
rect 24952 6316 25004 6322
rect 24952 6258 25004 6264
rect 24780 5302 24808 6258
rect 24952 6112 25004 6118
rect 24952 6054 25004 6060
rect 24964 5914 24992 6054
rect 24952 5908 25004 5914
rect 24952 5850 25004 5856
rect 24768 5296 24820 5302
rect 24768 5238 24820 5244
rect 24676 4480 24728 4486
rect 24676 4422 24728 4428
rect 24780 4282 24808 5238
rect 24860 5024 24912 5030
rect 24860 4966 24912 4972
rect 24872 4622 24900 4966
rect 25056 4826 25084 8622
rect 25320 8570 25372 8576
rect 25136 8492 25188 8498
rect 25136 8434 25188 8440
rect 25148 6798 25176 8434
rect 25700 8294 25728 9658
rect 26160 9489 26188 12406
rect 26240 12300 26292 12306
rect 26240 12242 26292 12248
rect 26252 12073 26280 12242
rect 26238 12064 26294 12073
rect 26238 11999 26294 12008
rect 26238 11792 26294 11801
rect 26238 11727 26240 11736
rect 26292 11727 26294 11736
rect 26240 11698 26292 11704
rect 26240 11076 26292 11082
rect 26240 11018 26292 11024
rect 26252 10674 26280 11018
rect 26240 10668 26292 10674
rect 26240 10610 26292 10616
rect 26146 9480 26202 9489
rect 26146 9415 26202 9424
rect 25780 8900 25832 8906
rect 25780 8842 25832 8848
rect 25228 8288 25280 8294
rect 25228 8230 25280 8236
rect 25608 8266 25728 8294
rect 25240 7886 25268 8230
rect 25228 7880 25280 7886
rect 25228 7822 25280 7828
rect 25412 7880 25464 7886
rect 25412 7822 25464 7828
rect 25424 7206 25452 7822
rect 25608 7546 25636 8266
rect 25792 8090 25820 8842
rect 25780 8084 25832 8090
rect 25780 8026 25832 8032
rect 25780 7948 25832 7954
rect 25780 7890 25832 7896
rect 25596 7540 25648 7546
rect 25596 7482 25648 7488
rect 25792 7410 25820 7890
rect 26148 7744 26200 7750
rect 26148 7686 26200 7692
rect 26160 7410 26188 7686
rect 25780 7404 25832 7410
rect 25780 7346 25832 7352
rect 26148 7404 26200 7410
rect 26148 7346 26200 7352
rect 26240 7336 26292 7342
rect 26240 7278 26292 7284
rect 25412 7200 25464 7206
rect 25412 7142 25464 7148
rect 25136 6792 25188 6798
rect 25136 6734 25188 6740
rect 25148 5846 25176 6734
rect 26056 6180 26108 6186
rect 26056 6122 26108 6128
rect 25136 5840 25188 5846
rect 25136 5782 25188 5788
rect 25148 5710 25176 5782
rect 25136 5704 25188 5710
rect 25136 5646 25188 5652
rect 25148 5234 25176 5646
rect 25964 5568 26016 5574
rect 25964 5510 26016 5516
rect 25976 5234 26004 5510
rect 25136 5228 25188 5234
rect 25136 5170 25188 5176
rect 25688 5228 25740 5234
rect 25688 5170 25740 5176
rect 25964 5228 26016 5234
rect 25964 5170 26016 5176
rect 25044 4820 25096 4826
rect 25044 4762 25096 4768
rect 24860 4616 24912 4622
rect 24860 4558 24912 4564
rect 24768 4276 24820 4282
rect 24768 4218 24820 4224
rect 25148 4214 25176 5170
rect 25596 4684 25648 4690
rect 25596 4626 25648 4632
rect 25136 4208 25188 4214
rect 25136 4150 25188 4156
rect 24490 3768 24546 3777
rect 24490 3703 24546 3712
rect 24308 3528 24360 3534
rect 24308 3470 24360 3476
rect 25136 3528 25188 3534
rect 25136 3470 25188 3476
rect 24032 2848 24084 2854
rect 23846 2816 23902 2825
rect 24032 2790 24084 2796
rect 23846 2751 23902 2760
rect 23756 2440 23808 2446
rect 23756 2382 23808 2388
rect 23768 800 23796 2382
rect 24044 800 24072 2790
rect 24320 800 24348 3470
rect 24860 2848 24912 2854
rect 24860 2790 24912 2796
rect 24584 2440 24636 2446
rect 24584 2382 24636 2388
rect 24596 800 24624 2382
rect 24872 800 24900 2790
rect 25148 800 25176 3470
rect 25412 2848 25464 2854
rect 25412 2790 25464 2796
rect 25424 800 25452 2790
rect 25608 2417 25636 4626
rect 25700 4622 25728 5170
rect 25780 5092 25832 5098
rect 25780 5034 25832 5040
rect 25688 4616 25740 4622
rect 25688 4558 25740 4564
rect 25792 4554 25820 5034
rect 25872 4616 25924 4622
rect 25872 4558 25924 4564
rect 25780 4548 25832 4554
rect 25780 4490 25832 4496
rect 25884 4282 25912 4558
rect 25872 4276 25924 4282
rect 25872 4218 25924 4224
rect 26068 4146 26096 6122
rect 26252 5778 26280 7278
rect 26240 5772 26292 5778
rect 26240 5714 26292 5720
rect 26148 5228 26200 5234
rect 26148 5170 26200 5176
rect 26056 4140 26108 4146
rect 26056 4082 26108 4088
rect 26160 3641 26188 5170
rect 26252 4146 26280 5714
rect 26344 5166 26372 12815
rect 26424 12786 26476 12792
rect 26436 11762 26464 12786
rect 26528 12782 26556 13398
rect 26516 12776 26568 12782
rect 26516 12718 26568 12724
rect 26606 12744 26662 12753
rect 26528 12442 26556 12718
rect 26606 12679 26662 12688
rect 26516 12436 26568 12442
rect 26516 12378 26568 12384
rect 26620 12374 26648 12679
rect 26608 12368 26660 12374
rect 26608 12310 26660 12316
rect 26424 11756 26476 11762
rect 26424 11698 26476 11704
rect 26804 11694 26832 13806
rect 26896 12442 26924 15438
rect 27528 14272 27580 14278
rect 27528 14214 27580 14220
rect 27540 13938 27568 14214
rect 27528 13932 27580 13938
rect 27528 13874 27580 13880
rect 27252 13796 27304 13802
rect 27252 13738 27304 13744
rect 27066 13288 27122 13297
rect 27066 13223 27122 13232
rect 27080 12782 27108 13223
rect 27068 12776 27120 12782
rect 27068 12718 27120 12724
rect 26884 12436 26936 12442
rect 26884 12378 26936 12384
rect 26700 11688 26752 11694
rect 26700 11630 26752 11636
rect 26792 11688 26844 11694
rect 26792 11630 26844 11636
rect 26424 10668 26476 10674
rect 26424 10610 26476 10616
rect 26436 10198 26464 10610
rect 26424 10192 26476 10198
rect 26424 10134 26476 10140
rect 26608 7268 26660 7274
rect 26608 7210 26660 7216
rect 26620 6866 26648 7210
rect 26608 6860 26660 6866
rect 26608 6802 26660 6808
rect 26516 5636 26568 5642
rect 26516 5578 26568 5584
rect 26528 5370 26556 5578
rect 26516 5364 26568 5370
rect 26516 5306 26568 5312
rect 26332 5160 26384 5166
rect 26332 5102 26384 5108
rect 26712 4593 26740 11630
rect 26804 10606 26832 11630
rect 26896 11082 26924 12378
rect 27160 11144 27212 11150
rect 27160 11086 27212 11092
rect 26884 11076 26936 11082
rect 26884 11018 26936 11024
rect 26792 10600 26844 10606
rect 26792 10542 26844 10548
rect 26804 9586 26832 10542
rect 27172 10538 27200 11086
rect 27160 10532 27212 10538
rect 27160 10474 27212 10480
rect 27172 10062 27200 10474
rect 27160 10056 27212 10062
rect 27160 9998 27212 10004
rect 26792 9580 26844 9586
rect 26792 9522 26844 9528
rect 27264 8974 27292 13738
rect 27540 13734 27568 13874
rect 27632 13870 27660 15438
rect 27620 13864 27672 13870
rect 27620 13806 27672 13812
rect 27528 13728 27580 13734
rect 27528 13670 27580 13676
rect 27436 13320 27488 13326
rect 27436 13262 27488 13268
rect 27448 13190 27476 13262
rect 27436 13184 27488 13190
rect 27436 13126 27488 13132
rect 27540 12918 27568 13670
rect 27528 12912 27580 12918
rect 27528 12854 27580 12860
rect 27344 12640 27396 12646
rect 27344 12582 27396 12588
rect 27252 8968 27304 8974
rect 27252 8910 27304 8916
rect 26976 7336 27028 7342
rect 26976 7278 27028 7284
rect 26988 7002 27016 7278
rect 27356 7206 27384 12582
rect 27724 11762 27752 16050
rect 27816 15706 27844 19110
rect 28080 18624 28132 18630
rect 28080 18566 28132 18572
rect 27988 16992 28040 16998
rect 27988 16934 28040 16940
rect 28000 16658 28028 16934
rect 27988 16652 28040 16658
rect 27988 16594 28040 16600
rect 28000 16114 28028 16594
rect 27988 16108 28040 16114
rect 27988 16050 28040 16056
rect 27804 15700 27856 15706
rect 27804 15642 27856 15648
rect 27816 15570 27844 15642
rect 27804 15564 27856 15570
rect 27804 15506 27856 15512
rect 28092 14822 28120 18566
rect 28368 17202 28396 19926
rect 28460 19378 28488 20334
rect 28816 19780 28868 19786
rect 28816 19722 28868 19728
rect 28632 19712 28684 19718
rect 28828 19689 28856 19722
rect 28632 19654 28684 19660
rect 28814 19680 28870 19689
rect 28644 19446 28672 19654
rect 28814 19615 28870 19624
rect 28632 19440 28684 19446
rect 28632 19382 28684 19388
rect 28448 19372 28500 19378
rect 28448 19314 28500 19320
rect 28460 18766 28488 19314
rect 28448 18760 28500 18766
rect 28448 18702 28500 18708
rect 28460 18222 28488 18702
rect 29000 18352 29052 18358
rect 29000 18294 29052 18300
rect 28448 18216 28500 18222
rect 28448 18158 28500 18164
rect 28460 17678 28488 18158
rect 28448 17672 28500 17678
rect 28448 17614 28500 17620
rect 28356 17196 28408 17202
rect 28356 17138 28408 17144
rect 28368 16590 28396 17138
rect 28460 16998 28488 17614
rect 29012 17338 29040 18294
rect 28540 17332 28592 17338
rect 28540 17274 28592 17280
rect 28632 17332 28684 17338
rect 28632 17274 28684 17280
rect 29000 17332 29052 17338
rect 29000 17274 29052 17280
rect 28448 16992 28500 16998
rect 28448 16934 28500 16940
rect 28552 16794 28580 17274
rect 28540 16788 28592 16794
rect 28540 16730 28592 16736
rect 28356 16584 28408 16590
rect 28356 16526 28408 16532
rect 28264 16516 28316 16522
rect 28264 16458 28316 16464
rect 28276 15434 28304 16458
rect 28540 16108 28592 16114
rect 28644 16096 28672 17274
rect 28908 17264 28960 17270
rect 28908 17206 28960 17212
rect 28920 16658 28948 17206
rect 28908 16652 28960 16658
rect 28908 16594 28960 16600
rect 28816 16584 28868 16590
rect 28816 16526 28868 16532
rect 28828 16114 28856 16526
rect 29472 16425 29500 23462
rect 29552 22772 29604 22778
rect 29552 22714 29604 22720
rect 29564 22681 29592 22714
rect 29550 22672 29606 22681
rect 29550 22607 29606 22616
rect 29656 22574 29684 23666
rect 29552 22568 29604 22574
rect 29552 22510 29604 22516
rect 29644 22568 29696 22574
rect 29644 22510 29696 22516
rect 29564 22098 29592 22510
rect 29552 22092 29604 22098
rect 29552 22034 29604 22040
rect 29552 20936 29604 20942
rect 29552 20878 29604 20884
rect 29564 20534 29592 20878
rect 29552 20528 29604 20534
rect 29552 20470 29604 20476
rect 29564 19514 29592 20470
rect 29656 19990 29684 22510
rect 29748 21962 29776 24550
rect 30288 24132 30340 24138
rect 30288 24074 30340 24080
rect 29920 24064 29972 24070
rect 29920 24006 29972 24012
rect 29828 23724 29880 23730
rect 29828 23666 29880 23672
rect 29840 23322 29868 23666
rect 29828 23316 29880 23322
rect 29828 23258 29880 23264
rect 29932 23118 29960 24006
rect 30300 23866 30328 24074
rect 30104 23860 30156 23866
rect 30104 23802 30156 23808
rect 30288 23860 30340 23866
rect 30288 23802 30340 23808
rect 29920 23112 29972 23118
rect 29920 23054 29972 23060
rect 29920 22976 29972 22982
rect 29920 22918 29972 22924
rect 30012 22976 30064 22982
rect 30012 22918 30064 22924
rect 29932 22166 29960 22918
rect 30024 22642 30052 22918
rect 30116 22642 30144 23802
rect 30472 23044 30524 23050
rect 30472 22986 30524 22992
rect 30012 22636 30064 22642
rect 30012 22578 30064 22584
rect 30104 22636 30156 22642
rect 30104 22578 30156 22584
rect 30288 22636 30340 22642
rect 30288 22578 30340 22584
rect 29920 22160 29972 22166
rect 29920 22102 29972 22108
rect 29932 22030 29960 22102
rect 30300 22030 30328 22578
rect 29920 22024 29972 22030
rect 29920 21966 29972 21972
rect 30288 22024 30340 22030
rect 30288 21966 30340 21972
rect 29736 21956 29788 21962
rect 29736 21898 29788 21904
rect 30484 21894 30512 22986
rect 30472 21888 30524 21894
rect 30472 21830 30524 21836
rect 30286 21584 30342 21593
rect 30484 21570 30512 21830
rect 30286 21519 30288 21528
rect 30340 21519 30342 21528
rect 30392 21542 30512 21570
rect 30288 21490 30340 21496
rect 30104 21412 30156 21418
rect 30104 21354 30156 21360
rect 29920 21140 29972 21146
rect 29920 21082 29972 21088
rect 29932 20942 29960 21082
rect 30116 20942 30144 21354
rect 29920 20936 29972 20942
rect 29920 20878 29972 20884
rect 30104 20936 30156 20942
rect 30104 20878 30156 20884
rect 30392 20874 30420 21542
rect 30472 21004 30524 21010
rect 30472 20946 30524 20952
rect 30380 20868 30432 20874
rect 30380 20810 30432 20816
rect 29736 20324 29788 20330
rect 29736 20266 29788 20272
rect 29748 19990 29776 20266
rect 30196 20256 30248 20262
rect 30196 20198 30248 20204
rect 29644 19984 29696 19990
rect 29644 19926 29696 19932
rect 29736 19984 29788 19990
rect 29736 19926 29788 19932
rect 30208 19854 30236 20198
rect 30288 19916 30340 19922
rect 30288 19858 30340 19864
rect 29736 19848 29788 19854
rect 29736 19790 29788 19796
rect 30196 19848 30248 19854
rect 30196 19790 30248 19796
rect 29552 19508 29604 19514
rect 29552 19450 29604 19456
rect 29644 18964 29696 18970
rect 29644 18906 29696 18912
rect 29552 18624 29604 18630
rect 29552 18566 29604 18572
rect 29564 18222 29592 18566
rect 29656 18358 29684 18906
rect 29644 18352 29696 18358
rect 29644 18294 29696 18300
rect 29552 18216 29604 18222
rect 29552 18158 29604 18164
rect 29458 16416 29514 16425
rect 29458 16351 29514 16360
rect 28592 16068 28672 16096
rect 28724 16108 28776 16114
rect 28540 16050 28592 16056
rect 28724 16050 28776 16056
rect 28816 16108 28868 16114
rect 28816 16050 28868 16056
rect 28356 15904 28408 15910
rect 28356 15846 28408 15852
rect 28264 15428 28316 15434
rect 28264 15370 28316 15376
rect 28276 15162 28304 15370
rect 28264 15156 28316 15162
rect 28264 15098 28316 15104
rect 28172 15020 28224 15026
rect 28172 14962 28224 14968
rect 28184 14822 28212 14962
rect 28080 14816 28132 14822
rect 28080 14758 28132 14764
rect 28172 14816 28224 14822
rect 28172 14758 28224 14764
rect 28368 14618 28396 15846
rect 28552 15502 28580 16050
rect 28736 15706 28764 16050
rect 29000 15972 29052 15978
rect 29000 15914 29052 15920
rect 28724 15700 28776 15706
rect 28724 15642 28776 15648
rect 28540 15496 28592 15502
rect 28540 15438 28592 15444
rect 29012 15434 29040 15914
rect 29656 15502 29684 18294
rect 29748 15638 29776 19790
rect 30104 19236 30156 19242
rect 30104 19178 30156 19184
rect 30012 18828 30064 18834
rect 30012 18770 30064 18776
rect 29828 18760 29880 18766
rect 29828 18702 29880 18708
rect 29840 18086 29868 18702
rect 29828 18080 29880 18086
rect 29828 18022 29880 18028
rect 29840 16504 29868 18022
rect 29920 17196 29972 17202
rect 29920 17138 29972 17144
rect 29932 16794 29960 17138
rect 29920 16788 29972 16794
rect 29920 16730 29972 16736
rect 30024 16561 30052 18770
rect 30116 16590 30144 19178
rect 30300 18970 30328 19858
rect 30484 19378 30512 20946
rect 30564 20868 30616 20874
rect 30564 20810 30616 20816
rect 30576 20058 30604 20810
rect 30564 20052 30616 20058
rect 30564 19994 30616 20000
rect 30668 19938 30696 25230
rect 32416 24682 32444 26318
rect 33232 26240 33284 26246
rect 33232 26182 33284 26188
rect 34060 26240 34112 26246
rect 34060 26182 34112 26188
rect 33244 25974 33272 26182
rect 34072 25974 34100 26182
rect 35176 26042 35204 26318
rect 35440 26308 35492 26314
rect 35440 26250 35492 26256
rect 35348 26240 35400 26246
rect 35348 26182 35400 26188
rect 34796 26036 34848 26042
rect 34796 25978 34848 25984
rect 35164 26036 35216 26042
rect 35164 25978 35216 25984
rect 33232 25968 33284 25974
rect 33232 25910 33284 25916
rect 34060 25968 34112 25974
rect 34060 25910 34112 25916
rect 33048 25832 33100 25838
rect 33048 25774 33100 25780
rect 32680 24744 32732 24750
rect 32680 24686 32732 24692
rect 32404 24676 32456 24682
rect 32404 24618 32456 24624
rect 32692 24410 32720 24686
rect 32772 24608 32824 24614
rect 32772 24550 32824 24556
rect 32680 24404 32732 24410
rect 32680 24346 32732 24352
rect 32784 24206 32812 24550
rect 31024 24200 31076 24206
rect 31024 24142 31076 24148
rect 32772 24200 32824 24206
rect 32772 24142 32824 24148
rect 30840 21344 30892 21350
rect 30840 21286 30892 21292
rect 30932 21344 30984 21350
rect 30932 21286 30984 21292
rect 30748 21004 30800 21010
rect 30748 20946 30800 20952
rect 30576 19910 30696 19938
rect 30472 19372 30524 19378
rect 30472 19314 30524 19320
rect 30288 18964 30340 18970
rect 30288 18906 30340 18912
rect 30380 18964 30432 18970
rect 30380 18906 30432 18912
rect 30392 18426 30420 18906
rect 30576 18902 30604 19910
rect 30656 19848 30708 19854
rect 30656 19790 30708 19796
rect 30564 18896 30616 18902
rect 30564 18838 30616 18844
rect 30380 18420 30432 18426
rect 30380 18362 30432 18368
rect 30196 18352 30248 18358
rect 30196 18294 30248 18300
rect 30208 18086 30236 18294
rect 30196 18080 30248 18086
rect 30196 18022 30248 18028
rect 30196 16720 30248 16726
rect 30196 16662 30248 16668
rect 30104 16584 30156 16590
rect 30010 16552 30066 16561
rect 29920 16516 29972 16522
rect 29840 16476 29920 16504
rect 30104 16526 30156 16532
rect 30010 16487 30066 16496
rect 29920 16458 29972 16464
rect 29736 15632 29788 15638
rect 29736 15574 29788 15580
rect 29644 15496 29696 15502
rect 29644 15438 29696 15444
rect 29000 15428 29052 15434
rect 29000 15370 29052 15376
rect 28630 15056 28686 15065
rect 28630 14991 28632 15000
rect 28684 14991 28686 15000
rect 28632 14962 28684 14968
rect 28356 14612 28408 14618
rect 28356 14554 28408 14560
rect 27804 14340 27856 14346
rect 27804 14282 27856 14288
rect 27816 13938 27844 14282
rect 27804 13932 27856 13938
rect 27804 13874 27856 13880
rect 27816 12434 27844 13874
rect 28172 13864 28224 13870
rect 28172 13806 28224 13812
rect 28540 13864 28592 13870
rect 28540 13806 28592 13812
rect 27988 13184 28040 13190
rect 27988 13126 28040 13132
rect 28000 12850 28028 13126
rect 27988 12844 28040 12850
rect 27988 12786 28040 12792
rect 27816 12406 27936 12434
rect 27436 11756 27488 11762
rect 27436 11698 27488 11704
rect 27712 11756 27764 11762
rect 27712 11698 27764 11704
rect 27448 10810 27476 11698
rect 27712 11552 27764 11558
rect 27712 11494 27764 11500
rect 27804 11552 27856 11558
rect 27804 11494 27856 11500
rect 27528 11076 27580 11082
rect 27528 11018 27580 11024
rect 27436 10804 27488 10810
rect 27436 10746 27488 10752
rect 27434 10160 27490 10169
rect 27434 10095 27436 10104
rect 27488 10095 27490 10104
rect 27436 10066 27488 10072
rect 27448 9722 27476 10066
rect 27436 9716 27488 9722
rect 27436 9658 27488 9664
rect 27540 8566 27568 11018
rect 27724 10742 27752 11494
rect 27712 10736 27764 10742
rect 27712 10678 27764 10684
rect 27712 9172 27764 9178
rect 27712 9114 27764 9120
rect 27528 8560 27580 8566
rect 27528 8502 27580 8508
rect 27724 8498 27752 9114
rect 27816 8906 27844 11494
rect 27804 8900 27856 8906
rect 27804 8842 27856 8848
rect 27712 8492 27764 8498
rect 27712 8434 27764 8440
rect 27804 8356 27856 8362
rect 27804 8298 27856 8304
rect 27344 7200 27396 7206
rect 27344 7142 27396 7148
rect 26976 6996 27028 7002
rect 26976 6938 27028 6944
rect 27712 6452 27764 6458
rect 27712 6394 27764 6400
rect 27620 6112 27672 6118
rect 27620 6054 27672 6060
rect 27632 5846 27660 6054
rect 27620 5840 27672 5846
rect 27620 5782 27672 5788
rect 26698 4584 26754 4593
rect 26698 4519 26754 4528
rect 27252 4548 27304 4554
rect 27252 4490 27304 4496
rect 27264 4146 27292 4490
rect 26240 4140 26292 4146
rect 26240 4082 26292 4088
rect 27252 4140 27304 4146
rect 27252 4082 27304 4088
rect 26146 3632 26202 3641
rect 26146 3567 26202 3576
rect 25964 3528 26016 3534
rect 25964 3470 26016 3476
rect 26792 3528 26844 3534
rect 26792 3470 26844 3476
rect 27620 3528 27672 3534
rect 27620 3470 27672 3476
rect 25688 2440 25740 2446
rect 25594 2408 25650 2417
rect 25688 2382 25740 2388
rect 25594 2343 25650 2352
rect 25700 800 25728 2382
rect 25976 800 26004 3470
rect 26240 2848 26292 2854
rect 26240 2790 26292 2796
rect 26252 800 26280 2790
rect 26516 2508 26568 2514
rect 26516 2450 26568 2456
rect 26528 800 26556 2450
rect 26804 800 26832 3470
rect 27068 2848 27120 2854
rect 27068 2790 27120 2796
rect 27080 800 27108 2790
rect 27344 2440 27396 2446
rect 27344 2382 27396 2388
rect 27356 800 27384 2382
rect 27632 800 27660 3470
rect 27724 2310 27752 6394
rect 27816 5234 27844 8298
rect 27908 6458 27936 12406
rect 28000 12374 28028 12786
rect 27988 12368 28040 12374
rect 27988 12310 28040 12316
rect 27988 12164 28040 12170
rect 27988 12106 28040 12112
rect 28000 11218 28028 12106
rect 28080 11552 28132 11558
rect 28078 11520 28080 11529
rect 28132 11520 28134 11529
rect 28078 11455 28134 11464
rect 27988 11212 28040 11218
rect 27988 11154 28040 11160
rect 27988 10668 28040 10674
rect 27988 10610 28040 10616
rect 28000 8362 28028 10610
rect 28092 10554 28120 11455
rect 28184 11218 28212 13806
rect 28552 13530 28580 13806
rect 28540 13524 28592 13530
rect 28540 13466 28592 13472
rect 28264 13320 28316 13326
rect 28264 13262 28316 13268
rect 28356 13320 28408 13326
rect 28552 13308 28580 13466
rect 28408 13280 28580 13308
rect 28356 13262 28408 13268
rect 28172 11212 28224 11218
rect 28172 11154 28224 11160
rect 28092 10526 28212 10554
rect 28080 10464 28132 10470
rect 28078 10432 28080 10441
rect 28132 10432 28134 10441
rect 28078 10367 28134 10376
rect 27988 8356 28040 8362
rect 27988 8298 28040 8304
rect 27896 6452 27948 6458
rect 27896 6394 27948 6400
rect 28080 6248 28132 6254
rect 28080 6190 28132 6196
rect 28092 5710 28120 6190
rect 28080 5704 28132 5710
rect 28080 5646 28132 5652
rect 28092 5302 28120 5646
rect 28080 5296 28132 5302
rect 28080 5238 28132 5244
rect 27804 5228 27856 5234
rect 27804 5170 27856 5176
rect 28184 4758 28212 10526
rect 28276 7342 28304 13262
rect 28356 12844 28408 12850
rect 28356 12786 28408 12792
rect 28368 10810 28396 12786
rect 28356 10804 28408 10810
rect 28356 10746 28408 10752
rect 28552 10062 28580 13280
rect 28644 12850 28672 14962
rect 28816 14816 28868 14822
rect 28816 14758 28868 14764
rect 28828 14550 28856 14758
rect 28816 14544 28868 14550
rect 28816 14486 28868 14492
rect 29012 14482 29040 15370
rect 29090 15328 29146 15337
rect 29090 15263 29146 15272
rect 29000 14476 29052 14482
rect 29000 14418 29052 14424
rect 28908 14272 28960 14278
rect 28960 14220 29040 14226
rect 28908 14214 29040 14220
rect 28920 14198 29040 14214
rect 29012 13954 29040 14198
rect 29104 14074 29132 15263
rect 29274 14240 29330 14249
rect 29274 14175 29330 14184
rect 29092 14068 29144 14074
rect 29092 14010 29144 14016
rect 29288 14006 29316 14175
rect 29276 14000 29328 14006
rect 29012 13926 29132 13954
rect 29276 13942 29328 13948
rect 29104 13802 29132 13926
rect 29184 13932 29236 13938
rect 29184 13874 29236 13880
rect 29552 13932 29604 13938
rect 29552 13874 29604 13880
rect 29092 13796 29144 13802
rect 29092 13738 29144 13744
rect 28722 13560 28778 13569
rect 28722 13495 28724 13504
rect 28776 13495 28778 13504
rect 28724 13466 28776 13472
rect 28632 12844 28684 12850
rect 28632 12786 28684 12792
rect 29104 12481 29132 13738
rect 29196 12850 29224 13874
rect 29460 13320 29512 13326
rect 29460 13262 29512 13268
rect 29368 12912 29420 12918
rect 29288 12872 29368 12900
rect 29184 12844 29236 12850
rect 29184 12786 29236 12792
rect 29090 12472 29146 12481
rect 29090 12407 29146 12416
rect 28632 12164 28684 12170
rect 28632 12106 28684 12112
rect 28644 11558 28672 12106
rect 28724 12096 28776 12102
rect 28724 12038 28776 12044
rect 29000 12096 29052 12102
rect 29000 12038 29052 12044
rect 28632 11552 28684 11558
rect 28632 11494 28684 11500
rect 28736 11354 28764 12038
rect 29012 11898 29040 12038
rect 29000 11892 29052 11898
rect 29000 11834 29052 11840
rect 28724 11348 28776 11354
rect 28724 11290 28776 11296
rect 28632 11212 28684 11218
rect 28632 11154 28684 11160
rect 28448 10056 28500 10062
rect 28448 9998 28500 10004
rect 28540 10056 28592 10062
rect 28540 9998 28592 10004
rect 28460 8838 28488 9998
rect 28448 8832 28500 8838
rect 28448 8774 28500 8780
rect 28460 7818 28488 8774
rect 28540 7948 28592 7954
rect 28644 7936 28672 11154
rect 29196 11014 29224 12786
rect 29288 11830 29316 12872
rect 29368 12854 29420 12860
rect 29472 12850 29500 13262
rect 29460 12844 29512 12850
rect 29460 12786 29512 12792
rect 29472 12730 29500 12786
rect 29380 12702 29500 12730
rect 29276 11824 29328 11830
rect 29276 11766 29328 11772
rect 29380 11014 29408 12702
rect 29460 12640 29512 12646
rect 29460 12582 29512 12588
rect 29472 12306 29500 12582
rect 29564 12322 29592 13874
rect 29644 13728 29696 13734
rect 29644 13670 29696 13676
rect 29656 13326 29684 13670
rect 29644 13320 29696 13326
rect 29644 13262 29696 13268
rect 29644 12776 29696 12782
rect 29644 12718 29696 12724
rect 29656 12434 29684 12718
rect 29748 12646 29776 15574
rect 29828 15496 29880 15502
rect 29828 15438 29880 15444
rect 29840 13802 29868 15438
rect 29932 14346 29960 16458
rect 30116 15994 30144 16526
rect 30024 15966 30144 15994
rect 30024 15910 30052 15966
rect 30012 15904 30064 15910
rect 30012 15846 30064 15852
rect 30104 15904 30156 15910
rect 30104 15846 30156 15852
rect 30012 15496 30064 15502
rect 30012 15438 30064 15444
rect 30024 15162 30052 15438
rect 30012 15156 30064 15162
rect 30012 15098 30064 15104
rect 30012 14952 30064 14958
rect 30012 14894 30064 14900
rect 29920 14340 29972 14346
rect 29920 14282 29972 14288
rect 29828 13796 29880 13802
rect 29828 13738 29880 13744
rect 29840 13530 29868 13738
rect 29828 13524 29880 13530
rect 29828 13466 29880 13472
rect 29932 13190 29960 14282
rect 29920 13184 29972 13190
rect 29920 13126 29972 13132
rect 29736 12640 29788 12646
rect 29736 12582 29788 12588
rect 29656 12406 29868 12434
rect 29460 12300 29512 12306
rect 29564 12294 29776 12322
rect 29840 12306 29868 12406
rect 29460 12242 29512 12248
rect 29472 11898 29500 12242
rect 29644 12232 29696 12238
rect 29644 12174 29696 12180
rect 29552 12164 29604 12170
rect 29552 12106 29604 12112
rect 29460 11892 29512 11898
rect 29460 11834 29512 11840
rect 29184 11008 29236 11014
rect 28722 10976 28778 10985
rect 29184 10950 29236 10956
rect 29368 11008 29420 11014
rect 29368 10950 29420 10956
rect 28722 10911 28778 10920
rect 28736 9994 28764 10911
rect 28908 10736 28960 10742
rect 28908 10678 28960 10684
rect 28816 10464 28868 10470
rect 28816 10406 28868 10412
rect 28828 10033 28856 10406
rect 28814 10024 28870 10033
rect 28724 9988 28776 9994
rect 28814 9959 28870 9968
rect 28724 9930 28776 9936
rect 28816 8832 28868 8838
rect 28920 8820 28948 10678
rect 29000 10056 29052 10062
rect 29000 9998 29052 10004
rect 29012 9178 29040 9998
rect 29196 9994 29224 10950
rect 29368 10668 29420 10674
rect 29368 10610 29420 10616
rect 29460 10668 29512 10674
rect 29460 10610 29512 10616
rect 29184 9988 29236 9994
rect 29184 9930 29236 9936
rect 29092 9580 29144 9586
rect 29092 9522 29144 9528
rect 29276 9580 29328 9586
rect 29276 9522 29328 9528
rect 29104 9450 29132 9522
rect 29092 9444 29144 9450
rect 29092 9386 29144 9392
rect 29000 9172 29052 9178
rect 29000 9114 29052 9120
rect 28868 8792 28948 8820
rect 28816 8774 28868 8780
rect 28724 8288 28776 8294
rect 28724 8230 28776 8236
rect 28592 7908 28672 7936
rect 28540 7890 28592 7896
rect 28356 7812 28408 7818
rect 28356 7754 28408 7760
rect 28448 7812 28500 7818
rect 28448 7754 28500 7760
rect 28264 7336 28316 7342
rect 28264 7278 28316 7284
rect 28264 6656 28316 6662
rect 28264 6598 28316 6604
rect 28276 6254 28304 6598
rect 28264 6248 28316 6254
rect 28264 6190 28316 6196
rect 28276 4758 28304 6190
rect 28368 6118 28396 7754
rect 28552 7206 28580 7890
rect 28540 7200 28592 7206
rect 28540 7142 28592 7148
rect 28552 6730 28580 7142
rect 28540 6724 28592 6730
rect 28540 6666 28592 6672
rect 28540 6316 28592 6322
rect 28540 6258 28592 6264
rect 28356 6112 28408 6118
rect 28356 6054 28408 6060
rect 28552 5914 28580 6258
rect 28540 5908 28592 5914
rect 28540 5850 28592 5856
rect 28540 5296 28592 5302
rect 28540 5238 28592 5244
rect 28172 4752 28224 4758
rect 28172 4694 28224 4700
rect 28264 4752 28316 4758
rect 28264 4694 28316 4700
rect 27804 4616 27856 4622
rect 27802 4584 27804 4593
rect 27856 4584 27858 4593
rect 27802 4519 27858 4528
rect 28552 4214 28580 5238
rect 28736 4826 28764 8230
rect 28828 6254 28856 8774
rect 29012 8378 29040 9114
rect 28920 8350 29040 8378
rect 28920 8090 28948 8350
rect 28908 8084 28960 8090
rect 28908 8026 28960 8032
rect 28908 7336 28960 7342
rect 28908 7278 28960 7284
rect 28920 6934 28948 7278
rect 28908 6928 28960 6934
rect 28908 6870 28960 6876
rect 29000 6316 29052 6322
rect 29104 6304 29132 9386
rect 29288 9178 29316 9522
rect 29276 9172 29328 9178
rect 29276 9114 29328 9120
rect 29380 8974 29408 10610
rect 29472 10266 29500 10610
rect 29460 10260 29512 10266
rect 29460 10202 29512 10208
rect 29368 8968 29420 8974
rect 29368 8910 29420 8916
rect 29184 8424 29236 8430
rect 29184 8366 29236 8372
rect 29196 7886 29224 8366
rect 29184 7880 29236 7886
rect 29184 7822 29236 7828
rect 29196 7002 29224 7822
rect 29564 7818 29592 12106
rect 29656 11898 29684 12174
rect 29644 11892 29696 11898
rect 29644 11834 29696 11840
rect 29748 11642 29776 12294
rect 29828 12300 29880 12306
rect 29828 12242 29880 12248
rect 29920 12232 29972 12238
rect 30024 12220 30052 14894
rect 29972 12192 30052 12220
rect 29920 12174 29972 12180
rect 29826 12064 29882 12073
rect 29826 11999 29882 12008
rect 29840 11762 29868 11999
rect 29828 11756 29880 11762
rect 29828 11698 29880 11704
rect 29656 11614 29776 11642
rect 29552 7812 29604 7818
rect 29552 7754 29604 7760
rect 29656 7206 29684 11614
rect 29736 11552 29788 11558
rect 29736 11494 29788 11500
rect 30012 11552 30064 11558
rect 30012 11494 30064 11500
rect 29748 11121 29776 11494
rect 29826 11384 29882 11393
rect 29826 11319 29882 11328
rect 29840 11286 29868 11319
rect 29828 11280 29880 11286
rect 29828 11222 29880 11228
rect 29734 11112 29790 11121
rect 29734 11047 29790 11056
rect 29920 11008 29972 11014
rect 29920 10950 29972 10956
rect 29932 10198 29960 10950
rect 29920 10192 29972 10198
rect 29920 10134 29972 10140
rect 29932 10062 29960 10134
rect 29920 10056 29972 10062
rect 29920 9998 29972 10004
rect 29828 9988 29880 9994
rect 29828 9930 29880 9936
rect 29736 9376 29788 9382
rect 29736 9318 29788 9324
rect 29748 7886 29776 9318
rect 29840 9110 29868 9930
rect 29920 9920 29972 9926
rect 29920 9862 29972 9868
rect 29828 9104 29880 9110
rect 29828 9046 29880 9052
rect 29932 8974 29960 9862
rect 29920 8968 29972 8974
rect 29920 8910 29972 8916
rect 29736 7880 29788 7886
rect 29736 7822 29788 7828
rect 29828 7744 29880 7750
rect 29828 7686 29880 7692
rect 29840 7410 29868 7686
rect 29828 7404 29880 7410
rect 29828 7346 29880 7352
rect 29644 7200 29696 7206
rect 29644 7142 29696 7148
rect 29656 7002 29684 7142
rect 29184 6996 29236 7002
rect 29184 6938 29236 6944
rect 29644 6996 29696 7002
rect 29644 6938 29696 6944
rect 29196 6322 29224 6938
rect 29052 6276 29132 6304
rect 29184 6316 29236 6322
rect 29000 6258 29052 6264
rect 29184 6258 29236 6264
rect 28816 6248 28868 6254
rect 28816 6190 28868 6196
rect 28816 5024 28868 5030
rect 28816 4966 28868 4972
rect 28724 4820 28776 4826
rect 28724 4762 28776 4768
rect 28632 4752 28684 4758
rect 28632 4694 28684 4700
rect 28644 4468 28672 4694
rect 28828 4622 28856 4966
rect 28908 4684 28960 4690
rect 28908 4626 28960 4632
rect 28816 4616 28868 4622
rect 28816 4558 28868 4564
rect 28920 4468 28948 4626
rect 29012 4622 29040 6258
rect 29656 5302 29684 6938
rect 29840 6798 29868 7346
rect 29828 6792 29880 6798
rect 29828 6734 29880 6740
rect 29644 5296 29696 5302
rect 29644 5238 29696 5244
rect 29920 5160 29972 5166
rect 29920 5102 29972 5108
rect 29932 4622 29960 5102
rect 29000 4616 29052 4622
rect 29000 4558 29052 4564
rect 29736 4616 29788 4622
rect 29736 4558 29788 4564
rect 29920 4616 29972 4622
rect 29920 4558 29972 4564
rect 28644 4440 28948 4468
rect 29748 4282 29776 4558
rect 29736 4276 29788 4282
rect 29736 4218 29788 4224
rect 28540 4208 28592 4214
rect 28540 4150 28592 4156
rect 30024 3942 30052 11494
rect 30116 10742 30144 15846
rect 30208 15502 30236 16662
rect 30293 16584 30345 16590
rect 30293 16526 30345 16532
rect 30196 15496 30248 15502
rect 30196 15438 30248 15444
rect 30300 15434 30328 16526
rect 30472 16040 30524 16046
rect 30472 15982 30524 15988
rect 30288 15428 30340 15434
rect 30288 15370 30340 15376
rect 30380 15360 30432 15366
rect 30208 15308 30380 15314
rect 30208 15302 30432 15308
rect 30208 15286 30420 15302
rect 30208 15094 30236 15286
rect 30196 15088 30248 15094
rect 30196 15030 30248 15036
rect 30288 15020 30340 15026
rect 30288 14962 30340 14968
rect 30196 14884 30248 14890
rect 30196 14826 30248 14832
rect 30208 14618 30236 14826
rect 30300 14618 30328 14962
rect 30196 14612 30248 14618
rect 30196 14554 30248 14560
rect 30288 14612 30340 14618
rect 30288 14554 30340 14560
rect 30208 13394 30236 14554
rect 30196 13388 30248 13394
rect 30196 13330 30248 13336
rect 30196 13252 30248 13258
rect 30196 13194 30248 13200
rect 30208 12238 30236 13194
rect 30196 12232 30248 12238
rect 30196 12174 30248 12180
rect 30380 12096 30432 12102
rect 30380 12038 30432 12044
rect 30392 11762 30420 12038
rect 30196 11756 30248 11762
rect 30196 11698 30248 11704
rect 30380 11756 30432 11762
rect 30380 11698 30432 11704
rect 30208 11558 30236 11698
rect 30196 11552 30248 11558
rect 30196 11494 30248 11500
rect 30286 11384 30342 11393
rect 30286 11319 30342 11328
rect 30196 11144 30248 11150
rect 30196 11086 30248 11092
rect 30300 11098 30328 11319
rect 30484 11218 30512 15982
rect 30564 15564 30616 15570
rect 30564 15506 30616 15512
rect 30472 11212 30524 11218
rect 30472 11154 30524 11160
rect 30104 10736 30156 10742
rect 30104 10678 30156 10684
rect 30208 8974 30236 11086
rect 30300 11070 30420 11098
rect 30392 10674 30420 11070
rect 30380 10668 30432 10674
rect 30380 10610 30432 10616
rect 30288 10464 30340 10470
rect 30288 10406 30340 10412
rect 30300 9654 30328 10406
rect 30576 9654 30604 15506
rect 30668 15162 30696 19790
rect 30760 18154 30788 20946
rect 30852 20942 30880 21286
rect 30840 20936 30892 20942
rect 30840 20878 30892 20884
rect 30944 20641 30972 21286
rect 30930 20632 30986 20641
rect 30930 20567 30986 20576
rect 30944 19854 30972 20567
rect 31036 19922 31064 24142
rect 32220 24132 32272 24138
rect 32220 24074 32272 24080
rect 32128 22432 32180 22438
rect 32128 22374 32180 22380
rect 32140 22030 32168 22374
rect 31668 22024 31720 22030
rect 31668 21966 31720 21972
rect 32128 22024 32180 22030
rect 32128 21966 32180 21972
rect 31680 20505 31708 21966
rect 32128 20936 32180 20942
rect 32128 20878 32180 20884
rect 31760 20800 31812 20806
rect 31760 20742 31812 20748
rect 31666 20496 31722 20505
rect 31666 20431 31722 20440
rect 31024 19916 31076 19922
rect 31024 19858 31076 19864
rect 30932 19848 30984 19854
rect 30932 19790 30984 19796
rect 31116 19712 31168 19718
rect 31116 19654 31168 19660
rect 31128 19378 31156 19654
rect 31116 19372 31168 19378
rect 31116 19314 31168 19320
rect 30748 18148 30800 18154
rect 30748 18090 30800 18096
rect 31128 17678 31156 19314
rect 31300 19304 31352 19310
rect 31300 19246 31352 19252
rect 31116 17672 31168 17678
rect 31116 17614 31168 17620
rect 31208 16992 31260 16998
rect 31208 16934 31260 16940
rect 31220 16590 31248 16934
rect 31208 16584 31260 16590
rect 31208 16526 31260 16532
rect 30840 16516 30892 16522
rect 30840 16458 30892 16464
rect 30852 15366 30880 16458
rect 31116 15564 31168 15570
rect 31116 15506 31168 15512
rect 31128 15434 31156 15506
rect 31116 15428 31168 15434
rect 31116 15370 31168 15376
rect 30840 15360 30892 15366
rect 30840 15302 30892 15308
rect 30656 15156 30708 15162
rect 30656 15098 30708 15104
rect 30656 15020 30708 15026
rect 30656 14962 30708 14968
rect 30668 14929 30696 14962
rect 30654 14920 30710 14929
rect 30654 14855 30710 14864
rect 30852 14346 30880 15302
rect 31022 15056 31078 15065
rect 31022 14991 31024 15000
rect 31076 14991 31078 15000
rect 31024 14962 31076 14968
rect 31220 14890 31248 16526
rect 31208 14884 31260 14890
rect 31208 14826 31260 14832
rect 31312 14770 31340 19246
rect 31484 17672 31536 17678
rect 31484 17614 31536 17620
rect 31496 17134 31524 17614
rect 31484 17128 31536 17134
rect 31484 17070 31536 17076
rect 31392 16788 31444 16794
rect 31392 16730 31444 16736
rect 31404 15026 31432 16730
rect 31496 15570 31524 17070
rect 31576 16652 31628 16658
rect 31576 16594 31628 16600
rect 31484 15564 31536 15570
rect 31484 15506 31536 15512
rect 31496 15162 31524 15506
rect 31484 15156 31536 15162
rect 31484 15098 31536 15104
rect 31392 15020 31444 15026
rect 31392 14962 31444 14968
rect 31220 14742 31340 14770
rect 31024 14408 31076 14414
rect 31024 14350 31076 14356
rect 30840 14340 30892 14346
rect 30840 14282 30892 14288
rect 31036 14074 31064 14350
rect 31024 14068 31076 14074
rect 31024 14010 31076 14016
rect 30656 13184 30708 13190
rect 30656 13126 30708 13132
rect 30668 12850 30696 13126
rect 30932 12912 30984 12918
rect 30932 12854 30984 12860
rect 30656 12844 30708 12850
rect 30656 12786 30708 12792
rect 30748 12844 30800 12850
rect 30748 12786 30800 12792
rect 30760 12434 30788 12786
rect 30668 12406 30788 12434
rect 30288 9648 30340 9654
rect 30288 9590 30340 9596
rect 30564 9648 30616 9654
rect 30564 9590 30616 9596
rect 30300 9450 30328 9590
rect 30288 9444 30340 9450
rect 30288 9386 30340 9392
rect 30196 8968 30248 8974
rect 30196 8910 30248 8916
rect 30668 7342 30696 12406
rect 30944 12306 30972 12854
rect 31116 12844 31168 12850
rect 31116 12786 31168 12792
rect 31128 12374 31156 12786
rect 31116 12368 31168 12374
rect 31116 12310 31168 12316
rect 30932 12300 30984 12306
rect 30932 12242 30984 12248
rect 31128 12073 31156 12310
rect 31114 12064 31170 12073
rect 31114 11999 31170 12008
rect 30838 10568 30894 10577
rect 30838 10503 30840 10512
rect 30892 10503 30894 10512
rect 30840 10474 30892 10480
rect 31116 10464 31168 10470
rect 31116 10406 31168 10412
rect 31128 9994 31156 10406
rect 31220 10169 31248 14742
rect 31404 14482 31432 14962
rect 31392 14476 31444 14482
rect 31392 14418 31444 14424
rect 31392 13456 31444 13462
rect 31390 13424 31392 13433
rect 31444 13424 31446 13433
rect 31390 13359 31446 13368
rect 31392 13320 31444 13326
rect 31392 13262 31444 13268
rect 31300 12640 31352 12646
rect 31298 12608 31300 12617
rect 31352 12608 31354 12617
rect 31298 12543 31354 12552
rect 31404 12442 31432 13262
rect 31392 12436 31444 12442
rect 31392 12378 31444 12384
rect 31404 12238 31432 12378
rect 31300 12232 31352 12238
rect 31300 12174 31352 12180
rect 31392 12232 31444 12238
rect 31392 12174 31444 12180
rect 31206 10160 31262 10169
rect 31206 10095 31262 10104
rect 31220 10062 31248 10095
rect 31208 10056 31260 10062
rect 31208 9998 31260 10004
rect 31116 9988 31168 9994
rect 31116 9930 31168 9936
rect 30748 9580 30800 9586
rect 30748 9522 30800 9528
rect 30760 9042 30788 9522
rect 31116 9512 31168 9518
rect 31116 9454 31168 9460
rect 30748 9036 30800 9042
rect 30748 8978 30800 8984
rect 30840 9036 30892 9042
rect 30840 8978 30892 8984
rect 30852 8634 30880 8978
rect 31128 8974 31156 9454
rect 31116 8968 31168 8974
rect 31116 8910 31168 8916
rect 31024 8900 31076 8906
rect 31024 8842 31076 8848
rect 30840 8628 30892 8634
rect 30840 8570 30892 8576
rect 31036 8090 31064 8842
rect 31024 8084 31076 8090
rect 31024 8026 31076 8032
rect 31036 7886 31064 8026
rect 31312 7954 31340 12174
rect 31588 12170 31616 16594
rect 31680 16017 31708 20431
rect 31772 19922 31800 20742
rect 32036 20460 32088 20466
rect 32036 20402 32088 20408
rect 31760 19916 31812 19922
rect 31760 19858 31812 19864
rect 31772 19310 31800 19858
rect 31852 19440 31904 19446
rect 31852 19382 31904 19388
rect 31760 19304 31812 19310
rect 31760 19246 31812 19252
rect 31864 18630 31892 19382
rect 32048 19174 32076 20402
rect 32140 20058 32168 20878
rect 32232 20262 32260 24074
rect 33060 23186 33088 25774
rect 34704 25696 34756 25702
rect 34704 25638 34756 25644
rect 34244 25356 34296 25362
rect 34244 25298 34296 25304
rect 33508 25220 33560 25226
rect 33508 25162 33560 25168
rect 33140 24812 33192 24818
rect 33140 24754 33192 24760
rect 33048 23180 33100 23186
rect 33048 23122 33100 23128
rect 32404 22024 32456 22030
rect 32404 21966 32456 21972
rect 32416 21554 32444 21966
rect 32496 21684 32548 21690
rect 32496 21626 32548 21632
rect 32312 21548 32364 21554
rect 32312 21490 32364 21496
rect 32404 21548 32456 21554
rect 32404 21490 32456 21496
rect 32324 20641 32352 21490
rect 32508 20942 32536 21626
rect 32956 21616 33008 21622
rect 32956 21558 33008 21564
rect 32772 21344 32824 21350
rect 32772 21286 32824 21292
rect 32496 20936 32548 20942
rect 32784 20913 32812 21286
rect 32496 20878 32548 20884
rect 32770 20904 32826 20913
rect 32770 20839 32826 20848
rect 32496 20800 32548 20806
rect 32496 20742 32548 20748
rect 32310 20632 32366 20641
rect 32310 20567 32366 20576
rect 32220 20256 32272 20262
rect 32220 20198 32272 20204
rect 32128 20052 32180 20058
rect 32128 19994 32180 20000
rect 32036 19168 32088 19174
rect 32036 19110 32088 19116
rect 31852 18624 31904 18630
rect 31852 18566 31904 18572
rect 32220 17740 32272 17746
rect 32324 17728 32352 20567
rect 32404 20528 32456 20534
rect 32404 20470 32456 20476
rect 32416 19718 32444 20470
rect 32508 20466 32536 20742
rect 32496 20460 32548 20466
rect 32496 20402 32548 20408
rect 32784 19854 32812 20839
rect 32968 20602 32996 21558
rect 33060 21554 33088 23122
rect 33048 21548 33100 21554
rect 33048 21490 33100 21496
rect 32956 20596 33008 20602
rect 32956 20538 33008 20544
rect 32772 19848 32824 19854
rect 32772 19790 32824 19796
rect 32404 19712 32456 19718
rect 32404 19654 32456 19660
rect 32588 19372 32640 19378
rect 32588 19314 32640 19320
rect 32496 19168 32548 19174
rect 32496 19110 32548 19116
rect 32404 18760 32456 18766
rect 32404 18702 32456 18708
rect 32272 17700 32352 17728
rect 32220 17682 32272 17688
rect 32232 17542 32260 17682
rect 32220 17536 32272 17542
rect 32220 17478 32272 17484
rect 31944 16788 31996 16794
rect 31944 16730 31996 16736
rect 31666 16008 31722 16017
rect 31666 15943 31722 15952
rect 31760 15496 31812 15502
rect 31760 15438 31812 15444
rect 31772 15162 31800 15438
rect 31760 15156 31812 15162
rect 31760 15098 31812 15104
rect 31668 14068 31720 14074
rect 31668 14010 31720 14016
rect 31680 13326 31708 14010
rect 31668 13320 31720 13326
rect 31668 13262 31720 13268
rect 31576 12164 31628 12170
rect 31576 12106 31628 12112
rect 31956 10742 31984 16730
rect 32128 15360 32180 15366
rect 32128 15302 32180 15308
rect 32140 15026 32168 15302
rect 32128 15020 32180 15026
rect 32128 14962 32180 14968
rect 32232 14498 32260 17478
rect 32416 16454 32444 18702
rect 32404 16448 32456 16454
rect 32404 16390 32456 16396
rect 32312 15020 32364 15026
rect 32312 14962 32364 14968
rect 32324 14618 32352 14962
rect 32312 14612 32364 14618
rect 32312 14554 32364 14560
rect 32232 14470 32352 14498
rect 32128 12232 32180 12238
rect 32128 12174 32180 12180
rect 31944 10736 31996 10742
rect 31944 10678 31996 10684
rect 31484 10668 31536 10674
rect 31484 10610 31536 10616
rect 31496 10266 31524 10610
rect 31760 10600 31812 10606
rect 31760 10542 31812 10548
rect 31484 10260 31536 10266
rect 31484 10202 31536 10208
rect 31772 10062 31800 10542
rect 32140 10538 32168 12174
rect 32220 12096 32272 12102
rect 32220 12038 32272 12044
rect 32232 11150 32260 12038
rect 32220 11144 32272 11150
rect 32220 11086 32272 11092
rect 32128 10532 32180 10538
rect 32128 10474 32180 10480
rect 32324 10441 32352 14470
rect 32508 14414 32536 19110
rect 32496 14408 32548 14414
rect 32496 14350 32548 14356
rect 32496 12300 32548 12306
rect 32496 12242 32548 12248
rect 32402 12200 32458 12209
rect 32402 12135 32404 12144
rect 32456 12135 32458 12144
rect 32404 12106 32456 12112
rect 32508 11150 32536 12242
rect 32496 11144 32548 11150
rect 32496 11086 32548 11092
rect 32310 10432 32366 10441
rect 32310 10367 32366 10376
rect 32036 10124 32088 10130
rect 32036 10066 32088 10072
rect 31760 10056 31812 10062
rect 31760 9998 31812 10004
rect 31482 9480 31538 9489
rect 31482 9415 31538 9424
rect 31496 8906 31524 9415
rect 31484 8900 31536 8906
rect 31484 8842 31536 8848
rect 31496 8634 31524 8842
rect 31484 8628 31536 8634
rect 31484 8570 31536 8576
rect 31576 8288 31628 8294
rect 31576 8230 31628 8236
rect 31588 7954 31616 8230
rect 31772 8090 31800 9998
rect 31944 9920 31996 9926
rect 31944 9862 31996 9868
rect 31852 9036 31904 9042
rect 31852 8978 31904 8984
rect 31864 8838 31892 8978
rect 31956 8974 31984 9862
rect 32048 9518 32076 10066
rect 32324 9761 32352 10367
rect 32600 10130 32628 19314
rect 33048 18760 33100 18766
rect 33152 18748 33180 24754
rect 33520 24614 33548 25162
rect 34256 24954 34284 25298
rect 34244 24948 34296 24954
rect 34244 24890 34296 24896
rect 33692 24812 33744 24818
rect 33692 24754 33744 24760
rect 34428 24812 34480 24818
rect 34428 24754 34480 24760
rect 33508 24608 33560 24614
rect 33508 24550 33560 24556
rect 33508 23248 33560 23254
rect 33508 23190 33560 23196
rect 33520 22681 33548 23190
rect 33600 22976 33652 22982
rect 33600 22918 33652 22924
rect 33506 22672 33562 22681
rect 33506 22607 33508 22616
rect 33560 22607 33562 22616
rect 33508 22578 33560 22584
rect 33612 21350 33640 22918
rect 33600 21344 33652 21350
rect 33600 21286 33652 21292
rect 33612 20942 33640 21286
rect 33704 21146 33732 24754
rect 34440 24410 34468 24754
rect 34716 24750 34744 25638
rect 34808 25430 34836 25978
rect 35360 25906 35388 26182
rect 35348 25900 35400 25906
rect 35348 25842 35400 25848
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 34796 25424 34848 25430
rect 34796 25366 34848 25372
rect 34808 24886 34836 25366
rect 35348 25288 35400 25294
rect 35348 25230 35400 25236
rect 34796 24880 34848 24886
rect 34796 24822 34848 24828
rect 34704 24744 34756 24750
rect 34704 24686 34756 24692
rect 34428 24404 34480 24410
rect 34428 24346 34480 24352
rect 34808 24274 34836 24822
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 35360 24410 35388 25230
rect 35452 25158 35480 26250
rect 35820 25702 35848 26318
rect 35808 25696 35860 25702
rect 35808 25638 35860 25644
rect 36096 25498 36124 26318
rect 37740 26308 37792 26314
rect 37740 26250 37792 26256
rect 36084 25492 36136 25498
rect 36084 25434 36136 25440
rect 35900 25288 35952 25294
rect 35900 25230 35952 25236
rect 35440 25152 35492 25158
rect 35440 25094 35492 25100
rect 35452 24614 35480 25094
rect 35440 24608 35492 24614
rect 35440 24550 35492 24556
rect 35348 24404 35400 24410
rect 35348 24346 35400 24352
rect 35452 24342 35480 24550
rect 35440 24336 35492 24342
rect 35440 24278 35492 24284
rect 34796 24268 34848 24274
rect 34796 24210 34848 24216
rect 34060 23724 34112 23730
rect 34060 23666 34112 23672
rect 33876 23656 33928 23662
rect 33876 23598 33928 23604
rect 33784 23520 33836 23526
rect 33784 23462 33836 23468
rect 33796 23118 33824 23462
rect 33784 23112 33836 23118
rect 33784 23054 33836 23060
rect 33796 22438 33824 23054
rect 33888 22642 33916 23598
rect 33968 23520 34020 23526
rect 33968 23462 34020 23468
rect 33980 23118 34008 23462
rect 34072 23322 34100 23666
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 34060 23316 34112 23322
rect 34060 23258 34112 23264
rect 33968 23112 34020 23118
rect 33968 23054 34020 23060
rect 33876 22636 33928 22642
rect 33876 22578 33928 22584
rect 33888 22506 33916 22578
rect 33876 22500 33928 22506
rect 33876 22442 33928 22448
rect 33784 22432 33836 22438
rect 33784 22374 33836 22380
rect 34072 21146 34100 23258
rect 35912 23118 35940 25230
rect 36728 25220 36780 25226
rect 36728 25162 36780 25168
rect 37464 25220 37516 25226
rect 37464 25162 37516 25168
rect 36740 24954 36768 25162
rect 36728 24948 36780 24954
rect 36728 24890 36780 24896
rect 37476 24818 37504 25162
rect 37752 24818 37780 26250
rect 37464 24812 37516 24818
rect 37464 24754 37516 24760
rect 37740 24812 37792 24818
rect 37740 24754 37792 24760
rect 38936 24812 38988 24818
rect 38936 24754 38988 24760
rect 36268 24744 36320 24750
rect 36268 24686 36320 24692
rect 38660 24744 38712 24750
rect 38660 24686 38712 24692
rect 36084 23316 36136 23322
rect 36084 23258 36136 23264
rect 34152 23112 34204 23118
rect 34152 23054 34204 23060
rect 35900 23112 35952 23118
rect 35900 23054 35952 23060
rect 34164 22982 34192 23054
rect 34428 23044 34480 23050
rect 34428 22986 34480 22992
rect 34796 23044 34848 23050
rect 34796 22986 34848 22992
rect 35624 23044 35676 23050
rect 35624 22986 35676 22992
rect 34152 22976 34204 22982
rect 34152 22918 34204 22924
rect 34164 22642 34192 22918
rect 34440 22642 34468 22986
rect 34808 22778 34836 22986
rect 34796 22772 34848 22778
rect 34796 22714 34848 22720
rect 34152 22636 34204 22642
rect 34152 22578 34204 22584
rect 34428 22636 34480 22642
rect 34428 22578 34480 22584
rect 34796 22636 34848 22642
rect 34796 22578 34848 22584
rect 35348 22636 35400 22642
rect 35348 22578 35400 22584
rect 34440 21554 34468 22578
rect 34808 22098 34836 22578
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 34796 22092 34848 22098
rect 34796 22034 34848 22040
rect 35360 21894 35388 22578
rect 35636 22506 35664 22986
rect 35808 22772 35860 22778
rect 35808 22714 35860 22720
rect 35624 22500 35676 22506
rect 35624 22442 35676 22448
rect 35440 22092 35492 22098
rect 35440 22034 35492 22040
rect 35348 21888 35400 21894
rect 35348 21830 35400 21836
rect 34428 21548 34480 21554
rect 34428 21490 34480 21496
rect 34704 21480 34756 21486
rect 34704 21422 34756 21428
rect 33692 21140 33744 21146
rect 33692 21082 33744 21088
rect 34060 21140 34112 21146
rect 34060 21082 34112 21088
rect 34336 21004 34388 21010
rect 34336 20946 34388 20952
rect 33324 20936 33376 20942
rect 33324 20878 33376 20884
rect 33600 20936 33652 20942
rect 33600 20878 33652 20884
rect 33692 20936 33744 20942
rect 33692 20878 33744 20884
rect 33336 19310 33364 20878
rect 33704 20466 33732 20878
rect 34348 20534 34376 20946
rect 34336 20528 34388 20534
rect 34336 20470 34388 20476
rect 33692 20460 33744 20466
rect 33692 20402 33744 20408
rect 33784 20392 33836 20398
rect 33784 20334 33836 20340
rect 34244 20392 34296 20398
rect 34244 20334 34296 20340
rect 33508 19848 33560 19854
rect 33508 19790 33560 19796
rect 33520 19378 33548 19790
rect 33796 19446 33824 20334
rect 34152 20256 34204 20262
rect 34152 20198 34204 20204
rect 34164 19922 34192 20198
rect 34256 20058 34284 20334
rect 34244 20052 34296 20058
rect 34244 19994 34296 20000
rect 34152 19916 34204 19922
rect 34152 19858 34204 19864
rect 33876 19848 33928 19854
rect 33876 19790 33928 19796
rect 33784 19440 33836 19446
rect 33784 19382 33836 19388
rect 33508 19372 33560 19378
rect 33508 19314 33560 19320
rect 33324 19304 33376 19310
rect 33324 19246 33376 19252
rect 33796 18766 33824 19382
rect 33100 18720 33180 18748
rect 33508 18760 33560 18766
rect 33048 18702 33100 18708
rect 33508 18702 33560 18708
rect 33784 18760 33836 18766
rect 33784 18702 33836 18708
rect 32680 18692 32732 18698
rect 32680 18634 32732 18640
rect 32692 17882 32720 18634
rect 33324 18624 33376 18630
rect 33324 18566 33376 18572
rect 32680 17876 32732 17882
rect 32680 17818 32732 17824
rect 33232 17808 33284 17814
rect 33232 17750 33284 17756
rect 32864 17536 32916 17542
rect 32864 17478 32916 17484
rect 32876 16794 32904 17478
rect 33244 17202 33272 17750
rect 33232 17196 33284 17202
rect 33232 17138 33284 17144
rect 32864 16788 32916 16794
rect 32864 16730 32916 16736
rect 33244 16454 33272 17138
rect 33336 16522 33364 18566
rect 33520 18306 33548 18702
rect 33600 18352 33652 18358
rect 33520 18300 33600 18306
rect 33520 18294 33652 18300
rect 33520 18278 33640 18294
rect 33416 17672 33468 17678
rect 33416 17614 33468 17620
rect 33324 16516 33376 16522
rect 33324 16458 33376 16464
rect 33232 16448 33284 16454
rect 33232 16390 33284 16396
rect 32864 16108 32916 16114
rect 32864 16050 32916 16056
rect 32876 15706 32904 16050
rect 32864 15700 32916 15706
rect 32864 15642 32916 15648
rect 32864 15020 32916 15026
rect 32864 14962 32916 14968
rect 32678 14920 32734 14929
rect 32678 14855 32680 14864
rect 32732 14855 32734 14864
rect 32680 14826 32732 14832
rect 32772 14816 32824 14822
rect 32772 14758 32824 14764
rect 32680 14476 32732 14482
rect 32680 14418 32732 14424
rect 32692 12434 32720 14418
rect 32784 14006 32812 14758
rect 32876 14385 32904 14962
rect 32862 14376 32918 14385
rect 33336 14346 33364 16458
rect 33428 15502 33456 17614
rect 33520 16114 33548 18278
rect 33888 18154 33916 19790
rect 34716 19718 34744 21422
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 35360 19786 35388 21830
rect 34796 19780 34848 19786
rect 34796 19722 34848 19728
rect 35348 19780 35400 19786
rect 35348 19722 35400 19728
rect 34704 19712 34756 19718
rect 34704 19654 34756 19660
rect 34612 19372 34664 19378
rect 34612 19314 34664 19320
rect 34624 18766 34652 19314
rect 34716 19310 34744 19654
rect 34808 19378 34836 19722
rect 34888 19712 34940 19718
rect 34886 19680 34888 19689
rect 34940 19680 34942 19689
rect 34886 19615 34942 19624
rect 34796 19372 34848 19378
rect 34796 19314 34848 19320
rect 34704 19304 34756 19310
rect 34704 19246 34756 19252
rect 34704 19168 34756 19174
rect 34704 19110 34756 19116
rect 34612 18760 34664 18766
rect 34612 18702 34664 18708
rect 33968 18692 34020 18698
rect 33968 18634 34020 18640
rect 33980 18426 34008 18634
rect 34612 18624 34664 18630
rect 34612 18566 34664 18572
rect 33968 18420 34020 18426
rect 33968 18362 34020 18368
rect 33980 18222 34008 18362
rect 33968 18216 34020 18222
rect 33968 18158 34020 18164
rect 33876 18148 33928 18154
rect 33876 18090 33928 18096
rect 34520 16992 34572 16998
rect 34520 16934 34572 16940
rect 33600 16584 33652 16590
rect 33600 16526 33652 16532
rect 33508 16108 33560 16114
rect 33508 16050 33560 16056
rect 33612 15910 33640 16526
rect 34532 16522 34560 16934
rect 33784 16516 33836 16522
rect 33784 16458 33836 16464
rect 34520 16516 34572 16522
rect 34520 16458 34572 16464
rect 33692 16040 33744 16046
rect 33692 15982 33744 15988
rect 33600 15904 33652 15910
rect 33600 15846 33652 15852
rect 33612 15502 33640 15846
rect 33416 15496 33468 15502
rect 33416 15438 33468 15444
rect 33600 15496 33652 15502
rect 33600 15438 33652 15444
rect 33704 15366 33732 15982
rect 33796 15366 33824 16458
rect 34532 15638 34560 16458
rect 34520 15632 34572 15638
rect 34520 15574 34572 15580
rect 33692 15360 33744 15366
rect 33692 15302 33744 15308
rect 33784 15360 33836 15366
rect 33784 15302 33836 15308
rect 33508 15088 33560 15094
rect 33508 15030 33560 15036
rect 32862 14311 32918 14320
rect 33140 14340 33192 14346
rect 33140 14282 33192 14288
rect 33324 14340 33376 14346
rect 33324 14282 33376 14288
rect 32772 14000 32824 14006
rect 32772 13942 32824 13948
rect 32692 12406 32904 12434
rect 32680 12232 32732 12238
rect 32680 12174 32732 12180
rect 32588 10124 32640 10130
rect 32588 10066 32640 10072
rect 32310 9752 32366 9761
rect 32310 9687 32366 9696
rect 32036 9512 32088 9518
rect 32036 9454 32088 9460
rect 31944 8968 31996 8974
rect 31944 8910 31996 8916
rect 31852 8832 31904 8838
rect 31852 8774 31904 8780
rect 32404 8832 32456 8838
rect 32404 8774 32456 8780
rect 32416 8566 32444 8774
rect 32404 8560 32456 8566
rect 32404 8502 32456 8508
rect 32128 8288 32180 8294
rect 32128 8230 32180 8236
rect 32140 8090 32168 8230
rect 31760 8084 31812 8090
rect 31760 8026 31812 8032
rect 32128 8084 32180 8090
rect 32128 8026 32180 8032
rect 31300 7948 31352 7954
rect 31300 7890 31352 7896
rect 31576 7948 31628 7954
rect 31576 7890 31628 7896
rect 31024 7880 31076 7886
rect 31024 7822 31076 7828
rect 31944 7744 31996 7750
rect 31944 7686 31996 7692
rect 30656 7336 30708 7342
rect 30656 7278 30708 7284
rect 30564 6860 30616 6866
rect 30564 6802 30616 6808
rect 30288 5296 30340 5302
rect 30288 5238 30340 5244
rect 30300 4826 30328 5238
rect 30576 5166 30604 6802
rect 30668 6798 30696 7278
rect 30932 7200 30984 7206
rect 30932 7142 30984 7148
rect 30944 6866 30972 7142
rect 31852 6996 31904 7002
rect 31852 6938 31904 6944
rect 30932 6860 30984 6866
rect 30932 6802 30984 6808
rect 30656 6792 30708 6798
rect 30656 6734 30708 6740
rect 30668 6458 30696 6734
rect 31668 6656 31720 6662
rect 31668 6598 31720 6604
rect 30656 6452 30708 6458
rect 30656 6394 30708 6400
rect 30668 5710 30696 6394
rect 31116 6248 31168 6254
rect 31116 6190 31168 6196
rect 30656 5704 30708 5710
rect 30656 5646 30708 5652
rect 31128 5370 31156 6190
rect 31680 5710 31708 6598
rect 31864 6458 31892 6938
rect 31956 6730 31984 7686
rect 32036 6792 32088 6798
rect 32036 6734 32088 6740
rect 32220 6792 32272 6798
rect 32220 6734 32272 6740
rect 31944 6724 31996 6730
rect 31944 6666 31996 6672
rect 32048 6458 32076 6734
rect 31852 6452 31904 6458
rect 31852 6394 31904 6400
rect 32036 6452 32088 6458
rect 32036 6394 32088 6400
rect 32232 5778 32260 6734
rect 32692 6322 32720 12174
rect 32876 11762 32904 12406
rect 33048 11892 33100 11898
rect 33048 11834 33100 11840
rect 32864 11756 32916 11762
rect 32864 11698 32916 11704
rect 32876 11558 32904 11698
rect 32864 11552 32916 11558
rect 32864 11494 32916 11500
rect 32876 11393 32904 11494
rect 32862 11384 32918 11393
rect 32862 11319 32918 11328
rect 32864 11280 32916 11286
rect 32862 11248 32864 11257
rect 32916 11248 32918 11257
rect 32862 11183 32918 11192
rect 33060 10810 33088 11834
rect 33048 10804 33100 10810
rect 33048 10746 33100 10752
rect 33152 10742 33180 14282
rect 33520 14006 33548 15030
rect 33796 14618 33824 15302
rect 33968 15088 34020 15094
rect 33968 15030 34020 15036
rect 33784 14612 33836 14618
rect 33784 14554 33836 14560
rect 33508 14000 33560 14006
rect 33508 13942 33560 13948
rect 33520 13410 33548 13942
rect 33428 13382 33548 13410
rect 33428 12866 33456 13382
rect 33508 13320 33560 13326
rect 33508 13262 33560 13268
rect 33336 12850 33456 12866
rect 33520 12850 33548 13262
rect 33876 13252 33928 13258
rect 33876 13194 33928 13200
rect 33324 12844 33456 12850
rect 33376 12838 33456 12844
rect 33508 12844 33560 12850
rect 33324 12786 33376 12792
rect 33508 12786 33560 12792
rect 33600 12300 33652 12306
rect 33600 12242 33652 12248
rect 33508 12164 33560 12170
rect 33508 12106 33560 12112
rect 33232 11144 33284 11150
rect 33232 11086 33284 11092
rect 33140 10736 33192 10742
rect 33140 10678 33192 10684
rect 33244 9450 33272 11086
rect 33416 11076 33468 11082
rect 33416 11018 33468 11024
rect 33322 10160 33378 10169
rect 33322 10095 33324 10104
rect 33376 10095 33378 10104
rect 33324 10066 33376 10072
rect 33322 9616 33378 9625
rect 33322 9551 33378 9560
rect 33232 9444 33284 9450
rect 33232 9386 33284 9392
rect 33336 9330 33364 9551
rect 33244 9302 33364 9330
rect 33244 8974 33272 9302
rect 33428 8974 33456 11018
rect 33520 10062 33548 12106
rect 33612 11762 33640 12242
rect 33888 12170 33916 13194
rect 33980 13190 34008 15030
rect 34624 14385 34652 18566
rect 34716 18086 34744 19110
rect 34808 18902 34836 19314
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 34796 18896 34848 18902
rect 34796 18838 34848 18844
rect 35072 18760 35124 18766
rect 35072 18702 35124 18708
rect 35084 18630 35112 18702
rect 35072 18624 35124 18630
rect 35072 18566 35124 18572
rect 35348 18624 35400 18630
rect 35348 18566 35400 18572
rect 35360 18358 35388 18566
rect 35348 18352 35400 18358
rect 35348 18294 35400 18300
rect 34704 18080 34756 18086
rect 34704 18022 34756 18028
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 35452 17542 35480 22034
rect 35532 21956 35584 21962
rect 35532 21898 35584 21904
rect 35544 21078 35572 21898
rect 35532 21072 35584 21078
rect 35532 21014 35584 21020
rect 35636 20806 35664 22442
rect 35820 22234 35848 22714
rect 35912 22710 35940 23054
rect 35900 22704 35952 22710
rect 35900 22646 35952 22652
rect 35808 22228 35860 22234
rect 35808 22170 35860 22176
rect 35820 22094 35848 22170
rect 35728 22066 35848 22094
rect 35728 21457 35756 22066
rect 35714 21448 35770 21457
rect 35714 21383 35770 21392
rect 35716 21004 35768 21010
rect 35716 20946 35768 20952
rect 35624 20800 35676 20806
rect 35624 20742 35676 20748
rect 35728 20602 35756 20946
rect 35808 20868 35860 20874
rect 35808 20810 35860 20816
rect 35716 20596 35768 20602
rect 35716 20538 35768 20544
rect 35820 20380 35848 20810
rect 35912 20534 35940 22646
rect 35992 22160 36044 22166
rect 35992 22102 36044 22108
rect 36004 21690 36032 22102
rect 35992 21684 36044 21690
rect 35992 21626 36044 21632
rect 36096 20942 36124 23258
rect 36084 20936 36136 20942
rect 36084 20878 36136 20884
rect 35992 20800 36044 20806
rect 35992 20742 36044 20748
rect 35900 20528 35952 20534
rect 35900 20470 35952 20476
rect 36004 20380 36032 20742
rect 35820 20352 36032 20380
rect 35912 18426 35940 20352
rect 36084 19916 36136 19922
rect 36084 19858 36136 19864
rect 35992 19440 36044 19446
rect 35992 19382 36044 19388
rect 36004 18698 36032 19382
rect 35992 18692 36044 18698
rect 35992 18634 36044 18640
rect 35900 18420 35952 18426
rect 35900 18362 35952 18368
rect 36096 18290 36124 19858
rect 36280 19378 36308 24686
rect 38672 24206 38700 24686
rect 38948 24206 38976 24754
rect 38660 24200 38712 24206
rect 38660 24142 38712 24148
rect 38936 24200 38988 24206
rect 38936 24142 38988 24148
rect 37924 24132 37976 24138
rect 37924 24074 37976 24080
rect 36452 24064 36504 24070
rect 36452 24006 36504 24012
rect 36464 23730 36492 24006
rect 37936 23866 37964 24074
rect 37924 23860 37976 23866
rect 37924 23802 37976 23808
rect 36452 23724 36504 23730
rect 36452 23666 36504 23672
rect 37280 23724 37332 23730
rect 37280 23666 37332 23672
rect 37648 23724 37700 23730
rect 37648 23666 37700 23672
rect 36464 22098 36492 23666
rect 36912 23044 36964 23050
rect 36912 22986 36964 22992
rect 36924 22778 36952 22986
rect 36912 22772 36964 22778
rect 36912 22714 36964 22720
rect 36636 22432 36688 22438
rect 36636 22374 36688 22380
rect 36452 22092 36504 22098
rect 36452 22034 36504 22040
rect 36544 21888 36596 21894
rect 36544 21830 36596 21836
rect 36360 21344 36412 21350
rect 36360 21286 36412 21292
rect 36372 20641 36400 21286
rect 36556 21010 36584 21830
rect 36544 21004 36596 21010
rect 36544 20946 36596 20952
rect 36358 20632 36414 20641
rect 36358 20567 36414 20576
rect 36268 19372 36320 19378
rect 36268 19314 36320 19320
rect 36280 19174 36308 19314
rect 36268 19168 36320 19174
rect 36268 19110 36320 19116
rect 36268 18896 36320 18902
rect 36268 18838 36320 18844
rect 36084 18284 36136 18290
rect 36084 18226 36136 18232
rect 35440 17536 35492 17542
rect 35440 17478 35492 17484
rect 35624 17536 35676 17542
rect 35624 17478 35676 17484
rect 35716 17536 35768 17542
rect 35716 17478 35768 17484
rect 35348 17196 35400 17202
rect 35348 17138 35400 17144
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 35360 16794 35388 17138
rect 34704 16788 34756 16794
rect 34704 16730 34756 16736
rect 35348 16788 35400 16794
rect 35348 16730 35400 16736
rect 34716 16590 34744 16730
rect 35636 16658 35664 17478
rect 35728 17270 35756 17478
rect 35716 17264 35768 17270
rect 35716 17206 35768 17212
rect 35728 16794 35756 17206
rect 36096 17202 36124 18226
rect 36280 17542 36308 18838
rect 36452 18692 36504 18698
rect 36452 18634 36504 18640
rect 36464 18086 36492 18634
rect 36452 18080 36504 18086
rect 36452 18022 36504 18028
rect 36268 17536 36320 17542
rect 36268 17478 36320 17484
rect 36084 17196 36136 17202
rect 36084 17138 36136 17144
rect 36084 16992 36136 16998
rect 36084 16934 36136 16940
rect 35716 16788 35768 16794
rect 35716 16730 35768 16736
rect 35992 16788 36044 16794
rect 35992 16730 36044 16736
rect 35624 16652 35676 16658
rect 35624 16594 35676 16600
rect 34704 16584 34756 16590
rect 34704 16526 34756 16532
rect 35532 16584 35584 16590
rect 35532 16526 35584 16532
rect 34716 16046 34744 16526
rect 35072 16176 35124 16182
rect 35072 16118 35124 16124
rect 34888 16108 34940 16114
rect 34888 16050 34940 16056
rect 34704 16040 34756 16046
rect 34900 15994 34928 16050
rect 35084 16046 35112 16118
rect 35544 16114 35572 16526
rect 35636 16153 35664 16594
rect 35622 16144 35678 16153
rect 35532 16108 35584 16114
rect 36004 16114 36032 16730
rect 36096 16425 36124 16934
rect 36082 16416 36138 16425
rect 36082 16351 36138 16360
rect 35622 16079 35678 16088
rect 35808 16108 35860 16114
rect 35532 16050 35584 16056
rect 34704 15982 34756 15988
rect 34716 14958 34744 15982
rect 34808 15966 34928 15994
rect 35072 16040 35124 16046
rect 35072 15982 35124 15988
rect 35348 16040 35400 16046
rect 35348 15982 35400 15988
rect 35440 16040 35492 16046
rect 35440 15982 35492 15988
rect 34808 15434 34836 15966
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 35360 15586 35388 15982
rect 35268 15558 35388 15586
rect 34796 15428 34848 15434
rect 34796 15370 34848 15376
rect 34808 15026 34836 15370
rect 34796 15020 34848 15026
rect 34796 14962 34848 14968
rect 35268 14958 35296 15558
rect 35348 15496 35400 15502
rect 35348 15438 35400 15444
rect 34704 14952 34756 14958
rect 34704 14894 34756 14900
rect 35256 14952 35308 14958
rect 35256 14894 35308 14900
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 34610 14376 34666 14385
rect 34520 14340 34572 14346
rect 34610 14311 34666 14320
rect 34520 14282 34572 14288
rect 34532 14006 34560 14282
rect 34520 14000 34572 14006
rect 34520 13942 34572 13948
rect 34152 13320 34204 13326
rect 34152 13262 34204 13268
rect 33968 13184 34020 13190
rect 33968 13126 34020 13132
rect 34164 12850 34192 13262
rect 34152 12844 34204 12850
rect 34152 12786 34204 12792
rect 33876 12164 33928 12170
rect 33876 12106 33928 12112
rect 34532 11898 34560 13942
rect 34624 12850 34652 14311
rect 35360 13938 35388 15438
rect 35452 15162 35480 15982
rect 35440 15156 35492 15162
rect 35440 15098 35492 15104
rect 35636 15042 35664 16079
rect 35992 16108 36044 16114
rect 35860 16068 35940 16096
rect 35808 16050 35860 16056
rect 35636 15014 35756 15042
rect 35532 14952 35584 14958
rect 35532 14894 35584 14900
rect 35440 14476 35492 14482
rect 35440 14418 35492 14424
rect 34704 13932 34756 13938
rect 34704 13874 34756 13880
rect 35348 13932 35400 13938
rect 35348 13874 35400 13880
rect 34716 12986 34744 13874
rect 34796 13728 34848 13734
rect 34796 13670 34848 13676
rect 34808 13394 34836 13670
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 34980 13524 35032 13530
rect 34980 13466 35032 13472
rect 34796 13388 34848 13394
rect 34796 13330 34848 13336
rect 34992 13326 35020 13466
rect 34980 13320 35032 13326
rect 34980 13262 35032 13268
rect 35256 13184 35308 13190
rect 35256 13126 35308 13132
rect 34704 12980 34756 12986
rect 34704 12922 34756 12928
rect 35268 12918 35296 13126
rect 35256 12912 35308 12918
rect 35256 12854 35308 12860
rect 34612 12844 34664 12850
rect 34612 12786 34664 12792
rect 34796 12640 34848 12646
rect 34796 12582 34848 12588
rect 34808 12170 34836 12582
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 35360 12238 35388 13874
rect 35452 13530 35480 14418
rect 35544 14414 35572 14894
rect 35532 14408 35584 14414
rect 35532 14350 35584 14356
rect 35544 14113 35572 14350
rect 35530 14104 35586 14113
rect 35530 14039 35586 14048
rect 35624 13932 35676 13938
rect 35624 13874 35676 13880
rect 35636 13530 35664 13874
rect 35440 13524 35492 13530
rect 35440 13466 35492 13472
rect 35624 13524 35676 13530
rect 35624 13466 35676 13472
rect 35728 12730 35756 15014
rect 35808 13456 35860 13462
rect 35808 13398 35860 13404
rect 35452 12702 35756 12730
rect 35348 12232 35400 12238
rect 35348 12174 35400 12180
rect 34796 12164 34848 12170
rect 34796 12106 34848 12112
rect 34520 11892 34572 11898
rect 34520 11834 34572 11840
rect 35360 11830 35388 12174
rect 35348 11824 35400 11830
rect 35348 11766 35400 11772
rect 33600 11756 33652 11762
rect 33600 11698 33652 11704
rect 34796 11756 34848 11762
rect 34796 11698 34848 11704
rect 33612 11218 33640 11698
rect 34520 11688 34572 11694
rect 34520 11630 34572 11636
rect 33600 11212 33652 11218
rect 33600 11154 33652 11160
rect 34428 11212 34480 11218
rect 34428 11154 34480 11160
rect 33968 11144 34020 11150
rect 33968 11086 34020 11092
rect 33600 10668 33652 10674
rect 33600 10610 33652 10616
rect 33508 10056 33560 10062
rect 33508 9998 33560 10004
rect 33508 9580 33560 9586
rect 33508 9522 33560 9528
rect 33520 9042 33548 9522
rect 33508 9036 33560 9042
rect 33508 8978 33560 8984
rect 33232 8968 33284 8974
rect 33232 8910 33284 8916
rect 33416 8968 33468 8974
rect 33416 8910 33468 8916
rect 33048 8832 33100 8838
rect 33048 8774 33100 8780
rect 33060 7886 33088 8774
rect 33048 7880 33100 7886
rect 33048 7822 33100 7828
rect 33244 7546 33272 8910
rect 33612 8498 33640 10610
rect 33784 10600 33836 10606
rect 33784 10542 33836 10548
rect 33692 10124 33744 10130
rect 33692 10066 33744 10072
rect 33704 9654 33732 10066
rect 33796 10062 33824 10542
rect 33784 10056 33836 10062
rect 33784 9998 33836 10004
rect 33876 9920 33928 9926
rect 33876 9862 33928 9868
rect 33692 9648 33744 9654
rect 33692 9590 33744 9596
rect 33888 9586 33916 9862
rect 33876 9580 33928 9586
rect 33876 9522 33928 9528
rect 33888 8974 33916 9522
rect 33876 8968 33928 8974
rect 33876 8910 33928 8916
rect 33980 8514 34008 11086
rect 34244 10464 34296 10470
rect 34244 10406 34296 10412
rect 34256 9586 34284 10406
rect 34440 9722 34468 11154
rect 34428 9716 34480 9722
rect 34428 9658 34480 9664
rect 34440 9586 34468 9658
rect 34244 9580 34296 9586
rect 34244 9522 34296 9528
rect 34428 9580 34480 9586
rect 34428 9522 34480 9528
rect 34060 8832 34112 8838
rect 34060 8774 34112 8780
rect 34072 8634 34100 8774
rect 34060 8628 34112 8634
rect 34060 8570 34112 8576
rect 33600 8492 33652 8498
rect 33600 8434 33652 8440
rect 33704 8486 34100 8514
rect 33508 8424 33560 8430
rect 33508 8366 33560 8372
rect 33520 8090 33548 8366
rect 33508 8084 33560 8090
rect 33508 8026 33560 8032
rect 33232 7540 33284 7546
rect 33232 7482 33284 7488
rect 33704 6390 33732 8486
rect 34072 8294 34100 8486
rect 34152 8492 34204 8498
rect 34152 8434 34204 8440
rect 34060 8288 34112 8294
rect 34060 8230 34112 8236
rect 34164 8090 34192 8434
rect 34256 8294 34284 9522
rect 34532 8906 34560 11630
rect 34612 11076 34664 11082
rect 34612 11018 34664 11024
rect 34520 8900 34572 8906
rect 34520 8842 34572 8848
rect 34624 8634 34652 11018
rect 34704 11008 34756 11014
rect 34704 10950 34756 10956
rect 34716 10742 34744 10950
rect 34704 10736 34756 10742
rect 34704 10678 34756 10684
rect 34808 10674 34836 11698
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 34978 11248 35034 11257
rect 35452 11234 35480 12702
rect 35820 12238 35848 13398
rect 35912 12918 35940 16068
rect 35992 16050 36044 16056
rect 36096 15194 36124 16351
rect 36464 16250 36492 18022
rect 36452 16244 36504 16250
rect 36452 16186 36504 16192
rect 36176 15904 36228 15910
rect 36176 15846 36228 15852
rect 36188 15502 36216 15846
rect 36176 15496 36228 15502
rect 36176 15438 36228 15444
rect 36004 15166 36124 15194
rect 35900 12912 35952 12918
rect 35900 12854 35952 12860
rect 35808 12232 35860 12238
rect 35808 12174 35860 12180
rect 35622 11928 35678 11937
rect 35622 11863 35624 11872
rect 35676 11863 35678 11872
rect 35624 11834 35676 11840
rect 35808 11824 35860 11830
rect 35808 11766 35860 11772
rect 34978 11183 35034 11192
rect 35360 11206 35480 11234
rect 34992 11150 35020 11183
rect 34980 11144 35032 11150
rect 34980 11086 35032 11092
rect 35164 11144 35216 11150
rect 35164 11086 35216 11092
rect 35176 10810 35204 11086
rect 35164 10804 35216 10810
rect 35164 10746 35216 10752
rect 34796 10668 34848 10674
rect 34796 10610 34848 10616
rect 34808 10266 34836 10610
rect 35360 10470 35388 11206
rect 35820 11150 35848 11766
rect 35808 11144 35860 11150
rect 35808 11086 35860 11092
rect 35440 11076 35492 11082
rect 35440 11018 35492 11024
rect 35348 10464 35400 10470
rect 35348 10406 35400 10412
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 34796 10260 34848 10266
rect 34796 10202 34848 10208
rect 34704 10056 34756 10062
rect 34704 9998 34756 10004
rect 34612 8628 34664 8634
rect 34612 8570 34664 8576
rect 34716 8566 34744 9998
rect 34796 9988 34848 9994
rect 34796 9930 34848 9936
rect 34704 8560 34756 8566
rect 34704 8502 34756 8508
rect 34244 8288 34296 8294
rect 34244 8230 34296 8236
rect 34152 8084 34204 8090
rect 34152 8026 34204 8032
rect 34520 8016 34572 8022
rect 34520 7958 34572 7964
rect 34532 7478 34560 7958
rect 34808 7750 34836 9930
rect 35072 9920 35124 9926
rect 35072 9862 35124 9868
rect 35084 9654 35112 9862
rect 35452 9654 35480 11018
rect 35820 10656 35848 11086
rect 35900 10668 35952 10674
rect 35820 10628 35900 10656
rect 35900 10610 35952 10616
rect 35808 10260 35860 10266
rect 36004 10248 36032 15166
rect 36648 15162 36676 22374
rect 37292 21962 37320 23666
rect 37464 23588 37516 23594
rect 37464 23530 37516 23536
rect 37372 22976 37424 22982
rect 37372 22918 37424 22924
rect 37384 22030 37412 22918
rect 37476 22030 37504 23530
rect 37660 23322 37688 23666
rect 37648 23316 37700 23322
rect 37648 23258 37700 23264
rect 38672 23118 38700 24142
rect 38660 23112 38712 23118
rect 38660 23054 38712 23060
rect 38672 22710 38700 23054
rect 38660 22704 38712 22710
rect 38660 22646 38712 22652
rect 38752 22636 38804 22642
rect 38752 22578 38804 22584
rect 38764 22098 38792 22578
rect 38752 22092 38804 22098
rect 38752 22034 38804 22040
rect 37372 22024 37424 22030
rect 37372 21966 37424 21972
rect 37464 22024 37516 22030
rect 37464 21966 37516 21972
rect 38384 22024 38436 22030
rect 38384 21966 38436 21972
rect 37280 21956 37332 21962
rect 37280 21898 37332 21904
rect 37292 21486 37320 21898
rect 37476 21554 37504 21966
rect 38200 21956 38252 21962
rect 38200 21898 38252 21904
rect 38212 21690 38240 21898
rect 38200 21684 38252 21690
rect 38200 21626 38252 21632
rect 37464 21548 37516 21554
rect 37464 21490 37516 21496
rect 37740 21548 37792 21554
rect 37740 21490 37792 21496
rect 37280 21480 37332 21486
rect 37280 21422 37332 21428
rect 37752 21146 37780 21490
rect 37832 21344 37884 21350
rect 37832 21286 37884 21292
rect 37740 21140 37792 21146
rect 37740 21082 37792 21088
rect 37648 20392 37700 20398
rect 37648 20334 37700 20340
rect 37372 20324 37424 20330
rect 37372 20266 37424 20272
rect 36728 19848 36780 19854
rect 36728 19790 36780 19796
rect 36740 18766 36768 19790
rect 37096 19780 37148 19786
rect 37096 19722 37148 19728
rect 37108 19514 37136 19722
rect 37384 19553 37412 20266
rect 37556 19848 37608 19854
rect 37556 19790 37608 19796
rect 37370 19544 37426 19553
rect 37096 19508 37148 19514
rect 37370 19479 37426 19488
rect 37096 19450 37148 19456
rect 36820 19440 36872 19446
rect 36820 19382 36872 19388
rect 36728 18760 36780 18766
rect 36728 18702 36780 18708
rect 36740 18290 36768 18702
rect 36728 18284 36780 18290
rect 36728 18226 36780 18232
rect 36636 15156 36688 15162
rect 36636 15098 36688 15104
rect 36648 13530 36676 15098
rect 36636 13524 36688 13530
rect 36636 13466 36688 13472
rect 36728 12844 36780 12850
rect 36728 12786 36780 12792
rect 36084 12776 36136 12782
rect 36084 12718 36136 12724
rect 36096 12442 36124 12718
rect 36084 12436 36136 12442
rect 36740 12434 36768 12786
rect 36084 12378 36136 12384
rect 36648 12406 36768 12434
rect 36648 11626 36676 12406
rect 36832 12322 36860 19382
rect 37384 19378 37412 19479
rect 37372 19372 37424 19378
rect 37372 19314 37424 19320
rect 37004 19168 37056 19174
rect 37004 19110 37056 19116
rect 37016 18766 37044 19110
rect 37568 18766 37596 19790
rect 37660 18970 37688 20334
rect 37740 20256 37792 20262
rect 37844 20244 37872 21286
rect 38016 21140 38068 21146
rect 38016 21082 38068 21088
rect 37924 20460 37976 20466
rect 37924 20402 37976 20408
rect 37792 20216 37872 20244
rect 37740 20198 37792 20204
rect 37752 19990 37780 20198
rect 37936 20058 37964 20402
rect 37924 20052 37976 20058
rect 37924 19994 37976 20000
rect 37740 19984 37792 19990
rect 37740 19926 37792 19932
rect 37648 18964 37700 18970
rect 37648 18906 37700 18912
rect 37004 18760 37056 18766
rect 37004 18702 37056 18708
rect 37556 18760 37608 18766
rect 37556 18702 37608 18708
rect 37568 18358 37596 18702
rect 37648 18624 37700 18630
rect 37648 18566 37700 18572
rect 37556 18352 37608 18358
rect 37556 18294 37608 18300
rect 37660 18290 37688 18566
rect 37648 18284 37700 18290
rect 37648 18226 37700 18232
rect 37752 18086 37780 19926
rect 37832 18284 37884 18290
rect 37832 18226 37884 18232
rect 37740 18080 37792 18086
rect 37740 18022 37792 18028
rect 37844 17762 37872 18226
rect 37752 17734 37872 17762
rect 37752 17678 37780 17734
rect 37740 17672 37792 17678
rect 37740 17614 37792 17620
rect 37648 17604 37700 17610
rect 37648 17546 37700 17552
rect 37188 17536 37240 17542
rect 37188 17478 37240 17484
rect 37464 17536 37516 17542
rect 37464 17478 37516 17484
rect 37200 16522 37228 17478
rect 37476 17202 37504 17478
rect 37280 17196 37332 17202
rect 37280 17138 37332 17144
rect 37464 17196 37516 17202
rect 37464 17138 37516 17144
rect 37556 17196 37608 17202
rect 37556 17138 37608 17144
rect 37292 16590 37320 17138
rect 37280 16584 37332 16590
rect 37280 16526 37332 16532
rect 37188 16516 37240 16522
rect 37188 16458 37240 16464
rect 37568 16454 37596 17138
rect 37372 16448 37424 16454
rect 37372 16390 37424 16396
rect 37556 16448 37608 16454
rect 37556 16390 37608 16396
rect 36912 15700 36964 15706
rect 36912 15642 36964 15648
rect 36924 15094 36952 15642
rect 37384 15094 37412 16390
rect 37660 16114 37688 17546
rect 37752 17338 37780 17614
rect 37832 17604 37884 17610
rect 37832 17546 37884 17552
rect 37844 17338 37872 17546
rect 37740 17332 37792 17338
rect 37740 17274 37792 17280
rect 37832 17332 37884 17338
rect 37832 17274 37884 17280
rect 37648 16108 37700 16114
rect 37648 16050 37700 16056
rect 37464 15904 37516 15910
rect 37464 15846 37516 15852
rect 36912 15088 36964 15094
rect 36912 15030 36964 15036
rect 37372 15088 37424 15094
rect 37372 15030 37424 15036
rect 37476 15026 37504 15846
rect 37660 15434 37688 16050
rect 37648 15428 37700 15434
rect 37648 15370 37700 15376
rect 37464 15020 37516 15026
rect 37464 14962 37516 14968
rect 37096 14816 37148 14822
rect 37096 14758 37148 14764
rect 37108 14346 37136 14758
rect 37752 14550 37780 17274
rect 37844 16726 37872 17274
rect 37832 16720 37884 16726
rect 37832 16662 37884 16668
rect 37924 16448 37976 16454
rect 37924 16390 37976 16396
rect 37936 16182 37964 16390
rect 37924 16176 37976 16182
rect 37924 16118 37976 16124
rect 37924 16040 37976 16046
rect 37924 15982 37976 15988
rect 37936 15366 37964 15982
rect 37924 15360 37976 15366
rect 37924 15302 37976 15308
rect 37936 14890 37964 15302
rect 37924 14884 37976 14890
rect 37924 14826 37976 14832
rect 37740 14544 37792 14550
rect 37740 14486 37792 14492
rect 37648 14408 37700 14414
rect 37648 14350 37700 14356
rect 36912 14340 36964 14346
rect 36912 14282 36964 14288
rect 37096 14340 37148 14346
rect 37096 14282 37148 14288
rect 36924 13326 36952 14282
rect 37108 14249 37136 14282
rect 37094 14240 37150 14249
rect 37094 14175 37150 14184
rect 37372 14068 37424 14074
rect 37372 14010 37424 14016
rect 37004 13524 37056 13530
rect 37004 13466 37056 13472
rect 36912 13320 36964 13326
rect 36912 13262 36964 13268
rect 36740 12294 36860 12322
rect 36636 11620 36688 11626
rect 36636 11562 36688 11568
rect 36084 11280 36136 11286
rect 36084 11222 36136 11228
rect 36096 11082 36124 11222
rect 36084 11076 36136 11082
rect 36084 11018 36136 11024
rect 36360 11076 36412 11082
rect 36360 11018 36412 11024
rect 36096 10985 36124 11018
rect 36082 10976 36138 10985
rect 36082 10911 36138 10920
rect 36372 10470 36400 11018
rect 36648 10674 36676 11562
rect 36636 10668 36688 10674
rect 36636 10610 36688 10616
rect 36360 10464 36412 10470
rect 36360 10406 36412 10412
rect 35860 10220 36032 10248
rect 35808 10202 35860 10208
rect 35072 9648 35124 9654
rect 35072 9590 35124 9596
rect 35440 9648 35492 9654
rect 35440 9590 35492 9596
rect 35820 9586 35848 10202
rect 36372 9586 36400 10406
rect 35164 9580 35216 9586
rect 35164 9522 35216 9528
rect 35808 9580 35860 9586
rect 35808 9522 35860 9528
rect 36360 9580 36412 9586
rect 36360 9522 36412 9528
rect 35176 9466 35204 9522
rect 35716 9512 35768 9518
rect 35176 9438 35388 9466
rect 35716 9454 35768 9460
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 35360 8634 35388 9438
rect 35532 9376 35584 9382
rect 35532 9318 35584 9324
rect 35348 8628 35400 8634
rect 35348 8570 35400 8576
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 34796 7744 34848 7750
rect 34796 7686 34848 7692
rect 34808 7546 34836 7686
rect 34796 7540 34848 7546
rect 34796 7482 34848 7488
rect 34520 7472 34572 7478
rect 34520 7414 34572 7420
rect 33784 6656 33836 6662
rect 33784 6598 33836 6604
rect 33692 6384 33744 6390
rect 33692 6326 33744 6332
rect 32680 6316 32732 6322
rect 32680 6258 32732 6264
rect 32956 6316 33008 6322
rect 32956 6258 33008 6264
rect 32772 5840 32824 5846
rect 32772 5782 32824 5788
rect 32220 5772 32272 5778
rect 32220 5714 32272 5720
rect 31668 5704 31720 5710
rect 31668 5646 31720 5652
rect 32588 5704 32640 5710
rect 32588 5646 32640 5652
rect 31116 5364 31168 5370
rect 31116 5306 31168 5312
rect 30564 5160 30616 5166
rect 30564 5102 30616 5108
rect 30288 4820 30340 4826
rect 30288 4762 30340 4768
rect 30288 4480 30340 4486
rect 30288 4422 30340 4428
rect 30300 4146 30328 4422
rect 30576 4214 30604 5102
rect 32128 4752 32180 4758
rect 32128 4694 32180 4700
rect 32140 4282 32168 4694
rect 32600 4622 32628 5646
rect 32784 5574 32812 5782
rect 32864 5704 32916 5710
rect 32864 5646 32916 5652
rect 32968 5658 32996 6258
rect 33048 6248 33100 6254
rect 33048 6190 33100 6196
rect 33060 5914 33088 6190
rect 33232 6112 33284 6118
rect 33232 6054 33284 6060
rect 33048 5908 33100 5914
rect 33048 5850 33100 5856
rect 33140 5704 33192 5710
rect 32968 5652 33140 5658
rect 32968 5646 33192 5652
rect 32876 5574 32904 5646
rect 32968 5630 33180 5646
rect 32772 5568 32824 5574
rect 32772 5510 32824 5516
rect 32864 5568 32916 5574
rect 32864 5510 32916 5516
rect 33244 5234 33272 6054
rect 33704 5778 33732 6326
rect 33796 6322 33824 6598
rect 33784 6316 33836 6322
rect 33784 6258 33836 6264
rect 34532 6254 34560 7414
rect 35544 7410 35572 9318
rect 35728 9110 35756 9454
rect 35820 9110 35848 9522
rect 36372 9178 36400 9522
rect 36360 9172 36412 9178
rect 36360 9114 36412 9120
rect 35716 9104 35768 9110
rect 35716 9046 35768 9052
rect 35808 9104 35860 9110
rect 35808 9046 35860 9052
rect 35716 8900 35768 8906
rect 35716 8842 35768 8848
rect 35728 7886 35756 8842
rect 36372 8566 36400 9114
rect 36360 8560 36412 8566
rect 36360 8502 36412 8508
rect 36542 8528 36598 8537
rect 36542 8463 36544 8472
rect 36596 8463 36598 8472
rect 36544 8434 36596 8440
rect 35808 8424 35860 8430
rect 35808 8366 35860 8372
rect 35820 8090 35848 8366
rect 35808 8084 35860 8090
rect 35808 8026 35860 8032
rect 35716 7880 35768 7886
rect 35716 7822 35768 7828
rect 35728 7478 35756 7822
rect 35716 7472 35768 7478
rect 35716 7414 35768 7420
rect 35532 7404 35584 7410
rect 35532 7346 35584 7352
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 34796 6792 34848 6798
rect 34796 6734 34848 6740
rect 34520 6248 34572 6254
rect 34520 6190 34572 6196
rect 33692 5772 33744 5778
rect 33692 5714 33744 5720
rect 34060 5704 34112 5710
rect 34060 5646 34112 5652
rect 34072 5574 34100 5646
rect 34060 5568 34112 5574
rect 34060 5510 34112 5516
rect 33232 5228 33284 5234
rect 33232 5170 33284 5176
rect 34532 4622 34560 6190
rect 34704 5568 34756 5574
rect 34704 5510 34756 5516
rect 34716 5234 34744 5510
rect 34808 5370 34836 6734
rect 36740 6390 36768 12294
rect 37016 12238 37044 13466
rect 37384 12646 37412 14010
rect 37660 13938 37688 14350
rect 37832 14272 37884 14278
rect 37832 14214 37884 14220
rect 37648 13932 37700 13938
rect 37648 13874 37700 13880
rect 37844 13920 37872 14214
rect 37924 13932 37976 13938
rect 37844 13892 37924 13920
rect 37740 13796 37792 13802
rect 37740 13738 37792 13744
rect 37752 13530 37780 13738
rect 37740 13524 37792 13530
rect 37740 13466 37792 13472
rect 37648 13252 37700 13258
rect 37648 13194 37700 13200
rect 37660 12850 37688 13194
rect 37844 12986 37872 13892
rect 37924 13874 37976 13880
rect 38028 12986 38056 21082
rect 38292 20936 38344 20942
rect 38292 20878 38344 20884
rect 38304 20602 38332 20878
rect 38292 20596 38344 20602
rect 38292 20538 38344 20544
rect 38108 20528 38160 20534
rect 38396 20505 38424 21966
rect 38108 20470 38160 20476
rect 38382 20496 38438 20505
rect 38120 15706 38148 20470
rect 38382 20431 38438 20440
rect 38200 19848 38252 19854
rect 38200 19790 38252 19796
rect 38212 19242 38240 19790
rect 38292 19780 38344 19786
rect 38292 19722 38344 19728
rect 38304 19378 38332 19722
rect 38292 19372 38344 19378
rect 38292 19314 38344 19320
rect 38200 19236 38252 19242
rect 38200 19178 38252 19184
rect 38108 15700 38160 15706
rect 38108 15642 38160 15648
rect 38212 13938 38240 19178
rect 38304 18970 38332 19314
rect 38292 18964 38344 18970
rect 38292 18906 38344 18912
rect 38396 18850 38424 20431
rect 38844 20392 38896 20398
rect 38844 20334 38896 20340
rect 38856 19922 38884 20334
rect 38844 19916 38896 19922
rect 38844 19858 38896 19864
rect 38304 18822 38424 18850
rect 38304 16794 38332 18822
rect 38752 18760 38804 18766
rect 38856 18748 38884 19858
rect 38804 18720 38884 18748
rect 38752 18702 38804 18708
rect 38856 18290 38884 18720
rect 38844 18284 38896 18290
rect 38844 18226 38896 18232
rect 38856 17202 38884 18226
rect 38844 17196 38896 17202
rect 38764 17156 38844 17184
rect 38292 16788 38344 16794
rect 38292 16730 38344 16736
rect 38200 13932 38252 13938
rect 38200 13874 38252 13880
rect 38212 13530 38240 13874
rect 38200 13524 38252 13530
rect 38200 13466 38252 13472
rect 37832 12980 37884 12986
rect 37832 12922 37884 12928
rect 38016 12980 38068 12986
rect 38016 12922 38068 12928
rect 37648 12844 37700 12850
rect 37648 12786 37700 12792
rect 37832 12844 37884 12850
rect 37832 12786 37884 12792
rect 37372 12640 37424 12646
rect 37372 12582 37424 12588
rect 36820 12232 36872 12238
rect 36820 12174 36872 12180
rect 37004 12232 37056 12238
rect 37004 12174 37056 12180
rect 37556 12232 37608 12238
rect 37556 12174 37608 12180
rect 36832 11354 36860 12174
rect 36912 11552 36964 11558
rect 36912 11494 36964 11500
rect 36820 11348 36872 11354
rect 36820 11290 36872 11296
rect 36924 11082 36952 11494
rect 37016 11257 37044 12174
rect 37280 12096 37332 12102
rect 37280 12038 37332 12044
rect 37002 11248 37058 11257
rect 37002 11183 37058 11192
rect 37292 11082 37320 12038
rect 37568 11762 37596 12174
rect 37556 11756 37608 11762
rect 37556 11698 37608 11704
rect 37372 11212 37424 11218
rect 37372 11154 37424 11160
rect 36912 11076 36964 11082
rect 36912 11018 36964 11024
rect 37280 11076 37332 11082
rect 37280 11018 37332 11024
rect 37188 10668 37240 10674
rect 37188 10610 37240 10616
rect 37200 9994 37228 10610
rect 37384 10554 37412 11154
rect 37292 10526 37412 10554
rect 37292 10062 37320 10526
rect 37568 10130 37596 11698
rect 37844 11558 37872 12786
rect 37924 12164 37976 12170
rect 37924 12106 37976 12112
rect 37832 11552 37884 11558
rect 37832 11494 37884 11500
rect 37936 10674 37964 12106
rect 37924 10668 37976 10674
rect 37924 10610 37976 10616
rect 37556 10124 37608 10130
rect 37556 10066 37608 10072
rect 37280 10056 37332 10062
rect 37280 9998 37332 10004
rect 37188 9988 37240 9994
rect 37188 9930 37240 9936
rect 37568 9586 37596 10066
rect 37936 9648 37964 10610
rect 38200 9920 38252 9926
rect 38304 9908 38332 16730
rect 38764 16114 38792 17156
rect 38844 17138 38896 17144
rect 38752 16108 38804 16114
rect 38752 16050 38804 16056
rect 39304 15496 39356 15502
rect 39304 15438 39356 15444
rect 38660 15428 38712 15434
rect 38660 15370 38712 15376
rect 38672 15162 38700 15370
rect 38660 15156 38712 15162
rect 38660 15098 38712 15104
rect 38384 15020 38436 15026
rect 38384 14962 38436 14968
rect 38396 14618 38424 14962
rect 39316 14822 39344 15438
rect 39304 14816 39356 14822
rect 39304 14758 39356 14764
rect 38384 14612 38436 14618
rect 38384 14554 38436 14560
rect 38384 12640 38436 12646
rect 38384 12582 38436 12588
rect 38660 12640 38712 12646
rect 38660 12582 38712 12588
rect 38396 12238 38424 12582
rect 38672 12306 38700 12582
rect 38660 12300 38712 12306
rect 38660 12242 38712 12248
rect 38384 12232 38436 12238
rect 38384 12174 38436 12180
rect 39028 12232 39080 12238
rect 39028 12174 39080 12180
rect 38252 9880 38332 9908
rect 38200 9862 38252 9868
rect 37936 9586 37967 9648
rect 38212 9586 38240 9862
rect 38396 9625 38424 12174
rect 39040 11150 39068 12174
rect 39028 11144 39080 11150
rect 39028 11086 39080 11092
rect 39040 10674 39068 11086
rect 39028 10668 39080 10674
rect 39028 10610 39080 10616
rect 39120 10668 39172 10674
rect 39120 10610 39172 10616
rect 39132 10266 39160 10610
rect 39120 10260 39172 10266
rect 39120 10202 39172 10208
rect 39304 9920 39356 9926
rect 39304 9862 39356 9868
rect 38382 9616 38438 9625
rect 37188 9580 37240 9586
rect 37188 9522 37240 9528
rect 37556 9580 37608 9586
rect 37556 9522 37608 9528
rect 37927 9580 37979 9586
rect 37927 9522 37979 9528
rect 38200 9580 38252 9586
rect 38382 9551 38438 9560
rect 38200 9522 38252 9528
rect 37096 9376 37148 9382
rect 37096 9318 37148 9324
rect 37108 7818 37136 9318
rect 37200 8974 37228 9522
rect 37188 8968 37240 8974
rect 37188 8910 37240 8916
rect 37372 8968 37424 8974
rect 37372 8910 37424 8916
rect 37200 8498 37228 8910
rect 37384 8634 37412 8910
rect 37936 8906 37964 9522
rect 38568 9512 38620 9518
rect 38568 9454 38620 9460
rect 38200 9036 38252 9042
rect 38200 8978 38252 8984
rect 37924 8900 37976 8906
rect 37844 8860 37924 8888
rect 37372 8628 37424 8634
rect 37372 8570 37424 8576
rect 37188 8492 37240 8498
rect 37760 8492 37812 8498
rect 37188 8434 37240 8440
rect 37752 8440 37760 8480
rect 37752 8434 37812 8440
rect 37752 8294 37780 8434
rect 37844 8362 37872 8860
rect 37924 8842 37976 8848
rect 38212 8566 38240 8978
rect 38200 8560 38252 8566
rect 38014 8528 38070 8537
rect 38200 8502 38252 8508
rect 38014 8463 38016 8472
rect 38068 8463 38070 8472
rect 38016 8434 38068 8440
rect 38580 8430 38608 9454
rect 39316 8906 39344 9862
rect 39304 8900 39356 8906
rect 39304 8842 39356 8848
rect 38660 8832 38712 8838
rect 38660 8774 38712 8780
rect 38672 8634 38700 8774
rect 38660 8628 38712 8634
rect 38660 8570 38712 8576
rect 37924 8424 37976 8430
rect 37924 8366 37976 8372
rect 38568 8424 38620 8430
rect 38568 8366 38620 8372
rect 37832 8356 37884 8362
rect 37832 8298 37884 8304
rect 37740 8288 37792 8294
rect 37740 8230 37792 8236
rect 37096 7812 37148 7818
rect 37096 7754 37148 7760
rect 37752 7546 37780 8230
rect 37936 7886 37964 8366
rect 38016 8288 38068 8294
rect 38016 8230 38068 8236
rect 38028 7886 38056 8230
rect 39316 8090 39344 8842
rect 39304 8084 39356 8090
rect 39304 8026 39356 8032
rect 37924 7880 37976 7886
rect 37924 7822 37976 7828
rect 38016 7880 38068 7886
rect 38016 7822 38068 7828
rect 37740 7540 37792 7546
rect 37740 7482 37792 7488
rect 36728 6384 36780 6390
rect 36728 6326 36780 6332
rect 39408 6322 39436 31726
rect 50294 31580 50602 31589
rect 50294 31578 50300 31580
rect 50356 31578 50380 31580
rect 50436 31578 50460 31580
rect 50516 31578 50540 31580
rect 50596 31578 50602 31580
rect 50356 31526 50358 31578
rect 50538 31526 50540 31578
rect 50294 31524 50300 31526
rect 50356 31524 50380 31526
rect 50436 31524 50460 31526
rect 50516 31524 50540 31526
rect 50596 31524 50602 31526
rect 50294 31515 50602 31524
rect 50294 30492 50602 30501
rect 50294 30490 50300 30492
rect 50356 30490 50380 30492
rect 50436 30490 50460 30492
rect 50516 30490 50540 30492
rect 50596 30490 50602 30492
rect 50356 30438 50358 30490
rect 50538 30438 50540 30490
rect 50294 30436 50300 30438
rect 50356 30436 50380 30438
rect 50436 30436 50460 30438
rect 50516 30436 50540 30438
rect 50596 30436 50602 30438
rect 50294 30427 50602 30436
rect 50294 29404 50602 29413
rect 50294 29402 50300 29404
rect 50356 29402 50380 29404
rect 50436 29402 50460 29404
rect 50516 29402 50540 29404
rect 50596 29402 50602 29404
rect 50356 29350 50358 29402
rect 50538 29350 50540 29402
rect 50294 29348 50300 29350
rect 50356 29348 50380 29350
rect 50436 29348 50460 29350
rect 50516 29348 50540 29350
rect 50596 29348 50602 29350
rect 50294 29339 50602 29348
rect 50294 28316 50602 28325
rect 50294 28314 50300 28316
rect 50356 28314 50380 28316
rect 50436 28314 50460 28316
rect 50516 28314 50540 28316
rect 50596 28314 50602 28316
rect 50356 28262 50358 28314
rect 50538 28262 50540 28314
rect 50294 28260 50300 28262
rect 50356 28260 50380 28262
rect 50436 28260 50460 28262
rect 50516 28260 50540 28262
rect 50596 28260 50602 28262
rect 50294 28251 50602 28260
rect 50294 27228 50602 27237
rect 50294 27226 50300 27228
rect 50356 27226 50380 27228
rect 50436 27226 50460 27228
rect 50516 27226 50540 27228
rect 50596 27226 50602 27228
rect 50356 27174 50358 27226
rect 50538 27174 50540 27226
rect 50294 27172 50300 27174
rect 50356 27172 50380 27174
rect 50436 27172 50460 27174
rect 50516 27172 50540 27174
rect 50596 27172 50602 27174
rect 50294 27163 50602 27172
rect 50294 26140 50602 26149
rect 50294 26138 50300 26140
rect 50356 26138 50380 26140
rect 50436 26138 50460 26140
rect 50516 26138 50540 26140
rect 50596 26138 50602 26140
rect 50356 26086 50358 26138
rect 50538 26086 50540 26138
rect 50294 26084 50300 26086
rect 50356 26084 50380 26086
rect 50436 26084 50460 26086
rect 50516 26084 50540 26086
rect 50596 26084 50602 26086
rect 50294 26075 50602 26084
rect 50294 25052 50602 25061
rect 50294 25050 50300 25052
rect 50356 25050 50380 25052
rect 50436 25050 50460 25052
rect 50516 25050 50540 25052
rect 50596 25050 50602 25052
rect 50356 24998 50358 25050
rect 50538 24998 50540 25050
rect 50294 24996 50300 24998
rect 50356 24996 50380 24998
rect 50436 24996 50460 24998
rect 50516 24996 50540 24998
rect 50596 24996 50602 24998
rect 50294 24987 50602 24996
rect 39948 24880 40000 24886
rect 39948 24822 40000 24828
rect 39960 24410 39988 24822
rect 43260 24812 43312 24818
rect 43260 24754 43312 24760
rect 41788 24744 41840 24750
rect 41788 24686 41840 24692
rect 42892 24744 42944 24750
rect 42892 24686 42944 24692
rect 41144 24608 41196 24614
rect 41144 24550 41196 24556
rect 39948 24404 40000 24410
rect 39948 24346 40000 24352
rect 41156 24206 41184 24550
rect 41800 24410 41828 24686
rect 41788 24404 41840 24410
rect 41788 24346 41840 24352
rect 42904 24206 42932 24686
rect 43272 24410 43300 24754
rect 56336 24614 56364 57190
rect 65654 57148 65962 57157
rect 65654 57146 65660 57148
rect 65716 57146 65740 57148
rect 65796 57146 65820 57148
rect 65876 57146 65900 57148
rect 65956 57146 65962 57148
rect 65716 57094 65718 57146
rect 65898 57094 65900 57146
rect 65654 57092 65660 57094
rect 65716 57092 65740 57094
rect 65796 57092 65820 57094
rect 65876 57092 65900 57094
rect 65956 57092 65962 57094
rect 65654 57083 65962 57092
rect 67640 56160 67692 56166
rect 67638 56128 67640 56137
rect 67692 56128 67694 56137
rect 65654 56060 65962 56069
rect 67638 56063 67694 56072
rect 65654 56058 65660 56060
rect 65716 56058 65740 56060
rect 65796 56058 65820 56060
rect 65876 56058 65900 56060
rect 65956 56058 65962 56060
rect 65716 56006 65718 56058
rect 65898 56006 65900 56058
rect 65654 56004 65660 56006
rect 65716 56004 65740 56006
rect 65796 56004 65820 56006
rect 65876 56004 65900 56006
rect 65956 56004 65962 56006
rect 65654 55995 65962 56004
rect 65654 54972 65962 54981
rect 65654 54970 65660 54972
rect 65716 54970 65740 54972
rect 65796 54970 65820 54972
rect 65876 54970 65900 54972
rect 65956 54970 65962 54972
rect 65716 54918 65718 54970
rect 65898 54918 65900 54970
rect 65654 54916 65660 54918
rect 65716 54916 65740 54918
rect 65796 54916 65820 54918
rect 65876 54916 65900 54918
rect 65956 54916 65962 54918
rect 65654 54907 65962 54916
rect 68100 54664 68152 54670
rect 68098 54632 68100 54641
rect 68152 54632 68154 54641
rect 68098 54567 68154 54576
rect 65654 53884 65962 53893
rect 65654 53882 65660 53884
rect 65716 53882 65740 53884
rect 65796 53882 65820 53884
rect 65876 53882 65900 53884
rect 65956 53882 65962 53884
rect 65716 53830 65718 53882
rect 65898 53830 65900 53882
rect 65654 53828 65660 53830
rect 65716 53828 65740 53830
rect 65796 53828 65820 53830
rect 65876 53828 65900 53830
rect 65956 53828 65962 53830
rect 65654 53819 65962 53828
rect 68100 53576 68152 53582
rect 68100 53518 68152 53524
rect 68112 53145 68140 53518
rect 68098 53136 68154 53145
rect 68098 53071 68154 53080
rect 65654 52796 65962 52805
rect 65654 52794 65660 52796
rect 65716 52794 65740 52796
rect 65796 52794 65820 52796
rect 65876 52794 65900 52796
rect 65956 52794 65962 52796
rect 65716 52742 65718 52794
rect 65898 52742 65900 52794
rect 65654 52740 65660 52742
rect 65716 52740 65740 52742
rect 65796 52740 65820 52742
rect 65876 52740 65900 52742
rect 65956 52740 65962 52742
rect 65654 52731 65962 52740
rect 67640 51808 67692 51814
rect 67640 51750 67692 51756
rect 65654 51708 65962 51717
rect 65654 51706 65660 51708
rect 65716 51706 65740 51708
rect 65796 51706 65820 51708
rect 65876 51706 65900 51708
rect 65956 51706 65962 51708
rect 65716 51654 65718 51706
rect 65898 51654 65900 51706
rect 65654 51652 65660 51654
rect 65716 51652 65740 51654
rect 65796 51652 65820 51654
rect 65876 51652 65900 51654
rect 65956 51652 65962 51654
rect 65654 51643 65962 51652
rect 67652 51649 67680 51750
rect 67638 51640 67694 51649
rect 67638 51575 67694 51584
rect 65654 50620 65962 50629
rect 65654 50618 65660 50620
rect 65716 50618 65740 50620
rect 65796 50618 65820 50620
rect 65876 50618 65900 50620
rect 65956 50618 65962 50620
rect 65716 50566 65718 50618
rect 65898 50566 65900 50618
rect 65654 50564 65660 50566
rect 65716 50564 65740 50566
rect 65796 50564 65820 50566
rect 65876 50564 65900 50566
rect 65956 50564 65962 50566
rect 65654 50555 65962 50564
rect 68100 50312 68152 50318
rect 68100 50254 68152 50260
rect 68112 50153 68140 50254
rect 68098 50144 68154 50153
rect 68098 50079 68154 50088
rect 65654 49532 65962 49541
rect 65654 49530 65660 49532
rect 65716 49530 65740 49532
rect 65796 49530 65820 49532
rect 65876 49530 65900 49532
rect 65956 49530 65962 49532
rect 65716 49478 65718 49530
rect 65898 49478 65900 49530
rect 65654 49476 65660 49478
rect 65716 49476 65740 49478
rect 65796 49476 65820 49478
rect 65876 49476 65900 49478
rect 65956 49476 65962 49478
rect 65654 49467 65962 49476
rect 67638 48648 67694 48657
rect 67638 48583 67640 48592
rect 67692 48583 67694 48592
rect 67640 48554 67692 48560
rect 65654 48444 65962 48453
rect 65654 48442 65660 48444
rect 65716 48442 65740 48444
rect 65796 48442 65820 48444
rect 65876 48442 65900 48444
rect 65956 48442 65962 48444
rect 65716 48390 65718 48442
rect 65898 48390 65900 48442
rect 65654 48388 65660 48390
rect 65716 48388 65740 48390
rect 65796 48388 65820 48390
rect 65876 48388 65900 48390
rect 65956 48388 65962 48390
rect 65654 48379 65962 48388
rect 67640 47456 67692 47462
rect 67640 47398 67692 47404
rect 65654 47356 65962 47365
rect 65654 47354 65660 47356
rect 65716 47354 65740 47356
rect 65796 47354 65820 47356
rect 65876 47354 65900 47356
rect 65956 47354 65962 47356
rect 65716 47302 65718 47354
rect 65898 47302 65900 47354
rect 65654 47300 65660 47302
rect 65716 47300 65740 47302
rect 65796 47300 65820 47302
rect 65876 47300 65900 47302
rect 65956 47300 65962 47302
rect 65654 47291 65962 47300
rect 67652 47161 67680 47398
rect 67638 47152 67694 47161
rect 67638 47087 67694 47096
rect 65654 46268 65962 46277
rect 65654 46266 65660 46268
rect 65716 46266 65740 46268
rect 65796 46266 65820 46268
rect 65876 46266 65900 46268
rect 65956 46266 65962 46268
rect 65716 46214 65718 46266
rect 65898 46214 65900 46266
rect 65654 46212 65660 46214
rect 65716 46212 65740 46214
rect 65796 46212 65820 46214
rect 65876 46212 65900 46214
rect 65956 46212 65962 46214
rect 65654 46203 65962 46212
rect 68100 45960 68152 45966
rect 68100 45902 68152 45908
rect 68112 45665 68140 45902
rect 68098 45656 68154 45665
rect 68098 45591 68154 45600
rect 65654 45180 65962 45189
rect 65654 45178 65660 45180
rect 65716 45178 65740 45180
rect 65796 45178 65820 45180
rect 65876 45178 65900 45180
rect 65956 45178 65962 45180
rect 65716 45126 65718 45178
rect 65898 45126 65900 45178
rect 65654 45124 65660 45126
rect 65716 45124 65740 45126
rect 65796 45124 65820 45126
rect 65876 45124 65900 45126
rect 65956 45124 65962 45126
rect 65654 45115 65962 45124
rect 67548 44192 67600 44198
rect 67546 44160 67548 44169
rect 67600 44160 67602 44169
rect 65654 44092 65962 44101
rect 67546 44095 67602 44104
rect 65654 44090 65660 44092
rect 65716 44090 65740 44092
rect 65796 44090 65820 44092
rect 65876 44090 65900 44092
rect 65956 44090 65962 44092
rect 65716 44038 65718 44090
rect 65898 44038 65900 44090
rect 65654 44036 65660 44038
rect 65716 44036 65740 44038
rect 65796 44036 65820 44038
rect 65876 44036 65900 44038
rect 65956 44036 65962 44038
rect 65654 44027 65962 44036
rect 65654 43004 65962 43013
rect 65654 43002 65660 43004
rect 65716 43002 65740 43004
rect 65796 43002 65820 43004
rect 65876 43002 65900 43004
rect 65956 43002 65962 43004
rect 65716 42950 65718 43002
rect 65898 42950 65900 43002
rect 65654 42948 65660 42950
rect 65716 42948 65740 42950
rect 65796 42948 65820 42950
rect 65876 42948 65900 42950
rect 65956 42948 65962 42950
rect 65654 42939 65962 42948
rect 68100 42696 68152 42702
rect 68098 42664 68100 42673
rect 68152 42664 68154 42673
rect 68098 42599 68154 42608
rect 65654 41916 65962 41925
rect 65654 41914 65660 41916
rect 65716 41914 65740 41916
rect 65796 41914 65820 41916
rect 65876 41914 65900 41916
rect 65956 41914 65962 41916
rect 65716 41862 65718 41914
rect 65898 41862 65900 41914
rect 65654 41860 65660 41862
rect 65716 41860 65740 41862
rect 65796 41860 65820 41862
rect 65876 41860 65900 41862
rect 65956 41860 65962 41862
rect 65654 41851 65962 41860
rect 68100 41608 68152 41614
rect 68100 41550 68152 41556
rect 68112 41177 68140 41550
rect 68098 41168 68154 41177
rect 68098 41103 68154 41112
rect 65654 40828 65962 40837
rect 65654 40826 65660 40828
rect 65716 40826 65740 40828
rect 65796 40826 65820 40828
rect 65876 40826 65900 40828
rect 65956 40826 65962 40828
rect 65716 40774 65718 40826
rect 65898 40774 65900 40826
rect 65654 40772 65660 40774
rect 65716 40772 65740 40774
rect 65796 40772 65820 40774
rect 65876 40772 65900 40774
rect 65956 40772 65962 40774
rect 65654 40763 65962 40772
rect 67640 39840 67692 39846
rect 67640 39782 67692 39788
rect 65654 39740 65962 39749
rect 65654 39738 65660 39740
rect 65716 39738 65740 39740
rect 65796 39738 65820 39740
rect 65876 39738 65900 39740
rect 65956 39738 65962 39740
rect 65716 39686 65718 39738
rect 65898 39686 65900 39738
rect 65654 39684 65660 39686
rect 65716 39684 65740 39686
rect 65796 39684 65820 39686
rect 65876 39684 65900 39686
rect 65956 39684 65962 39686
rect 65654 39675 65962 39684
rect 67652 39681 67680 39782
rect 67638 39672 67694 39681
rect 67638 39607 67694 39616
rect 65654 38652 65962 38661
rect 65654 38650 65660 38652
rect 65716 38650 65740 38652
rect 65796 38650 65820 38652
rect 65876 38650 65900 38652
rect 65956 38650 65962 38652
rect 65716 38598 65718 38650
rect 65898 38598 65900 38650
rect 65654 38596 65660 38598
rect 65716 38596 65740 38598
rect 65796 38596 65820 38598
rect 65876 38596 65900 38598
rect 65956 38596 65962 38598
rect 65654 38587 65962 38596
rect 68100 38344 68152 38350
rect 68100 38286 68152 38292
rect 68112 38185 68140 38286
rect 68098 38176 68154 38185
rect 68098 38111 68154 38120
rect 65654 37564 65962 37573
rect 65654 37562 65660 37564
rect 65716 37562 65740 37564
rect 65796 37562 65820 37564
rect 65876 37562 65900 37564
rect 65956 37562 65962 37564
rect 65716 37510 65718 37562
rect 65898 37510 65900 37562
rect 65654 37508 65660 37510
rect 65716 37508 65740 37510
rect 65796 37508 65820 37510
rect 65876 37508 65900 37510
rect 65956 37508 65962 37510
rect 65654 37499 65962 37508
rect 67638 36680 67694 36689
rect 67638 36615 67640 36624
rect 67692 36615 67694 36624
rect 67640 36586 67692 36592
rect 65654 36476 65962 36485
rect 65654 36474 65660 36476
rect 65716 36474 65740 36476
rect 65796 36474 65820 36476
rect 65876 36474 65900 36476
rect 65956 36474 65962 36476
rect 65716 36422 65718 36474
rect 65898 36422 65900 36474
rect 65654 36420 65660 36422
rect 65716 36420 65740 36422
rect 65796 36420 65820 36422
rect 65876 36420 65900 36422
rect 65956 36420 65962 36422
rect 65654 36411 65962 36420
rect 67640 35488 67692 35494
rect 67640 35430 67692 35436
rect 65654 35388 65962 35397
rect 65654 35386 65660 35388
rect 65716 35386 65740 35388
rect 65796 35386 65820 35388
rect 65876 35386 65900 35388
rect 65956 35386 65962 35388
rect 65716 35334 65718 35386
rect 65898 35334 65900 35386
rect 65654 35332 65660 35334
rect 65716 35332 65740 35334
rect 65796 35332 65820 35334
rect 65876 35332 65900 35334
rect 65956 35332 65962 35334
rect 65654 35323 65962 35332
rect 67652 35193 67680 35430
rect 67638 35184 67694 35193
rect 67638 35119 67694 35128
rect 65654 34300 65962 34309
rect 65654 34298 65660 34300
rect 65716 34298 65740 34300
rect 65796 34298 65820 34300
rect 65876 34298 65900 34300
rect 65956 34298 65962 34300
rect 65716 34246 65718 34298
rect 65898 34246 65900 34298
rect 65654 34244 65660 34246
rect 65716 34244 65740 34246
rect 65796 34244 65820 34246
rect 65876 34244 65900 34246
rect 65956 34244 65962 34246
rect 65654 34235 65962 34244
rect 68100 33992 68152 33998
rect 68100 33934 68152 33940
rect 68112 33697 68140 33934
rect 68098 33688 68154 33697
rect 68098 33623 68154 33632
rect 65654 33212 65962 33221
rect 65654 33210 65660 33212
rect 65716 33210 65740 33212
rect 65796 33210 65820 33212
rect 65876 33210 65900 33212
rect 65956 33210 65962 33212
rect 65716 33158 65718 33210
rect 65898 33158 65900 33210
rect 65654 33156 65660 33158
rect 65716 33156 65740 33158
rect 65796 33156 65820 33158
rect 65876 33156 65900 33158
rect 65956 33156 65962 33158
rect 65654 33147 65962 33156
rect 67640 32224 67692 32230
rect 67638 32192 67640 32201
rect 67692 32192 67694 32201
rect 65654 32124 65962 32133
rect 67638 32127 67694 32136
rect 65654 32122 65660 32124
rect 65716 32122 65740 32124
rect 65796 32122 65820 32124
rect 65876 32122 65900 32124
rect 65956 32122 65962 32124
rect 65716 32070 65718 32122
rect 65898 32070 65900 32122
rect 65654 32068 65660 32070
rect 65716 32068 65740 32070
rect 65796 32068 65820 32070
rect 65876 32068 65900 32070
rect 65956 32068 65962 32070
rect 65654 32059 65962 32068
rect 65654 31036 65962 31045
rect 65654 31034 65660 31036
rect 65716 31034 65740 31036
rect 65796 31034 65820 31036
rect 65876 31034 65900 31036
rect 65956 31034 65962 31036
rect 65716 30982 65718 31034
rect 65898 30982 65900 31034
rect 65654 30980 65660 30982
rect 65716 30980 65740 30982
rect 65796 30980 65820 30982
rect 65876 30980 65900 30982
rect 65956 30980 65962 30982
rect 65654 30971 65962 30980
rect 68100 30728 68152 30734
rect 68098 30696 68100 30705
rect 68152 30696 68154 30705
rect 68098 30631 68154 30640
rect 65654 29948 65962 29957
rect 65654 29946 65660 29948
rect 65716 29946 65740 29948
rect 65796 29946 65820 29948
rect 65876 29946 65900 29948
rect 65956 29946 65962 29948
rect 65716 29894 65718 29946
rect 65898 29894 65900 29946
rect 65654 29892 65660 29894
rect 65716 29892 65740 29894
rect 65796 29892 65820 29894
rect 65876 29892 65900 29894
rect 65956 29892 65962 29894
rect 65654 29883 65962 29892
rect 68100 29640 68152 29646
rect 68100 29582 68152 29588
rect 68112 29209 68140 29582
rect 68098 29200 68154 29209
rect 68098 29135 68154 29144
rect 65654 28860 65962 28869
rect 65654 28858 65660 28860
rect 65716 28858 65740 28860
rect 65796 28858 65820 28860
rect 65876 28858 65900 28860
rect 65956 28858 65962 28860
rect 65716 28806 65718 28858
rect 65898 28806 65900 28858
rect 65654 28804 65660 28806
rect 65716 28804 65740 28806
rect 65796 28804 65820 28806
rect 65876 28804 65900 28806
rect 65956 28804 65962 28806
rect 65654 28795 65962 28804
rect 67640 27872 67692 27878
rect 67640 27814 67692 27820
rect 65654 27772 65962 27781
rect 65654 27770 65660 27772
rect 65716 27770 65740 27772
rect 65796 27770 65820 27772
rect 65876 27770 65900 27772
rect 65956 27770 65962 27772
rect 65716 27718 65718 27770
rect 65898 27718 65900 27770
rect 65654 27716 65660 27718
rect 65716 27716 65740 27718
rect 65796 27716 65820 27718
rect 65876 27716 65900 27718
rect 65956 27716 65962 27718
rect 65654 27707 65962 27716
rect 67652 27713 67680 27814
rect 67638 27704 67694 27713
rect 67638 27639 67694 27648
rect 65654 26684 65962 26693
rect 65654 26682 65660 26684
rect 65716 26682 65740 26684
rect 65796 26682 65820 26684
rect 65876 26682 65900 26684
rect 65956 26682 65962 26684
rect 65716 26630 65718 26682
rect 65898 26630 65900 26682
rect 65654 26628 65660 26630
rect 65716 26628 65740 26630
rect 65796 26628 65820 26630
rect 65876 26628 65900 26630
rect 65956 26628 65962 26630
rect 65654 26619 65962 26628
rect 68100 26376 68152 26382
rect 68100 26318 68152 26324
rect 68112 26217 68140 26318
rect 68098 26208 68154 26217
rect 68098 26143 68154 26152
rect 65654 25596 65962 25605
rect 65654 25594 65660 25596
rect 65716 25594 65740 25596
rect 65796 25594 65820 25596
rect 65876 25594 65900 25596
rect 65956 25594 65962 25596
rect 65716 25542 65718 25594
rect 65898 25542 65900 25594
rect 65654 25540 65660 25542
rect 65716 25540 65740 25542
rect 65796 25540 65820 25542
rect 65876 25540 65900 25542
rect 65956 25540 65962 25542
rect 65654 25531 65962 25540
rect 67638 24712 67694 24721
rect 67638 24647 67640 24656
rect 67692 24647 67694 24656
rect 67640 24618 67692 24624
rect 56324 24608 56376 24614
rect 56324 24550 56376 24556
rect 65654 24508 65962 24517
rect 65654 24506 65660 24508
rect 65716 24506 65740 24508
rect 65796 24506 65820 24508
rect 65876 24506 65900 24508
rect 65956 24506 65962 24508
rect 65716 24454 65718 24506
rect 65898 24454 65900 24506
rect 65654 24452 65660 24454
rect 65716 24452 65740 24454
rect 65796 24452 65820 24454
rect 65876 24452 65900 24454
rect 65956 24452 65962 24454
rect 65654 24443 65962 24452
rect 43260 24404 43312 24410
rect 43260 24346 43312 24352
rect 40040 24200 40092 24206
rect 40040 24142 40092 24148
rect 41144 24200 41196 24206
rect 41144 24142 41196 24148
rect 42524 24200 42576 24206
rect 42524 24142 42576 24148
rect 42892 24200 42944 24206
rect 42892 24142 42944 24148
rect 43260 24200 43312 24206
rect 43260 24142 43312 24148
rect 39856 23112 39908 23118
rect 39856 23054 39908 23060
rect 39868 22098 39896 23054
rect 40052 22642 40080 24142
rect 42432 24064 42484 24070
rect 42432 24006 42484 24012
rect 42444 23730 42472 24006
rect 42432 23724 42484 23730
rect 42432 23666 42484 23672
rect 41604 23656 41656 23662
rect 41604 23598 41656 23604
rect 41616 23322 41644 23598
rect 41696 23520 41748 23526
rect 41696 23462 41748 23468
rect 41604 23316 41656 23322
rect 41604 23258 41656 23264
rect 40132 23044 40184 23050
rect 40132 22986 40184 22992
rect 40144 22778 40172 22986
rect 40132 22772 40184 22778
rect 40132 22714 40184 22720
rect 40040 22636 40092 22642
rect 40040 22578 40092 22584
rect 39856 22092 39908 22098
rect 39856 22034 39908 22040
rect 41616 21554 41644 23258
rect 41708 22642 41736 23462
rect 42444 22642 42472 23666
rect 41696 22636 41748 22642
rect 41696 22578 41748 22584
rect 41880 22636 41932 22642
rect 41880 22578 41932 22584
rect 42432 22636 42484 22642
rect 42432 22578 42484 22584
rect 41788 21888 41840 21894
rect 41788 21830 41840 21836
rect 41236 21548 41288 21554
rect 41236 21490 41288 21496
rect 41604 21548 41656 21554
rect 41604 21490 41656 21496
rect 40132 21004 40184 21010
rect 40132 20946 40184 20952
rect 39488 20256 39540 20262
rect 39488 20198 39540 20204
rect 39500 19786 39528 20198
rect 40144 19854 40172 20946
rect 40224 20392 40276 20398
rect 40224 20334 40276 20340
rect 40236 20058 40264 20334
rect 41248 20058 41276 21490
rect 41420 21480 41472 21486
rect 41616 21434 41644 21490
rect 41420 21422 41472 21428
rect 41432 21078 41460 21422
rect 41524 21406 41644 21434
rect 41420 21072 41472 21078
rect 41420 21014 41472 21020
rect 41328 20800 41380 20806
rect 41328 20742 41380 20748
rect 41340 20602 41368 20742
rect 41328 20596 41380 20602
rect 41328 20538 41380 20544
rect 41432 20534 41460 21014
rect 41524 20942 41552 21406
rect 41604 21344 41656 21350
rect 41604 21286 41656 21292
rect 41616 20942 41644 21286
rect 41696 21004 41748 21010
rect 41696 20946 41748 20952
rect 41512 20936 41564 20942
rect 41512 20878 41564 20884
rect 41604 20936 41656 20942
rect 41604 20878 41656 20884
rect 41420 20528 41472 20534
rect 41420 20470 41472 20476
rect 41708 20398 41736 20946
rect 41800 20874 41828 21830
rect 41892 21350 41920 22578
rect 42064 22432 42116 22438
rect 42064 22374 42116 22380
rect 42076 22030 42104 22374
rect 42064 22024 42116 22030
rect 42064 21966 42116 21972
rect 42536 21894 42564 24142
rect 42800 23860 42852 23866
rect 42800 23802 42852 23808
rect 42812 22642 42840 23802
rect 42904 22778 42932 24142
rect 43272 23866 43300 24142
rect 50294 23964 50602 23973
rect 50294 23962 50300 23964
rect 50356 23962 50380 23964
rect 50436 23962 50460 23964
rect 50516 23962 50540 23964
rect 50596 23962 50602 23964
rect 50356 23910 50358 23962
rect 50538 23910 50540 23962
rect 50294 23908 50300 23910
rect 50356 23908 50380 23910
rect 50436 23908 50460 23910
rect 50516 23908 50540 23910
rect 50596 23908 50602 23910
rect 50294 23899 50602 23908
rect 43260 23860 43312 23866
rect 43260 23802 43312 23808
rect 67548 23520 67600 23526
rect 67548 23462 67600 23468
rect 65654 23420 65962 23429
rect 65654 23418 65660 23420
rect 65716 23418 65740 23420
rect 65796 23418 65820 23420
rect 65876 23418 65900 23420
rect 65956 23418 65962 23420
rect 65716 23366 65718 23418
rect 65898 23366 65900 23418
rect 65654 23364 65660 23366
rect 65716 23364 65740 23366
rect 65796 23364 65820 23366
rect 65876 23364 65900 23366
rect 65956 23364 65962 23366
rect 65654 23355 65962 23364
rect 67560 23225 67588 23462
rect 67546 23216 67602 23225
rect 67546 23151 67602 23160
rect 43352 23112 43404 23118
rect 43352 23054 43404 23060
rect 43628 23112 43680 23118
rect 43628 23054 43680 23060
rect 42892 22772 42944 22778
rect 42892 22714 42944 22720
rect 42616 22636 42668 22642
rect 42616 22578 42668 22584
rect 42800 22636 42852 22642
rect 42800 22578 42852 22584
rect 42524 21888 42576 21894
rect 42524 21830 42576 21836
rect 42536 21622 42564 21830
rect 42628 21690 42656 22578
rect 43364 21690 43392 23054
rect 43640 22778 43668 23054
rect 50294 22876 50602 22885
rect 50294 22874 50300 22876
rect 50356 22874 50380 22876
rect 50436 22874 50460 22876
rect 50516 22874 50540 22876
rect 50596 22874 50602 22876
rect 50356 22822 50358 22874
rect 50538 22822 50540 22874
rect 50294 22820 50300 22822
rect 50356 22820 50380 22822
rect 50436 22820 50460 22822
rect 50516 22820 50540 22822
rect 50596 22820 50602 22822
rect 50294 22811 50602 22820
rect 43628 22772 43680 22778
rect 43628 22714 43680 22720
rect 65654 22332 65962 22341
rect 65654 22330 65660 22332
rect 65716 22330 65740 22332
rect 65796 22330 65820 22332
rect 65876 22330 65900 22332
rect 65956 22330 65962 22332
rect 65716 22278 65718 22330
rect 65898 22278 65900 22330
rect 65654 22276 65660 22278
rect 65716 22276 65740 22278
rect 65796 22276 65820 22278
rect 65876 22276 65900 22278
rect 65956 22276 65962 22278
rect 65654 22267 65962 22276
rect 68100 22160 68152 22166
rect 68100 22102 68152 22108
rect 50294 21788 50602 21797
rect 50294 21786 50300 21788
rect 50356 21786 50380 21788
rect 50436 21786 50460 21788
rect 50516 21786 50540 21788
rect 50596 21786 50602 21788
rect 50356 21734 50358 21786
rect 50538 21734 50540 21786
rect 50294 21732 50300 21734
rect 50356 21732 50380 21734
rect 50436 21732 50460 21734
rect 50516 21732 50540 21734
rect 50596 21732 50602 21734
rect 50294 21723 50602 21732
rect 68112 21729 68140 22102
rect 68098 21720 68154 21729
rect 42616 21684 42668 21690
rect 42616 21626 42668 21632
rect 43352 21684 43404 21690
rect 68098 21655 68154 21664
rect 43352 21626 43404 21632
rect 42524 21616 42576 21622
rect 42524 21558 42576 21564
rect 42432 21548 42484 21554
rect 42432 21490 42484 21496
rect 42800 21548 42852 21554
rect 42800 21490 42852 21496
rect 41880 21344 41932 21350
rect 41880 21286 41932 21292
rect 42444 21146 42472 21490
rect 42432 21140 42484 21146
rect 42432 21082 42484 21088
rect 41788 20868 41840 20874
rect 41788 20810 41840 20816
rect 41800 20466 41828 20810
rect 42812 20602 42840 21490
rect 65654 21244 65962 21253
rect 65654 21242 65660 21244
rect 65716 21242 65740 21244
rect 65796 21242 65820 21244
rect 65876 21242 65900 21244
rect 65956 21242 65962 21244
rect 65716 21190 65718 21242
rect 65898 21190 65900 21242
rect 65654 21188 65660 21190
rect 65716 21188 65740 21190
rect 65796 21188 65820 21190
rect 65876 21188 65900 21190
rect 65956 21188 65962 21190
rect 65654 21179 65962 21188
rect 50294 20700 50602 20709
rect 50294 20698 50300 20700
rect 50356 20698 50380 20700
rect 50436 20698 50460 20700
rect 50516 20698 50540 20700
rect 50596 20698 50602 20700
rect 50356 20646 50358 20698
rect 50538 20646 50540 20698
rect 50294 20644 50300 20646
rect 50356 20644 50380 20646
rect 50436 20644 50460 20646
rect 50516 20644 50540 20646
rect 50596 20644 50602 20646
rect 50294 20635 50602 20644
rect 42800 20596 42852 20602
rect 42800 20538 42852 20544
rect 41788 20460 41840 20466
rect 41788 20402 41840 20408
rect 42432 20460 42484 20466
rect 42432 20402 42484 20408
rect 41696 20392 41748 20398
rect 41696 20334 41748 20340
rect 41800 20346 41828 20402
rect 40224 20052 40276 20058
rect 40224 19994 40276 20000
rect 41236 20052 41288 20058
rect 41236 19994 41288 20000
rect 40132 19848 40184 19854
rect 40132 19790 40184 19796
rect 39488 19780 39540 19786
rect 39488 19722 39540 19728
rect 39500 19446 39528 19722
rect 40236 19446 40264 19994
rect 39488 19440 39540 19446
rect 39488 19382 39540 19388
rect 40224 19440 40276 19446
rect 40224 19382 40276 19388
rect 40236 18970 40264 19382
rect 41328 19168 41380 19174
rect 41328 19110 41380 19116
rect 40224 18964 40276 18970
rect 40224 18906 40276 18912
rect 40236 18426 40264 18906
rect 41340 18834 41368 19110
rect 41328 18828 41380 18834
rect 41328 18770 41380 18776
rect 41420 18760 41472 18766
rect 41420 18702 41472 18708
rect 40224 18420 40276 18426
rect 40224 18362 40276 18368
rect 40040 17740 40092 17746
rect 40040 17682 40092 17688
rect 40052 16250 40080 17682
rect 40040 16244 40092 16250
rect 40040 16186 40092 16192
rect 41432 15162 41460 18702
rect 41420 15156 41472 15162
rect 41420 15098 41472 15104
rect 39856 14816 39908 14822
rect 39856 14758 39908 14764
rect 39868 13326 39896 14758
rect 39948 13864 40000 13870
rect 39948 13806 40000 13812
rect 39960 13326 39988 13806
rect 39856 13320 39908 13326
rect 39856 13262 39908 13268
rect 39948 13320 40000 13326
rect 39948 13262 40000 13268
rect 39868 12238 39896 13262
rect 41708 12986 41736 20334
rect 41800 20318 41920 20346
rect 41788 20256 41840 20262
rect 41788 20198 41840 20204
rect 41800 18902 41828 20198
rect 41892 20058 41920 20318
rect 41880 20052 41932 20058
rect 41880 19994 41932 20000
rect 41788 18896 41840 18902
rect 41788 18838 41840 18844
rect 41696 12980 41748 12986
rect 41696 12922 41748 12928
rect 41236 12844 41288 12850
rect 41236 12786 41288 12792
rect 41248 12442 41276 12786
rect 41236 12436 41288 12442
rect 41236 12378 41288 12384
rect 39856 12232 39908 12238
rect 39856 12174 39908 12180
rect 40408 11348 40460 11354
rect 40408 11290 40460 11296
rect 40420 10810 40448 11290
rect 42444 10810 42472 20402
rect 67640 20256 67692 20262
rect 67638 20224 67640 20233
rect 67692 20224 67694 20233
rect 65654 20156 65962 20165
rect 67638 20159 67694 20168
rect 65654 20154 65660 20156
rect 65716 20154 65740 20156
rect 65796 20154 65820 20156
rect 65876 20154 65900 20156
rect 65956 20154 65962 20156
rect 65716 20102 65718 20154
rect 65898 20102 65900 20154
rect 65654 20100 65660 20102
rect 65716 20100 65740 20102
rect 65796 20100 65820 20102
rect 65876 20100 65900 20102
rect 65956 20100 65962 20102
rect 65654 20091 65962 20100
rect 50294 19612 50602 19621
rect 50294 19610 50300 19612
rect 50356 19610 50380 19612
rect 50436 19610 50460 19612
rect 50516 19610 50540 19612
rect 50596 19610 50602 19612
rect 50356 19558 50358 19610
rect 50538 19558 50540 19610
rect 50294 19556 50300 19558
rect 50356 19556 50380 19558
rect 50436 19556 50460 19558
rect 50516 19556 50540 19558
rect 50596 19556 50602 19558
rect 50294 19547 50602 19556
rect 65654 19068 65962 19077
rect 65654 19066 65660 19068
rect 65716 19066 65740 19068
rect 65796 19066 65820 19068
rect 65876 19066 65900 19068
rect 65956 19066 65962 19068
rect 65716 19014 65718 19066
rect 65898 19014 65900 19066
rect 65654 19012 65660 19014
rect 65716 19012 65740 19014
rect 65796 19012 65820 19014
rect 65876 19012 65900 19014
rect 65956 19012 65962 19014
rect 65654 19003 65962 19012
rect 68100 18760 68152 18766
rect 68098 18728 68100 18737
rect 68152 18728 68154 18737
rect 68098 18663 68154 18672
rect 50294 18524 50602 18533
rect 50294 18522 50300 18524
rect 50356 18522 50380 18524
rect 50436 18522 50460 18524
rect 50516 18522 50540 18524
rect 50596 18522 50602 18524
rect 50356 18470 50358 18522
rect 50538 18470 50540 18522
rect 50294 18468 50300 18470
rect 50356 18468 50380 18470
rect 50436 18468 50460 18470
rect 50516 18468 50540 18470
rect 50596 18468 50602 18470
rect 50294 18459 50602 18468
rect 65654 17980 65962 17989
rect 65654 17978 65660 17980
rect 65716 17978 65740 17980
rect 65796 17978 65820 17980
rect 65876 17978 65900 17980
rect 65956 17978 65962 17980
rect 65716 17926 65718 17978
rect 65898 17926 65900 17978
rect 65654 17924 65660 17926
rect 65716 17924 65740 17926
rect 65796 17924 65820 17926
rect 65876 17924 65900 17926
rect 65956 17924 65962 17926
rect 65654 17915 65962 17924
rect 68100 17672 68152 17678
rect 68100 17614 68152 17620
rect 50294 17436 50602 17445
rect 50294 17434 50300 17436
rect 50356 17434 50380 17436
rect 50436 17434 50460 17436
rect 50516 17434 50540 17436
rect 50596 17434 50602 17436
rect 50356 17382 50358 17434
rect 50538 17382 50540 17434
rect 50294 17380 50300 17382
rect 50356 17380 50380 17382
rect 50436 17380 50460 17382
rect 50516 17380 50540 17382
rect 50596 17380 50602 17382
rect 50294 17371 50602 17380
rect 68112 17241 68140 17614
rect 68098 17232 68154 17241
rect 68098 17167 68154 17176
rect 65654 16892 65962 16901
rect 65654 16890 65660 16892
rect 65716 16890 65740 16892
rect 65796 16890 65820 16892
rect 65876 16890 65900 16892
rect 65956 16890 65962 16892
rect 65716 16838 65718 16890
rect 65898 16838 65900 16890
rect 65654 16836 65660 16838
rect 65716 16836 65740 16838
rect 65796 16836 65820 16838
rect 65876 16836 65900 16838
rect 65956 16836 65962 16838
rect 65654 16827 65962 16836
rect 50294 16348 50602 16357
rect 50294 16346 50300 16348
rect 50356 16346 50380 16348
rect 50436 16346 50460 16348
rect 50516 16346 50540 16348
rect 50596 16346 50602 16348
rect 50356 16294 50358 16346
rect 50538 16294 50540 16346
rect 50294 16292 50300 16294
rect 50356 16292 50380 16294
rect 50436 16292 50460 16294
rect 50516 16292 50540 16294
rect 50596 16292 50602 16294
rect 50294 16283 50602 16292
rect 67640 15904 67692 15910
rect 67640 15846 67692 15852
rect 65654 15804 65962 15813
rect 65654 15802 65660 15804
rect 65716 15802 65740 15804
rect 65796 15802 65820 15804
rect 65876 15802 65900 15804
rect 65956 15802 65962 15804
rect 65716 15750 65718 15802
rect 65898 15750 65900 15802
rect 65654 15748 65660 15750
rect 65716 15748 65740 15750
rect 65796 15748 65820 15750
rect 65876 15748 65900 15750
rect 65956 15748 65962 15750
rect 65654 15739 65962 15748
rect 67652 15745 67680 15846
rect 67638 15736 67694 15745
rect 67638 15671 67694 15680
rect 50294 15260 50602 15269
rect 50294 15258 50300 15260
rect 50356 15258 50380 15260
rect 50436 15258 50460 15260
rect 50516 15258 50540 15260
rect 50596 15258 50602 15260
rect 50356 15206 50358 15258
rect 50538 15206 50540 15258
rect 50294 15204 50300 15206
rect 50356 15204 50380 15206
rect 50436 15204 50460 15206
rect 50516 15204 50540 15206
rect 50596 15204 50602 15206
rect 50294 15195 50602 15204
rect 65654 14716 65962 14725
rect 65654 14714 65660 14716
rect 65716 14714 65740 14716
rect 65796 14714 65820 14716
rect 65876 14714 65900 14716
rect 65956 14714 65962 14716
rect 65716 14662 65718 14714
rect 65898 14662 65900 14714
rect 65654 14660 65660 14662
rect 65716 14660 65740 14662
rect 65796 14660 65820 14662
rect 65876 14660 65900 14662
rect 65956 14660 65962 14662
rect 65654 14651 65962 14660
rect 68100 14408 68152 14414
rect 68100 14350 68152 14356
rect 68112 14249 68140 14350
rect 68098 14240 68154 14249
rect 50294 14172 50602 14181
rect 68098 14175 68154 14184
rect 50294 14170 50300 14172
rect 50356 14170 50380 14172
rect 50436 14170 50460 14172
rect 50516 14170 50540 14172
rect 50596 14170 50602 14172
rect 50356 14118 50358 14170
rect 50538 14118 50540 14170
rect 50294 14116 50300 14118
rect 50356 14116 50380 14118
rect 50436 14116 50460 14118
rect 50516 14116 50540 14118
rect 50596 14116 50602 14118
rect 50294 14107 50602 14116
rect 65654 13628 65962 13637
rect 65654 13626 65660 13628
rect 65716 13626 65740 13628
rect 65796 13626 65820 13628
rect 65876 13626 65900 13628
rect 65956 13626 65962 13628
rect 65716 13574 65718 13626
rect 65898 13574 65900 13626
rect 65654 13572 65660 13574
rect 65716 13572 65740 13574
rect 65796 13572 65820 13574
rect 65876 13572 65900 13574
rect 65956 13572 65962 13574
rect 65654 13563 65962 13572
rect 50294 13084 50602 13093
rect 50294 13082 50300 13084
rect 50356 13082 50380 13084
rect 50436 13082 50460 13084
rect 50516 13082 50540 13084
rect 50596 13082 50602 13084
rect 50356 13030 50358 13082
rect 50538 13030 50540 13082
rect 50294 13028 50300 13030
rect 50356 13028 50380 13030
rect 50436 13028 50460 13030
rect 50516 13028 50540 13030
rect 50596 13028 50602 13030
rect 50294 13019 50602 13028
rect 67638 12744 67694 12753
rect 67638 12679 67640 12688
rect 67692 12679 67694 12688
rect 67640 12650 67692 12656
rect 65654 12540 65962 12549
rect 65654 12538 65660 12540
rect 65716 12538 65740 12540
rect 65796 12538 65820 12540
rect 65876 12538 65900 12540
rect 65956 12538 65962 12540
rect 65716 12486 65718 12538
rect 65898 12486 65900 12538
rect 65654 12484 65660 12486
rect 65716 12484 65740 12486
rect 65796 12484 65820 12486
rect 65876 12484 65900 12486
rect 65956 12484 65962 12486
rect 65654 12475 65962 12484
rect 50294 11996 50602 12005
rect 50294 11994 50300 11996
rect 50356 11994 50380 11996
rect 50436 11994 50460 11996
rect 50516 11994 50540 11996
rect 50596 11994 50602 11996
rect 50356 11942 50358 11994
rect 50538 11942 50540 11994
rect 50294 11940 50300 11942
rect 50356 11940 50380 11942
rect 50436 11940 50460 11942
rect 50516 11940 50540 11942
rect 50596 11940 50602 11942
rect 50294 11931 50602 11940
rect 67640 11552 67692 11558
rect 67640 11494 67692 11500
rect 65654 11452 65962 11461
rect 65654 11450 65660 11452
rect 65716 11450 65740 11452
rect 65796 11450 65820 11452
rect 65876 11450 65900 11452
rect 65956 11450 65962 11452
rect 65716 11398 65718 11450
rect 65898 11398 65900 11450
rect 65654 11396 65660 11398
rect 65716 11396 65740 11398
rect 65796 11396 65820 11398
rect 65876 11396 65900 11398
rect 65956 11396 65962 11398
rect 65654 11387 65962 11396
rect 67652 11257 67680 11494
rect 67638 11248 67694 11257
rect 67638 11183 67694 11192
rect 50294 10908 50602 10917
rect 50294 10906 50300 10908
rect 50356 10906 50380 10908
rect 50436 10906 50460 10908
rect 50516 10906 50540 10908
rect 50596 10906 50602 10908
rect 50356 10854 50358 10906
rect 50538 10854 50540 10906
rect 50294 10852 50300 10854
rect 50356 10852 50380 10854
rect 50436 10852 50460 10854
rect 50516 10852 50540 10854
rect 50596 10852 50602 10854
rect 50294 10843 50602 10852
rect 40408 10804 40460 10810
rect 40408 10746 40460 10752
rect 42432 10804 42484 10810
rect 42432 10746 42484 10752
rect 39856 10668 39908 10674
rect 39856 10610 39908 10616
rect 39868 9926 39896 10610
rect 40960 10600 41012 10606
rect 40960 10542 41012 10548
rect 40868 10464 40920 10470
rect 40868 10406 40920 10412
rect 39856 9920 39908 9926
rect 39856 9862 39908 9868
rect 40880 9382 40908 10406
rect 40868 9376 40920 9382
rect 40868 9318 40920 9324
rect 40972 8498 41000 10542
rect 65654 10364 65962 10373
rect 65654 10362 65660 10364
rect 65716 10362 65740 10364
rect 65796 10362 65820 10364
rect 65876 10362 65900 10364
rect 65956 10362 65962 10364
rect 65716 10310 65718 10362
rect 65898 10310 65900 10362
rect 65654 10308 65660 10310
rect 65716 10308 65740 10310
rect 65796 10308 65820 10310
rect 65876 10308 65900 10310
rect 65956 10308 65962 10310
rect 65654 10299 65962 10308
rect 68100 10056 68152 10062
rect 68100 9998 68152 10004
rect 50294 9820 50602 9829
rect 50294 9818 50300 9820
rect 50356 9818 50380 9820
rect 50436 9818 50460 9820
rect 50516 9818 50540 9820
rect 50596 9818 50602 9820
rect 50356 9766 50358 9818
rect 50538 9766 50540 9818
rect 50294 9764 50300 9766
rect 50356 9764 50380 9766
rect 50436 9764 50460 9766
rect 50516 9764 50540 9766
rect 50596 9764 50602 9766
rect 50294 9755 50602 9764
rect 68112 9761 68140 9998
rect 68098 9752 68154 9761
rect 68098 9687 68154 9696
rect 65654 9276 65962 9285
rect 65654 9274 65660 9276
rect 65716 9274 65740 9276
rect 65796 9274 65820 9276
rect 65876 9274 65900 9276
rect 65956 9274 65962 9276
rect 65716 9222 65718 9274
rect 65898 9222 65900 9274
rect 65654 9220 65660 9222
rect 65716 9220 65740 9222
rect 65796 9220 65820 9222
rect 65876 9220 65900 9222
rect 65956 9220 65962 9222
rect 65654 9211 65962 9220
rect 50294 8732 50602 8741
rect 50294 8730 50300 8732
rect 50356 8730 50380 8732
rect 50436 8730 50460 8732
rect 50516 8730 50540 8732
rect 50596 8730 50602 8732
rect 50356 8678 50358 8730
rect 50538 8678 50540 8730
rect 50294 8676 50300 8678
rect 50356 8676 50380 8678
rect 50436 8676 50460 8678
rect 50516 8676 50540 8678
rect 50596 8676 50602 8678
rect 50294 8667 50602 8676
rect 40960 8492 41012 8498
rect 40960 8434 41012 8440
rect 67548 8356 67600 8362
rect 67548 8298 67600 8304
rect 67560 8265 67588 8298
rect 67546 8256 67602 8265
rect 65654 8188 65962 8197
rect 67546 8191 67602 8200
rect 65654 8186 65660 8188
rect 65716 8186 65740 8188
rect 65796 8186 65820 8188
rect 65876 8186 65900 8188
rect 65956 8186 65962 8188
rect 65716 8134 65718 8186
rect 65898 8134 65900 8186
rect 65654 8132 65660 8134
rect 65716 8132 65740 8134
rect 65796 8132 65820 8134
rect 65876 8132 65900 8134
rect 65956 8132 65962 8134
rect 65654 8123 65962 8132
rect 50294 7644 50602 7653
rect 50294 7642 50300 7644
rect 50356 7642 50380 7644
rect 50436 7642 50460 7644
rect 50516 7642 50540 7644
rect 50596 7642 50602 7644
rect 50356 7590 50358 7642
rect 50538 7590 50540 7642
rect 50294 7588 50300 7590
rect 50356 7588 50380 7590
rect 50436 7588 50460 7590
rect 50516 7588 50540 7590
rect 50596 7588 50602 7590
rect 50294 7579 50602 7588
rect 65654 7100 65962 7109
rect 65654 7098 65660 7100
rect 65716 7098 65740 7100
rect 65796 7098 65820 7100
rect 65876 7098 65900 7100
rect 65956 7098 65962 7100
rect 65716 7046 65718 7098
rect 65898 7046 65900 7098
rect 65654 7044 65660 7046
rect 65716 7044 65740 7046
rect 65796 7044 65820 7046
rect 65876 7044 65900 7046
rect 65956 7044 65962 7046
rect 65654 7035 65962 7044
rect 68100 6792 68152 6798
rect 68098 6760 68100 6769
rect 68152 6760 68154 6769
rect 68098 6695 68154 6704
rect 50294 6556 50602 6565
rect 50294 6554 50300 6556
rect 50356 6554 50380 6556
rect 50436 6554 50460 6556
rect 50516 6554 50540 6556
rect 50596 6554 50602 6556
rect 50356 6502 50358 6554
rect 50538 6502 50540 6554
rect 50294 6500 50300 6502
rect 50356 6500 50380 6502
rect 50436 6500 50460 6502
rect 50516 6500 50540 6502
rect 50596 6500 50602 6502
rect 50294 6491 50602 6500
rect 37740 6316 37792 6322
rect 37740 6258 37792 6264
rect 39396 6316 39448 6322
rect 39396 6258 39448 6264
rect 36268 6248 36320 6254
rect 36268 6190 36320 6196
rect 36280 6118 36308 6190
rect 36268 6112 36320 6118
rect 36268 6054 36320 6060
rect 36728 6112 36780 6118
rect 36728 6054 36780 6060
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 36280 5914 36308 6054
rect 36268 5908 36320 5914
rect 36268 5850 36320 5856
rect 36268 5704 36320 5710
rect 36268 5646 36320 5652
rect 36452 5704 36504 5710
rect 36452 5646 36504 5652
rect 36176 5636 36228 5642
rect 36176 5578 36228 5584
rect 36188 5370 36216 5578
rect 34796 5364 34848 5370
rect 34796 5306 34848 5312
rect 36176 5364 36228 5370
rect 36176 5306 36228 5312
rect 36280 5234 36308 5646
rect 34704 5228 34756 5234
rect 34704 5170 34756 5176
rect 36176 5228 36228 5234
rect 36176 5170 36228 5176
rect 36268 5228 36320 5234
rect 36268 5170 36320 5176
rect 34612 5024 34664 5030
rect 34612 4966 34664 4972
rect 32588 4616 32640 4622
rect 32588 4558 32640 4564
rect 34520 4616 34572 4622
rect 34520 4558 34572 4564
rect 32128 4276 32180 4282
rect 32128 4218 32180 4224
rect 34532 4214 34560 4558
rect 30564 4208 30616 4214
rect 30564 4150 30616 4156
rect 34520 4208 34572 4214
rect 34520 4150 34572 4156
rect 30288 4140 30340 4146
rect 30288 4082 30340 4088
rect 34624 4078 34652 4966
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 36188 4690 36216 5170
rect 36280 4758 36308 5170
rect 36464 4826 36492 5646
rect 36740 5302 36768 6054
rect 37752 5914 37780 6258
rect 65654 6012 65962 6021
rect 65654 6010 65660 6012
rect 65716 6010 65740 6012
rect 65796 6010 65820 6012
rect 65876 6010 65900 6012
rect 65956 6010 65962 6012
rect 65716 5958 65718 6010
rect 65898 5958 65900 6010
rect 65654 5956 65660 5958
rect 65716 5956 65740 5958
rect 65796 5956 65820 5958
rect 65876 5956 65900 5958
rect 65956 5956 65962 5958
rect 65654 5947 65962 5956
rect 37740 5908 37792 5914
rect 37740 5850 37792 5856
rect 68100 5704 68152 5710
rect 68100 5646 68152 5652
rect 50294 5468 50602 5477
rect 50294 5466 50300 5468
rect 50356 5466 50380 5468
rect 50436 5466 50460 5468
rect 50516 5466 50540 5468
rect 50596 5466 50602 5468
rect 50356 5414 50358 5466
rect 50538 5414 50540 5466
rect 50294 5412 50300 5414
rect 50356 5412 50380 5414
rect 50436 5412 50460 5414
rect 50516 5412 50540 5414
rect 50596 5412 50602 5414
rect 50294 5403 50602 5412
rect 36728 5296 36780 5302
rect 68112 5273 68140 5646
rect 36728 5238 36780 5244
rect 68098 5264 68154 5273
rect 68098 5199 68154 5208
rect 58808 5160 58860 5166
rect 58808 5102 58860 5108
rect 58716 5024 58768 5030
rect 58716 4966 58768 4972
rect 36452 4820 36504 4826
rect 36452 4762 36504 4768
rect 36268 4752 36320 4758
rect 36268 4694 36320 4700
rect 57244 4752 57296 4758
rect 57244 4694 57296 4700
rect 58256 4752 58308 4758
rect 58256 4694 58308 4700
rect 36176 4684 36228 4690
rect 36176 4626 36228 4632
rect 36912 4616 36964 4622
rect 36912 4558 36964 4564
rect 57152 4616 57204 4622
rect 57152 4558 57204 4564
rect 36924 4282 36952 4558
rect 50294 4380 50602 4389
rect 50294 4378 50300 4380
rect 50356 4378 50380 4380
rect 50436 4378 50460 4380
rect 50516 4378 50540 4380
rect 50596 4378 50602 4380
rect 50356 4326 50358 4378
rect 50538 4326 50540 4378
rect 50294 4324 50300 4326
rect 50356 4324 50380 4326
rect 50436 4324 50460 4326
rect 50516 4324 50540 4326
rect 50596 4324 50602 4326
rect 50294 4315 50602 4324
rect 36912 4276 36964 4282
rect 36912 4218 36964 4224
rect 34612 4072 34664 4078
rect 34612 4014 34664 4020
rect 30012 3936 30064 3942
rect 30012 3878 30064 3884
rect 56140 3936 56192 3942
rect 56140 3878 56192 3884
rect 56324 3936 56376 3942
rect 56324 3878 56376 3884
rect 56968 3936 57020 3942
rect 56968 3878 57020 3884
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 41144 3664 41196 3670
rect 41144 3606 41196 3612
rect 28724 3528 28776 3534
rect 28724 3470 28776 3476
rect 29828 3528 29880 3534
rect 29828 3470 29880 3476
rect 30656 3528 30708 3534
rect 30656 3470 30708 3476
rect 31484 3528 31536 3534
rect 31484 3470 31536 3476
rect 32312 3528 32364 3534
rect 32312 3470 32364 3476
rect 33140 3528 33192 3534
rect 33140 3470 33192 3476
rect 39212 3528 39264 3534
rect 39212 3470 39264 3476
rect 40040 3528 40092 3534
rect 40040 3470 40092 3476
rect 40868 3528 40920 3534
rect 40868 3470 40920 3476
rect 27896 2848 27948 2854
rect 27896 2790 27948 2796
rect 28448 2848 28500 2854
rect 28448 2790 28500 2796
rect 27712 2304 27764 2310
rect 27712 2246 27764 2252
rect 27908 800 27936 2790
rect 28172 2440 28224 2446
rect 28172 2382 28224 2388
rect 28184 800 28212 2382
rect 28460 800 28488 2790
rect 28736 800 28764 3470
rect 29276 2848 29328 2854
rect 29276 2790 29328 2796
rect 29000 2576 29052 2582
rect 29000 2518 29052 2524
rect 29012 800 29040 2518
rect 29288 800 29316 2790
rect 29552 2440 29604 2446
rect 29552 2382 29604 2388
rect 29564 800 29592 2382
rect 29840 800 29868 3470
rect 30104 2848 30156 2854
rect 30104 2790 30156 2796
rect 30380 2848 30432 2854
rect 30380 2790 30432 2796
rect 30116 800 30144 2790
rect 30392 800 30420 2790
rect 30668 800 30696 3470
rect 31208 2848 31260 2854
rect 31208 2790 31260 2796
rect 30932 2576 30984 2582
rect 30932 2518 30984 2524
rect 30944 800 30972 2518
rect 31220 800 31248 2790
rect 31496 800 31524 3470
rect 32036 2848 32088 2854
rect 32036 2790 32088 2796
rect 31760 2372 31812 2378
rect 31760 2314 31812 2320
rect 31772 800 31800 2314
rect 32048 800 32076 2790
rect 32324 800 32352 3470
rect 32864 2848 32916 2854
rect 32864 2790 32916 2796
rect 32588 2440 32640 2446
rect 32588 2382 32640 2388
rect 32600 800 32628 2382
rect 32876 800 32904 2790
rect 33152 800 33180 3470
rect 37280 2984 37332 2990
rect 37280 2926 37332 2932
rect 33692 2848 33744 2854
rect 33692 2790 33744 2796
rect 34244 2848 34296 2854
rect 34244 2790 34296 2796
rect 34520 2848 34572 2854
rect 34520 2790 34572 2796
rect 35348 2848 35400 2854
rect 35348 2790 35400 2796
rect 36176 2848 36228 2854
rect 36176 2790 36228 2796
rect 36728 2848 36780 2854
rect 36728 2790 36780 2796
rect 33416 2440 33468 2446
rect 33416 2382 33468 2388
rect 33428 800 33456 2382
rect 33704 800 33732 2790
rect 33968 2440 34020 2446
rect 33968 2382 34020 2388
rect 33980 800 34008 2382
rect 34256 800 34284 2790
rect 34532 800 34560 2790
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 34796 2440 34848 2446
rect 34796 2382 34848 2388
rect 35072 2440 35124 2446
rect 35072 2382 35124 2388
rect 34808 800 34836 2382
rect 35084 800 35112 2382
rect 35360 800 35388 2790
rect 35624 2440 35676 2446
rect 35624 2382 35676 2388
rect 35900 2440 35952 2446
rect 35900 2382 35952 2388
rect 35636 800 35664 2382
rect 35912 800 35940 2382
rect 36188 800 36216 2790
rect 36452 2440 36504 2446
rect 36452 2382 36504 2388
rect 36464 800 36492 2382
rect 36740 800 36768 2790
rect 37004 2508 37056 2514
rect 37004 2450 37056 2456
rect 37016 800 37044 2450
rect 37292 800 37320 2926
rect 38384 2916 38436 2922
rect 38384 2858 38436 2864
rect 37832 2848 37884 2854
rect 37832 2790 37884 2796
rect 37556 2440 37608 2446
rect 37556 2382 37608 2388
rect 37568 800 37596 2382
rect 37844 800 37872 2790
rect 38108 2508 38160 2514
rect 38108 2450 38160 2456
rect 38120 800 38148 2450
rect 38396 800 38424 2858
rect 38936 2848 38988 2854
rect 38936 2790 38988 2796
rect 38660 2440 38712 2446
rect 38660 2382 38712 2388
rect 38672 800 38700 2382
rect 38948 800 38976 2790
rect 39224 800 39252 3470
rect 39764 2916 39816 2922
rect 39764 2858 39816 2864
rect 39488 2372 39540 2378
rect 39488 2314 39540 2320
rect 39500 800 39528 2314
rect 39776 800 39804 2858
rect 40052 800 40080 3470
rect 40316 2848 40368 2854
rect 40316 2790 40368 2796
rect 40328 800 40356 2790
rect 40592 2576 40644 2582
rect 40592 2518 40644 2524
rect 40604 800 40632 2518
rect 40880 800 40908 3470
rect 41156 800 41184 3606
rect 55772 3596 55824 3602
rect 55772 3538 55824 3544
rect 42524 3528 42576 3534
rect 42524 3470 42576 3476
rect 43076 3528 43128 3534
rect 43076 3470 43128 3476
rect 45008 3528 45060 3534
rect 45008 3470 45060 3476
rect 45284 3528 45336 3534
rect 45284 3470 45336 3476
rect 46112 3528 46164 3534
rect 46112 3470 46164 3476
rect 46940 3528 46992 3534
rect 46940 3470 46992 3476
rect 47768 3528 47820 3534
rect 47768 3470 47820 3476
rect 48872 3528 48924 3534
rect 48872 3470 48924 3476
rect 50160 3528 50212 3534
rect 50160 3470 50212 3476
rect 50804 3528 50856 3534
rect 50804 3470 50856 3476
rect 51356 3528 51408 3534
rect 51356 3470 51408 3476
rect 52736 3528 52788 3534
rect 52736 3470 52788 3476
rect 53012 3528 53064 3534
rect 53012 3470 53064 3476
rect 54668 3528 54720 3534
rect 54668 3470 54720 3476
rect 55496 3528 55548 3534
rect 55496 3470 55548 3476
rect 42248 2916 42300 2922
rect 42248 2858 42300 2864
rect 41696 2848 41748 2854
rect 41696 2790 41748 2796
rect 41420 2508 41472 2514
rect 41420 2450 41472 2456
rect 41432 800 41460 2450
rect 41708 800 41736 2790
rect 41972 2440 42024 2446
rect 41972 2382 42024 2388
rect 41984 800 42012 2382
rect 42260 800 42288 2858
rect 42536 800 42564 3470
rect 42800 2848 42852 2854
rect 42800 2790 42852 2796
rect 42812 800 42840 2790
rect 43088 800 43116 3470
rect 44732 2984 44784 2990
rect 44732 2926 44784 2932
rect 43628 2916 43680 2922
rect 43628 2858 43680 2864
rect 43352 2508 43404 2514
rect 43352 2450 43404 2456
rect 43364 800 43392 2450
rect 43640 800 43668 2858
rect 44180 2848 44232 2854
rect 44180 2790 44232 2796
rect 43904 2372 43956 2378
rect 43904 2314 43956 2320
rect 43916 800 43944 2314
rect 44192 800 44220 2790
rect 44456 2576 44508 2582
rect 44456 2518 44508 2524
rect 44468 800 44496 2518
rect 44744 800 44772 2926
rect 45020 800 45048 3470
rect 45296 800 45324 3470
rect 45560 2848 45612 2854
rect 45560 2790 45612 2796
rect 45572 800 45600 2790
rect 45836 2440 45888 2446
rect 45836 2382 45888 2388
rect 45848 800 45876 2382
rect 46124 800 46152 3470
rect 46664 2848 46716 2854
rect 46664 2790 46716 2796
rect 46388 2508 46440 2514
rect 46388 2450 46440 2456
rect 46400 800 46428 2450
rect 46676 800 46704 2790
rect 46952 800 46980 3470
rect 47492 2916 47544 2922
rect 47492 2858 47544 2864
rect 47216 2372 47268 2378
rect 47216 2314 47268 2320
rect 47228 800 47256 2314
rect 47504 800 47532 2858
rect 47780 800 47808 3470
rect 48596 2984 48648 2990
rect 48596 2926 48648 2932
rect 48044 2848 48096 2854
rect 48044 2790 48096 2796
rect 48056 800 48084 2790
rect 48320 2576 48372 2582
rect 48320 2518 48372 2524
rect 48332 800 48360 2518
rect 48608 800 48636 2926
rect 48884 800 48912 3470
rect 49424 2916 49476 2922
rect 49424 2858 49476 2864
rect 49148 2508 49200 2514
rect 49148 2450 49200 2456
rect 49160 800 49188 2450
rect 49436 800 49464 2858
rect 49976 2848 50028 2854
rect 49976 2790 50028 2796
rect 49700 2440 49752 2446
rect 49700 2382 49752 2388
rect 49712 800 49740 2382
rect 49988 800 50016 2790
rect 50172 1850 50200 3470
rect 50294 3292 50602 3301
rect 50294 3290 50300 3292
rect 50356 3290 50380 3292
rect 50436 3290 50460 3292
rect 50516 3290 50540 3292
rect 50596 3290 50602 3292
rect 50356 3238 50358 3290
rect 50538 3238 50540 3290
rect 50294 3236 50300 3238
rect 50356 3236 50380 3238
rect 50436 3236 50460 3238
rect 50516 3236 50540 3238
rect 50596 3236 50602 3238
rect 50294 3227 50602 3236
rect 50620 2916 50672 2922
rect 50620 2858 50672 2864
rect 50294 2204 50602 2213
rect 50294 2202 50300 2204
rect 50356 2202 50380 2204
rect 50436 2202 50460 2204
rect 50516 2202 50540 2204
rect 50596 2202 50602 2204
rect 50356 2150 50358 2202
rect 50538 2150 50540 2202
rect 50294 2148 50300 2150
rect 50356 2148 50380 2150
rect 50436 2148 50460 2150
rect 50516 2148 50540 2150
rect 50596 2148 50602 2150
rect 50294 2139 50602 2148
rect 50172 1822 50292 1850
rect 50264 800 50292 1822
rect 50632 1442 50660 2858
rect 50540 1414 50660 1442
rect 50540 800 50568 1414
rect 50816 800 50844 3470
rect 51080 2508 51132 2514
rect 51080 2450 51132 2456
rect 51092 800 51120 2450
rect 51368 800 51396 3470
rect 52460 2984 52512 2990
rect 52460 2926 52512 2932
rect 51908 2848 51960 2854
rect 51908 2790 51960 2796
rect 51632 2440 51684 2446
rect 51632 2382 51684 2388
rect 51644 800 51672 2382
rect 51920 800 51948 2790
rect 52184 2576 52236 2582
rect 52184 2518 52236 2524
rect 52196 800 52224 2518
rect 52472 800 52500 2926
rect 52748 800 52776 3470
rect 53024 800 53052 3470
rect 53564 2984 53616 2990
rect 53564 2926 53616 2932
rect 53288 2916 53340 2922
rect 53288 2858 53340 2864
rect 53300 800 53328 2858
rect 53576 800 53604 2926
rect 54392 2916 54444 2922
rect 54392 2858 54444 2864
rect 53840 2848 53892 2854
rect 53840 2790 53892 2796
rect 53852 800 53880 2790
rect 54116 2372 54168 2378
rect 54116 2314 54168 2320
rect 54128 800 54156 2314
rect 54404 800 54432 2858
rect 54680 800 54708 3470
rect 55220 2984 55272 2990
rect 55220 2926 55272 2932
rect 55232 2650 55260 2926
rect 55404 2848 55456 2854
rect 55404 2790 55456 2796
rect 55220 2644 55272 2650
rect 55220 2586 55272 2592
rect 54944 2508 54996 2514
rect 54944 2450 54996 2456
rect 54956 800 54984 2450
rect 55416 1442 55444 2790
rect 55232 1414 55444 1442
rect 55232 800 55260 1414
rect 55508 800 55536 3470
rect 55680 2916 55732 2922
rect 55680 2858 55732 2864
rect 55692 800 55720 2858
rect 55784 800 55812 3538
rect 55956 3188 56008 3194
rect 55956 3130 56008 3136
rect 55864 2576 55916 2582
rect 55864 2518 55916 2524
rect 55876 800 55904 2518
rect 55968 800 55996 3130
rect 56048 2848 56100 2854
rect 56048 2790 56100 2796
rect 56060 800 56088 2790
rect 56152 800 56180 3878
rect 56232 3528 56284 3534
rect 56232 3470 56284 3476
rect 56244 800 56272 3470
rect 56336 800 56364 3878
rect 56508 3664 56560 3670
rect 56508 3606 56560 3612
rect 56416 2440 56468 2446
rect 56416 2382 56468 2388
rect 56428 800 56456 2382
rect 56520 800 56548 3606
rect 56784 3596 56836 3602
rect 56784 3538 56836 3544
rect 56692 2984 56744 2990
rect 56692 2926 56744 2932
rect 56704 1442 56732 2926
rect 56612 1414 56732 1442
rect 56612 800 56640 1414
rect 56796 1306 56824 3538
rect 56876 2304 56928 2310
rect 56876 2246 56928 2252
rect 56704 1278 56824 1306
rect 56704 800 56732 1278
rect 56784 1216 56836 1222
rect 56784 1158 56836 1164
rect 56796 800 56824 1158
rect 56888 800 56916 2246
rect 56980 800 57008 3878
rect 57060 2916 57112 2922
rect 57060 2858 57112 2864
rect 57072 1222 57100 2858
rect 57060 1216 57112 1222
rect 57060 1158 57112 1164
rect 57060 1080 57112 1086
rect 57060 1022 57112 1028
rect 57072 800 57100 1022
rect 57164 800 57192 4558
rect 57256 800 57284 4694
rect 57612 4616 57664 4622
rect 57612 4558 57664 4564
rect 57520 4004 57572 4010
rect 57520 3946 57572 3952
rect 57336 3528 57388 3534
rect 57336 3470 57388 3476
rect 57348 800 57376 3470
rect 57428 2644 57480 2650
rect 57428 2586 57480 2592
rect 57440 800 57468 2586
rect 57532 800 57560 3946
rect 57624 800 57652 4558
rect 57980 4140 58032 4146
rect 57980 4082 58032 4088
rect 57796 3732 57848 3738
rect 57796 3674 57848 3680
rect 57704 3120 57756 3126
rect 57704 3062 57756 3068
rect 57716 800 57744 3062
rect 57808 800 57836 3674
rect 57886 3224 57942 3233
rect 57886 3159 57942 3168
rect 57900 800 57928 3159
rect 57992 800 58020 4082
rect 58072 3936 58124 3942
rect 58072 3878 58124 3884
rect 58084 3738 58112 3878
rect 58072 3732 58124 3738
rect 58072 3674 58124 3680
rect 58072 3188 58124 3194
rect 58072 3130 58124 3136
rect 58084 2582 58112 3130
rect 58164 3052 58216 3058
rect 58164 2994 58216 3000
rect 58072 2576 58124 2582
rect 58072 2518 58124 2524
rect 58072 2100 58124 2106
rect 58072 2042 58124 2048
rect 58084 800 58112 2042
rect 58176 800 58204 2994
rect 58268 800 58296 4694
rect 58624 4004 58676 4010
rect 58624 3946 58676 3952
rect 58348 3664 58400 3670
rect 58348 3606 58400 3612
rect 58360 800 58388 3606
rect 58440 2984 58492 2990
rect 58440 2926 58492 2932
rect 58452 800 58480 2926
rect 58532 1964 58584 1970
rect 58532 1906 58584 1912
rect 58544 800 58572 1906
rect 58636 800 58664 3946
rect 58728 800 58756 4966
rect 58820 800 58848 5102
rect 59268 5092 59320 5098
rect 59268 5034 59320 5040
rect 58900 4684 58952 4690
rect 58900 4626 58952 4632
rect 58912 800 58940 4626
rect 59176 4072 59228 4078
rect 59176 4014 59228 4020
rect 58992 3596 59044 3602
rect 58992 3538 59044 3544
rect 59004 800 59032 3538
rect 59084 2032 59136 2038
rect 59084 1974 59136 1980
rect 59096 800 59124 1974
rect 59188 800 59216 4014
rect 59280 800 59308 5034
rect 65654 4924 65962 4933
rect 65654 4922 65660 4924
rect 65716 4922 65740 4924
rect 65796 4922 65820 4924
rect 65876 4922 65900 4924
rect 65956 4922 65962 4924
rect 65716 4870 65718 4922
rect 65898 4870 65900 4922
rect 65654 4868 65660 4870
rect 65716 4868 65740 4870
rect 65796 4868 65820 4870
rect 65876 4868 65900 4870
rect 65956 4868 65962 4870
rect 65654 4859 65962 4868
rect 67640 3936 67692 3942
rect 67640 3878 67692 3884
rect 65654 3836 65962 3845
rect 65654 3834 65660 3836
rect 65716 3834 65740 3836
rect 65796 3834 65820 3836
rect 65876 3834 65900 3836
rect 65956 3834 65962 3836
rect 65716 3782 65718 3834
rect 65898 3782 65900 3834
rect 65654 3780 65660 3782
rect 65716 3780 65740 3782
rect 65796 3780 65820 3782
rect 65876 3780 65900 3782
rect 65956 3780 65962 3782
rect 65654 3771 65962 3780
rect 67652 3777 67680 3878
rect 67638 3768 67694 3777
rect 67638 3703 67694 3712
rect 60464 3528 60516 3534
rect 60464 3470 60516 3476
rect 60476 3233 60504 3470
rect 60462 3224 60518 3233
rect 60462 3159 60518 3168
rect 60464 3120 60516 3126
rect 60464 3062 60516 3068
rect 59360 2916 59412 2922
rect 59360 2858 59412 2864
rect 59372 800 59400 2858
rect 60476 2854 60504 3062
rect 59452 2848 59504 2854
rect 59452 2790 59504 2796
rect 60464 2848 60516 2854
rect 60464 2790 60516 2796
rect 59464 1086 59492 2790
rect 65654 2748 65962 2757
rect 65654 2746 65660 2748
rect 65716 2746 65740 2748
rect 65796 2746 65820 2748
rect 65876 2746 65900 2748
rect 65956 2746 65962 2748
rect 65716 2694 65718 2746
rect 65898 2694 65900 2746
rect 65654 2692 65660 2694
rect 65716 2692 65740 2694
rect 65796 2692 65820 2694
rect 65876 2692 65900 2694
rect 65956 2692 65962 2694
rect 65654 2683 65962 2692
rect 63684 2508 63736 2514
rect 63684 2450 63736 2456
rect 61752 2440 61804 2446
rect 61752 2382 61804 2388
rect 63040 2440 63092 2446
rect 63040 2382 63092 2388
rect 61764 2106 61792 2382
rect 61752 2100 61804 2106
rect 61752 2042 61804 2048
rect 63052 1970 63080 2382
rect 63696 2038 63724 2450
rect 67640 2440 67692 2446
rect 67640 2382 67692 2388
rect 67652 2281 67680 2382
rect 67638 2272 67694 2281
rect 67638 2207 67694 2216
rect 63684 2032 63736 2038
rect 63684 1974 63736 1980
rect 63040 1964 63092 1970
rect 63040 1906 63092 1912
rect 59452 1080 59504 1086
rect 59452 1022 59504 1028
rect 10598 0 10654 800
rect 10690 0 10746 800
rect 10782 0 10838 800
rect 10874 0 10930 800
rect 10966 0 11022 800
rect 11058 0 11114 800
rect 11150 0 11206 800
rect 11242 0 11298 800
rect 11334 0 11390 800
rect 11426 0 11482 800
rect 11518 0 11574 800
rect 11610 0 11666 800
rect 11702 0 11758 800
rect 11794 0 11850 800
rect 11886 0 11942 800
rect 11978 0 12034 800
rect 12070 0 12126 800
rect 12162 0 12218 800
rect 12254 0 12310 800
rect 12346 0 12402 800
rect 12438 0 12494 800
rect 12530 0 12586 800
rect 12622 0 12678 800
rect 12714 0 12770 800
rect 12806 0 12862 800
rect 12898 0 12954 800
rect 12990 0 13046 800
rect 13082 0 13138 800
rect 13174 0 13230 800
rect 13266 0 13322 800
rect 13358 0 13414 800
rect 13450 0 13506 800
rect 13542 0 13598 800
rect 13634 0 13690 800
rect 13726 0 13782 800
rect 13818 0 13874 800
rect 13910 0 13966 800
rect 14002 0 14058 800
rect 14094 0 14150 800
rect 14186 0 14242 800
rect 14278 0 14334 800
rect 14370 0 14426 800
rect 14462 0 14518 800
rect 14554 0 14610 800
rect 14646 0 14702 800
rect 14738 0 14794 800
rect 14830 0 14886 800
rect 14922 0 14978 800
rect 15014 0 15070 800
rect 15106 0 15162 800
rect 15198 0 15254 800
rect 15290 0 15346 800
rect 15382 0 15438 800
rect 15474 0 15530 800
rect 15566 0 15622 800
rect 15658 0 15714 800
rect 15750 0 15806 800
rect 15842 0 15898 800
rect 15934 0 15990 800
rect 16026 0 16082 800
rect 16118 0 16174 800
rect 16210 0 16266 800
rect 16302 0 16358 800
rect 16394 0 16450 800
rect 16486 0 16542 800
rect 16578 0 16634 800
rect 16670 0 16726 800
rect 16762 0 16818 800
rect 16854 0 16910 800
rect 16946 0 17002 800
rect 17038 0 17094 800
rect 17130 0 17186 800
rect 17222 0 17278 800
rect 17314 0 17370 800
rect 17406 0 17462 800
rect 17498 0 17554 800
rect 17590 0 17646 800
rect 17682 0 17738 800
rect 17774 0 17830 800
rect 17866 0 17922 800
rect 17958 0 18014 800
rect 18050 0 18106 800
rect 18142 0 18198 800
rect 18234 0 18290 800
rect 18326 0 18382 800
rect 18418 0 18474 800
rect 18510 0 18566 800
rect 18602 0 18658 800
rect 18694 0 18750 800
rect 18786 0 18842 800
rect 18878 0 18934 800
rect 18970 0 19026 800
rect 19062 0 19118 800
rect 19154 0 19210 800
rect 19246 0 19302 800
rect 19338 0 19394 800
rect 19430 0 19486 800
rect 19522 0 19578 800
rect 19614 0 19670 800
rect 19706 0 19762 800
rect 19798 0 19854 800
rect 19890 0 19946 800
rect 19982 0 20038 800
rect 20074 0 20130 800
rect 20166 0 20222 800
rect 20258 0 20314 800
rect 20350 0 20406 800
rect 20442 0 20498 800
rect 20534 0 20590 800
rect 20626 0 20682 800
rect 20718 0 20774 800
rect 20810 0 20866 800
rect 20902 0 20958 800
rect 20994 0 21050 800
rect 21086 0 21142 800
rect 21178 0 21234 800
rect 21270 0 21326 800
rect 21362 0 21418 800
rect 21454 0 21510 800
rect 21546 0 21602 800
rect 21638 0 21694 800
rect 21730 0 21786 800
rect 21822 0 21878 800
rect 21914 0 21970 800
rect 22006 0 22062 800
rect 22098 0 22154 800
rect 22190 0 22246 800
rect 22282 0 22338 800
rect 22374 0 22430 800
rect 22466 0 22522 800
rect 22558 0 22614 800
rect 22650 0 22706 800
rect 22742 0 22798 800
rect 22834 0 22890 800
rect 22926 0 22982 800
rect 23018 0 23074 800
rect 23110 0 23166 800
rect 23202 0 23258 800
rect 23294 0 23350 800
rect 23386 0 23442 800
rect 23478 0 23534 800
rect 23570 0 23626 800
rect 23662 0 23718 800
rect 23754 0 23810 800
rect 23846 0 23902 800
rect 23938 0 23994 800
rect 24030 0 24086 800
rect 24122 0 24178 800
rect 24214 0 24270 800
rect 24306 0 24362 800
rect 24398 0 24454 800
rect 24490 0 24546 800
rect 24582 0 24638 800
rect 24674 0 24730 800
rect 24766 0 24822 800
rect 24858 0 24914 800
rect 24950 0 25006 800
rect 25042 0 25098 800
rect 25134 0 25190 800
rect 25226 0 25282 800
rect 25318 0 25374 800
rect 25410 0 25466 800
rect 25502 0 25558 800
rect 25594 0 25650 800
rect 25686 0 25742 800
rect 25778 0 25834 800
rect 25870 0 25926 800
rect 25962 0 26018 800
rect 26054 0 26110 800
rect 26146 0 26202 800
rect 26238 0 26294 800
rect 26330 0 26386 800
rect 26422 0 26478 800
rect 26514 0 26570 800
rect 26606 0 26662 800
rect 26698 0 26754 800
rect 26790 0 26846 800
rect 26882 0 26938 800
rect 26974 0 27030 800
rect 27066 0 27122 800
rect 27158 0 27214 800
rect 27250 0 27306 800
rect 27342 0 27398 800
rect 27434 0 27490 800
rect 27526 0 27582 800
rect 27618 0 27674 800
rect 27710 0 27766 800
rect 27802 0 27858 800
rect 27894 0 27950 800
rect 27986 0 28042 800
rect 28078 0 28134 800
rect 28170 0 28226 800
rect 28262 0 28318 800
rect 28354 0 28410 800
rect 28446 0 28502 800
rect 28538 0 28594 800
rect 28630 0 28686 800
rect 28722 0 28778 800
rect 28814 0 28870 800
rect 28906 0 28962 800
rect 28998 0 29054 800
rect 29090 0 29146 800
rect 29182 0 29238 800
rect 29274 0 29330 800
rect 29366 0 29422 800
rect 29458 0 29514 800
rect 29550 0 29606 800
rect 29642 0 29698 800
rect 29734 0 29790 800
rect 29826 0 29882 800
rect 29918 0 29974 800
rect 30010 0 30066 800
rect 30102 0 30158 800
rect 30194 0 30250 800
rect 30286 0 30342 800
rect 30378 0 30434 800
rect 30470 0 30526 800
rect 30562 0 30618 800
rect 30654 0 30710 800
rect 30746 0 30802 800
rect 30838 0 30894 800
rect 30930 0 30986 800
rect 31022 0 31078 800
rect 31114 0 31170 800
rect 31206 0 31262 800
rect 31298 0 31354 800
rect 31390 0 31446 800
rect 31482 0 31538 800
rect 31574 0 31630 800
rect 31666 0 31722 800
rect 31758 0 31814 800
rect 31850 0 31906 800
rect 31942 0 31998 800
rect 32034 0 32090 800
rect 32126 0 32182 800
rect 32218 0 32274 800
rect 32310 0 32366 800
rect 32402 0 32458 800
rect 32494 0 32550 800
rect 32586 0 32642 800
rect 32678 0 32734 800
rect 32770 0 32826 800
rect 32862 0 32918 800
rect 32954 0 33010 800
rect 33046 0 33102 800
rect 33138 0 33194 800
rect 33230 0 33286 800
rect 33322 0 33378 800
rect 33414 0 33470 800
rect 33506 0 33562 800
rect 33598 0 33654 800
rect 33690 0 33746 800
rect 33782 0 33838 800
rect 33874 0 33930 800
rect 33966 0 34022 800
rect 34058 0 34114 800
rect 34150 0 34206 800
rect 34242 0 34298 800
rect 34334 0 34390 800
rect 34426 0 34482 800
rect 34518 0 34574 800
rect 34610 0 34666 800
rect 34702 0 34758 800
rect 34794 0 34850 800
rect 34886 0 34942 800
rect 34978 0 35034 800
rect 35070 0 35126 800
rect 35162 0 35218 800
rect 35254 0 35310 800
rect 35346 0 35402 800
rect 35438 0 35494 800
rect 35530 0 35586 800
rect 35622 0 35678 800
rect 35714 0 35770 800
rect 35806 0 35862 800
rect 35898 0 35954 800
rect 35990 0 36046 800
rect 36082 0 36138 800
rect 36174 0 36230 800
rect 36266 0 36322 800
rect 36358 0 36414 800
rect 36450 0 36506 800
rect 36542 0 36598 800
rect 36634 0 36690 800
rect 36726 0 36782 800
rect 36818 0 36874 800
rect 36910 0 36966 800
rect 37002 0 37058 800
rect 37094 0 37150 800
rect 37186 0 37242 800
rect 37278 0 37334 800
rect 37370 0 37426 800
rect 37462 0 37518 800
rect 37554 0 37610 800
rect 37646 0 37702 800
rect 37738 0 37794 800
rect 37830 0 37886 800
rect 37922 0 37978 800
rect 38014 0 38070 800
rect 38106 0 38162 800
rect 38198 0 38254 800
rect 38290 0 38346 800
rect 38382 0 38438 800
rect 38474 0 38530 800
rect 38566 0 38622 800
rect 38658 0 38714 800
rect 38750 0 38806 800
rect 38842 0 38898 800
rect 38934 0 38990 800
rect 39026 0 39082 800
rect 39118 0 39174 800
rect 39210 0 39266 800
rect 39302 0 39358 800
rect 39394 0 39450 800
rect 39486 0 39542 800
rect 39578 0 39634 800
rect 39670 0 39726 800
rect 39762 0 39818 800
rect 39854 0 39910 800
rect 39946 0 40002 800
rect 40038 0 40094 800
rect 40130 0 40186 800
rect 40222 0 40278 800
rect 40314 0 40370 800
rect 40406 0 40462 800
rect 40498 0 40554 800
rect 40590 0 40646 800
rect 40682 0 40738 800
rect 40774 0 40830 800
rect 40866 0 40922 800
rect 40958 0 41014 800
rect 41050 0 41106 800
rect 41142 0 41198 800
rect 41234 0 41290 800
rect 41326 0 41382 800
rect 41418 0 41474 800
rect 41510 0 41566 800
rect 41602 0 41658 800
rect 41694 0 41750 800
rect 41786 0 41842 800
rect 41878 0 41934 800
rect 41970 0 42026 800
rect 42062 0 42118 800
rect 42154 0 42210 800
rect 42246 0 42302 800
rect 42338 0 42394 800
rect 42430 0 42486 800
rect 42522 0 42578 800
rect 42614 0 42670 800
rect 42706 0 42762 800
rect 42798 0 42854 800
rect 42890 0 42946 800
rect 42982 0 43038 800
rect 43074 0 43130 800
rect 43166 0 43222 800
rect 43258 0 43314 800
rect 43350 0 43406 800
rect 43442 0 43498 800
rect 43534 0 43590 800
rect 43626 0 43682 800
rect 43718 0 43774 800
rect 43810 0 43866 800
rect 43902 0 43958 800
rect 43994 0 44050 800
rect 44086 0 44142 800
rect 44178 0 44234 800
rect 44270 0 44326 800
rect 44362 0 44418 800
rect 44454 0 44510 800
rect 44546 0 44602 800
rect 44638 0 44694 800
rect 44730 0 44786 800
rect 44822 0 44878 800
rect 44914 0 44970 800
rect 45006 0 45062 800
rect 45098 0 45154 800
rect 45190 0 45246 800
rect 45282 0 45338 800
rect 45374 0 45430 800
rect 45466 0 45522 800
rect 45558 0 45614 800
rect 45650 0 45706 800
rect 45742 0 45798 800
rect 45834 0 45890 800
rect 45926 0 45982 800
rect 46018 0 46074 800
rect 46110 0 46166 800
rect 46202 0 46258 800
rect 46294 0 46350 800
rect 46386 0 46442 800
rect 46478 0 46534 800
rect 46570 0 46626 800
rect 46662 0 46718 800
rect 46754 0 46810 800
rect 46846 0 46902 800
rect 46938 0 46994 800
rect 47030 0 47086 800
rect 47122 0 47178 800
rect 47214 0 47270 800
rect 47306 0 47362 800
rect 47398 0 47454 800
rect 47490 0 47546 800
rect 47582 0 47638 800
rect 47674 0 47730 800
rect 47766 0 47822 800
rect 47858 0 47914 800
rect 47950 0 48006 800
rect 48042 0 48098 800
rect 48134 0 48190 800
rect 48226 0 48282 800
rect 48318 0 48374 800
rect 48410 0 48466 800
rect 48502 0 48558 800
rect 48594 0 48650 800
rect 48686 0 48742 800
rect 48778 0 48834 800
rect 48870 0 48926 800
rect 48962 0 49018 800
rect 49054 0 49110 800
rect 49146 0 49202 800
rect 49238 0 49294 800
rect 49330 0 49386 800
rect 49422 0 49478 800
rect 49514 0 49570 800
rect 49606 0 49662 800
rect 49698 0 49754 800
rect 49790 0 49846 800
rect 49882 0 49938 800
rect 49974 0 50030 800
rect 50066 0 50122 800
rect 50158 0 50214 800
rect 50250 0 50306 800
rect 50342 0 50398 800
rect 50434 0 50490 800
rect 50526 0 50582 800
rect 50618 0 50674 800
rect 50710 0 50766 800
rect 50802 0 50858 800
rect 50894 0 50950 800
rect 50986 0 51042 800
rect 51078 0 51134 800
rect 51170 0 51226 800
rect 51262 0 51318 800
rect 51354 0 51410 800
rect 51446 0 51502 800
rect 51538 0 51594 800
rect 51630 0 51686 800
rect 51722 0 51778 800
rect 51814 0 51870 800
rect 51906 0 51962 800
rect 51998 0 52054 800
rect 52090 0 52146 800
rect 52182 0 52238 800
rect 52274 0 52330 800
rect 52366 0 52422 800
rect 52458 0 52514 800
rect 52550 0 52606 800
rect 52642 0 52698 800
rect 52734 0 52790 800
rect 52826 0 52882 800
rect 52918 0 52974 800
rect 53010 0 53066 800
rect 53102 0 53158 800
rect 53194 0 53250 800
rect 53286 0 53342 800
rect 53378 0 53434 800
rect 53470 0 53526 800
rect 53562 0 53618 800
rect 53654 0 53710 800
rect 53746 0 53802 800
rect 53838 0 53894 800
rect 53930 0 53986 800
rect 54022 0 54078 800
rect 54114 0 54170 800
rect 54206 0 54262 800
rect 54298 0 54354 800
rect 54390 0 54446 800
rect 54482 0 54538 800
rect 54574 0 54630 800
rect 54666 0 54722 800
rect 54758 0 54814 800
rect 54850 0 54906 800
rect 54942 0 54998 800
rect 55034 0 55090 800
rect 55126 0 55182 800
rect 55218 0 55274 800
rect 55310 0 55366 800
rect 55402 0 55458 800
rect 55494 0 55550 800
rect 55586 0 55642 800
rect 55678 0 55734 800
rect 55770 0 55826 800
rect 55862 0 55918 800
rect 55954 0 56010 800
rect 56046 0 56102 800
rect 56138 0 56194 800
rect 56230 0 56286 800
rect 56322 0 56378 800
rect 56414 0 56470 800
rect 56506 0 56562 800
rect 56598 0 56654 800
rect 56690 0 56746 800
rect 56782 0 56838 800
rect 56874 0 56930 800
rect 56966 0 57022 800
rect 57058 0 57114 800
rect 57150 0 57206 800
rect 57242 0 57298 800
rect 57334 0 57390 800
rect 57426 0 57482 800
rect 57518 0 57574 800
rect 57610 0 57666 800
rect 57702 0 57758 800
rect 57794 0 57850 800
rect 57886 0 57942 800
rect 57978 0 58034 800
rect 58070 0 58126 800
rect 58162 0 58218 800
rect 58254 0 58310 800
rect 58346 0 58402 800
rect 58438 0 58494 800
rect 58530 0 58586 800
rect 58622 0 58678 800
rect 58714 0 58770 800
rect 58806 0 58862 800
rect 58898 0 58954 800
rect 58990 0 59046 800
rect 59082 0 59138 800
rect 59174 0 59230 800
rect 59266 0 59322 800
rect 59358 0 59414 800
<< via2 >>
rect 19580 57690 19636 57692
rect 19660 57690 19716 57692
rect 19740 57690 19796 57692
rect 19820 57690 19876 57692
rect 19580 57638 19626 57690
rect 19626 57638 19636 57690
rect 19660 57638 19690 57690
rect 19690 57638 19702 57690
rect 19702 57638 19716 57690
rect 19740 57638 19754 57690
rect 19754 57638 19766 57690
rect 19766 57638 19796 57690
rect 19820 57638 19830 57690
rect 19830 57638 19876 57690
rect 19580 57636 19636 57638
rect 19660 57636 19716 57638
rect 19740 57636 19796 57638
rect 19820 57636 19876 57638
rect 50300 57690 50356 57692
rect 50380 57690 50436 57692
rect 50460 57690 50516 57692
rect 50540 57690 50596 57692
rect 50300 57638 50346 57690
rect 50346 57638 50356 57690
rect 50380 57638 50410 57690
rect 50410 57638 50422 57690
rect 50422 57638 50436 57690
rect 50460 57638 50474 57690
rect 50474 57638 50486 57690
rect 50486 57638 50516 57690
rect 50540 57638 50550 57690
rect 50550 57638 50596 57690
rect 50300 57636 50356 57638
rect 50380 57636 50436 57638
rect 50460 57636 50516 57638
rect 50540 57636 50596 57638
rect 67638 57568 67694 57624
rect 4220 57146 4276 57148
rect 4300 57146 4356 57148
rect 4380 57146 4436 57148
rect 4460 57146 4516 57148
rect 4220 57094 4266 57146
rect 4266 57094 4276 57146
rect 4300 57094 4330 57146
rect 4330 57094 4342 57146
rect 4342 57094 4356 57146
rect 4380 57094 4394 57146
rect 4394 57094 4406 57146
rect 4406 57094 4436 57146
rect 4460 57094 4470 57146
rect 4470 57094 4516 57146
rect 4220 57092 4276 57094
rect 4300 57092 4356 57094
rect 4380 57092 4436 57094
rect 4460 57092 4516 57094
rect 19580 56602 19636 56604
rect 19660 56602 19716 56604
rect 19740 56602 19796 56604
rect 19820 56602 19876 56604
rect 19580 56550 19626 56602
rect 19626 56550 19636 56602
rect 19660 56550 19690 56602
rect 19690 56550 19702 56602
rect 19702 56550 19716 56602
rect 19740 56550 19754 56602
rect 19754 56550 19766 56602
rect 19766 56550 19796 56602
rect 19820 56550 19830 56602
rect 19830 56550 19876 56602
rect 19580 56548 19636 56550
rect 19660 56548 19716 56550
rect 19740 56548 19796 56550
rect 19820 56548 19876 56550
rect 4220 56058 4276 56060
rect 4300 56058 4356 56060
rect 4380 56058 4436 56060
rect 4460 56058 4516 56060
rect 4220 56006 4266 56058
rect 4266 56006 4276 56058
rect 4300 56006 4330 56058
rect 4330 56006 4342 56058
rect 4342 56006 4356 56058
rect 4380 56006 4394 56058
rect 4394 56006 4406 56058
rect 4406 56006 4436 56058
rect 4460 56006 4470 56058
rect 4470 56006 4516 56058
rect 4220 56004 4276 56006
rect 4300 56004 4356 56006
rect 4380 56004 4436 56006
rect 4460 56004 4516 56006
rect 19580 55514 19636 55516
rect 19660 55514 19716 55516
rect 19740 55514 19796 55516
rect 19820 55514 19876 55516
rect 19580 55462 19626 55514
rect 19626 55462 19636 55514
rect 19660 55462 19690 55514
rect 19690 55462 19702 55514
rect 19702 55462 19716 55514
rect 19740 55462 19754 55514
rect 19754 55462 19766 55514
rect 19766 55462 19796 55514
rect 19820 55462 19830 55514
rect 19830 55462 19876 55514
rect 19580 55460 19636 55462
rect 19660 55460 19716 55462
rect 19740 55460 19796 55462
rect 19820 55460 19876 55462
rect 4220 54970 4276 54972
rect 4300 54970 4356 54972
rect 4380 54970 4436 54972
rect 4460 54970 4516 54972
rect 4220 54918 4266 54970
rect 4266 54918 4276 54970
rect 4300 54918 4330 54970
rect 4330 54918 4342 54970
rect 4342 54918 4356 54970
rect 4380 54918 4394 54970
rect 4394 54918 4406 54970
rect 4406 54918 4436 54970
rect 4460 54918 4470 54970
rect 4470 54918 4516 54970
rect 4220 54916 4276 54918
rect 4300 54916 4356 54918
rect 4380 54916 4436 54918
rect 4460 54916 4516 54918
rect 19580 54426 19636 54428
rect 19660 54426 19716 54428
rect 19740 54426 19796 54428
rect 19820 54426 19876 54428
rect 19580 54374 19626 54426
rect 19626 54374 19636 54426
rect 19660 54374 19690 54426
rect 19690 54374 19702 54426
rect 19702 54374 19716 54426
rect 19740 54374 19754 54426
rect 19754 54374 19766 54426
rect 19766 54374 19796 54426
rect 19820 54374 19830 54426
rect 19830 54374 19876 54426
rect 19580 54372 19636 54374
rect 19660 54372 19716 54374
rect 19740 54372 19796 54374
rect 19820 54372 19876 54374
rect 4220 53882 4276 53884
rect 4300 53882 4356 53884
rect 4380 53882 4436 53884
rect 4460 53882 4516 53884
rect 4220 53830 4266 53882
rect 4266 53830 4276 53882
rect 4300 53830 4330 53882
rect 4330 53830 4342 53882
rect 4342 53830 4356 53882
rect 4380 53830 4394 53882
rect 4394 53830 4406 53882
rect 4406 53830 4436 53882
rect 4460 53830 4470 53882
rect 4470 53830 4516 53882
rect 4220 53828 4276 53830
rect 4300 53828 4356 53830
rect 4380 53828 4436 53830
rect 4460 53828 4516 53830
rect 19580 53338 19636 53340
rect 19660 53338 19716 53340
rect 19740 53338 19796 53340
rect 19820 53338 19876 53340
rect 19580 53286 19626 53338
rect 19626 53286 19636 53338
rect 19660 53286 19690 53338
rect 19690 53286 19702 53338
rect 19702 53286 19716 53338
rect 19740 53286 19754 53338
rect 19754 53286 19766 53338
rect 19766 53286 19796 53338
rect 19820 53286 19830 53338
rect 19830 53286 19876 53338
rect 19580 53284 19636 53286
rect 19660 53284 19716 53286
rect 19740 53284 19796 53286
rect 19820 53284 19876 53286
rect 4220 52794 4276 52796
rect 4300 52794 4356 52796
rect 4380 52794 4436 52796
rect 4460 52794 4516 52796
rect 4220 52742 4266 52794
rect 4266 52742 4276 52794
rect 4300 52742 4330 52794
rect 4330 52742 4342 52794
rect 4342 52742 4356 52794
rect 4380 52742 4394 52794
rect 4394 52742 4406 52794
rect 4406 52742 4436 52794
rect 4460 52742 4470 52794
rect 4470 52742 4516 52794
rect 4220 52740 4276 52742
rect 4300 52740 4356 52742
rect 4380 52740 4436 52742
rect 4460 52740 4516 52742
rect 19580 52250 19636 52252
rect 19660 52250 19716 52252
rect 19740 52250 19796 52252
rect 19820 52250 19876 52252
rect 19580 52198 19626 52250
rect 19626 52198 19636 52250
rect 19660 52198 19690 52250
rect 19690 52198 19702 52250
rect 19702 52198 19716 52250
rect 19740 52198 19754 52250
rect 19754 52198 19766 52250
rect 19766 52198 19796 52250
rect 19820 52198 19830 52250
rect 19830 52198 19876 52250
rect 19580 52196 19636 52198
rect 19660 52196 19716 52198
rect 19740 52196 19796 52198
rect 19820 52196 19876 52198
rect 4220 51706 4276 51708
rect 4300 51706 4356 51708
rect 4380 51706 4436 51708
rect 4460 51706 4516 51708
rect 4220 51654 4266 51706
rect 4266 51654 4276 51706
rect 4300 51654 4330 51706
rect 4330 51654 4342 51706
rect 4342 51654 4356 51706
rect 4380 51654 4394 51706
rect 4394 51654 4406 51706
rect 4406 51654 4436 51706
rect 4460 51654 4470 51706
rect 4470 51654 4516 51706
rect 4220 51652 4276 51654
rect 4300 51652 4356 51654
rect 4380 51652 4436 51654
rect 4460 51652 4516 51654
rect 19580 51162 19636 51164
rect 19660 51162 19716 51164
rect 19740 51162 19796 51164
rect 19820 51162 19876 51164
rect 19580 51110 19626 51162
rect 19626 51110 19636 51162
rect 19660 51110 19690 51162
rect 19690 51110 19702 51162
rect 19702 51110 19716 51162
rect 19740 51110 19754 51162
rect 19754 51110 19766 51162
rect 19766 51110 19796 51162
rect 19820 51110 19830 51162
rect 19830 51110 19876 51162
rect 19580 51108 19636 51110
rect 19660 51108 19716 51110
rect 19740 51108 19796 51110
rect 19820 51108 19876 51110
rect 4220 50618 4276 50620
rect 4300 50618 4356 50620
rect 4380 50618 4436 50620
rect 4460 50618 4516 50620
rect 4220 50566 4266 50618
rect 4266 50566 4276 50618
rect 4300 50566 4330 50618
rect 4330 50566 4342 50618
rect 4342 50566 4356 50618
rect 4380 50566 4394 50618
rect 4394 50566 4406 50618
rect 4406 50566 4436 50618
rect 4460 50566 4470 50618
rect 4470 50566 4516 50618
rect 4220 50564 4276 50566
rect 4300 50564 4356 50566
rect 4380 50564 4436 50566
rect 4460 50564 4516 50566
rect 19580 50074 19636 50076
rect 19660 50074 19716 50076
rect 19740 50074 19796 50076
rect 19820 50074 19876 50076
rect 19580 50022 19626 50074
rect 19626 50022 19636 50074
rect 19660 50022 19690 50074
rect 19690 50022 19702 50074
rect 19702 50022 19716 50074
rect 19740 50022 19754 50074
rect 19754 50022 19766 50074
rect 19766 50022 19796 50074
rect 19820 50022 19830 50074
rect 19830 50022 19876 50074
rect 19580 50020 19636 50022
rect 19660 50020 19716 50022
rect 19740 50020 19796 50022
rect 19820 50020 19876 50022
rect 4220 49530 4276 49532
rect 4300 49530 4356 49532
rect 4380 49530 4436 49532
rect 4460 49530 4516 49532
rect 4220 49478 4266 49530
rect 4266 49478 4276 49530
rect 4300 49478 4330 49530
rect 4330 49478 4342 49530
rect 4342 49478 4356 49530
rect 4380 49478 4394 49530
rect 4394 49478 4406 49530
rect 4406 49478 4436 49530
rect 4460 49478 4470 49530
rect 4470 49478 4516 49530
rect 4220 49476 4276 49478
rect 4300 49476 4356 49478
rect 4380 49476 4436 49478
rect 4460 49476 4516 49478
rect 19580 48986 19636 48988
rect 19660 48986 19716 48988
rect 19740 48986 19796 48988
rect 19820 48986 19876 48988
rect 19580 48934 19626 48986
rect 19626 48934 19636 48986
rect 19660 48934 19690 48986
rect 19690 48934 19702 48986
rect 19702 48934 19716 48986
rect 19740 48934 19754 48986
rect 19754 48934 19766 48986
rect 19766 48934 19796 48986
rect 19820 48934 19830 48986
rect 19830 48934 19876 48986
rect 19580 48932 19636 48934
rect 19660 48932 19716 48934
rect 19740 48932 19796 48934
rect 19820 48932 19876 48934
rect 4220 48442 4276 48444
rect 4300 48442 4356 48444
rect 4380 48442 4436 48444
rect 4460 48442 4516 48444
rect 4220 48390 4266 48442
rect 4266 48390 4276 48442
rect 4300 48390 4330 48442
rect 4330 48390 4342 48442
rect 4342 48390 4356 48442
rect 4380 48390 4394 48442
rect 4394 48390 4406 48442
rect 4406 48390 4436 48442
rect 4460 48390 4470 48442
rect 4470 48390 4516 48442
rect 4220 48388 4276 48390
rect 4300 48388 4356 48390
rect 4380 48388 4436 48390
rect 4460 48388 4516 48390
rect 19580 47898 19636 47900
rect 19660 47898 19716 47900
rect 19740 47898 19796 47900
rect 19820 47898 19876 47900
rect 19580 47846 19626 47898
rect 19626 47846 19636 47898
rect 19660 47846 19690 47898
rect 19690 47846 19702 47898
rect 19702 47846 19716 47898
rect 19740 47846 19754 47898
rect 19754 47846 19766 47898
rect 19766 47846 19796 47898
rect 19820 47846 19830 47898
rect 19830 47846 19876 47898
rect 19580 47844 19636 47846
rect 19660 47844 19716 47846
rect 19740 47844 19796 47846
rect 19820 47844 19876 47846
rect 4220 47354 4276 47356
rect 4300 47354 4356 47356
rect 4380 47354 4436 47356
rect 4460 47354 4516 47356
rect 4220 47302 4266 47354
rect 4266 47302 4276 47354
rect 4300 47302 4330 47354
rect 4330 47302 4342 47354
rect 4342 47302 4356 47354
rect 4380 47302 4394 47354
rect 4394 47302 4406 47354
rect 4406 47302 4436 47354
rect 4460 47302 4470 47354
rect 4470 47302 4516 47354
rect 4220 47300 4276 47302
rect 4300 47300 4356 47302
rect 4380 47300 4436 47302
rect 4460 47300 4516 47302
rect 19580 46810 19636 46812
rect 19660 46810 19716 46812
rect 19740 46810 19796 46812
rect 19820 46810 19876 46812
rect 19580 46758 19626 46810
rect 19626 46758 19636 46810
rect 19660 46758 19690 46810
rect 19690 46758 19702 46810
rect 19702 46758 19716 46810
rect 19740 46758 19754 46810
rect 19754 46758 19766 46810
rect 19766 46758 19796 46810
rect 19820 46758 19830 46810
rect 19830 46758 19876 46810
rect 19580 46756 19636 46758
rect 19660 46756 19716 46758
rect 19740 46756 19796 46758
rect 19820 46756 19876 46758
rect 4220 46266 4276 46268
rect 4300 46266 4356 46268
rect 4380 46266 4436 46268
rect 4460 46266 4516 46268
rect 4220 46214 4266 46266
rect 4266 46214 4276 46266
rect 4300 46214 4330 46266
rect 4330 46214 4342 46266
rect 4342 46214 4356 46266
rect 4380 46214 4394 46266
rect 4394 46214 4406 46266
rect 4406 46214 4436 46266
rect 4460 46214 4470 46266
rect 4470 46214 4516 46266
rect 4220 46212 4276 46214
rect 4300 46212 4356 46214
rect 4380 46212 4436 46214
rect 4460 46212 4516 46214
rect 19580 45722 19636 45724
rect 19660 45722 19716 45724
rect 19740 45722 19796 45724
rect 19820 45722 19876 45724
rect 19580 45670 19626 45722
rect 19626 45670 19636 45722
rect 19660 45670 19690 45722
rect 19690 45670 19702 45722
rect 19702 45670 19716 45722
rect 19740 45670 19754 45722
rect 19754 45670 19766 45722
rect 19766 45670 19796 45722
rect 19820 45670 19830 45722
rect 19830 45670 19876 45722
rect 19580 45668 19636 45670
rect 19660 45668 19716 45670
rect 19740 45668 19796 45670
rect 19820 45668 19876 45670
rect 4220 45178 4276 45180
rect 4300 45178 4356 45180
rect 4380 45178 4436 45180
rect 4460 45178 4516 45180
rect 4220 45126 4266 45178
rect 4266 45126 4276 45178
rect 4300 45126 4330 45178
rect 4330 45126 4342 45178
rect 4342 45126 4356 45178
rect 4380 45126 4394 45178
rect 4394 45126 4406 45178
rect 4406 45126 4436 45178
rect 4460 45126 4470 45178
rect 4470 45126 4516 45178
rect 4220 45124 4276 45126
rect 4300 45124 4356 45126
rect 4380 45124 4436 45126
rect 4460 45124 4516 45126
rect 19580 44634 19636 44636
rect 19660 44634 19716 44636
rect 19740 44634 19796 44636
rect 19820 44634 19876 44636
rect 19580 44582 19626 44634
rect 19626 44582 19636 44634
rect 19660 44582 19690 44634
rect 19690 44582 19702 44634
rect 19702 44582 19716 44634
rect 19740 44582 19754 44634
rect 19754 44582 19766 44634
rect 19766 44582 19796 44634
rect 19820 44582 19830 44634
rect 19830 44582 19876 44634
rect 19580 44580 19636 44582
rect 19660 44580 19716 44582
rect 19740 44580 19796 44582
rect 19820 44580 19876 44582
rect 4220 44090 4276 44092
rect 4300 44090 4356 44092
rect 4380 44090 4436 44092
rect 4460 44090 4516 44092
rect 4220 44038 4266 44090
rect 4266 44038 4276 44090
rect 4300 44038 4330 44090
rect 4330 44038 4342 44090
rect 4342 44038 4356 44090
rect 4380 44038 4394 44090
rect 4394 44038 4406 44090
rect 4406 44038 4436 44090
rect 4460 44038 4470 44090
rect 4470 44038 4516 44090
rect 4220 44036 4276 44038
rect 4300 44036 4356 44038
rect 4380 44036 4436 44038
rect 4460 44036 4516 44038
rect 19580 43546 19636 43548
rect 19660 43546 19716 43548
rect 19740 43546 19796 43548
rect 19820 43546 19876 43548
rect 19580 43494 19626 43546
rect 19626 43494 19636 43546
rect 19660 43494 19690 43546
rect 19690 43494 19702 43546
rect 19702 43494 19716 43546
rect 19740 43494 19754 43546
rect 19754 43494 19766 43546
rect 19766 43494 19796 43546
rect 19820 43494 19830 43546
rect 19830 43494 19876 43546
rect 19580 43492 19636 43494
rect 19660 43492 19716 43494
rect 19740 43492 19796 43494
rect 19820 43492 19876 43494
rect 4220 43002 4276 43004
rect 4300 43002 4356 43004
rect 4380 43002 4436 43004
rect 4460 43002 4516 43004
rect 4220 42950 4266 43002
rect 4266 42950 4276 43002
rect 4300 42950 4330 43002
rect 4330 42950 4342 43002
rect 4342 42950 4356 43002
rect 4380 42950 4394 43002
rect 4394 42950 4406 43002
rect 4406 42950 4436 43002
rect 4460 42950 4470 43002
rect 4470 42950 4516 43002
rect 4220 42948 4276 42950
rect 4300 42948 4356 42950
rect 4380 42948 4436 42950
rect 4460 42948 4516 42950
rect 19580 42458 19636 42460
rect 19660 42458 19716 42460
rect 19740 42458 19796 42460
rect 19820 42458 19876 42460
rect 19580 42406 19626 42458
rect 19626 42406 19636 42458
rect 19660 42406 19690 42458
rect 19690 42406 19702 42458
rect 19702 42406 19716 42458
rect 19740 42406 19754 42458
rect 19754 42406 19766 42458
rect 19766 42406 19796 42458
rect 19820 42406 19830 42458
rect 19830 42406 19876 42458
rect 19580 42404 19636 42406
rect 19660 42404 19716 42406
rect 19740 42404 19796 42406
rect 19820 42404 19876 42406
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 19580 41370 19636 41372
rect 19660 41370 19716 41372
rect 19740 41370 19796 41372
rect 19820 41370 19876 41372
rect 19580 41318 19626 41370
rect 19626 41318 19636 41370
rect 19660 41318 19690 41370
rect 19690 41318 19702 41370
rect 19702 41318 19716 41370
rect 19740 41318 19754 41370
rect 19754 41318 19766 41370
rect 19766 41318 19796 41370
rect 19820 41318 19830 41370
rect 19830 41318 19876 41370
rect 19580 41316 19636 41318
rect 19660 41316 19716 41318
rect 19740 41316 19796 41318
rect 19820 41316 19876 41318
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 19580 40282 19636 40284
rect 19660 40282 19716 40284
rect 19740 40282 19796 40284
rect 19820 40282 19876 40284
rect 19580 40230 19626 40282
rect 19626 40230 19636 40282
rect 19660 40230 19690 40282
rect 19690 40230 19702 40282
rect 19702 40230 19716 40282
rect 19740 40230 19754 40282
rect 19754 40230 19766 40282
rect 19766 40230 19796 40282
rect 19820 40230 19830 40282
rect 19830 40230 19876 40282
rect 19580 40228 19636 40230
rect 19660 40228 19716 40230
rect 19740 40228 19796 40230
rect 19820 40228 19876 40230
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 19580 39194 19636 39196
rect 19660 39194 19716 39196
rect 19740 39194 19796 39196
rect 19820 39194 19876 39196
rect 19580 39142 19626 39194
rect 19626 39142 19636 39194
rect 19660 39142 19690 39194
rect 19690 39142 19702 39194
rect 19702 39142 19716 39194
rect 19740 39142 19754 39194
rect 19754 39142 19766 39194
rect 19766 39142 19796 39194
rect 19820 39142 19830 39194
rect 19830 39142 19876 39194
rect 19580 39140 19636 39142
rect 19660 39140 19716 39142
rect 19740 39140 19796 39142
rect 19820 39140 19876 39142
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 19580 38106 19636 38108
rect 19660 38106 19716 38108
rect 19740 38106 19796 38108
rect 19820 38106 19876 38108
rect 19580 38054 19626 38106
rect 19626 38054 19636 38106
rect 19660 38054 19690 38106
rect 19690 38054 19702 38106
rect 19702 38054 19716 38106
rect 19740 38054 19754 38106
rect 19754 38054 19766 38106
rect 19766 38054 19796 38106
rect 19820 38054 19830 38106
rect 19830 38054 19876 38106
rect 19580 38052 19636 38054
rect 19660 38052 19716 38054
rect 19740 38052 19796 38054
rect 19820 38052 19876 38054
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 2502 22616 2558 22672
rect 4342 23860 4398 23896
rect 4342 23840 4344 23860
rect 4344 23840 4396 23860
rect 4396 23840 4398 23860
rect 4894 23724 4950 23760
rect 4894 23704 4896 23724
rect 4896 23704 4948 23724
rect 4948 23704 4950 23724
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 5906 22636 5962 22672
rect 5906 22616 5908 22636
rect 5908 22616 5960 22636
rect 5960 22616 5962 22636
rect 5538 20460 5594 20496
rect 5538 20440 5540 20460
rect 5540 20440 5592 20460
rect 5592 20440 5594 20460
rect 6550 21140 6606 21176
rect 6550 21120 6552 21140
rect 6552 21120 6604 21140
rect 6604 21120 6606 21140
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 5446 14864 5502 14920
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4618 12708 4674 12744
rect 4618 12688 4620 12708
rect 4620 12688 4672 12708
rect 4672 12688 4674 12708
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 3422 12144 3478 12200
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4710 10512 4766 10568
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 5722 7812 5778 7848
rect 5722 7792 5724 7812
rect 5724 7792 5776 7812
rect 5776 7792 5778 7812
rect 6090 9868 6092 9888
rect 6092 9868 6144 9888
rect 6144 9868 6146 9888
rect 6090 9832 6146 9868
rect 5906 6976 5962 7032
rect 5630 5752 5686 5808
rect 3974 5072 4030 5128
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4986 4140 5042 4176
rect 4986 4120 4988 4140
rect 4988 4120 5040 4140
rect 5040 4120 5042 4140
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4618 3712 4674 3768
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 8574 23840 8630 23896
rect 8482 23724 8538 23760
rect 8482 23704 8484 23724
rect 8484 23704 8536 23724
rect 8536 23704 8538 23724
rect 8114 20984 8170 21040
rect 6274 9696 6330 9752
rect 7746 13912 7802 13968
rect 7286 8780 7288 8800
rect 7288 8780 7340 8800
rect 7340 8780 7342 8800
rect 7286 8744 7342 8780
rect 8022 13776 8078 13832
rect 8114 9696 8170 9752
rect 8758 21140 8814 21176
rect 8758 21120 8760 21140
rect 8760 21120 8812 21140
rect 8812 21120 8814 21140
rect 9678 21428 9680 21448
rect 9680 21428 9732 21448
rect 9732 21428 9734 21448
rect 9678 21392 9734 21428
rect 9586 17040 9642 17096
rect 7838 8744 7894 8800
rect 6458 3168 6514 3224
rect 7930 8336 7986 8392
rect 8390 8336 8446 8392
rect 7286 5072 7342 5128
rect 7654 4004 7710 4040
rect 7654 3984 7656 4004
rect 7656 3984 7708 4004
rect 7708 3984 7710 4004
rect 10598 15408 10654 15464
rect 10414 14048 10470 14104
rect 9494 10668 9550 10704
rect 9494 10648 9496 10668
rect 9496 10648 9548 10668
rect 9548 10648 9550 10668
rect 9126 10512 9182 10568
rect 8114 4664 8170 4720
rect 9218 6196 9220 6216
rect 9220 6196 9272 6216
rect 9272 6196 9274 6216
rect 9218 6160 9274 6196
rect 8942 4156 8944 4176
rect 8944 4156 8996 4176
rect 8996 4156 8998 4176
rect 8942 4120 8998 4156
rect 8666 3168 8722 3224
rect 7930 2624 7986 2680
rect 6458 2080 6514 2136
rect 6734 1944 6790 2000
rect 10046 9832 10102 9888
rect 9770 4528 9826 4584
rect 9954 4528 10010 4584
rect 9310 3440 9366 3496
rect 9586 2760 9642 2816
rect 10046 2352 10102 2408
rect 9034 1808 9090 1864
rect 10782 10668 10838 10704
rect 10782 10648 10784 10668
rect 10784 10648 10836 10668
rect 10836 10648 10838 10668
rect 10322 3984 10378 4040
rect 10598 3984 10654 4040
rect 10506 3848 10562 3904
rect 10874 6024 10930 6080
rect 11702 21392 11758 21448
rect 11978 18128 12034 18184
rect 11426 16532 11428 16552
rect 11428 16532 11480 16552
rect 11480 16532 11482 16552
rect 11426 16496 11482 16532
rect 11886 15544 11942 15600
rect 11242 13232 11298 13288
rect 11058 11500 11060 11520
rect 11060 11500 11112 11520
rect 11112 11500 11114 11520
rect 11058 11464 11114 11500
rect 12622 16496 12678 16552
rect 13082 24404 13138 24440
rect 13082 24384 13084 24404
rect 13084 24384 13136 24404
rect 13136 24384 13138 24404
rect 12898 21392 12954 21448
rect 12898 13640 12954 13696
rect 12898 13368 12954 13424
rect 12530 12844 12586 12880
rect 12530 12824 12532 12844
rect 12532 12824 12584 12844
rect 12584 12824 12586 12844
rect 12806 12144 12862 12200
rect 11058 8880 11114 8936
rect 11150 8780 11152 8800
rect 11152 8780 11204 8800
rect 11204 8780 11206 8800
rect 11150 8744 11206 8780
rect 11702 7404 11758 7440
rect 11702 7384 11704 7404
rect 11704 7384 11756 7404
rect 11756 7384 11758 7404
rect 11058 6976 11114 7032
rect 11426 6840 11482 6896
rect 11978 6840 12034 6896
rect 11058 5888 11114 5944
rect 10966 4004 11022 4040
rect 10966 3984 10968 4004
rect 10968 3984 11020 4004
rect 11020 3984 11022 4004
rect 10874 3576 10930 3632
rect 10874 2080 10930 2136
rect 11334 4664 11390 4720
rect 11426 4120 11482 4176
rect 11334 3848 11390 3904
rect 11702 5092 11758 5128
rect 11702 5072 11704 5092
rect 11704 5072 11756 5092
rect 11756 5072 11758 5092
rect 11978 4936 12034 4992
rect 12162 5888 12218 5944
rect 12162 5344 12218 5400
rect 11518 2896 11574 2952
rect 11886 2760 11942 2816
rect 12622 6160 12678 6216
rect 12162 3576 12218 3632
rect 12070 2796 12072 2816
rect 12072 2796 12124 2816
rect 12124 2796 12126 2816
rect 12070 2760 12126 2796
rect 12714 1264 12770 1320
rect 12898 1264 12954 1320
rect 14186 15136 14242 15192
rect 15198 18400 15254 18456
rect 14646 14864 14702 14920
rect 14738 13912 14794 13968
rect 14646 13252 14702 13288
rect 14646 13232 14648 13252
rect 14648 13232 14700 13252
rect 14700 13232 14702 13252
rect 14922 12180 14924 12200
rect 14924 12180 14976 12200
rect 14976 12180 14978 12200
rect 14922 12144 14978 12180
rect 15106 11872 15162 11928
rect 15750 20304 15806 20360
rect 15474 17620 15476 17640
rect 15476 17620 15528 17640
rect 15528 17620 15530 17640
rect 15474 17584 15530 17620
rect 13450 6024 13506 6080
rect 15474 11736 15530 11792
rect 14094 3712 14150 3768
rect 14094 2896 14150 2952
rect 14922 5480 14978 5536
rect 15106 3612 15108 3632
rect 15108 3612 15160 3632
rect 15160 3612 15162 3632
rect 15106 3576 15162 3612
rect 15198 2896 15254 2952
rect 15382 5752 15438 5808
rect 16762 24384 16818 24440
rect 16210 18400 16266 18456
rect 16118 18284 16174 18320
rect 16118 18264 16120 18284
rect 16120 18264 16172 18284
rect 16172 18264 16174 18284
rect 16394 17584 16450 17640
rect 16026 13368 16082 13424
rect 16118 12280 16174 12336
rect 15842 7792 15898 7848
rect 16854 21140 16910 21176
rect 16854 21120 16856 21140
rect 16856 21120 16908 21140
rect 16908 21120 16910 21140
rect 17222 21120 17278 21176
rect 16670 17040 16726 17096
rect 16578 13640 16634 13696
rect 16486 13388 16542 13424
rect 16486 13368 16488 13388
rect 16488 13368 16540 13388
rect 16540 13368 16542 13388
rect 18142 21936 18198 21992
rect 16854 15444 16856 15464
rect 16856 15444 16908 15464
rect 16908 15444 16910 15464
rect 16854 15408 16910 15444
rect 17222 17040 17278 17096
rect 17038 14048 17094 14104
rect 17222 15544 17278 15600
rect 17682 16088 17738 16144
rect 18326 16496 18382 16552
rect 17406 14456 17462 14512
rect 16486 11212 16542 11248
rect 16486 11192 16488 11212
rect 16488 11192 16540 11212
rect 16540 11192 16542 11212
rect 15934 4936 15990 4992
rect 15658 3032 15714 3088
rect 15658 2080 15714 2136
rect 15842 1808 15898 1864
rect 16210 5344 16266 5400
rect 16302 3848 16358 3904
rect 16762 12008 16818 12064
rect 16762 11092 16764 11112
rect 16764 11092 16816 11112
rect 16816 11092 16818 11112
rect 16762 11056 16818 11092
rect 17130 9580 17186 9616
rect 17406 12552 17462 12608
rect 17314 11328 17370 11384
rect 17130 9560 17132 9580
rect 17132 9560 17184 9580
rect 17184 9560 17186 9580
rect 17866 12144 17922 12200
rect 17866 12044 17868 12064
rect 17868 12044 17920 12064
rect 17920 12044 17922 12064
rect 17866 12008 17922 12044
rect 18418 15036 18420 15056
rect 18420 15036 18472 15056
rect 18472 15036 18474 15056
rect 18418 15000 18474 15036
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 18878 21120 18934 21176
rect 18786 18284 18842 18320
rect 18786 18264 18788 18284
rect 18788 18264 18840 18284
rect 18840 18264 18842 18284
rect 18694 18128 18750 18184
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19614 16496 19670 16552
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19338 15136 19394 15192
rect 18510 11872 18566 11928
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19062 13232 19118 13288
rect 19154 12144 19210 12200
rect 18234 9968 18290 10024
rect 16854 6840 16910 6896
rect 17406 5480 17462 5536
rect 17314 5072 17370 5128
rect 18234 2644 18290 2680
rect 18234 2624 18236 2644
rect 18236 2624 18288 2644
rect 18288 2624 18290 2644
rect 18970 10512 19026 10568
rect 19890 13776 19946 13832
rect 19706 13504 19762 13560
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 34940 57146 34996 57148
rect 35020 57146 35076 57148
rect 35100 57146 35156 57148
rect 35180 57146 35236 57148
rect 34940 57094 34986 57146
rect 34986 57094 34996 57146
rect 35020 57094 35050 57146
rect 35050 57094 35062 57146
rect 35062 57094 35076 57146
rect 35100 57094 35114 57146
rect 35114 57094 35126 57146
rect 35126 57094 35156 57146
rect 35180 57094 35190 57146
rect 35190 57094 35236 57146
rect 34940 57092 34996 57094
rect 35020 57092 35076 57094
rect 35100 57092 35156 57094
rect 35180 57092 35236 57094
rect 34940 56058 34996 56060
rect 35020 56058 35076 56060
rect 35100 56058 35156 56060
rect 35180 56058 35236 56060
rect 34940 56006 34986 56058
rect 34986 56006 34996 56058
rect 35020 56006 35050 56058
rect 35050 56006 35062 56058
rect 35062 56006 35076 56058
rect 35100 56006 35114 56058
rect 35114 56006 35126 56058
rect 35126 56006 35156 56058
rect 35180 56006 35190 56058
rect 35190 56006 35236 56058
rect 34940 56004 34996 56006
rect 35020 56004 35076 56006
rect 35100 56004 35156 56006
rect 35180 56004 35236 56006
rect 34940 54970 34996 54972
rect 35020 54970 35076 54972
rect 35100 54970 35156 54972
rect 35180 54970 35236 54972
rect 34940 54918 34986 54970
rect 34986 54918 34996 54970
rect 35020 54918 35050 54970
rect 35050 54918 35062 54970
rect 35062 54918 35076 54970
rect 35100 54918 35114 54970
rect 35114 54918 35126 54970
rect 35126 54918 35156 54970
rect 35180 54918 35190 54970
rect 35190 54918 35236 54970
rect 34940 54916 34996 54918
rect 35020 54916 35076 54918
rect 35100 54916 35156 54918
rect 35180 54916 35236 54918
rect 34940 53882 34996 53884
rect 35020 53882 35076 53884
rect 35100 53882 35156 53884
rect 35180 53882 35236 53884
rect 34940 53830 34986 53882
rect 34986 53830 34996 53882
rect 35020 53830 35050 53882
rect 35050 53830 35062 53882
rect 35062 53830 35076 53882
rect 35100 53830 35114 53882
rect 35114 53830 35126 53882
rect 35126 53830 35156 53882
rect 35180 53830 35190 53882
rect 35190 53830 35236 53882
rect 34940 53828 34996 53830
rect 35020 53828 35076 53830
rect 35100 53828 35156 53830
rect 35180 53828 35236 53830
rect 34940 52794 34996 52796
rect 35020 52794 35076 52796
rect 35100 52794 35156 52796
rect 35180 52794 35236 52796
rect 34940 52742 34986 52794
rect 34986 52742 34996 52794
rect 35020 52742 35050 52794
rect 35050 52742 35062 52794
rect 35062 52742 35076 52794
rect 35100 52742 35114 52794
rect 35114 52742 35126 52794
rect 35126 52742 35156 52794
rect 35180 52742 35190 52794
rect 35190 52742 35236 52794
rect 34940 52740 34996 52742
rect 35020 52740 35076 52742
rect 35100 52740 35156 52742
rect 35180 52740 35236 52742
rect 34940 51706 34996 51708
rect 35020 51706 35076 51708
rect 35100 51706 35156 51708
rect 35180 51706 35236 51708
rect 34940 51654 34986 51706
rect 34986 51654 34996 51706
rect 35020 51654 35050 51706
rect 35050 51654 35062 51706
rect 35062 51654 35076 51706
rect 35100 51654 35114 51706
rect 35114 51654 35126 51706
rect 35126 51654 35156 51706
rect 35180 51654 35190 51706
rect 35190 51654 35236 51706
rect 34940 51652 34996 51654
rect 35020 51652 35076 51654
rect 35100 51652 35156 51654
rect 35180 51652 35236 51654
rect 34940 50618 34996 50620
rect 35020 50618 35076 50620
rect 35100 50618 35156 50620
rect 35180 50618 35236 50620
rect 34940 50566 34986 50618
rect 34986 50566 34996 50618
rect 35020 50566 35050 50618
rect 35050 50566 35062 50618
rect 35062 50566 35076 50618
rect 35100 50566 35114 50618
rect 35114 50566 35126 50618
rect 35126 50566 35156 50618
rect 35180 50566 35190 50618
rect 35190 50566 35236 50618
rect 34940 50564 34996 50566
rect 35020 50564 35076 50566
rect 35100 50564 35156 50566
rect 35180 50564 35236 50566
rect 34940 49530 34996 49532
rect 35020 49530 35076 49532
rect 35100 49530 35156 49532
rect 35180 49530 35236 49532
rect 34940 49478 34986 49530
rect 34986 49478 34996 49530
rect 35020 49478 35050 49530
rect 35050 49478 35062 49530
rect 35062 49478 35076 49530
rect 35100 49478 35114 49530
rect 35114 49478 35126 49530
rect 35126 49478 35156 49530
rect 35180 49478 35190 49530
rect 35190 49478 35236 49530
rect 34940 49476 34996 49478
rect 35020 49476 35076 49478
rect 35100 49476 35156 49478
rect 35180 49476 35236 49478
rect 34940 48442 34996 48444
rect 35020 48442 35076 48444
rect 35100 48442 35156 48444
rect 35180 48442 35236 48444
rect 34940 48390 34986 48442
rect 34986 48390 34996 48442
rect 35020 48390 35050 48442
rect 35050 48390 35062 48442
rect 35062 48390 35076 48442
rect 35100 48390 35114 48442
rect 35114 48390 35126 48442
rect 35126 48390 35156 48442
rect 35180 48390 35190 48442
rect 35190 48390 35236 48442
rect 34940 48388 34996 48390
rect 35020 48388 35076 48390
rect 35100 48388 35156 48390
rect 35180 48388 35236 48390
rect 34940 47354 34996 47356
rect 35020 47354 35076 47356
rect 35100 47354 35156 47356
rect 35180 47354 35236 47356
rect 34940 47302 34986 47354
rect 34986 47302 34996 47354
rect 35020 47302 35050 47354
rect 35050 47302 35062 47354
rect 35062 47302 35076 47354
rect 35100 47302 35114 47354
rect 35114 47302 35126 47354
rect 35126 47302 35156 47354
rect 35180 47302 35190 47354
rect 35190 47302 35236 47354
rect 34940 47300 34996 47302
rect 35020 47300 35076 47302
rect 35100 47300 35156 47302
rect 35180 47300 35236 47302
rect 34940 46266 34996 46268
rect 35020 46266 35076 46268
rect 35100 46266 35156 46268
rect 35180 46266 35236 46268
rect 34940 46214 34986 46266
rect 34986 46214 34996 46266
rect 35020 46214 35050 46266
rect 35050 46214 35062 46266
rect 35062 46214 35076 46266
rect 35100 46214 35114 46266
rect 35114 46214 35126 46266
rect 35126 46214 35156 46266
rect 35180 46214 35190 46266
rect 35190 46214 35236 46266
rect 34940 46212 34996 46214
rect 35020 46212 35076 46214
rect 35100 46212 35156 46214
rect 35180 46212 35236 46214
rect 34940 45178 34996 45180
rect 35020 45178 35076 45180
rect 35100 45178 35156 45180
rect 35180 45178 35236 45180
rect 34940 45126 34986 45178
rect 34986 45126 34996 45178
rect 35020 45126 35050 45178
rect 35050 45126 35062 45178
rect 35062 45126 35076 45178
rect 35100 45126 35114 45178
rect 35114 45126 35126 45178
rect 35126 45126 35156 45178
rect 35180 45126 35190 45178
rect 35190 45126 35236 45178
rect 34940 45124 34996 45126
rect 35020 45124 35076 45126
rect 35100 45124 35156 45126
rect 35180 45124 35236 45126
rect 34940 44090 34996 44092
rect 35020 44090 35076 44092
rect 35100 44090 35156 44092
rect 35180 44090 35236 44092
rect 34940 44038 34986 44090
rect 34986 44038 34996 44090
rect 35020 44038 35050 44090
rect 35050 44038 35062 44090
rect 35062 44038 35076 44090
rect 35100 44038 35114 44090
rect 35114 44038 35126 44090
rect 35126 44038 35156 44090
rect 35180 44038 35190 44090
rect 35190 44038 35236 44090
rect 34940 44036 34996 44038
rect 35020 44036 35076 44038
rect 35100 44036 35156 44038
rect 35180 44036 35236 44038
rect 34940 43002 34996 43004
rect 35020 43002 35076 43004
rect 35100 43002 35156 43004
rect 35180 43002 35236 43004
rect 34940 42950 34986 43002
rect 34986 42950 34996 43002
rect 35020 42950 35050 43002
rect 35050 42950 35062 43002
rect 35062 42950 35076 43002
rect 35100 42950 35114 43002
rect 35114 42950 35126 43002
rect 35126 42950 35156 43002
rect 35180 42950 35190 43002
rect 35190 42950 35236 43002
rect 34940 42948 34996 42950
rect 35020 42948 35076 42950
rect 35100 42948 35156 42950
rect 35180 42948 35236 42950
rect 34940 41914 34996 41916
rect 35020 41914 35076 41916
rect 35100 41914 35156 41916
rect 35180 41914 35236 41916
rect 34940 41862 34986 41914
rect 34986 41862 34996 41914
rect 35020 41862 35050 41914
rect 35050 41862 35062 41914
rect 35062 41862 35076 41914
rect 35100 41862 35114 41914
rect 35114 41862 35126 41914
rect 35126 41862 35156 41914
rect 35180 41862 35190 41914
rect 35190 41862 35236 41914
rect 34940 41860 34996 41862
rect 35020 41860 35076 41862
rect 35100 41860 35156 41862
rect 35180 41860 35236 41862
rect 34940 40826 34996 40828
rect 35020 40826 35076 40828
rect 35100 40826 35156 40828
rect 35180 40826 35236 40828
rect 34940 40774 34986 40826
rect 34986 40774 34996 40826
rect 35020 40774 35050 40826
rect 35050 40774 35062 40826
rect 35062 40774 35076 40826
rect 35100 40774 35114 40826
rect 35114 40774 35126 40826
rect 35126 40774 35156 40826
rect 35180 40774 35190 40826
rect 35190 40774 35236 40826
rect 34940 40772 34996 40774
rect 35020 40772 35076 40774
rect 35100 40772 35156 40774
rect 35180 40772 35236 40774
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 20902 20848 20958 20904
rect 20258 13932 20314 13968
rect 20258 13912 20260 13932
rect 20260 13912 20312 13932
rect 20312 13912 20314 13932
rect 20534 20576 20590 20632
rect 23478 27648 23534 27704
rect 22006 21392 22062 21448
rect 22006 18148 22062 18184
rect 22006 18128 22008 18148
rect 22008 18128 22060 18148
rect 22060 18128 22062 18148
rect 20442 14456 20498 14512
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19062 1944 19118 2000
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 20810 12960 20866 13016
rect 20626 10240 20682 10296
rect 19430 3984 19486 4040
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 20442 3848 20498 3904
rect 22742 20304 22798 20360
rect 22926 21800 22982 21856
rect 23386 24656 23442 24712
rect 23570 22208 23626 22264
rect 23386 21120 23442 21176
rect 22558 16108 22614 16144
rect 22558 16088 22560 16108
rect 22560 16088 22612 16108
rect 22612 16088 22614 16108
rect 22374 12688 22430 12744
rect 21914 12144 21970 12200
rect 21822 11600 21878 11656
rect 21178 8900 21234 8936
rect 21178 8880 21180 8900
rect 21180 8880 21232 8900
rect 21232 8880 21234 8900
rect 20810 3984 20866 4040
rect 22926 12044 22928 12064
rect 22928 12044 22980 12064
rect 22980 12044 22982 12064
rect 22926 12008 22982 12044
rect 23570 15000 23626 15056
rect 23294 11736 23350 11792
rect 23478 12960 23534 13016
rect 23478 12688 23534 12744
rect 22834 4664 22890 4720
rect 24030 20712 24086 20768
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 25042 23044 25098 23080
rect 25042 23024 25044 23044
rect 25044 23024 25096 23044
rect 25096 23024 25098 23044
rect 24398 21936 24454 21992
rect 24490 21836 24492 21856
rect 24492 21836 24544 21856
rect 24544 21836 24546 21856
rect 24490 21800 24546 21836
rect 24306 20984 24362 21040
rect 24674 20440 24730 20496
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 50300 56602 50356 56604
rect 50380 56602 50436 56604
rect 50460 56602 50516 56604
rect 50540 56602 50596 56604
rect 50300 56550 50346 56602
rect 50346 56550 50356 56602
rect 50380 56550 50410 56602
rect 50410 56550 50422 56602
rect 50422 56550 50436 56602
rect 50460 56550 50474 56602
rect 50474 56550 50486 56602
rect 50486 56550 50516 56602
rect 50540 56550 50550 56602
rect 50550 56550 50596 56602
rect 50300 56548 50356 56550
rect 50380 56548 50436 56550
rect 50460 56548 50516 56550
rect 50540 56548 50596 56550
rect 50300 55514 50356 55516
rect 50380 55514 50436 55516
rect 50460 55514 50516 55516
rect 50540 55514 50596 55516
rect 50300 55462 50346 55514
rect 50346 55462 50356 55514
rect 50380 55462 50410 55514
rect 50410 55462 50422 55514
rect 50422 55462 50436 55514
rect 50460 55462 50474 55514
rect 50474 55462 50486 55514
rect 50486 55462 50516 55514
rect 50540 55462 50550 55514
rect 50550 55462 50596 55514
rect 50300 55460 50356 55462
rect 50380 55460 50436 55462
rect 50460 55460 50516 55462
rect 50540 55460 50596 55462
rect 50300 54426 50356 54428
rect 50380 54426 50436 54428
rect 50460 54426 50516 54428
rect 50540 54426 50596 54428
rect 50300 54374 50346 54426
rect 50346 54374 50356 54426
rect 50380 54374 50410 54426
rect 50410 54374 50422 54426
rect 50422 54374 50436 54426
rect 50460 54374 50474 54426
rect 50474 54374 50486 54426
rect 50486 54374 50516 54426
rect 50540 54374 50550 54426
rect 50550 54374 50596 54426
rect 50300 54372 50356 54374
rect 50380 54372 50436 54374
rect 50460 54372 50516 54374
rect 50540 54372 50596 54374
rect 50300 53338 50356 53340
rect 50380 53338 50436 53340
rect 50460 53338 50516 53340
rect 50540 53338 50596 53340
rect 50300 53286 50346 53338
rect 50346 53286 50356 53338
rect 50380 53286 50410 53338
rect 50410 53286 50422 53338
rect 50422 53286 50436 53338
rect 50460 53286 50474 53338
rect 50474 53286 50486 53338
rect 50486 53286 50516 53338
rect 50540 53286 50550 53338
rect 50550 53286 50596 53338
rect 50300 53284 50356 53286
rect 50380 53284 50436 53286
rect 50460 53284 50516 53286
rect 50540 53284 50596 53286
rect 50300 52250 50356 52252
rect 50380 52250 50436 52252
rect 50460 52250 50516 52252
rect 50540 52250 50596 52252
rect 50300 52198 50346 52250
rect 50346 52198 50356 52250
rect 50380 52198 50410 52250
rect 50410 52198 50422 52250
rect 50422 52198 50436 52250
rect 50460 52198 50474 52250
rect 50474 52198 50486 52250
rect 50486 52198 50516 52250
rect 50540 52198 50550 52250
rect 50550 52198 50596 52250
rect 50300 52196 50356 52198
rect 50380 52196 50436 52198
rect 50460 52196 50516 52198
rect 50540 52196 50596 52198
rect 50300 51162 50356 51164
rect 50380 51162 50436 51164
rect 50460 51162 50516 51164
rect 50540 51162 50596 51164
rect 50300 51110 50346 51162
rect 50346 51110 50356 51162
rect 50380 51110 50410 51162
rect 50410 51110 50422 51162
rect 50422 51110 50436 51162
rect 50460 51110 50474 51162
rect 50474 51110 50486 51162
rect 50486 51110 50516 51162
rect 50540 51110 50550 51162
rect 50550 51110 50596 51162
rect 50300 51108 50356 51110
rect 50380 51108 50436 51110
rect 50460 51108 50516 51110
rect 50540 51108 50596 51110
rect 50300 50074 50356 50076
rect 50380 50074 50436 50076
rect 50460 50074 50516 50076
rect 50540 50074 50596 50076
rect 50300 50022 50346 50074
rect 50346 50022 50356 50074
rect 50380 50022 50410 50074
rect 50410 50022 50422 50074
rect 50422 50022 50436 50074
rect 50460 50022 50474 50074
rect 50474 50022 50486 50074
rect 50486 50022 50516 50074
rect 50540 50022 50550 50074
rect 50550 50022 50596 50074
rect 50300 50020 50356 50022
rect 50380 50020 50436 50022
rect 50460 50020 50516 50022
rect 50540 50020 50596 50022
rect 50300 48986 50356 48988
rect 50380 48986 50436 48988
rect 50460 48986 50516 48988
rect 50540 48986 50596 48988
rect 50300 48934 50346 48986
rect 50346 48934 50356 48986
rect 50380 48934 50410 48986
rect 50410 48934 50422 48986
rect 50422 48934 50436 48986
rect 50460 48934 50474 48986
rect 50474 48934 50486 48986
rect 50486 48934 50516 48986
rect 50540 48934 50550 48986
rect 50550 48934 50596 48986
rect 50300 48932 50356 48934
rect 50380 48932 50436 48934
rect 50460 48932 50516 48934
rect 50540 48932 50596 48934
rect 50300 47898 50356 47900
rect 50380 47898 50436 47900
rect 50460 47898 50516 47900
rect 50540 47898 50596 47900
rect 50300 47846 50346 47898
rect 50346 47846 50356 47898
rect 50380 47846 50410 47898
rect 50410 47846 50422 47898
rect 50422 47846 50436 47898
rect 50460 47846 50474 47898
rect 50474 47846 50486 47898
rect 50486 47846 50516 47898
rect 50540 47846 50550 47898
rect 50550 47846 50596 47898
rect 50300 47844 50356 47846
rect 50380 47844 50436 47846
rect 50460 47844 50516 47846
rect 50540 47844 50596 47846
rect 50300 46810 50356 46812
rect 50380 46810 50436 46812
rect 50460 46810 50516 46812
rect 50540 46810 50596 46812
rect 50300 46758 50346 46810
rect 50346 46758 50356 46810
rect 50380 46758 50410 46810
rect 50410 46758 50422 46810
rect 50422 46758 50436 46810
rect 50460 46758 50474 46810
rect 50474 46758 50486 46810
rect 50486 46758 50516 46810
rect 50540 46758 50550 46810
rect 50550 46758 50596 46810
rect 50300 46756 50356 46758
rect 50380 46756 50436 46758
rect 50460 46756 50516 46758
rect 50540 46756 50596 46758
rect 50300 45722 50356 45724
rect 50380 45722 50436 45724
rect 50460 45722 50516 45724
rect 50540 45722 50596 45724
rect 50300 45670 50346 45722
rect 50346 45670 50356 45722
rect 50380 45670 50410 45722
rect 50410 45670 50422 45722
rect 50422 45670 50436 45722
rect 50460 45670 50474 45722
rect 50474 45670 50486 45722
rect 50486 45670 50516 45722
rect 50540 45670 50550 45722
rect 50550 45670 50596 45722
rect 50300 45668 50356 45670
rect 50380 45668 50436 45670
rect 50460 45668 50516 45670
rect 50540 45668 50596 45670
rect 50300 44634 50356 44636
rect 50380 44634 50436 44636
rect 50460 44634 50516 44636
rect 50540 44634 50596 44636
rect 50300 44582 50346 44634
rect 50346 44582 50356 44634
rect 50380 44582 50410 44634
rect 50410 44582 50422 44634
rect 50422 44582 50436 44634
rect 50460 44582 50474 44634
rect 50474 44582 50486 44634
rect 50486 44582 50516 44634
rect 50540 44582 50550 44634
rect 50550 44582 50596 44634
rect 50300 44580 50356 44582
rect 50380 44580 50436 44582
rect 50460 44580 50516 44582
rect 50540 44580 50596 44582
rect 50300 43546 50356 43548
rect 50380 43546 50436 43548
rect 50460 43546 50516 43548
rect 50540 43546 50596 43548
rect 50300 43494 50346 43546
rect 50346 43494 50356 43546
rect 50380 43494 50410 43546
rect 50410 43494 50422 43546
rect 50422 43494 50436 43546
rect 50460 43494 50474 43546
rect 50474 43494 50486 43546
rect 50486 43494 50516 43546
rect 50540 43494 50550 43546
rect 50550 43494 50596 43546
rect 50300 43492 50356 43494
rect 50380 43492 50436 43494
rect 50460 43492 50516 43494
rect 50540 43492 50596 43494
rect 50300 42458 50356 42460
rect 50380 42458 50436 42460
rect 50460 42458 50516 42460
rect 50540 42458 50596 42460
rect 50300 42406 50346 42458
rect 50346 42406 50356 42458
rect 50380 42406 50410 42458
rect 50410 42406 50422 42458
rect 50422 42406 50436 42458
rect 50460 42406 50474 42458
rect 50474 42406 50486 42458
rect 50486 42406 50516 42458
rect 50540 42406 50550 42458
rect 50550 42406 50596 42458
rect 50300 42404 50356 42406
rect 50380 42404 50436 42406
rect 50460 42404 50516 42406
rect 50540 42404 50596 42406
rect 50300 41370 50356 41372
rect 50380 41370 50436 41372
rect 50460 41370 50516 41372
rect 50540 41370 50596 41372
rect 50300 41318 50346 41370
rect 50346 41318 50356 41370
rect 50380 41318 50410 41370
rect 50410 41318 50422 41370
rect 50422 41318 50436 41370
rect 50460 41318 50474 41370
rect 50474 41318 50486 41370
rect 50486 41318 50516 41370
rect 50540 41318 50550 41370
rect 50550 41318 50596 41370
rect 50300 41316 50356 41318
rect 50380 41316 50436 41318
rect 50460 41316 50516 41318
rect 50540 41316 50596 41318
rect 50300 40282 50356 40284
rect 50380 40282 50436 40284
rect 50460 40282 50516 40284
rect 50540 40282 50596 40284
rect 50300 40230 50346 40282
rect 50346 40230 50356 40282
rect 50380 40230 50410 40282
rect 50410 40230 50422 40282
rect 50422 40230 50436 40282
rect 50460 40230 50474 40282
rect 50474 40230 50486 40282
rect 50486 40230 50516 40282
rect 50540 40230 50550 40282
rect 50550 40230 50596 40282
rect 50300 40228 50356 40230
rect 50380 40228 50436 40230
rect 50460 40228 50516 40230
rect 50540 40228 50596 40230
rect 50300 39194 50356 39196
rect 50380 39194 50436 39196
rect 50460 39194 50516 39196
rect 50540 39194 50596 39196
rect 50300 39142 50346 39194
rect 50346 39142 50356 39194
rect 50380 39142 50410 39194
rect 50410 39142 50422 39194
rect 50422 39142 50436 39194
rect 50460 39142 50474 39194
rect 50474 39142 50486 39194
rect 50486 39142 50516 39194
rect 50540 39142 50550 39194
rect 50550 39142 50596 39194
rect 50300 39140 50356 39142
rect 50380 39140 50436 39142
rect 50460 39140 50516 39142
rect 50540 39140 50596 39142
rect 50300 38106 50356 38108
rect 50380 38106 50436 38108
rect 50460 38106 50516 38108
rect 50540 38106 50596 38108
rect 50300 38054 50346 38106
rect 50346 38054 50356 38106
rect 50380 38054 50410 38106
rect 50410 38054 50422 38106
rect 50422 38054 50436 38106
rect 50460 38054 50474 38106
rect 50474 38054 50486 38106
rect 50486 38054 50516 38106
rect 50540 38054 50550 38106
rect 50550 38054 50596 38106
rect 50300 38052 50356 38054
rect 50380 38052 50436 38054
rect 50460 38052 50516 38054
rect 50540 38052 50596 38054
rect 50300 37018 50356 37020
rect 50380 37018 50436 37020
rect 50460 37018 50516 37020
rect 50540 37018 50596 37020
rect 50300 36966 50346 37018
rect 50346 36966 50356 37018
rect 50380 36966 50410 37018
rect 50410 36966 50422 37018
rect 50422 36966 50436 37018
rect 50460 36966 50474 37018
rect 50474 36966 50486 37018
rect 50486 36966 50516 37018
rect 50540 36966 50550 37018
rect 50550 36966 50596 37018
rect 50300 36964 50356 36966
rect 50380 36964 50436 36966
rect 50460 36964 50516 36966
rect 50540 36964 50596 36966
rect 50300 35930 50356 35932
rect 50380 35930 50436 35932
rect 50460 35930 50516 35932
rect 50540 35930 50596 35932
rect 50300 35878 50346 35930
rect 50346 35878 50356 35930
rect 50380 35878 50410 35930
rect 50410 35878 50422 35930
rect 50422 35878 50436 35930
rect 50460 35878 50474 35930
rect 50474 35878 50486 35930
rect 50486 35878 50516 35930
rect 50540 35878 50550 35930
rect 50550 35878 50596 35930
rect 50300 35876 50356 35878
rect 50380 35876 50436 35878
rect 50460 35876 50516 35878
rect 50540 35876 50596 35878
rect 50300 34842 50356 34844
rect 50380 34842 50436 34844
rect 50460 34842 50516 34844
rect 50540 34842 50596 34844
rect 50300 34790 50346 34842
rect 50346 34790 50356 34842
rect 50380 34790 50410 34842
rect 50410 34790 50422 34842
rect 50422 34790 50436 34842
rect 50460 34790 50474 34842
rect 50474 34790 50486 34842
rect 50486 34790 50516 34842
rect 50540 34790 50550 34842
rect 50550 34790 50596 34842
rect 50300 34788 50356 34790
rect 50380 34788 50436 34790
rect 50460 34788 50516 34790
rect 50540 34788 50596 34790
rect 50300 33754 50356 33756
rect 50380 33754 50436 33756
rect 50460 33754 50516 33756
rect 50540 33754 50596 33756
rect 50300 33702 50346 33754
rect 50346 33702 50356 33754
rect 50380 33702 50410 33754
rect 50410 33702 50422 33754
rect 50422 33702 50436 33754
rect 50460 33702 50474 33754
rect 50474 33702 50486 33754
rect 50486 33702 50516 33754
rect 50540 33702 50550 33754
rect 50550 33702 50596 33754
rect 50300 33700 50356 33702
rect 50380 33700 50436 33702
rect 50460 33700 50516 33702
rect 50540 33700 50596 33702
rect 50300 32666 50356 32668
rect 50380 32666 50436 32668
rect 50460 32666 50516 32668
rect 50540 32666 50596 32668
rect 50300 32614 50346 32666
rect 50346 32614 50356 32666
rect 50380 32614 50410 32666
rect 50410 32614 50422 32666
rect 50422 32614 50436 32666
rect 50460 32614 50474 32666
rect 50474 32614 50486 32666
rect 50486 32614 50516 32666
rect 50540 32614 50550 32666
rect 50550 32614 50596 32666
rect 50300 32612 50356 32614
rect 50380 32612 50436 32614
rect 50460 32612 50516 32614
rect 50540 32612 50596 32614
rect 25778 22752 25834 22808
rect 27618 23060 27620 23080
rect 27620 23060 27672 23080
rect 27672 23060 27674 23080
rect 25318 20440 25374 20496
rect 24490 19488 24546 19544
rect 25042 16532 25044 16552
rect 25044 16532 25096 16552
rect 25096 16532 25098 16552
rect 25042 16496 25098 16532
rect 24398 15000 24454 15056
rect 24214 14900 24216 14920
rect 24216 14900 24268 14920
rect 24268 14900 24270 14920
rect 24214 14864 24270 14900
rect 23754 13268 23756 13288
rect 23756 13268 23808 13288
rect 23808 13268 23810 13288
rect 23754 13232 23810 13268
rect 24122 11600 24178 11656
rect 24674 15272 24730 15328
rect 24766 13232 24822 13288
rect 24674 12824 24730 12880
rect 24766 11872 24822 11928
rect 23754 3032 23810 3088
rect 25134 14320 25190 14376
rect 25134 12008 25190 12064
rect 25134 11772 25136 11792
rect 25136 11772 25188 11792
rect 25188 11772 25190 11792
rect 25134 11736 25190 11772
rect 25410 12980 25466 13016
rect 25410 12960 25412 12980
rect 25412 12960 25464 12980
rect 25464 12960 25466 12980
rect 25318 12416 25374 12472
rect 25410 12316 25412 12336
rect 25412 12316 25464 12336
rect 25464 12316 25466 12336
rect 25410 12280 25466 12316
rect 25870 16088 25926 16144
rect 25962 15952 26018 16008
rect 26238 14864 26294 14920
rect 27158 16360 27214 16416
rect 27618 23024 27674 23060
rect 27342 21120 27398 21176
rect 27894 21564 27896 21584
rect 27896 21564 27948 21584
rect 27948 21564 27950 21584
rect 27894 21528 27950 21564
rect 28906 22772 28962 22808
rect 28906 22752 28908 22772
rect 28908 22752 28960 22772
rect 28960 22752 28962 22772
rect 28998 21548 29054 21584
rect 28998 21528 29000 21548
rect 29000 21528 29052 21548
rect 29052 21528 29054 21548
rect 27250 16088 27306 16144
rect 29090 20576 29146 20632
rect 26146 12980 26202 13016
rect 26146 12960 26148 12980
rect 26148 12960 26200 12980
rect 26200 12960 26202 12980
rect 26330 12824 26386 12880
rect 26238 12008 26294 12064
rect 26238 11756 26294 11792
rect 26238 11736 26240 11756
rect 26240 11736 26292 11756
rect 26292 11736 26294 11756
rect 26146 9424 26202 9480
rect 24490 3712 24546 3768
rect 23846 2760 23902 2816
rect 26606 12688 26662 12744
rect 27066 13232 27122 13288
rect 28814 19624 28870 19680
rect 29550 22616 29606 22672
rect 30286 21548 30342 21584
rect 30286 21528 30288 21548
rect 30288 21528 30340 21548
rect 30340 21528 30342 21548
rect 29458 16360 29514 16416
rect 30010 16496 30066 16552
rect 28630 15020 28686 15056
rect 28630 15000 28632 15020
rect 28632 15000 28684 15020
rect 28684 15000 28686 15020
rect 27434 10124 27490 10160
rect 27434 10104 27436 10124
rect 27436 10104 27488 10124
rect 27488 10104 27490 10124
rect 26698 4528 26754 4584
rect 26146 3576 26202 3632
rect 25594 2352 25650 2408
rect 28078 11500 28080 11520
rect 28080 11500 28132 11520
rect 28132 11500 28134 11520
rect 28078 11464 28134 11500
rect 28078 10412 28080 10432
rect 28080 10412 28132 10432
rect 28132 10412 28134 10432
rect 28078 10376 28134 10412
rect 29090 15272 29146 15328
rect 29274 14184 29330 14240
rect 28722 13524 28778 13560
rect 28722 13504 28724 13524
rect 28724 13504 28776 13524
rect 28776 13504 28778 13524
rect 29090 12416 29146 12472
rect 28722 10920 28778 10976
rect 28814 9968 28870 10024
rect 27802 4564 27804 4584
rect 27804 4564 27856 4584
rect 27856 4564 27858 4584
rect 27802 4528 27858 4564
rect 29826 12008 29882 12064
rect 29826 11328 29882 11384
rect 29734 11056 29790 11112
rect 30286 11328 30342 11384
rect 30930 20576 30986 20632
rect 31666 20440 31722 20496
rect 30654 14864 30710 14920
rect 31022 15020 31078 15056
rect 31022 15000 31024 15020
rect 31024 15000 31076 15020
rect 31076 15000 31078 15020
rect 31114 12008 31170 12064
rect 30838 10532 30894 10568
rect 30838 10512 30840 10532
rect 30840 10512 30892 10532
rect 30892 10512 30894 10532
rect 31390 13404 31392 13424
rect 31392 13404 31444 13424
rect 31444 13404 31446 13424
rect 31390 13368 31446 13404
rect 31298 12588 31300 12608
rect 31300 12588 31352 12608
rect 31352 12588 31354 12608
rect 31298 12552 31354 12588
rect 31206 10104 31262 10160
rect 32770 20848 32826 20904
rect 32310 20576 32366 20632
rect 31666 15952 31722 16008
rect 32402 12164 32458 12200
rect 32402 12144 32404 12164
rect 32404 12144 32456 12164
rect 32456 12144 32458 12164
rect 32310 10376 32366 10432
rect 31482 9424 31538 9480
rect 33506 22636 33562 22672
rect 33506 22616 33508 22636
rect 33508 22616 33560 22636
rect 33560 22616 33562 22636
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 32678 14884 32734 14920
rect 32678 14864 32680 14884
rect 32680 14864 32732 14884
rect 32732 14864 32734 14884
rect 32862 14320 32918 14376
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34886 19660 34888 19680
rect 34888 19660 34940 19680
rect 34940 19660 34942 19680
rect 34886 19624 34942 19660
rect 32310 9696 32366 9752
rect 32862 11328 32918 11384
rect 32862 11228 32864 11248
rect 32864 11228 32916 11248
rect 32916 11228 32918 11248
rect 32862 11192 32918 11228
rect 33322 10124 33378 10160
rect 33322 10104 33324 10124
rect 33324 10104 33376 10124
rect 33376 10104 33378 10124
rect 33322 9560 33378 9616
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 35714 21392 35770 21448
rect 36358 20576 36414 20632
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 35622 16088 35678 16144
rect 36082 16360 36138 16416
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34610 14320 34666 14376
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 35530 14048 35586 14104
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34978 11192 35034 11248
rect 35622 11892 35678 11928
rect 35622 11872 35624 11892
rect 35624 11872 35676 11892
rect 35676 11872 35678 11892
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 37370 19488 37426 19544
rect 37094 14184 37150 14240
rect 36082 10920 36138 10976
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 36542 8492 36598 8528
rect 36542 8472 36544 8492
rect 36544 8472 36596 8492
rect 36596 8472 36598 8492
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 38382 20440 38438 20496
rect 37002 11192 37058 11248
rect 38382 9560 38438 9616
rect 38014 8492 38070 8528
rect 38014 8472 38016 8492
rect 38016 8472 38068 8492
rect 38068 8472 38070 8492
rect 50300 31578 50356 31580
rect 50380 31578 50436 31580
rect 50460 31578 50516 31580
rect 50540 31578 50596 31580
rect 50300 31526 50346 31578
rect 50346 31526 50356 31578
rect 50380 31526 50410 31578
rect 50410 31526 50422 31578
rect 50422 31526 50436 31578
rect 50460 31526 50474 31578
rect 50474 31526 50486 31578
rect 50486 31526 50516 31578
rect 50540 31526 50550 31578
rect 50550 31526 50596 31578
rect 50300 31524 50356 31526
rect 50380 31524 50436 31526
rect 50460 31524 50516 31526
rect 50540 31524 50596 31526
rect 50300 30490 50356 30492
rect 50380 30490 50436 30492
rect 50460 30490 50516 30492
rect 50540 30490 50596 30492
rect 50300 30438 50346 30490
rect 50346 30438 50356 30490
rect 50380 30438 50410 30490
rect 50410 30438 50422 30490
rect 50422 30438 50436 30490
rect 50460 30438 50474 30490
rect 50474 30438 50486 30490
rect 50486 30438 50516 30490
rect 50540 30438 50550 30490
rect 50550 30438 50596 30490
rect 50300 30436 50356 30438
rect 50380 30436 50436 30438
rect 50460 30436 50516 30438
rect 50540 30436 50596 30438
rect 50300 29402 50356 29404
rect 50380 29402 50436 29404
rect 50460 29402 50516 29404
rect 50540 29402 50596 29404
rect 50300 29350 50346 29402
rect 50346 29350 50356 29402
rect 50380 29350 50410 29402
rect 50410 29350 50422 29402
rect 50422 29350 50436 29402
rect 50460 29350 50474 29402
rect 50474 29350 50486 29402
rect 50486 29350 50516 29402
rect 50540 29350 50550 29402
rect 50550 29350 50596 29402
rect 50300 29348 50356 29350
rect 50380 29348 50436 29350
rect 50460 29348 50516 29350
rect 50540 29348 50596 29350
rect 50300 28314 50356 28316
rect 50380 28314 50436 28316
rect 50460 28314 50516 28316
rect 50540 28314 50596 28316
rect 50300 28262 50346 28314
rect 50346 28262 50356 28314
rect 50380 28262 50410 28314
rect 50410 28262 50422 28314
rect 50422 28262 50436 28314
rect 50460 28262 50474 28314
rect 50474 28262 50486 28314
rect 50486 28262 50516 28314
rect 50540 28262 50550 28314
rect 50550 28262 50596 28314
rect 50300 28260 50356 28262
rect 50380 28260 50436 28262
rect 50460 28260 50516 28262
rect 50540 28260 50596 28262
rect 50300 27226 50356 27228
rect 50380 27226 50436 27228
rect 50460 27226 50516 27228
rect 50540 27226 50596 27228
rect 50300 27174 50346 27226
rect 50346 27174 50356 27226
rect 50380 27174 50410 27226
rect 50410 27174 50422 27226
rect 50422 27174 50436 27226
rect 50460 27174 50474 27226
rect 50474 27174 50486 27226
rect 50486 27174 50516 27226
rect 50540 27174 50550 27226
rect 50550 27174 50596 27226
rect 50300 27172 50356 27174
rect 50380 27172 50436 27174
rect 50460 27172 50516 27174
rect 50540 27172 50596 27174
rect 50300 26138 50356 26140
rect 50380 26138 50436 26140
rect 50460 26138 50516 26140
rect 50540 26138 50596 26140
rect 50300 26086 50346 26138
rect 50346 26086 50356 26138
rect 50380 26086 50410 26138
rect 50410 26086 50422 26138
rect 50422 26086 50436 26138
rect 50460 26086 50474 26138
rect 50474 26086 50486 26138
rect 50486 26086 50516 26138
rect 50540 26086 50550 26138
rect 50550 26086 50596 26138
rect 50300 26084 50356 26086
rect 50380 26084 50436 26086
rect 50460 26084 50516 26086
rect 50540 26084 50596 26086
rect 50300 25050 50356 25052
rect 50380 25050 50436 25052
rect 50460 25050 50516 25052
rect 50540 25050 50596 25052
rect 50300 24998 50346 25050
rect 50346 24998 50356 25050
rect 50380 24998 50410 25050
rect 50410 24998 50422 25050
rect 50422 24998 50436 25050
rect 50460 24998 50474 25050
rect 50474 24998 50486 25050
rect 50486 24998 50516 25050
rect 50540 24998 50550 25050
rect 50550 24998 50596 25050
rect 50300 24996 50356 24998
rect 50380 24996 50436 24998
rect 50460 24996 50516 24998
rect 50540 24996 50596 24998
rect 65660 57146 65716 57148
rect 65740 57146 65796 57148
rect 65820 57146 65876 57148
rect 65900 57146 65956 57148
rect 65660 57094 65706 57146
rect 65706 57094 65716 57146
rect 65740 57094 65770 57146
rect 65770 57094 65782 57146
rect 65782 57094 65796 57146
rect 65820 57094 65834 57146
rect 65834 57094 65846 57146
rect 65846 57094 65876 57146
rect 65900 57094 65910 57146
rect 65910 57094 65956 57146
rect 65660 57092 65716 57094
rect 65740 57092 65796 57094
rect 65820 57092 65876 57094
rect 65900 57092 65956 57094
rect 67638 56108 67640 56128
rect 67640 56108 67692 56128
rect 67692 56108 67694 56128
rect 67638 56072 67694 56108
rect 65660 56058 65716 56060
rect 65740 56058 65796 56060
rect 65820 56058 65876 56060
rect 65900 56058 65956 56060
rect 65660 56006 65706 56058
rect 65706 56006 65716 56058
rect 65740 56006 65770 56058
rect 65770 56006 65782 56058
rect 65782 56006 65796 56058
rect 65820 56006 65834 56058
rect 65834 56006 65846 56058
rect 65846 56006 65876 56058
rect 65900 56006 65910 56058
rect 65910 56006 65956 56058
rect 65660 56004 65716 56006
rect 65740 56004 65796 56006
rect 65820 56004 65876 56006
rect 65900 56004 65956 56006
rect 65660 54970 65716 54972
rect 65740 54970 65796 54972
rect 65820 54970 65876 54972
rect 65900 54970 65956 54972
rect 65660 54918 65706 54970
rect 65706 54918 65716 54970
rect 65740 54918 65770 54970
rect 65770 54918 65782 54970
rect 65782 54918 65796 54970
rect 65820 54918 65834 54970
rect 65834 54918 65846 54970
rect 65846 54918 65876 54970
rect 65900 54918 65910 54970
rect 65910 54918 65956 54970
rect 65660 54916 65716 54918
rect 65740 54916 65796 54918
rect 65820 54916 65876 54918
rect 65900 54916 65956 54918
rect 68098 54612 68100 54632
rect 68100 54612 68152 54632
rect 68152 54612 68154 54632
rect 68098 54576 68154 54612
rect 65660 53882 65716 53884
rect 65740 53882 65796 53884
rect 65820 53882 65876 53884
rect 65900 53882 65956 53884
rect 65660 53830 65706 53882
rect 65706 53830 65716 53882
rect 65740 53830 65770 53882
rect 65770 53830 65782 53882
rect 65782 53830 65796 53882
rect 65820 53830 65834 53882
rect 65834 53830 65846 53882
rect 65846 53830 65876 53882
rect 65900 53830 65910 53882
rect 65910 53830 65956 53882
rect 65660 53828 65716 53830
rect 65740 53828 65796 53830
rect 65820 53828 65876 53830
rect 65900 53828 65956 53830
rect 68098 53080 68154 53136
rect 65660 52794 65716 52796
rect 65740 52794 65796 52796
rect 65820 52794 65876 52796
rect 65900 52794 65956 52796
rect 65660 52742 65706 52794
rect 65706 52742 65716 52794
rect 65740 52742 65770 52794
rect 65770 52742 65782 52794
rect 65782 52742 65796 52794
rect 65820 52742 65834 52794
rect 65834 52742 65846 52794
rect 65846 52742 65876 52794
rect 65900 52742 65910 52794
rect 65910 52742 65956 52794
rect 65660 52740 65716 52742
rect 65740 52740 65796 52742
rect 65820 52740 65876 52742
rect 65900 52740 65956 52742
rect 65660 51706 65716 51708
rect 65740 51706 65796 51708
rect 65820 51706 65876 51708
rect 65900 51706 65956 51708
rect 65660 51654 65706 51706
rect 65706 51654 65716 51706
rect 65740 51654 65770 51706
rect 65770 51654 65782 51706
rect 65782 51654 65796 51706
rect 65820 51654 65834 51706
rect 65834 51654 65846 51706
rect 65846 51654 65876 51706
rect 65900 51654 65910 51706
rect 65910 51654 65956 51706
rect 65660 51652 65716 51654
rect 65740 51652 65796 51654
rect 65820 51652 65876 51654
rect 65900 51652 65956 51654
rect 67638 51584 67694 51640
rect 65660 50618 65716 50620
rect 65740 50618 65796 50620
rect 65820 50618 65876 50620
rect 65900 50618 65956 50620
rect 65660 50566 65706 50618
rect 65706 50566 65716 50618
rect 65740 50566 65770 50618
rect 65770 50566 65782 50618
rect 65782 50566 65796 50618
rect 65820 50566 65834 50618
rect 65834 50566 65846 50618
rect 65846 50566 65876 50618
rect 65900 50566 65910 50618
rect 65910 50566 65956 50618
rect 65660 50564 65716 50566
rect 65740 50564 65796 50566
rect 65820 50564 65876 50566
rect 65900 50564 65956 50566
rect 68098 50088 68154 50144
rect 65660 49530 65716 49532
rect 65740 49530 65796 49532
rect 65820 49530 65876 49532
rect 65900 49530 65956 49532
rect 65660 49478 65706 49530
rect 65706 49478 65716 49530
rect 65740 49478 65770 49530
rect 65770 49478 65782 49530
rect 65782 49478 65796 49530
rect 65820 49478 65834 49530
rect 65834 49478 65846 49530
rect 65846 49478 65876 49530
rect 65900 49478 65910 49530
rect 65910 49478 65956 49530
rect 65660 49476 65716 49478
rect 65740 49476 65796 49478
rect 65820 49476 65876 49478
rect 65900 49476 65956 49478
rect 67638 48612 67694 48648
rect 67638 48592 67640 48612
rect 67640 48592 67692 48612
rect 67692 48592 67694 48612
rect 65660 48442 65716 48444
rect 65740 48442 65796 48444
rect 65820 48442 65876 48444
rect 65900 48442 65956 48444
rect 65660 48390 65706 48442
rect 65706 48390 65716 48442
rect 65740 48390 65770 48442
rect 65770 48390 65782 48442
rect 65782 48390 65796 48442
rect 65820 48390 65834 48442
rect 65834 48390 65846 48442
rect 65846 48390 65876 48442
rect 65900 48390 65910 48442
rect 65910 48390 65956 48442
rect 65660 48388 65716 48390
rect 65740 48388 65796 48390
rect 65820 48388 65876 48390
rect 65900 48388 65956 48390
rect 65660 47354 65716 47356
rect 65740 47354 65796 47356
rect 65820 47354 65876 47356
rect 65900 47354 65956 47356
rect 65660 47302 65706 47354
rect 65706 47302 65716 47354
rect 65740 47302 65770 47354
rect 65770 47302 65782 47354
rect 65782 47302 65796 47354
rect 65820 47302 65834 47354
rect 65834 47302 65846 47354
rect 65846 47302 65876 47354
rect 65900 47302 65910 47354
rect 65910 47302 65956 47354
rect 65660 47300 65716 47302
rect 65740 47300 65796 47302
rect 65820 47300 65876 47302
rect 65900 47300 65956 47302
rect 67638 47096 67694 47152
rect 65660 46266 65716 46268
rect 65740 46266 65796 46268
rect 65820 46266 65876 46268
rect 65900 46266 65956 46268
rect 65660 46214 65706 46266
rect 65706 46214 65716 46266
rect 65740 46214 65770 46266
rect 65770 46214 65782 46266
rect 65782 46214 65796 46266
rect 65820 46214 65834 46266
rect 65834 46214 65846 46266
rect 65846 46214 65876 46266
rect 65900 46214 65910 46266
rect 65910 46214 65956 46266
rect 65660 46212 65716 46214
rect 65740 46212 65796 46214
rect 65820 46212 65876 46214
rect 65900 46212 65956 46214
rect 68098 45600 68154 45656
rect 65660 45178 65716 45180
rect 65740 45178 65796 45180
rect 65820 45178 65876 45180
rect 65900 45178 65956 45180
rect 65660 45126 65706 45178
rect 65706 45126 65716 45178
rect 65740 45126 65770 45178
rect 65770 45126 65782 45178
rect 65782 45126 65796 45178
rect 65820 45126 65834 45178
rect 65834 45126 65846 45178
rect 65846 45126 65876 45178
rect 65900 45126 65910 45178
rect 65910 45126 65956 45178
rect 65660 45124 65716 45126
rect 65740 45124 65796 45126
rect 65820 45124 65876 45126
rect 65900 45124 65956 45126
rect 67546 44140 67548 44160
rect 67548 44140 67600 44160
rect 67600 44140 67602 44160
rect 67546 44104 67602 44140
rect 65660 44090 65716 44092
rect 65740 44090 65796 44092
rect 65820 44090 65876 44092
rect 65900 44090 65956 44092
rect 65660 44038 65706 44090
rect 65706 44038 65716 44090
rect 65740 44038 65770 44090
rect 65770 44038 65782 44090
rect 65782 44038 65796 44090
rect 65820 44038 65834 44090
rect 65834 44038 65846 44090
rect 65846 44038 65876 44090
rect 65900 44038 65910 44090
rect 65910 44038 65956 44090
rect 65660 44036 65716 44038
rect 65740 44036 65796 44038
rect 65820 44036 65876 44038
rect 65900 44036 65956 44038
rect 65660 43002 65716 43004
rect 65740 43002 65796 43004
rect 65820 43002 65876 43004
rect 65900 43002 65956 43004
rect 65660 42950 65706 43002
rect 65706 42950 65716 43002
rect 65740 42950 65770 43002
rect 65770 42950 65782 43002
rect 65782 42950 65796 43002
rect 65820 42950 65834 43002
rect 65834 42950 65846 43002
rect 65846 42950 65876 43002
rect 65900 42950 65910 43002
rect 65910 42950 65956 43002
rect 65660 42948 65716 42950
rect 65740 42948 65796 42950
rect 65820 42948 65876 42950
rect 65900 42948 65956 42950
rect 68098 42644 68100 42664
rect 68100 42644 68152 42664
rect 68152 42644 68154 42664
rect 68098 42608 68154 42644
rect 65660 41914 65716 41916
rect 65740 41914 65796 41916
rect 65820 41914 65876 41916
rect 65900 41914 65956 41916
rect 65660 41862 65706 41914
rect 65706 41862 65716 41914
rect 65740 41862 65770 41914
rect 65770 41862 65782 41914
rect 65782 41862 65796 41914
rect 65820 41862 65834 41914
rect 65834 41862 65846 41914
rect 65846 41862 65876 41914
rect 65900 41862 65910 41914
rect 65910 41862 65956 41914
rect 65660 41860 65716 41862
rect 65740 41860 65796 41862
rect 65820 41860 65876 41862
rect 65900 41860 65956 41862
rect 68098 41112 68154 41168
rect 65660 40826 65716 40828
rect 65740 40826 65796 40828
rect 65820 40826 65876 40828
rect 65900 40826 65956 40828
rect 65660 40774 65706 40826
rect 65706 40774 65716 40826
rect 65740 40774 65770 40826
rect 65770 40774 65782 40826
rect 65782 40774 65796 40826
rect 65820 40774 65834 40826
rect 65834 40774 65846 40826
rect 65846 40774 65876 40826
rect 65900 40774 65910 40826
rect 65910 40774 65956 40826
rect 65660 40772 65716 40774
rect 65740 40772 65796 40774
rect 65820 40772 65876 40774
rect 65900 40772 65956 40774
rect 65660 39738 65716 39740
rect 65740 39738 65796 39740
rect 65820 39738 65876 39740
rect 65900 39738 65956 39740
rect 65660 39686 65706 39738
rect 65706 39686 65716 39738
rect 65740 39686 65770 39738
rect 65770 39686 65782 39738
rect 65782 39686 65796 39738
rect 65820 39686 65834 39738
rect 65834 39686 65846 39738
rect 65846 39686 65876 39738
rect 65900 39686 65910 39738
rect 65910 39686 65956 39738
rect 65660 39684 65716 39686
rect 65740 39684 65796 39686
rect 65820 39684 65876 39686
rect 65900 39684 65956 39686
rect 67638 39616 67694 39672
rect 65660 38650 65716 38652
rect 65740 38650 65796 38652
rect 65820 38650 65876 38652
rect 65900 38650 65956 38652
rect 65660 38598 65706 38650
rect 65706 38598 65716 38650
rect 65740 38598 65770 38650
rect 65770 38598 65782 38650
rect 65782 38598 65796 38650
rect 65820 38598 65834 38650
rect 65834 38598 65846 38650
rect 65846 38598 65876 38650
rect 65900 38598 65910 38650
rect 65910 38598 65956 38650
rect 65660 38596 65716 38598
rect 65740 38596 65796 38598
rect 65820 38596 65876 38598
rect 65900 38596 65956 38598
rect 68098 38120 68154 38176
rect 65660 37562 65716 37564
rect 65740 37562 65796 37564
rect 65820 37562 65876 37564
rect 65900 37562 65956 37564
rect 65660 37510 65706 37562
rect 65706 37510 65716 37562
rect 65740 37510 65770 37562
rect 65770 37510 65782 37562
rect 65782 37510 65796 37562
rect 65820 37510 65834 37562
rect 65834 37510 65846 37562
rect 65846 37510 65876 37562
rect 65900 37510 65910 37562
rect 65910 37510 65956 37562
rect 65660 37508 65716 37510
rect 65740 37508 65796 37510
rect 65820 37508 65876 37510
rect 65900 37508 65956 37510
rect 67638 36644 67694 36680
rect 67638 36624 67640 36644
rect 67640 36624 67692 36644
rect 67692 36624 67694 36644
rect 65660 36474 65716 36476
rect 65740 36474 65796 36476
rect 65820 36474 65876 36476
rect 65900 36474 65956 36476
rect 65660 36422 65706 36474
rect 65706 36422 65716 36474
rect 65740 36422 65770 36474
rect 65770 36422 65782 36474
rect 65782 36422 65796 36474
rect 65820 36422 65834 36474
rect 65834 36422 65846 36474
rect 65846 36422 65876 36474
rect 65900 36422 65910 36474
rect 65910 36422 65956 36474
rect 65660 36420 65716 36422
rect 65740 36420 65796 36422
rect 65820 36420 65876 36422
rect 65900 36420 65956 36422
rect 65660 35386 65716 35388
rect 65740 35386 65796 35388
rect 65820 35386 65876 35388
rect 65900 35386 65956 35388
rect 65660 35334 65706 35386
rect 65706 35334 65716 35386
rect 65740 35334 65770 35386
rect 65770 35334 65782 35386
rect 65782 35334 65796 35386
rect 65820 35334 65834 35386
rect 65834 35334 65846 35386
rect 65846 35334 65876 35386
rect 65900 35334 65910 35386
rect 65910 35334 65956 35386
rect 65660 35332 65716 35334
rect 65740 35332 65796 35334
rect 65820 35332 65876 35334
rect 65900 35332 65956 35334
rect 67638 35128 67694 35184
rect 65660 34298 65716 34300
rect 65740 34298 65796 34300
rect 65820 34298 65876 34300
rect 65900 34298 65956 34300
rect 65660 34246 65706 34298
rect 65706 34246 65716 34298
rect 65740 34246 65770 34298
rect 65770 34246 65782 34298
rect 65782 34246 65796 34298
rect 65820 34246 65834 34298
rect 65834 34246 65846 34298
rect 65846 34246 65876 34298
rect 65900 34246 65910 34298
rect 65910 34246 65956 34298
rect 65660 34244 65716 34246
rect 65740 34244 65796 34246
rect 65820 34244 65876 34246
rect 65900 34244 65956 34246
rect 68098 33632 68154 33688
rect 65660 33210 65716 33212
rect 65740 33210 65796 33212
rect 65820 33210 65876 33212
rect 65900 33210 65956 33212
rect 65660 33158 65706 33210
rect 65706 33158 65716 33210
rect 65740 33158 65770 33210
rect 65770 33158 65782 33210
rect 65782 33158 65796 33210
rect 65820 33158 65834 33210
rect 65834 33158 65846 33210
rect 65846 33158 65876 33210
rect 65900 33158 65910 33210
rect 65910 33158 65956 33210
rect 65660 33156 65716 33158
rect 65740 33156 65796 33158
rect 65820 33156 65876 33158
rect 65900 33156 65956 33158
rect 67638 32172 67640 32192
rect 67640 32172 67692 32192
rect 67692 32172 67694 32192
rect 67638 32136 67694 32172
rect 65660 32122 65716 32124
rect 65740 32122 65796 32124
rect 65820 32122 65876 32124
rect 65900 32122 65956 32124
rect 65660 32070 65706 32122
rect 65706 32070 65716 32122
rect 65740 32070 65770 32122
rect 65770 32070 65782 32122
rect 65782 32070 65796 32122
rect 65820 32070 65834 32122
rect 65834 32070 65846 32122
rect 65846 32070 65876 32122
rect 65900 32070 65910 32122
rect 65910 32070 65956 32122
rect 65660 32068 65716 32070
rect 65740 32068 65796 32070
rect 65820 32068 65876 32070
rect 65900 32068 65956 32070
rect 65660 31034 65716 31036
rect 65740 31034 65796 31036
rect 65820 31034 65876 31036
rect 65900 31034 65956 31036
rect 65660 30982 65706 31034
rect 65706 30982 65716 31034
rect 65740 30982 65770 31034
rect 65770 30982 65782 31034
rect 65782 30982 65796 31034
rect 65820 30982 65834 31034
rect 65834 30982 65846 31034
rect 65846 30982 65876 31034
rect 65900 30982 65910 31034
rect 65910 30982 65956 31034
rect 65660 30980 65716 30982
rect 65740 30980 65796 30982
rect 65820 30980 65876 30982
rect 65900 30980 65956 30982
rect 68098 30676 68100 30696
rect 68100 30676 68152 30696
rect 68152 30676 68154 30696
rect 68098 30640 68154 30676
rect 65660 29946 65716 29948
rect 65740 29946 65796 29948
rect 65820 29946 65876 29948
rect 65900 29946 65956 29948
rect 65660 29894 65706 29946
rect 65706 29894 65716 29946
rect 65740 29894 65770 29946
rect 65770 29894 65782 29946
rect 65782 29894 65796 29946
rect 65820 29894 65834 29946
rect 65834 29894 65846 29946
rect 65846 29894 65876 29946
rect 65900 29894 65910 29946
rect 65910 29894 65956 29946
rect 65660 29892 65716 29894
rect 65740 29892 65796 29894
rect 65820 29892 65876 29894
rect 65900 29892 65956 29894
rect 68098 29144 68154 29200
rect 65660 28858 65716 28860
rect 65740 28858 65796 28860
rect 65820 28858 65876 28860
rect 65900 28858 65956 28860
rect 65660 28806 65706 28858
rect 65706 28806 65716 28858
rect 65740 28806 65770 28858
rect 65770 28806 65782 28858
rect 65782 28806 65796 28858
rect 65820 28806 65834 28858
rect 65834 28806 65846 28858
rect 65846 28806 65876 28858
rect 65900 28806 65910 28858
rect 65910 28806 65956 28858
rect 65660 28804 65716 28806
rect 65740 28804 65796 28806
rect 65820 28804 65876 28806
rect 65900 28804 65956 28806
rect 65660 27770 65716 27772
rect 65740 27770 65796 27772
rect 65820 27770 65876 27772
rect 65900 27770 65956 27772
rect 65660 27718 65706 27770
rect 65706 27718 65716 27770
rect 65740 27718 65770 27770
rect 65770 27718 65782 27770
rect 65782 27718 65796 27770
rect 65820 27718 65834 27770
rect 65834 27718 65846 27770
rect 65846 27718 65876 27770
rect 65900 27718 65910 27770
rect 65910 27718 65956 27770
rect 65660 27716 65716 27718
rect 65740 27716 65796 27718
rect 65820 27716 65876 27718
rect 65900 27716 65956 27718
rect 67638 27648 67694 27704
rect 65660 26682 65716 26684
rect 65740 26682 65796 26684
rect 65820 26682 65876 26684
rect 65900 26682 65956 26684
rect 65660 26630 65706 26682
rect 65706 26630 65716 26682
rect 65740 26630 65770 26682
rect 65770 26630 65782 26682
rect 65782 26630 65796 26682
rect 65820 26630 65834 26682
rect 65834 26630 65846 26682
rect 65846 26630 65876 26682
rect 65900 26630 65910 26682
rect 65910 26630 65956 26682
rect 65660 26628 65716 26630
rect 65740 26628 65796 26630
rect 65820 26628 65876 26630
rect 65900 26628 65956 26630
rect 68098 26152 68154 26208
rect 65660 25594 65716 25596
rect 65740 25594 65796 25596
rect 65820 25594 65876 25596
rect 65900 25594 65956 25596
rect 65660 25542 65706 25594
rect 65706 25542 65716 25594
rect 65740 25542 65770 25594
rect 65770 25542 65782 25594
rect 65782 25542 65796 25594
rect 65820 25542 65834 25594
rect 65834 25542 65846 25594
rect 65846 25542 65876 25594
rect 65900 25542 65910 25594
rect 65910 25542 65956 25594
rect 65660 25540 65716 25542
rect 65740 25540 65796 25542
rect 65820 25540 65876 25542
rect 65900 25540 65956 25542
rect 67638 24676 67694 24712
rect 67638 24656 67640 24676
rect 67640 24656 67692 24676
rect 67692 24656 67694 24676
rect 65660 24506 65716 24508
rect 65740 24506 65796 24508
rect 65820 24506 65876 24508
rect 65900 24506 65956 24508
rect 65660 24454 65706 24506
rect 65706 24454 65716 24506
rect 65740 24454 65770 24506
rect 65770 24454 65782 24506
rect 65782 24454 65796 24506
rect 65820 24454 65834 24506
rect 65834 24454 65846 24506
rect 65846 24454 65876 24506
rect 65900 24454 65910 24506
rect 65910 24454 65956 24506
rect 65660 24452 65716 24454
rect 65740 24452 65796 24454
rect 65820 24452 65876 24454
rect 65900 24452 65956 24454
rect 50300 23962 50356 23964
rect 50380 23962 50436 23964
rect 50460 23962 50516 23964
rect 50540 23962 50596 23964
rect 50300 23910 50346 23962
rect 50346 23910 50356 23962
rect 50380 23910 50410 23962
rect 50410 23910 50422 23962
rect 50422 23910 50436 23962
rect 50460 23910 50474 23962
rect 50474 23910 50486 23962
rect 50486 23910 50516 23962
rect 50540 23910 50550 23962
rect 50550 23910 50596 23962
rect 50300 23908 50356 23910
rect 50380 23908 50436 23910
rect 50460 23908 50516 23910
rect 50540 23908 50596 23910
rect 65660 23418 65716 23420
rect 65740 23418 65796 23420
rect 65820 23418 65876 23420
rect 65900 23418 65956 23420
rect 65660 23366 65706 23418
rect 65706 23366 65716 23418
rect 65740 23366 65770 23418
rect 65770 23366 65782 23418
rect 65782 23366 65796 23418
rect 65820 23366 65834 23418
rect 65834 23366 65846 23418
rect 65846 23366 65876 23418
rect 65900 23366 65910 23418
rect 65910 23366 65956 23418
rect 65660 23364 65716 23366
rect 65740 23364 65796 23366
rect 65820 23364 65876 23366
rect 65900 23364 65956 23366
rect 67546 23160 67602 23216
rect 50300 22874 50356 22876
rect 50380 22874 50436 22876
rect 50460 22874 50516 22876
rect 50540 22874 50596 22876
rect 50300 22822 50346 22874
rect 50346 22822 50356 22874
rect 50380 22822 50410 22874
rect 50410 22822 50422 22874
rect 50422 22822 50436 22874
rect 50460 22822 50474 22874
rect 50474 22822 50486 22874
rect 50486 22822 50516 22874
rect 50540 22822 50550 22874
rect 50550 22822 50596 22874
rect 50300 22820 50356 22822
rect 50380 22820 50436 22822
rect 50460 22820 50516 22822
rect 50540 22820 50596 22822
rect 65660 22330 65716 22332
rect 65740 22330 65796 22332
rect 65820 22330 65876 22332
rect 65900 22330 65956 22332
rect 65660 22278 65706 22330
rect 65706 22278 65716 22330
rect 65740 22278 65770 22330
rect 65770 22278 65782 22330
rect 65782 22278 65796 22330
rect 65820 22278 65834 22330
rect 65834 22278 65846 22330
rect 65846 22278 65876 22330
rect 65900 22278 65910 22330
rect 65910 22278 65956 22330
rect 65660 22276 65716 22278
rect 65740 22276 65796 22278
rect 65820 22276 65876 22278
rect 65900 22276 65956 22278
rect 50300 21786 50356 21788
rect 50380 21786 50436 21788
rect 50460 21786 50516 21788
rect 50540 21786 50596 21788
rect 50300 21734 50346 21786
rect 50346 21734 50356 21786
rect 50380 21734 50410 21786
rect 50410 21734 50422 21786
rect 50422 21734 50436 21786
rect 50460 21734 50474 21786
rect 50474 21734 50486 21786
rect 50486 21734 50516 21786
rect 50540 21734 50550 21786
rect 50550 21734 50596 21786
rect 50300 21732 50356 21734
rect 50380 21732 50436 21734
rect 50460 21732 50516 21734
rect 50540 21732 50596 21734
rect 68098 21664 68154 21720
rect 65660 21242 65716 21244
rect 65740 21242 65796 21244
rect 65820 21242 65876 21244
rect 65900 21242 65956 21244
rect 65660 21190 65706 21242
rect 65706 21190 65716 21242
rect 65740 21190 65770 21242
rect 65770 21190 65782 21242
rect 65782 21190 65796 21242
rect 65820 21190 65834 21242
rect 65834 21190 65846 21242
rect 65846 21190 65876 21242
rect 65900 21190 65910 21242
rect 65910 21190 65956 21242
rect 65660 21188 65716 21190
rect 65740 21188 65796 21190
rect 65820 21188 65876 21190
rect 65900 21188 65956 21190
rect 50300 20698 50356 20700
rect 50380 20698 50436 20700
rect 50460 20698 50516 20700
rect 50540 20698 50596 20700
rect 50300 20646 50346 20698
rect 50346 20646 50356 20698
rect 50380 20646 50410 20698
rect 50410 20646 50422 20698
rect 50422 20646 50436 20698
rect 50460 20646 50474 20698
rect 50474 20646 50486 20698
rect 50486 20646 50516 20698
rect 50540 20646 50550 20698
rect 50550 20646 50596 20698
rect 50300 20644 50356 20646
rect 50380 20644 50436 20646
rect 50460 20644 50516 20646
rect 50540 20644 50596 20646
rect 67638 20204 67640 20224
rect 67640 20204 67692 20224
rect 67692 20204 67694 20224
rect 67638 20168 67694 20204
rect 65660 20154 65716 20156
rect 65740 20154 65796 20156
rect 65820 20154 65876 20156
rect 65900 20154 65956 20156
rect 65660 20102 65706 20154
rect 65706 20102 65716 20154
rect 65740 20102 65770 20154
rect 65770 20102 65782 20154
rect 65782 20102 65796 20154
rect 65820 20102 65834 20154
rect 65834 20102 65846 20154
rect 65846 20102 65876 20154
rect 65900 20102 65910 20154
rect 65910 20102 65956 20154
rect 65660 20100 65716 20102
rect 65740 20100 65796 20102
rect 65820 20100 65876 20102
rect 65900 20100 65956 20102
rect 50300 19610 50356 19612
rect 50380 19610 50436 19612
rect 50460 19610 50516 19612
rect 50540 19610 50596 19612
rect 50300 19558 50346 19610
rect 50346 19558 50356 19610
rect 50380 19558 50410 19610
rect 50410 19558 50422 19610
rect 50422 19558 50436 19610
rect 50460 19558 50474 19610
rect 50474 19558 50486 19610
rect 50486 19558 50516 19610
rect 50540 19558 50550 19610
rect 50550 19558 50596 19610
rect 50300 19556 50356 19558
rect 50380 19556 50436 19558
rect 50460 19556 50516 19558
rect 50540 19556 50596 19558
rect 65660 19066 65716 19068
rect 65740 19066 65796 19068
rect 65820 19066 65876 19068
rect 65900 19066 65956 19068
rect 65660 19014 65706 19066
rect 65706 19014 65716 19066
rect 65740 19014 65770 19066
rect 65770 19014 65782 19066
rect 65782 19014 65796 19066
rect 65820 19014 65834 19066
rect 65834 19014 65846 19066
rect 65846 19014 65876 19066
rect 65900 19014 65910 19066
rect 65910 19014 65956 19066
rect 65660 19012 65716 19014
rect 65740 19012 65796 19014
rect 65820 19012 65876 19014
rect 65900 19012 65956 19014
rect 68098 18708 68100 18728
rect 68100 18708 68152 18728
rect 68152 18708 68154 18728
rect 68098 18672 68154 18708
rect 50300 18522 50356 18524
rect 50380 18522 50436 18524
rect 50460 18522 50516 18524
rect 50540 18522 50596 18524
rect 50300 18470 50346 18522
rect 50346 18470 50356 18522
rect 50380 18470 50410 18522
rect 50410 18470 50422 18522
rect 50422 18470 50436 18522
rect 50460 18470 50474 18522
rect 50474 18470 50486 18522
rect 50486 18470 50516 18522
rect 50540 18470 50550 18522
rect 50550 18470 50596 18522
rect 50300 18468 50356 18470
rect 50380 18468 50436 18470
rect 50460 18468 50516 18470
rect 50540 18468 50596 18470
rect 65660 17978 65716 17980
rect 65740 17978 65796 17980
rect 65820 17978 65876 17980
rect 65900 17978 65956 17980
rect 65660 17926 65706 17978
rect 65706 17926 65716 17978
rect 65740 17926 65770 17978
rect 65770 17926 65782 17978
rect 65782 17926 65796 17978
rect 65820 17926 65834 17978
rect 65834 17926 65846 17978
rect 65846 17926 65876 17978
rect 65900 17926 65910 17978
rect 65910 17926 65956 17978
rect 65660 17924 65716 17926
rect 65740 17924 65796 17926
rect 65820 17924 65876 17926
rect 65900 17924 65956 17926
rect 50300 17434 50356 17436
rect 50380 17434 50436 17436
rect 50460 17434 50516 17436
rect 50540 17434 50596 17436
rect 50300 17382 50346 17434
rect 50346 17382 50356 17434
rect 50380 17382 50410 17434
rect 50410 17382 50422 17434
rect 50422 17382 50436 17434
rect 50460 17382 50474 17434
rect 50474 17382 50486 17434
rect 50486 17382 50516 17434
rect 50540 17382 50550 17434
rect 50550 17382 50596 17434
rect 50300 17380 50356 17382
rect 50380 17380 50436 17382
rect 50460 17380 50516 17382
rect 50540 17380 50596 17382
rect 68098 17176 68154 17232
rect 65660 16890 65716 16892
rect 65740 16890 65796 16892
rect 65820 16890 65876 16892
rect 65900 16890 65956 16892
rect 65660 16838 65706 16890
rect 65706 16838 65716 16890
rect 65740 16838 65770 16890
rect 65770 16838 65782 16890
rect 65782 16838 65796 16890
rect 65820 16838 65834 16890
rect 65834 16838 65846 16890
rect 65846 16838 65876 16890
rect 65900 16838 65910 16890
rect 65910 16838 65956 16890
rect 65660 16836 65716 16838
rect 65740 16836 65796 16838
rect 65820 16836 65876 16838
rect 65900 16836 65956 16838
rect 50300 16346 50356 16348
rect 50380 16346 50436 16348
rect 50460 16346 50516 16348
rect 50540 16346 50596 16348
rect 50300 16294 50346 16346
rect 50346 16294 50356 16346
rect 50380 16294 50410 16346
rect 50410 16294 50422 16346
rect 50422 16294 50436 16346
rect 50460 16294 50474 16346
rect 50474 16294 50486 16346
rect 50486 16294 50516 16346
rect 50540 16294 50550 16346
rect 50550 16294 50596 16346
rect 50300 16292 50356 16294
rect 50380 16292 50436 16294
rect 50460 16292 50516 16294
rect 50540 16292 50596 16294
rect 65660 15802 65716 15804
rect 65740 15802 65796 15804
rect 65820 15802 65876 15804
rect 65900 15802 65956 15804
rect 65660 15750 65706 15802
rect 65706 15750 65716 15802
rect 65740 15750 65770 15802
rect 65770 15750 65782 15802
rect 65782 15750 65796 15802
rect 65820 15750 65834 15802
rect 65834 15750 65846 15802
rect 65846 15750 65876 15802
rect 65900 15750 65910 15802
rect 65910 15750 65956 15802
rect 65660 15748 65716 15750
rect 65740 15748 65796 15750
rect 65820 15748 65876 15750
rect 65900 15748 65956 15750
rect 67638 15680 67694 15736
rect 50300 15258 50356 15260
rect 50380 15258 50436 15260
rect 50460 15258 50516 15260
rect 50540 15258 50596 15260
rect 50300 15206 50346 15258
rect 50346 15206 50356 15258
rect 50380 15206 50410 15258
rect 50410 15206 50422 15258
rect 50422 15206 50436 15258
rect 50460 15206 50474 15258
rect 50474 15206 50486 15258
rect 50486 15206 50516 15258
rect 50540 15206 50550 15258
rect 50550 15206 50596 15258
rect 50300 15204 50356 15206
rect 50380 15204 50436 15206
rect 50460 15204 50516 15206
rect 50540 15204 50596 15206
rect 65660 14714 65716 14716
rect 65740 14714 65796 14716
rect 65820 14714 65876 14716
rect 65900 14714 65956 14716
rect 65660 14662 65706 14714
rect 65706 14662 65716 14714
rect 65740 14662 65770 14714
rect 65770 14662 65782 14714
rect 65782 14662 65796 14714
rect 65820 14662 65834 14714
rect 65834 14662 65846 14714
rect 65846 14662 65876 14714
rect 65900 14662 65910 14714
rect 65910 14662 65956 14714
rect 65660 14660 65716 14662
rect 65740 14660 65796 14662
rect 65820 14660 65876 14662
rect 65900 14660 65956 14662
rect 68098 14184 68154 14240
rect 50300 14170 50356 14172
rect 50380 14170 50436 14172
rect 50460 14170 50516 14172
rect 50540 14170 50596 14172
rect 50300 14118 50346 14170
rect 50346 14118 50356 14170
rect 50380 14118 50410 14170
rect 50410 14118 50422 14170
rect 50422 14118 50436 14170
rect 50460 14118 50474 14170
rect 50474 14118 50486 14170
rect 50486 14118 50516 14170
rect 50540 14118 50550 14170
rect 50550 14118 50596 14170
rect 50300 14116 50356 14118
rect 50380 14116 50436 14118
rect 50460 14116 50516 14118
rect 50540 14116 50596 14118
rect 65660 13626 65716 13628
rect 65740 13626 65796 13628
rect 65820 13626 65876 13628
rect 65900 13626 65956 13628
rect 65660 13574 65706 13626
rect 65706 13574 65716 13626
rect 65740 13574 65770 13626
rect 65770 13574 65782 13626
rect 65782 13574 65796 13626
rect 65820 13574 65834 13626
rect 65834 13574 65846 13626
rect 65846 13574 65876 13626
rect 65900 13574 65910 13626
rect 65910 13574 65956 13626
rect 65660 13572 65716 13574
rect 65740 13572 65796 13574
rect 65820 13572 65876 13574
rect 65900 13572 65956 13574
rect 50300 13082 50356 13084
rect 50380 13082 50436 13084
rect 50460 13082 50516 13084
rect 50540 13082 50596 13084
rect 50300 13030 50346 13082
rect 50346 13030 50356 13082
rect 50380 13030 50410 13082
rect 50410 13030 50422 13082
rect 50422 13030 50436 13082
rect 50460 13030 50474 13082
rect 50474 13030 50486 13082
rect 50486 13030 50516 13082
rect 50540 13030 50550 13082
rect 50550 13030 50596 13082
rect 50300 13028 50356 13030
rect 50380 13028 50436 13030
rect 50460 13028 50516 13030
rect 50540 13028 50596 13030
rect 67638 12708 67694 12744
rect 67638 12688 67640 12708
rect 67640 12688 67692 12708
rect 67692 12688 67694 12708
rect 65660 12538 65716 12540
rect 65740 12538 65796 12540
rect 65820 12538 65876 12540
rect 65900 12538 65956 12540
rect 65660 12486 65706 12538
rect 65706 12486 65716 12538
rect 65740 12486 65770 12538
rect 65770 12486 65782 12538
rect 65782 12486 65796 12538
rect 65820 12486 65834 12538
rect 65834 12486 65846 12538
rect 65846 12486 65876 12538
rect 65900 12486 65910 12538
rect 65910 12486 65956 12538
rect 65660 12484 65716 12486
rect 65740 12484 65796 12486
rect 65820 12484 65876 12486
rect 65900 12484 65956 12486
rect 50300 11994 50356 11996
rect 50380 11994 50436 11996
rect 50460 11994 50516 11996
rect 50540 11994 50596 11996
rect 50300 11942 50346 11994
rect 50346 11942 50356 11994
rect 50380 11942 50410 11994
rect 50410 11942 50422 11994
rect 50422 11942 50436 11994
rect 50460 11942 50474 11994
rect 50474 11942 50486 11994
rect 50486 11942 50516 11994
rect 50540 11942 50550 11994
rect 50550 11942 50596 11994
rect 50300 11940 50356 11942
rect 50380 11940 50436 11942
rect 50460 11940 50516 11942
rect 50540 11940 50596 11942
rect 65660 11450 65716 11452
rect 65740 11450 65796 11452
rect 65820 11450 65876 11452
rect 65900 11450 65956 11452
rect 65660 11398 65706 11450
rect 65706 11398 65716 11450
rect 65740 11398 65770 11450
rect 65770 11398 65782 11450
rect 65782 11398 65796 11450
rect 65820 11398 65834 11450
rect 65834 11398 65846 11450
rect 65846 11398 65876 11450
rect 65900 11398 65910 11450
rect 65910 11398 65956 11450
rect 65660 11396 65716 11398
rect 65740 11396 65796 11398
rect 65820 11396 65876 11398
rect 65900 11396 65956 11398
rect 67638 11192 67694 11248
rect 50300 10906 50356 10908
rect 50380 10906 50436 10908
rect 50460 10906 50516 10908
rect 50540 10906 50596 10908
rect 50300 10854 50346 10906
rect 50346 10854 50356 10906
rect 50380 10854 50410 10906
rect 50410 10854 50422 10906
rect 50422 10854 50436 10906
rect 50460 10854 50474 10906
rect 50474 10854 50486 10906
rect 50486 10854 50516 10906
rect 50540 10854 50550 10906
rect 50550 10854 50596 10906
rect 50300 10852 50356 10854
rect 50380 10852 50436 10854
rect 50460 10852 50516 10854
rect 50540 10852 50596 10854
rect 65660 10362 65716 10364
rect 65740 10362 65796 10364
rect 65820 10362 65876 10364
rect 65900 10362 65956 10364
rect 65660 10310 65706 10362
rect 65706 10310 65716 10362
rect 65740 10310 65770 10362
rect 65770 10310 65782 10362
rect 65782 10310 65796 10362
rect 65820 10310 65834 10362
rect 65834 10310 65846 10362
rect 65846 10310 65876 10362
rect 65900 10310 65910 10362
rect 65910 10310 65956 10362
rect 65660 10308 65716 10310
rect 65740 10308 65796 10310
rect 65820 10308 65876 10310
rect 65900 10308 65956 10310
rect 50300 9818 50356 9820
rect 50380 9818 50436 9820
rect 50460 9818 50516 9820
rect 50540 9818 50596 9820
rect 50300 9766 50346 9818
rect 50346 9766 50356 9818
rect 50380 9766 50410 9818
rect 50410 9766 50422 9818
rect 50422 9766 50436 9818
rect 50460 9766 50474 9818
rect 50474 9766 50486 9818
rect 50486 9766 50516 9818
rect 50540 9766 50550 9818
rect 50550 9766 50596 9818
rect 50300 9764 50356 9766
rect 50380 9764 50436 9766
rect 50460 9764 50516 9766
rect 50540 9764 50596 9766
rect 68098 9696 68154 9752
rect 65660 9274 65716 9276
rect 65740 9274 65796 9276
rect 65820 9274 65876 9276
rect 65900 9274 65956 9276
rect 65660 9222 65706 9274
rect 65706 9222 65716 9274
rect 65740 9222 65770 9274
rect 65770 9222 65782 9274
rect 65782 9222 65796 9274
rect 65820 9222 65834 9274
rect 65834 9222 65846 9274
rect 65846 9222 65876 9274
rect 65900 9222 65910 9274
rect 65910 9222 65956 9274
rect 65660 9220 65716 9222
rect 65740 9220 65796 9222
rect 65820 9220 65876 9222
rect 65900 9220 65956 9222
rect 50300 8730 50356 8732
rect 50380 8730 50436 8732
rect 50460 8730 50516 8732
rect 50540 8730 50596 8732
rect 50300 8678 50346 8730
rect 50346 8678 50356 8730
rect 50380 8678 50410 8730
rect 50410 8678 50422 8730
rect 50422 8678 50436 8730
rect 50460 8678 50474 8730
rect 50474 8678 50486 8730
rect 50486 8678 50516 8730
rect 50540 8678 50550 8730
rect 50550 8678 50596 8730
rect 50300 8676 50356 8678
rect 50380 8676 50436 8678
rect 50460 8676 50516 8678
rect 50540 8676 50596 8678
rect 67546 8200 67602 8256
rect 65660 8186 65716 8188
rect 65740 8186 65796 8188
rect 65820 8186 65876 8188
rect 65900 8186 65956 8188
rect 65660 8134 65706 8186
rect 65706 8134 65716 8186
rect 65740 8134 65770 8186
rect 65770 8134 65782 8186
rect 65782 8134 65796 8186
rect 65820 8134 65834 8186
rect 65834 8134 65846 8186
rect 65846 8134 65876 8186
rect 65900 8134 65910 8186
rect 65910 8134 65956 8186
rect 65660 8132 65716 8134
rect 65740 8132 65796 8134
rect 65820 8132 65876 8134
rect 65900 8132 65956 8134
rect 50300 7642 50356 7644
rect 50380 7642 50436 7644
rect 50460 7642 50516 7644
rect 50540 7642 50596 7644
rect 50300 7590 50346 7642
rect 50346 7590 50356 7642
rect 50380 7590 50410 7642
rect 50410 7590 50422 7642
rect 50422 7590 50436 7642
rect 50460 7590 50474 7642
rect 50474 7590 50486 7642
rect 50486 7590 50516 7642
rect 50540 7590 50550 7642
rect 50550 7590 50596 7642
rect 50300 7588 50356 7590
rect 50380 7588 50436 7590
rect 50460 7588 50516 7590
rect 50540 7588 50596 7590
rect 65660 7098 65716 7100
rect 65740 7098 65796 7100
rect 65820 7098 65876 7100
rect 65900 7098 65956 7100
rect 65660 7046 65706 7098
rect 65706 7046 65716 7098
rect 65740 7046 65770 7098
rect 65770 7046 65782 7098
rect 65782 7046 65796 7098
rect 65820 7046 65834 7098
rect 65834 7046 65846 7098
rect 65846 7046 65876 7098
rect 65900 7046 65910 7098
rect 65910 7046 65956 7098
rect 65660 7044 65716 7046
rect 65740 7044 65796 7046
rect 65820 7044 65876 7046
rect 65900 7044 65956 7046
rect 68098 6740 68100 6760
rect 68100 6740 68152 6760
rect 68152 6740 68154 6760
rect 68098 6704 68154 6740
rect 50300 6554 50356 6556
rect 50380 6554 50436 6556
rect 50460 6554 50516 6556
rect 50540 6554 50596 6556
rect 50300 6502 50346 6554
rect 50346 6502 50356 6554
rect 50380 6502 50410 6554
rect 50410 6502 50422 6554
rect 50422 6502 50436 6554
rect 50460 6502 50474 6554
rect 50474 6502 50486 6554
rect 50486 6502 50516 6554
rect 50540 6502 50550 6554
rect 50550 6502 50596 6554
rect 50300 6500 50356 6502
rect 50380 6500 50436 6502
rect 50460 6500 50516 6502
rect 50540 6500 50596 6502
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 65660 6010 65716 6012
rect 65740 6010 65796 6012
rect 65820 6010 65876 6012
rect 65900 6010 65956 6012
rect 65660 5958 65706 6010
rect 65706 5958 65716 6010
rect 65740 5958 65770 6010
rect 65770 5958 65782 6010
rect 65782 5958 65796 6010
rect 65820 5958 65834 6010
rect 65834 5958 65846 6010
rect 65846 5958 65876 6010
rect 65900 5958 65910 6010
rect 65910 5958 65956 6010
rect 65660 5956 65716 5958
rect 65740 5956 65796 5958
rect 65820 5956 65876 5958
rect 65900 5956 65956 5958
rect 50300 5466 50356 5468
rect 50380 5466 50436 5468
rect 50460 5466 50516 5468
rect 50540 5466 50596 5468
rect 50300 5414 50346 5466
rect 50346 5414 50356 5466
rect 50380 5414 50410 5466
rect 50410 5414 50422 5466
rect 50422 5414 50436 5466
rect 50460 5414 50474 5466
rect 50474 5414 50486 5466
rect 50486 5414 50516 5466
rect 50540 5414 50550 5466
rect 50550 5414 50596 5466
rect 50300 5412 50356 5414
rect 50380 5412 50436 5414
rect 50460 5412 50516 5414
rect 50540 5412 50596 5414
rect 68098 5208 68154 5264
rect 50300 4378 50356 4380
rect 50380 4378 50436 4380
rect 50460 4378 50516 4380
rect 50540 4378 50596 4380
rect 50300 4326 50346 4378
rect 50346 4326 50356 4378
rect 50380 4326 50410 4378
rect 50410 4326 50422 4378
rect 50422 4326 50436 4378
rect 50460 4326 50474 4378
rect 50474 4326 50486 4378
rect 50486 4326 50516 4378
rect 50540 4326 50550 4378
rect 50550 4326 50596 4378
rect 50300 4324 50356 4326
rect 50380 4324 50436 4326
rect 50460 4324 50516 4326
rect 50540 4324 50596 4326
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 50300 3290 50356 3292
rect 50380 3290 50436 3292
rect 50460 3290 50516 3292
rect 50540 3290 50596 3292
rect 50300 3238 50346 3290
rect 50346 3238 50356 3290
rect 50380 3238 50410 3290
rect 50410 3238 50422 3290
rect 50422 3238 50436 3290
rect 50460 3238 50474 3290
rect 50474 3238 50486 3290
rect 50486 3238 50516 3290
rect 50540 3238 50550 3290
rect 50550 3238 50596 3290
rect 50300 3236 50356 3238
rect 50380 3236 50436 3238
rect 50460 3236 50516 3238
rect 50540 3236 50596 3238
rect 50300 2202 50356 2204
rect 50380 2202 50436 2204
rect 50460 2202 50516 2204
rect 50540 2202 50596 2204
rect 50300 2150 50346 2202
rect 50346 2150 50356 2202
rect 50380 2150 50410 2202
rect 50410 2150 50422 2202
rect 50422 2150 50436 2202
rect 50460 2150 50474 2202
rect 50474 2150 50486 2202
rect 50486 2150 50516 2202
rect 50540 2150 50550 2202
rect 50550 2150 50596 2202
rect 50300 2148 50356 2150
rect 50380 2148 50436 2150
rect 50460 2148 50516 2150
rect 50540 2148 50596 2150
rect 57886 3168 57942 3224
rect 65660 4922 65716 4924
rect 65740 4922 65796 4924
rect 65820 4922 65876 4924
rect 65900 4922 65956 4924
rect 65660 4870 65706 4922
rect 65706 4870 65716 4922
rect 65740 4870 65770 4922
rect 65770 4870 65782 4922
rect 65782 4870 65796 4922
rect 65820 4870 65834 4922
rect 65834 4870 65846 4922
rect 65846 4870 65876 4922
rect 65900 4870 65910 4922
rect 65910 4870 65956 4922
rect 65660 4868 65716 4870
rect 65740 4868 65796 4870
rect 65820 4868 65876 4870
rect 65900 4868 65956 4870
rect 65660 3834 65716 3836
rect 65740 3834 65796 3836
rect 65820 3834 65876 3836
rect 65900 3834 65956 3836
rect 65660 3782 65706 3834
rect 65706 3782 65716 3834
rect 65740 3782 65770 3834
rect 65770 3782 65782 3834
rect 65782 3782 65796 3834
rect 65820 3782 65834 3834
rect 65834 3782 65846 3834
rect 65846 3782 65876 3834
rect 65900 3782 65910 3834
rect 65910 3782 65956 3834
rect 65660 3780 65716 3782
rect 65740 3780 65796 3782
rect 65820 3780 65876 3782
rect 65900 3780 65956 3782
rect 67638 3712 67694 3768
rect 60462 3168 60518 3224
rect 65660 2746 65716 2748
rect 65740 2746 65796 2748
rect 65820 2746 65876 2748
rect 65900 2746 65956 2748
rect 65660 2694 65706 2746
rect 65706 2694 65716 2746
rect 65740 2694 65770 2746
rect 65770 2694 65782 2746
rect 65782 2694 65796 2746
rect 65820 2694 65834 2746
rect 65834 2694 65846 2746
rect 65846 2694 65876 2746
rect 65900 2694 65910 2746
rect 65910 2694 65956 2746
rect 65660 2692 65716 2694
rect 65740 2692 65796 2694
rect 65820 2692 65876 2694
rect 65900 2692 65956 2694
rect 67638 2216 67694 2272
<< metal3 >>
rect 19570 57696 19886 57697
rect 0 57536 800 57656
rect 19570 57632 19576 57696
rect 19640 57632 19656 57696
rect 19720 57632 19736 57696
rect 19800 57632 19816 57696
rect 19880 57632 19886 57696
rect 19570 57631 19886 57632
rect 50290 57696 50606 57697
rect 50290 57632 50296 57696
rect 50360 57632 50376 57696
rect 50440 57632 50456 57696
rect 50520 57632 50536 57696
rect 50600 57632 50606 57696
rect 50290 57631 50606 57632
rect 67633 57626 67699 57629
rect 69200 57626 70000 57656
rect 67633 57624 70000 57626
rect 67633 57568 67638 57624
rect 67694 57568 70000 57624
rect 67633 57566 70000 57568
rect 67633 57563 67699 57566
rect 69200 57536 70000 57566
rect 4210 57152 4526 57153
rect 4210 57088 4216 57152
rect 4280 57088 4296 57152
rect 4360 57088 4376 57152
rect 4440 57088 4456 57152
rect 4520 57088 4526 57152
rect 4210 57087 4526 57088
rect 34930 57152 35246 57153
rect 34930 57088 34936 57152
rect 35000 57088 35016 57152
rect 35080 57088 35096 57152
rect 35160 57088 35176 57152
rect 35240 57088 35246 57152
rect 34930 57087 35246 57088
rect 65650 57152 65966 57153
rect 65650 57088 65656 57152
rect 65720 57088 65736 57152
rect 65800 57088 65816 57152
rect 65880 57088 65896 57152
rect 65960 57088 65966 57152
rect 65650 57087 65966 57088
rect 19570 56608 19886 56609
rect 19570 56544 19576 56608
rect 19640 56544 19656 56608
rect 19720 56544 19736 56608
rect 19800 56544 19816 56608
rect 19880 56544 19886 56608
rect 19570 56543 19886 56544
rect 50290 56608 50606 56609
rect 50290 56544 50296 56608
rect 50360 56544 50376 56608
rect 50440 56544 50456 56608
rect 50520 56544 50536 56608
rect 50600 56544 50606 56608
rect 50290 56543 50606 56544
rect 0 56040 800 56160
rect 67633 56130 67699 56133
rect 69200 56130 70000 56160
rect 67633 56128 70000 56130
rect 67633 56072 67638 56128
rect 67694 56072 70000 56128
rect 67633 56070 70000 56072
rect 67633 56067 67699 56070
rect 4210 56064 4526 56065
rect 4210 56000 4216 56064
rect 4280 56000 4296 56064
rect 4360 56000 4376 56064
rect 4440 56000 4456 56064
rect 4520 56000 4526 56064
rect 4210 55999 4526 56000
rect 34930 56064 35246 56065
rect 34930 56000 34936 56064
rect 35000 56000 35016 56064
rect 35080 56000 35096 56064
rect 35160 56000 35176 56064
rect 35240 56000 35246 56064
rect 34930 55999 35246 56000
rect 65650 56064 65966 56065
rect 65650 56000 65656 56064
rect 65720 56000 65736 56064
rect 65800 56000 65816 56064
rect 65880 56000 65896 56064
rect 65960 56000 65966 56064
rect 69200 56040 70000 56070
rect 65650 55999 65966 56000
rect 19570 55520 19886 55521
rect 19570 55456 19576 55520
rect 19640 55456 19656 55520
rect 19720 55456 19736 55520
rect 19800 55456 19816 55520
rect 19880 55456 19886 55520
rect 19570 55455 19886 55456
rect 50290 55520 50606 55521
rect 50290 55456 50296 55520
rect 50360 55456 50376 55520
rect 50440 55456 50456 55520
rect 50520 55456 50536 55520
rect 50600 55456 50606 55520
rect 50290 55455 50606 55456
rect 4210 54976 4526 54977
rect 4210 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4526 54976
rect 4210 54911 4526 54912
rect 34930 54976 35246 54977
rect 34930 54912 34936 54976
rect 35000 54912 35016 54976
rect 35080 54912 35096 54976
rect 35160 54912 35176 54976
rect 35240 54912 35246 54976
rect 34930 54911 35246 54912
rect 65650 54976 65966 54977
rect 65650 54912 65656 54976
rect 65720 54912 65736 54976
rect 65800 54912 65816 54976
rect 65880 54912 65896 54976
rect 65960 54912 65966 54976
rect 65650 54911 65966 54912
rect 0 54544 800 54664
rect 68093 54634 68159 54637
rect 69200 54634 70000 54664
rect 68093 54632 70000 54634
rect 68093 54576 68098 54632
rect 68154 54576 70000 54632
rect 68093 54574 70000 54576
rect 68093 54571 68159 54574
rect 69200 54544 70000 54574
rect 19570 54432 19886 54433
rect 19570 54368 19576 54432
rect 19640 54368 19656 54432
rect 19720 54368 19736 54432
rect 19800 54368 19816 54432
rect 19880 54368 19886 54432
rect 19570 54367 19886 54368
rect 50290 54432 50606 54433
rect 50290 54368 50296 54432
rect 50360 54368 50376 54432
rect 50440 54368 50456 54432
rect 50520 54368 50536 54432
rect 50600 54368 50606 54432
rect 50290 54367 50606 54368
rect 4210 53888 4526 53889
rect 4210 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4526 53888
rect 4210 53823 4526 53824
rect 34930 53888 35246 53889
rect 34930 53824 34936 53888
rect 35000 53824 35016 53888
rect 35080 53824 35096 53888
rect 35160 53824 35176 53888
rect 35240 53824 35246 53888
rect 34930 53823 35246 53824
rect 65650 53888 65966 53889
rect 65650 53824 65656 53888
rect 65720 53824 65736 53888
rect 65800 53824 65816 53888
rect 65880 53824 65896 53888
rect 65960 53824 65966 53888
rect 65650 53823 65966 53824
rect 19570 53344 19886 53345
rect 19570 53280 19576 53344
rect 19640 53280 19656 53344
rect 19720 53280 19736 53344
rect 19800 53280 19816 53344
rect 19880 53280 19886 53344
rect 19570 53279 19886 53280
rect 50290 53344 50606 53345
rect 50290 53280 50296 53344
rect 50360 53280 50376 53344
rect 50440 53280 50456 53344
rect 50520 53280 50536 53344
rect 50600 53280 50606 53344
rect 50290 53279 50606 53280
rect 0 53048 800 53168
rect 68093 53138 68159 53141
rect 69200 53138 70000 53168
rect 68093 53136 70000 53138
rect 68093 53080 68098 53136
rect 68154 53080 70000 53136
rect 68093 53078 70000 53080
rect 68093 53075 68159 53078
rect 69200 53048 70000 53078
rect 4210 52800 4526 52801
rect 4210 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4526 52800
rect 4210 52735 4526 52736
rect 34930 52800 35246 52801
rect 34930 52736 34936 52800
rect 35000 52736 35016 52800
rect 35080 52736 35096 52800
rect 35160 52736 35176 52800
rect 35240 52736 35246 52800
rect 34930 52735 35246 52736
rect 65650 52800 65966 52801
rect 65650 52736 65656 52800
rect 65720 52736 65736 52800
rect 65800 52736 65816 52800
rect 65880 52736 65896 52800
rect 65960 52736 65966 52800
rect 65650 52735 65966 52736
rect 19570 52256 19886 52257
rect 19570 52192 19576 52256
rect 19640 52192 19656 52256
rect 19720 52192 19736 52256
rect 19800 52192 19816 52256
rect 19880 52192 19886 52256
rect 19570 52191 19886 52192
rect 50290 52256 50606 52257
rect 50290 52192 50296 52256
rect 50360 52192 50376 52256
rect 50440 52192 50456 52256
rect 50520 52192 50536 52256
rect 50600 52192 50606 52256
rect 50290 52191 50606 52192
rect 4210 51712 4526 51713
rect 0 51552 800 51672
rect 4210 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4526 51712
rect 4210 51647 4526 51648
rect 34930 51712 35246 51713
rect 34930 51648 34936 51712
rect 35000 51648 35016 51712
rect 35080 51648 35096 51712
rect 35160 51648 35176 51712
rect 35240 51648 35246 51712
rect 34930 51647 35246 51648
rect 65650 51712 65966 51713
rect 65650 51648 65656 51712
rect 65720 51648 65736 51712
rect 65800 51648 65816 51712
rect 65880 51648 65896 51712
rect 65960 51648 65966 51712
rect 65650 51647 65966 51648
rect 67633 51642 67699 51645
rect 69200 51642 70000 51672
rect 67633 51640 70000 51642
rect 67633 51584 67638 51640
rect 67694 51584 70000 51640
rect 67633 51582 70000 51584
rect 67633 51579 67699 51582
rect 69200 51552 70000 51582
rect 19570 51168 19886 51169
rect 19570 51104 19576 51168
rect 19640 51104 19656 51168
rect 19720 51104 19736 51168
rect 19800 51104 19816 51168
rect 19880 51104 19886 51168
rect 19570 51103 19886 51104
rect 50290 51168 50606 51169
rect 50290 51104 50296 51168
rect 50360 51104 50376 51168
rect 50440 51104 50456 51168
rect 50520 51104 50536 51168
rect 50600 51104 50606 51168
rect 50290 51103 50606 51104
rect 4210 50624 4526 50625
rect 4210 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4526 50624
rect 4210 50559 4526 50560
rect 34930 50624 35246 50625
rect 34930 50560 34936 50624
rect 35000 50560 35016 50624
rect 35080 50560 35096 50624
rect 35160 50560 35176 50624
rect 35240 50560 35246 50624
rect 34930 50559 35246 50560
rect 65650 50624 65966 50625
rect 65650 50560 65656 50624
rect 65720 50560 65736 50624
rect 65800 50560 65816 50624
rect 65880 50560 65896 50624
rect 65960 50560 65966 50624
rect 65650 50559 65966 50560
rect 0 50056 800 50176
rect 68093 50146 68159 50149
rect 69200 50146 70000 50176
rect 68093 50144 70000 50146
rect 68093 50088 68098 50144
rect 68154 50088 70000 50144
rect 68093 50086 70000 50088
rect 68093 50083 68159 50086
rect 19570 50080 19886 50081
rect 19570 50016 19576 50080
rect 19640 50016 19656 50080
rect 19720 50016 19736 50080
rect 19800 50016 19816 50080
rect 19880 50016 19886 50080
rect 19570 50015 19886 50016
rect 50290 50080 50606 50081
rect 50290 50016 50296 50080
rect 50360 50016 50376 50080
rect 50440 50016 50456 50080
rect 50520 50016 50536 50080
rect 50600 50016 50606 50080
rect 69200 50056 70000 50086
rect 50290 50015 50606 50016
rect 4210 49536 4526 49537
rect 4210 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4526 49536
rect 4210 49471 4526 49472
rect 34930 49536 35246 49537
rect 34930 49472 34936 49536
rect 35000 49472 35016 49536
rect 35080 49472 35096 49536
rect 35160 49472 35176 49536
rect 35240 49472 35246 49536
rect 34930 49471 35246 49472
rect 65650 49536 65966 49537
rect 65650 49472 65656 49536
rect 65720 49472 65736 49536
rect 65800 49472 65816 49536
rect 65880 49472 65896 49536
rect 65960 49472 65966 49536
rect 65650 49471 65966 49472
rect 19570 48992 19886 48993
rect 19570 48928 19576 48992
rect 19640 48928 19656 48992
rect 19720 48928 19736 48992
rect 19800 48928 19816 48992
rect 19880 48928 19886 48992
rect 19570 48927 19886 48928
rect 50290 48992 50606 48993
rect 50290 48928 50296 48992
rect 50360 48928 50376 48992
rect 50440 48928 50456 48992
rect 50520 48928 50536 48992
rect 50600 48928 50606 48992
rect 50290 48927 50606 48928
rect 0 48560 800 48680
rect 67633 48650 67699 48653
rect 69200 48650 70000 48680
rect 67633 48648 70000 48650
rect 67633 48592 67638 48648
rect 67694 48592 70000 48648
rect 67633 48590 70000 48592
rect 67633 48587 67699 48590
rect 69200 48560 70000 48590
rect 4210 48448 4526 48449
rect 4210 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4526 48448
rect 4210 48383 4526 48384
rect 34930 48448 35246 48449
rect 34930 48384 34936 48448
rect 35000 48384 35016 48448
rect 35080 48384 35096 48448
rect 35160 48384 35176 48448
rect 35240 48384 35246 48448
rect 34930 48383 35246 48384
rect 65650 48448 65966 48449
rect 65650 48384 65656 48448
rect 65720 48384 65736 48448
rect 65800 48384 65816 48448
rect 65880 48384 65896 48448
rect 65960 48384 65966 48448
rect 65650 48383 65966 48384
rect 19570 47904 19886 47905
rect 19570 47840 19576 47904
rect 19640 47840 19656 47904
rect 19720 47840 19736 47904
rect 19800 47840 19816 47904
rect 19880 47840 19886 47904
rect 19570 47839 19886 47840
rect 50290 47904 50606 47905
rect 50290 47840 50296 47904
rect 50360 47840 50376 47904
rect 50440 47840 50456 47904
rect 50520 47840 50536 47904
rect 50600 47840 50606 47904
rect 50290 47839 50606 47840
rect 4210 47360 4526 47361
rect 4210 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4526 47360
rect 4210 47295 4526 47296
rect 34930 47360 35246 47361
rect 34930 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35246 47360
rect 34930 47295 35246 47296
rect 65650 47360 65966 47361
rect 65650 47296 65656 47360
rect 65720 47296 65736 47360
rect 65800 47296 65816 47360
rect 65880 47296 65896 47360
rect 65960 47296 65966 47360
rect 65650 47295 65966 47296
rect 0 47064 800 47184
rect 67633 47154 67699 47157
rect 69200 47154 70000 47184
rect 67633 47152 70000 47154
rect 67633 47096 67638 47152
rect 67694 47096 70000 47152
rect 67633 47094 70000 47096
rect 67633 47091 67699 47094
rect 69200 47064 70000 47094
rect 19570 46816 19886 46817
rect 19570 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19886 46816
rect 19570 46751 19886 46752
rect 50290 46816 50606 46817
rect 50290 46752 50296 46816
rect 50360 46752 50376 46816
rect 50440 46752 50456 46816
rect 50520 46752 50536 46816
rect 50600 46752 50606 46816
rect 50290 46751 50606 46752
rect 4210 46272 4526 46273
rect 4210 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4526 46272
rect 4210 46207 4526 46208
rect 34930 46272 35246 46273
rect 34930 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35246 46272
rect 34930 46207 35246 46208
rect 65650 46272 65966 46273
rect 65650 46208 65656 46272
rect 65720 46208 65736 46272
rect 65800 46208 65816 46272
rect 65880 46208 65896 46272
rect 65960 46208 65966 46272
rect 65650 46207 65966 46208
rect 19570 45728 19886 45729
rect 0 45568 800 45688
rect 19570 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19886 45728
rect 19570 45663 19886 45664
rect 50290 45728 50606 45729
rect 50290 45664 50296 45728
rect 50360 45664 50376 45728
rect 50440 45664 50456 45728
rect 50520 45664 50536 45728
rect 50600 45664 50606 45728
rect 50290 45663 50606 45664
rect 68093 45658 68159 45661
rect 69200 45658 70000 45688
rect 68093 45656 70000 45658
rect 68093 45600 68098 45656
rect 68154 45600 70000 45656
rect 68093 45598 70000 45600
rect 68093 45595 68159 45598
rect 69200 45568 70000 45598
rect 4210 45184 4526 45185
rect 4210 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4526 45184
rect 4210 45119 4526 45120
rect 34930 45184 35246 45185
rect 34930 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35246 45184
rect 34930 45119 35246 45120
rect 65650 45184 65966 45185
rect 65650 45120 65656 45184
rect 65720 45120 65736 45184
rect 65800 45120 65816 45184
rect 65880 45120 65896 45184
rect 65960 45120 65966 45184
rect 65650 45119 65966 45120
rect 19570 44640 19886 44641
rect 19570 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19886 44640
rect 19570 44575 19886 44576
rect 50290 44640 50606 44641
rect 50290 44576 50296 44640
rect 50360 44576 50376 44640
rect 50440 44576 50456 44640
rect 50520 44576 50536 44640
rect 50600 44576 50606 44640
rect 50290 44575 50606 44576
rect 0 44072 800 44192
rect 67541 44162 67607 44165
rect 69200 44162 70000 44192
rect 67541 44160 70000 44162
rect 67541 44104 67546 44160
rect 67602 44104 70000 44160
rect 67541 44102 70000 44104
rect 67541 44099 67607 44102
rect 4210 44096 4526 44097
rect 4210 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4526 44096
rect 4210 44031 4526 44032
rect 34930 44096 35246 44097
rect 34930 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35246 44096
rect 34930 44031 35246 44032
rect 65650 44096 65966 44097
rect 65650 44032 65656 44096
rect 65720 44032 65736 44096
rect 65800 44032 65816 44096
rect 65880 44032 65896 44096
rect 65960 44032 65966 44096
rect 69200 44072 70000 44102
rect 65650 44031 65966 44032
rect 19570 43552 19886 43553
rect 19570 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19886 43552
rect 19570 43487 19886 43488
rect 50290 43552 50606 43553
rect 50290 43488 50296 43552
rect 50360 43488 50376 43552
rect 50440 43488 50456 43552
rect 50520 43488 50536 43552
rect 50600 43488 50606 43552
rect 50290 43487 50606 43488
rect 4210 43008 4526 43009
rect 4210 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4526 43008
rect 4210 42943 4526 42944
rect 34930 43008 35246 43009
rect 34930 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35246 43008
rect 34930 42943 35246 42944
rect 65650 43008 65966 43009
rect 65650 42944 65656 43008
rect 65720 42944 65736 43008
rect 65800 42944 65816 43008
rect 65880 42944 65896 43008
rect 65960 42944 65966 43008
rect 65650 42943 65966 42944
rect 0 42576 800 42696
rect 68093 42666 68159 42669
rect 69200 42666 70000 42696
rect 68093 42664 70000 42666
rect 68093 42608 68098 42664
rect 68154 42608 70000 42664
rect 68093 42606 70000 42608
rect 68093 42603 68159 42606
rect 69200 42576 70000 42606
rect 19570 42464 19886 42465
rect 19570 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19886 42464
rect 19570 42399 19886 42400
rect 50290 42464 50606 42465
rect 50290 42400 50296 42464
rect 50360 42400 50376 42464
rect 50440 42400 50456 42464
rect 50520 42400 50536 42464
rect 50600 42400 50606 42464
rect 50290 42399 50606 42400
rect 4210 41920 4526 41921
rect 4210 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4526 41920
rect 4210 41855 4526 41856
rect 34930 41920 35246 41921
rect 34930 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35246 41920
rect 34930 41855 35246 41856
rect 65650 41920 65966 41921
rect 65650 41856 65656 41920
rect 65720 41856 65736 41920
rect 65800 41856 65816 41920
rect 65880 41856 65896 41920
rect 65960 41856 65966 41920
rect 65650 41855 65966 41856
rect 19570 41376 19886 41377
rect 19570 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19886 41376
rect 19570 41311 19886 41312
rect 50290 41376 50606 41377
rect 50290 41312 50296 41376
rect 50360 41312 50376 41376
rect 50440 41312 50456 41376
rect 50520 41312 50536 41376
rect 50600 41312 50606 41376
rect 50290 41311 50606 41312
rect 0 41080 800 41200
rect 68093 41170 68159 41173
rect 69200 41170 70000 41200
rect 68093 41168 70000 41170
rect 68093 41112 68098 41168
rect 68154 41112 70000 41168
rect 68093 41110 70000 41112
rect 68093 41107 68159 41110
rect 69200 41080 70000 41110
rect 4210 40832 4526 40833
rect 4210 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4526 40832
rect 4210 40767 4526 40768
rect 34930 40832 35246 40833
rect 34930 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35246 40832
rect 34930 40767 35246 40768
rect 65650 40832 65966 40833
rect 65650 40768 65656 40832
rect 65720 40768 65736 40832
rect 65800 40768 65816 40832
rect 65880 40768 65896 40832
rect 65960 40768 65966 40832
rect 65650 40767 65966 40768
rect 19570 40288 19886 40289
rect 19570 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19886 40288
rect 19570 40223 19886 40224
rect 50290 40288 50606 40289
rect 50290 40224 50296 40288
rect 50360 40224 50376 40288
rect 50440 40224 50456 40288
rect 50520 40224 50536 40288
rect 50600 40224 50606 40288
rect 50290 40223 50606 40224
rect 4210 39744 4526 39745
rect 0 39584 800 39704
rect 4210 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4526 39744
rect 4210 39679 4526 39680
rect 34930 39744 35246 39745
rect 34930 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35246 39744
rect 34930 39679 35246 39680
rect 65650 39744 65966 39745
rect 65650 39680 65656 39744
rect 65720 39680 65736 39744
rect 65800 39680 65816 39744
rect 65880 39680 65896 39744
rect 65960 39680 65966 39744
rect 65650 39679 65966 39680
rect 67633 39674 67699 39677
rect 69200 39674 70000 39704
rect 67633 39672 70000 39674
rect 67633 39616 67638 39672
rect 67694 39616 70000 39672
rect 67633 39614 70000 39616
rect 67633 39611 67699 39614
rect 69200 39584 70000 39614
rect 19570 39200 19886 39201
rect 19570 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19886 39200
rect 19570 39135 19886 39136
rect 50290 39200 50606 39201
rect 50290 39136 50296 39200
rect 50360 39136 50376 39200
rect 50440 39136 50456 39200
rect 50520 39136 50536 39200
rect 50600 39136 50606 39200
rect 50290 39135 50606 39136
rect 4210 38656 4526 38657
rect 4210 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4526 38656
rect 4210 38591 4526 38592
rect 34930 38656 35246 38657
rect 34930 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35246 38656
rect 34930 38591 35246 38592
rect 65650 38656 65966 38657
rect 65650 38592 65656 38656
rect 65720 38592 65736 38656
rect 65800 38592 65816 38656
rect 65880 38592 65896 38656
rect 65960 38592 65966 38656
rect 65650 38591 65966 38592
rect 0 38088 800 38208
rect 68093 38178 68159 38181
rect 69200 38178 70000 38208
rect 68093 38176 70000 38178
rect 68093 38120 68098 38176
rect 68154 38120 70000 38176
rect 68093 38118 70000 38120
rect 68093 38115 68159 38118
rect 19570 38112 19886 38113
rect 19570 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19886 38112
rect 19570 38047 19886 38048
rect 50290 38112 50606 38113
rect 50290 38048 50296 38112
rect 50360 38048 50376 38112
rect 50440 38048 50456 38112
rect 50520 38048 50536 38112
rect 50600 38048 50606 38112
rect 69200 38088 70000 38118
rect 50290 38047 50606 38048
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 65650 37568 65966 37569
rect 65650 37504 65656 37568
rect 65720 37504 65736 37568
rect 65800 37504 65816 37568
rect 65880 37504 65896 37568
rect 65960 37504 65966 37568
rect 65650 37503 65966 37504
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 50290 37024 50606 37025
rect 50290 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50606 37024
rect 50290 36959 50606 36960
rect 0 36592 800 36712
rect 67633 36682 67699 36685
rect 69200 36682 70000 36712
rect 67633 36680 70000 36682
rect 67633 36624 67638 36680
rect 67694 36624 70000 36680
rect 67633 36622 70000 36624
rect 67633 36619 67699 36622
rect 69200 36592 70000 36622
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 65650 36480 65966 36481
rect 65650 36416 65656 36480
rect 65720 36416 65736 36480
rect 65800 36416 65816 36480
rect 65880 36416 65896 36480
rect 65960 36416 65966 36480
rect 65650 36415 65966 36416
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 50290 35936 50606 35937
rect 50290 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50606 35936
rect 50290 35871 50606 35872
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 65650 35392 65966 35393
rect 65650 35328 65656 35392
rect 65720 35328 65736 35392
rect 65800 35328 65816 35392
rect 65880 35328 65896 35392
rect 65960 35328 65966 35392
rect 65650 35327 65966 35328
rect 0 35096 800 35216
rect 67633 35186 67699 35189
rect 69200 35186 70000 35216
rect 67633 35184 70000 35186
rect 67633 35128 67638 35184
rect 67694 35128 70000 35184
rect 67633 35126 70000 35128
rect 67633 35123 67699 35126
rect 69200 35096 70000 35126
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 50290 34848 50606 34849
rect 50290 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50606 34848
rect 50290 34783 50606 34784
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 65650 34304 65966 34305
rect 65650 34240 65656 34304
rect 65720 34240 65736 34304
rect 65800 34240 65816 34304
rect 65880 34240 65896 34304
rect 65960 34240 65966 34304
rect 65650 34239 65966 34240
rect 19570 33760 19886 33761
rect 0 33600 800 33720
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 50290 33760 50606 33761
rect 50290 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50606 33760
rect 50290 33695 50606 33696
rect 68093 33690 68159 33693
rect 69200 33690 70000 33720
rect 68093 33688 70000 33690
rect 68093 33632 68098 33688
rect 68154 33632 70000 33688
rect 68093 33630 70000 33632
rect 68093 33627 68159 33630
rect 69200 33600 70000 33630
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 65650 33216 65966 33217
rect 65650 33152 65656 33216
rect 65720 33152 65736 33216
rect 65800 33152 65816 33216
rect 65880 33152 65896 33216
rect 65960 33152 65966 33216
rect 65650 33151 65966 33152
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 19570 32607 19886 32608
rect 50290 32672 50606 32673
rect 50290 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50606 32672
rect 50290 32607 50606 32608
rect 0 32104 800 32224
rect 67633 32194 67699 32197
rect 69200 32194 70000 32224
rect 67633 32192 70000 32194
rect 67633 32136 67638 32192
rect 67694 32136 70000 32192
rect 67633 32134 70000 32136
rect 67633 32131 67699 32134
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 65650 32128 65966 32129
rect 65650 32064 65656 32128
rect 65720 32064 65736 32128
rect 65800 32064 65816 32128
rect 65880 32064 65896 32128
rect 65960 32064 65966 32128
rect 69200 32104 70000 32134
rect 65650 32063 65966 32064
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 50290 31584 50606 31585
rect 50290 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50606 31584
rect 50290 31519 50606 31520
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 65650 31040 65966 31041
rect 65650 30976 65656 31040
rect 65720 30976 65736 31040
rect 65800 30976 65816 31040
rect 65880 30976 65896 31040
rect 65960 30976 65966 31040
rect 65650 30975 65966 30976
rect 0 30608 800 30728
rect 68093 30698 68159 30701
rect 69200 30698 70000 30728
rect 68093 30696 70000 30698
rect 68093 30640 68098 30696
rect 68154 30640 70000 30696
rect 68093 30638 70000 30640
rect 68093 30635 68159 30638
rect 69200 30608 70000 30638
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 50290 30496 50606 30497
rect 50290 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50606 30496
rect 50290 30431 50606 30432
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 65650 29952 65966 29953
rect 65650 29888 65656 29952
rect 65720 29888 65736 29952
rect 65800 29888 65816 29952
rect 65880 29888 65896 29952
rect 65960 29888 65966 29952
rect 65650 29887 65966 29888
rect 19570 29408 19886 29409
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 50290 29408 50606 29409
rect 50290 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50606 29408
rect 50290 29343 50606 29344
rect 0 29112 800 29232
rect 68093 29202 68159 29205
rect 69200 29202 70000 29232
rect 68093 29200 70000 29202
rect 68093 29144 68098 29200
rect 68154 29144 70000 29200
rect 68093 29142 70000 29144
rect 68093 29139 68159 29142
rect 69200 29112 70000 29142
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 65650 28864 65966 28865
rect 65650 28800 65656 28864
rect 65720 28800 65736 28864
rect 65800 28800 65816 28864
rect 65880 28800 65896 28864
rect 65960 28800 65966 28864
rect 65650 28799 65966 28800
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 50290 28320 50606 28321
rect 50290 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50606 28320
rect 50290 28255 50606 28256
rect 4210 27776 4526 27777
rect 0 27616 800 27736
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 65650 27776 65966 27777
rect 65650 27712 65656 27776
rect 65720 27712 65736 27776
rect 65800 27712 65816 27776
rect 65880 27712 65896 27776
rect 65960 27712 65966 27776
rect 65650 27711 65966 27712
rect 23473 27708 23539 27709
rect 23422 27706 23428 27708
rect 23382 27646 23428 27706
rect 23492 27704 23539 27708
rect 23534 27648 23539 27704
rect 23422 27644 23428 27646
rect 23492 27644 23539 27648
rect 23473 27643 23539 27644
rect 67633 27706 67699 27709
rect 69200 27706 70000 27736
rect 67633 27704 70000 27706
rect 67633 27648 67638 27704
rect 67694 27648 70000 27704
rect 67633 27646 70000 27648
rect 67633 27643 67699 27646
rect 69200 27616 70000 27646
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 19570 27167 19886 27168
rect 50290 27232 50606 27233
rect 50290 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50606 27232
rect 50290 27167 50606 27168
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 65650 26688 65966 26689
rect 65650 26624 65656 26688
rect 65720 26624 65736 26688
rect 65800 26624 65816 26688
rect 65880 26624 65896 26688
rect 65960 26624 65966 26688
rect 65650 26623 65966 26624
rect 0 26120 800 26240
rect 68093 26210 68159 26213
rect 69200 26210 70000 26240
rect 68093 26208 70000 26210
rect 68093 26152 68098 26208
rect 68154 26152 70000 26208
rect 68093 26150 70000 26152
rect 68093 26147 68159 26150
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 50290 26144 50606 26145
rect 50290 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50606 26144
rect 69200 26120 70000 26150
rect 50290 26079 50606 26080
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 65650 25600 65966 25601
rect 65650 25536 65656 25600
rect 65720 25536 65736 25600
rect 65800 25536 65816 25600
rect 65880 25536 65896 25600
rect 65960 25536 65966 25600
rect 65650 25535 65966 25536
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 50290 25056 50606 25057
rect 50290 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50606 25056
rect 50290 24991 50606 24992
rect 0 24624 800 24744
rect 23381 24716 23447 24717
rect 23381 24714 23428 24716
rect 23336 24712 23428 24714
rect 23336 24656 23386 24712
rect 23336 24654 23428 24656
rect 23381 24652 23428 24654
rect 23492 24652 23498 24716
rect 67633 24714 67699 24717
rect 69200 24714 70000 24744
rect 67633 24712 70000 24714
rect 67633 24656 67638 24712
rect 67694 24656 70000 24712
rect 67633 24654 70000 24656
rect 23381 24651 23447 24652
rect 67633 24651 67699 24654
rect 69200 24624 70000 24654
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 65650 24512 65966 24513
rect 65650 24448 65656 24512
rect 65720 24448 65736 24512
rect 65800 24448 65816 24512
rect 65880 24448 65896 24512
rect 65960 24448 65966 24512
rect 65650 24447 65966 24448
rect 13077 24442 13143 24445
rect 16757 24442 16823 24445
rect 13077 24440 16823 24442
rect 13077 24384 13082 24440
rect 13138 24384 16762 24440
rect 16818 24384 16823 24440
rect 13077 24382 16823 24384
rect 13077 24379 13143 24382
rect 16757 24379 16823 24382
rect 19570 23968 19886 23969
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 50290 23968 50606 23969
rect 50290 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50606 23968
rect 50290 23903 50606 23904
rect 4337 23898 4403 23901
rect 8569 23898 8635 23901
rect 4337 23896 8635 23898
rect 4337 23840 4342 23896
rect 4398 23840 8574 23896
rect 8630 23840 8635 23896
rect 4337 23838 8635 23840
rect 4337 23835 4403 23838
rect 8569 23835 8635 23838
rect 4889 23762 4955 23765
rect 8477 23762 8543 23765
rect 4889 23760 8543 23762
rect 4889 23704 4894 23760
rect 4950 23704 8482 23760
rect 8538 23704 8543 23760
rect 4889 23702 8543 23704
rect 4889 23699 4955 23702
rect 8477 23699 8543 23702
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 65650 23424 65966 23425
rect 65650 23360 65656 23424
rect 65720 23360 65736 23424
rect 65800 23360 65816 23424
rect 65880 23360 65896 23424
rect 65960 23360 65966 23424
rect 65650 23359 65966 23360
rect 0 23128 800 23248
rect 67541 23218 67607 23221
rect 69200 23218 70000 23248
rect 67541 23216 70000 23218
rect 67541 23160 67546 23216
rect 67602 23160 70000 23216
rect 67541 23158 70000 23160
rect 67541 23155 67607 23158
rect 69200 23128 70000 23158
rect 25037 23082 25103 23085
rect 27613 23082 27679 23085
rect 25037 23080 27679 23082
rect 25037 23024 25042 23080
rect 25098 23024 27618 23080
rect 27674 23024 27679 23080
rect 25037 23022 27679 23024
rect 25037 23019 25103 23022
rect 27613 23019 27679 23022
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 50290 22880 50606 22881
rect 50290 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50606 22880
rect 50290 22815 50606 22816
rect 25773 22810 25839 22813
rect 28901 22810 28967 22813
rect 25773 22808 28967 22810
rect 25773 22752 25778 22808
rect 25834 22752 28906 22808
rect 28962 22752 28967 22808
rect 25773 22750 28967 22752
rect 25773 22747 25839 22750
rect 28901 22747 28967 22750
rect 2497 22674 2563 22677
rect 5901 22674 5967 22677
rect 2497 22672 5967 22674
rect 2497 22616 2502 22672
rect 2558 22616 5906 22672
rect 5962 22616 5967 22672
rect 2497 22614 5967 22616
rect 2497 22611 2563 22614
rect 5901 22611 5967 22614
rect 29545 22674 29611 22677
rect 33501 22674 33567 22677
rect 29545 22672 33567 22674
rect 29545 22616 29550 22672
rect 29606 22616 33506 22672
rect 33562 22616 33567 22672
rect 29545 22614 33567 22616
rect 29545 22611 29611 22614
rect 33501 22611 33567 22614
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 65650 22336 65966 22337
rect 65650 22272 65656 22336
rect 65720 22272 65736 22336
rect 65800 22272 65816 22336
rect 65880 22272 65896 22336
rect 65960 22272 65966 22336
rect 65650 22271 65966 22272
rect 23565 22268 23631 22269
rect 23565 22264 23612 22268
rect 23676 22266 23682 22268
rect 23565 22208 23570 22264
rect 23565 22204 23612 22208
rect 23676 22206 23722 22266
rect 23676 22204 23682 22206
rect 23565 22203 23631 22204
rect 18137 21994 18203 21997
rect 24393 21994 24459 21997
rect 18137 21992 24459 21994
rect 18137 21936 18142 21992
rect 18198 21936 24398 21992
rect 24454 21936 24459 21992
rect 18137 21934 24459 21936
rect 18137 21931 18203 21934
rect 24393 21931 24459 21934
rect 22921 21858 22987 21861
rect 24485 21858 24551 21861
rect 22921 21856 24551 21858
rect 22921 21800 22926 21856
rect 22982 21800 24490 21856
rect 24546 21800 24551 21856
rect 22921 21798 24551 21800
rect 22921 21795 22987 21798
rect 24485 21795 24551 21798
rect 19570 21792 19886 21793
rect 0 21632 800 21752
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 19570 21727 19886 21728
rect 50290 21792 50606 21793
rect 50290 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50606 21792
rect 50290 21727 50606 21728
rect 68093 21722 68159 21725
rect 69200 21722 70000 21752
rect 68093 21720 70000 21722
rect 68093 21664 68098 21720
rect 68154 21664 70000 21720
rect 68093 21662 70000 21664
rect 68093 21659 68159 21662
rect 69200 21632 70000 21662
rect 27889 21586 27955 21589
rect 28993 21586 29059 21589
rect 30281 21586 30347 21589
rect 27889 21584 30347 21586
rect 27889 21528 27894 21584
rect 27950 21528 28998 21584
rect 29054 21528 30286 21584
rect 30342 21528 30347 21584
rect 27889 21526 30347 21528
rect 27889 21523 27955 21526
rect 28993 21523 29059 21526
rect 30281 21523 30347 21526
rect 9673 21450 9739 21453
rect 11697 21450 11763 21453
rect 12893 21450 12959 21453
rect 9673 21448 12959 21450
rect 9673 21392 9678 21448
rect 9734 21392 11702 21448
rect 11758 21392 12898 21448
rect 12954 21392 12959 21448
rect 9673 21390 12959 21392
rect 9673 21387 9739 21390
rect 11697 21387 11763 21390
rect 12893 21387 12959 21390
rect 22001 21450 22067 21453
rect 35709 21450 35775 21453
rect 22001 21448 35775 21450
rect 22001 21392 22006 21448
rect 22062 21392 35714 21448
rect 35770 21392 35775 21448
rect 22001 21390 35775 21392
rect 22001 21387 22067 21390
rect 35709 21387 35775 21390
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 65650 21248 65966 21249
rect 65650 21184 65656 21248
rect 65720 21184 65736 21248
rect 65800 21184 65816 21248
rect 65880 21184 65896 21248
rect 65960 21184 65966 21248
rect 65650 21183 65966 21184
rect 6545 21178 6611 21181
rect 8753 21178 8819 21181
rect 6545 21176 8819 21178
rect 6545 21120 6550 21176
rect 6606 21120 8758 21176
rect 8814 21120 8819 21176
rect 6545 21118 8819 21120
rect 6545 21115 6611 21118
rect 8753 21115 8819 21118
rect 16849 21178 16915 21181
rect 17217 21178 17283 21181
rect 18873 21178 18939 21181
rect 16849 21176 18939 21178
rect 16849 21120 16854 21176
rect 16910 21120 17222 21176
rect 17278 21120 18878 21176
rect 18934 21120 18939 21176
rect 16849 21118 18939 21120
rect 16849 21115 16915 21118
rect 17217 21115 17283 21118
rect 18873 21115 18939 21118
rect 23381 21178 23447 21181
rect 27337 21178 27403 21181
rect 23381 21176 27403 21178
rect 23381 21120 23386 21176
rect 23442 21120 27342 21176
rect 27398 21120 27403 21176
rect 23381 21118 27403 21120
rect 23381 21115 23447 21118
rect 27337 21115 27403 21118
rect 8109 21042 8175 21045
rect 24301 21042 24367 21045
rect 8109 21040 24367 21042
rect 8109 20984 8114 21040
rect 8170 20984 24306 21040
rect 24362 20984 24367 21040
rect 8109 20982 24367 20984
rect 8109 20979 8175 20982
rect 24301 20979 24367 20982
rect 20897 20906 20963 20909
rect 32765 20906 32831 20909
rect 20897 20904 32831 20906
rect 20897 20848 20902 20904
rect 20958 20848 32770 20904
rect 32826 20848 32831 20904
rect 20897 20846 32831 20848
rect 20897 20843 20963 20846
rect 32765 20843 32831 20846
rect 24025 20770 24091 20773
rect 24158 20770 24164 20772
rect 24025 20768 24164 20770
rect 24025 20712 24030 20768
rect 24086 20712 24164 20768
rect 24025 20710 24164 20712
rect 24025 20707 24091 20710
rect 24158 20708 24164 20710
rect 24228 20708 24234 20772
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 50290 20704 50606 20705
rect 50290 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50606 20704
rect 50290 20639 50606 20640
rect 20529 20634 20595 20637
rect 29085 20634 29151 20637
rect 30925 20634 30991 20637
rect 20529 20632 30991 20634
rect 20529 20576 20534 20632
rect 20590 20576 29090 20632
rect 29146 20576 30930 20632
rect 30986 20576 30991 20632
rect 20529 20574 30991 20576
rect 20529 20571 20595 20574
rect 29085 20571 29151 20574
rect 30925 20571 30991 20574
rect 32305 20634 32371 20637
rect 36353 20634 36419 20637
rect 32305 20632 36419 20634
rect 32305 20576 32310 20632
rect 32366 20576 36358 20632
rect 36414 20576 36419 20632
rect 32305 20574 36419 20576
rect 32305 20571 32371 20574
rect 36353 20571 36419 20574
rect 5533 20498 5599 20501
rect 24669 20498 24735 20501
rect 25313 20498 25379 20501
rect 5533 20496 25379 20498
rect 5533 20440 5538 20496
rect 5594 20440 24674 20496
rect 24730 20440 25318 20496
rect 25374 20440 25379 20496
rect 5533 20438 25379 20440
rect 5533 20435 5599 20438
rect 24669 20435 24735 20438
rect 25313 20435 25379 20438
rect 31661 20498 31727 20501
rect 38377 20498 38443 20501
rect 31661 20496 38443 20498
rect 31661 20440 31666 20496
rect 31722 20440 38382 20496
rect 38438 20440 38443 20496
rect 31661 20438 38443 20440
rect 31661 20435 31727 20438
rect 38377 20435 38443 20438
rect 15745 20362 15811 20365
rect 22737 20362 22803 20365
rect 15745 20360 22803 20362
rect 15745 20304 15750 20360
rect 15806 20304 22742 20360
rect 22798 20304 22803 20360
rect 15745 20302 22803 20304
rect 15745 20299 15811 20302
rect 22737 20299 22803 20302
rect 0 20136 800 20256
rect 67633 20226 67699 20229
rect 69200 20226 70000 20256
rect 67633 20224 70000 20226
rect 67633 20168 67638 20224
rect 67694 20168 70000 20224
rect 67633 20166 70000 20168
rect 67633 20163 67699 20166
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 65650 20160 65966 20161
rect 65650 20096 65656 20160
rect 65720 20096 65736 20160
rect 65800 20096 65816 20160
rect 65880 20096 65896 20160
rect 65960 20096 65966 20160
rect 69200 20136 70000 20166
rect 65650 20095 65966 20096
rect 28809 19682 28875 19685
rect 34881 19682 34947 19685
rect 28809 19680 34947 19682
rect 28809 19624 28814 19680
rect 28870 19624 34886 19680
rect 34942 19624 34947 19680
rect 28809 19622 34947 19624
rect 28809 19619 28875 19622
rect 34881 19619 34947 19622
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 50290 19616 50606 19617
rect 50290 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50606 19616
rect 50290 19551 50606 19552
rect 24485 19546 24551 19549
rect 37365 19546 37431 19549
rect 24485 19544 37431 19546
rect 24485 19488 24490 19544
rect 24546 19488 37370 19544
rect 37426 19488 37431 19544
rect 24485 19486 37431 19488
rect 24485 19483 24551 19486
rect 37365 19483 37431 19486
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 65650 19072 65966 19073
rect 65650 19008 65656 19072
rect 65720 19008 65736 19072
rect 65800 19008 65816 19072
rect 65880 19008 65896 19072
rect 65960 19008 65966 19072
rect 65650 19007 65966 19008
rect 0 18640 800 18760
rect 68093 18730 68159 18733
rect 69200 18730 70000 18760
rect 68093 18728 70000 18730
rect 68093 18672 68098 18728
rect 68154 18672 70000 18728
rect 68093 18670 70000 18672
rect 68093 18667 68159 18670
rect 69200 18640 70000 18670
rect 19570 18528 19886 18529
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 50290 18528 50606 18529
rect 50290 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50606 18528
rect 50290 18463 50606 18464
rect 15193 18458 15259 18461
rect 16205 18458 16271 18461
rect 15193 18456 16271 18458
rect 15193 18400 15198 18456
rect 15254 18400 16210 18456
rect 16266 18400 16271 18456
rect 15193 18398 16271 18400
rect 15193 18395 15259 18398
rect 16205 18395 16271 18398
rect 16113 18322 16179 18325
rect 18781 18322 18847 18325
rect 16113 18320 18847 18322
rect 16113 18264 16118 18320
rect 16174 18264 18786 18320
rect 18842 18264 18847 18320
rect 16113 18262 18847 18264
rect 16113 18259 16179 18262
rect 18781 18259 18847 18262
rect 11973 18186 12039 18189
rect 18689 18186 18755 18189
rect 22001 18188 22067 18189
rect 21950 18186 21956 18188
rect 11973 18184 18755 18186
rect 11973 18128 11978 18184
rect 12034 18128 18694 18184
rect 18750 18128 18755 18184
rect 11973 18126 18755 18128
rect 21910 18126 21956 18186
rect 22020 18184 22067 18188
rect 22062 18128 22067 18184
rect 11973 18123 12039 18126
rect 18689 18123 18755 18126
rect 21950 18124 21956 18126
rect 22020 18124 22067 18128
rect 22001 18123 22067 18124
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 65650 17984 65966 17985
rect 65650 17920 65656 17984
rect 65720 17920 65736 17984
rect 65800 17920 65816 17984
rect 65880 17920 65896 17984
rect 65960 17920 65966 17984
rect 65650 17919 65966 17920
rect 15469 17642 15535 17645
rect 16389 17642 16455 17645
rect 15469 17640 16455 17642
rect 15469 17584 15474 17640
rect 15530 17584 16394 17640
rect 16450 17584 16455 17640
rect 15469 17582 16455 17584
rect 15469 17579 15535 17582
rect 16389 17579 16455 17582
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 50290 17440 50606 17441
rect 50290 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50606 17440
rect 50290 17375 50606 17376
rect 0 17144 800 17264
rect 68093 17234 68159 17237
rect 69200 17234 70000 17264
rect 68093 17232 70000 17234
rect 68093 17176 68098 17232
rect 68154 17176 70000 17232
rect 68093 17174 70000 17176
rect 68093 17171 68159 17174
rect 69200 17144 70000 17174
rect 9581 17098 9647 17101
rect 16665 17098 16731 17101
rect 17217 17098 17283 17101
rect 9581 17096 17283 17098
rect 9581 17040 9586 17096
rect 9642 17040 16670 17096
rect 16726 17040 17222 17096
rect 17278 17040 17283 17096
rect 9581 17038 17283 17040
rect 9581 17035 9647 17038
rect 16665 17035 16731 17038
rect 17217 17035 17283 17038
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 65650 16896 65966 16897
rect 65650 16832 65656 16896
rect 65720 16832 65736 16896
rect 65800 16832 65816 16896
rect 65880 16832 65896 16896
rect 65960 16832 65966 16896
rect 65650 16831 65966 16832
rect 11421 16554 11487 16557
rect 12617 16554 12683 16557
rect 18321 16554 18387 16557
rect 19609 16554 19675 16557
rect 11421 16552 19675 16554
rect 11421 16496 11426 16552
rect 11482 16496 12622 16552
rect 12678 16496 18326 16552
rect 18382 16496 19614 16552
rect 19670 16496 19675 16552
rect 11421 16494 19675 16496
rect 11421 16491 11487 16494
rect 12617 16491 12683 16494
rect 18321 16491 18387 16494
rect 19609 16491 19675 16494
rect 25037 16554 25103 16557
rect 30005 16554 30071 16557
rect 25037 16552 30071 16554
rect 25037 16496 25042 16552
rect 25098 16496 30010 16552
rect 30066 16496 30071 16552
rect 25037 16494 30071 16496
rect 25037 16491 25103 16494
rect 30005 16491 30071 16494
rect 27153 16418 27219 16421
rect 29453 16418 29519 16421
rect 36077 16418 36143 16421
rect 27153 16416 36143 16418
rect 27153 16360 27158 16416
rect 27214 16360 29458 16416
rect 29514 16360 36082 16416
rect 36138 16360 36143 16416
rect 27153 16358 36143 16360
rect 27153 16355 27219 16358
rect 29453 16355 29519 16358
rect 36077 16355 36143 16358
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 50290 16352 50606 16353
rect 50290 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50606 16352
rect 50290 16287 50606 16288
rect 17677 16146 17743 16149
rect 22553 16146 22619 16149
rect 17677 16144 22619 16146
rect 17677 16088 17682 16144
rect 17738 16088 22558 16144
rect 22614 16088 22619 16144
rect 17677 16086 22619 16088
rect 17677 16083 17743 16086
rect 22553 16083 22619 16086
rect 25865 16146 25931 16149
rect 27245 16146 27311 16149
rect 35617 16146 35683 16149
rect 25865 16144 35683 16146
rect 25865 16088 25870 16144
rect 25926 16088 27250 16144
rect 27306 16088 35622 16144
rect 35678 16088 35683 16144
rect 25865 16086 35683 16088
rect 25865 16083 25931 16086
rect 27245 16083 27311 16086
rect 35617 16083 35683 16086
rect 25957 16010 26023 16013
rect 31661 16010 31727 16013
rect 25957 16008 31727 16010
rect 25957 15952 25962 16008
rect 26018 15952 31666 16008
rect 31722 15952 31727 16008
rect 25957 15950 31727 15952
rect 25957 15947 26023 15950
rect 31661 15947 31727 15950
rect 4210 15808 4526 15809
rect 0 15648 800 15768
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 65650 15808 65966 15809
rect 65650 15744 65656 15808
rect 65720 15744 65736 15808
rect 65800 15744 65816 15808
rect 65880 15744 65896 15808
rect 65960 15744 65966 15808
rect 65650 15743 65966 15744
rect 67633 15738 67699 15741
rect 69200 15738 70000 15768
rect 67633 15736 70000 15738
rect 67633 15680 67638 15736
rect 67694 15680 70000 15736
rect 67633 15678 70000 15680
rect 67633 15675 67699 15678
rect 69200 15648 70000 15678
rect 11881 15602 11947 15605
rect 17217 15602 17283 15605
rect 11881 15600 17283 15602
rect 11881 15544 11886 15600
rect 11942 15544 17222 15600
rect 17278 15544 17283 15600
rect 11881 15542 17283 15544
rect 11881 15539 11947 15542
rect 17217 15539 17283 15542
rect 10593 15466 10659 15469
rect 16849 15466 16915 15469
rect 10593 15464 16915 15466
rect 10593 15408 10598 15464
rect 10654 15408 16854 15464
rect 16910 15408 16915 15464
rect 10593 15406 16915 15408
rect 10593 15403 10659 15406
rect 16849 15403 16915 15406
rect 24669 15330 24735 15333
rect 29085 15330 29151 15333
rect 24669 15328 29151 15330
rect 24669 15272 24674 15328
rect 24730 15272 29090 15328
rect 29146 15272 29151 15328
rect 24669 15270 29151 15272
rect 24669 15267 24735 15270
rect 29085 15267 29151 15270
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 50290 15264 50606 15265
rect 50290 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50606 15264
rect 50290 15199 50606 15200
rect 14181 15194 14247 15197
rect 19333 15194 19399 15197
rect 14181 15192 19399 15194
rect 14181 15136 14186 15192
rect 14242 15136 19338 15192
rect 19394 15136 19399 15192
rect 14181 15134 19399 15136
rect 14181 15131 14247 15134
rect 19333 15131 19399 15134
rect 18413 15058 18479 15061
rect 23565 15058 23631 15061
rect 24393 15058 24459 15061
rect 18413 15056 24459 15058
rect 18413 15000 18418 15056
rect 18474 15000 23570 15056
rect 23626 15000 24398 15056
rect 24454 15000 24459 15056
rect 18413 14998 24459 15000
rect 18413 14995 18479 14998
rect 23565 14995 23631 14998
rect 24393 14995 24459 14998
rect 28625 15058 28691 15061
rect 31017 15058 31083 15061
rect 28625 15056 31083 15058
rect 28625 15000 28630 15056
rect 28686 15000 31022 15056
rect 31078 15000 31083 15056
rect 28625 14998 31083 15000
rect 28625 14995 28691 14998
rect 31017 14995 31083 14998
rect 5441 14922 5507 14925
rect 14641 14922 14707 14925
rect 5441 14920 14707 14922
rect 5441 14864 5446 14920
rect 5502 14864 14646 14920
rect 14702 14864 14707 14920
rect 5441 14862 14707 14864
rect 5441 14859 5507 14862
rect 14641 14859 14707 14862
rect 24209 14922 24275 14925
rect 26233 14922 26299 14925
rect 24209 14920 26299 14922
rect 24209 14864 24214 14920
rect 24270 14864 26238 14920
rect 26294 14864 26299 14920
rect 24209 14862 26299 14864
rect 24209 14859 24275 14862
rect 26233 14859 26299 14862
rect 30649 14922 30715 14925
rect 32673 14922 32739 14925
rect 30649 14920 32739 14922
rect 30649 14864 30654 14920
rect 30710 14864 32678 14920
rect 32734 14864 32739 14920
rect 30649 14862 32739 14864
rect 30649 14859 30715 14862
rect 32673 14859 32739 14862
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 65650 14720 65966 14721
rect 65650 14656 65656 14720
rect 65720 14656 65736 14720
rect 65800 14656 65816 14720
rect 65880 14656 65896 14720
rect 65960 14656 65966 14720
rect 65650 14655 65966 14656
rect 17401 14514 17467 14517
rect 20437 14514 20503 14517
rect 17401 14512 20503 14514
rect 17401 14456 17406 14512
rect 17462 14456 20442 14512
rect 20498 14456 20503 14512
rect 17401 14454 20503 14456
rect 17401 14451 17467 14454
rect 20437 14451 20503 14454
rect 25129 14378 25195 14381
rect 32857 14378 32923 14381
rect 34605 14378 34671 14381
rect 25129 14376 34671 14378
rect 25129 14320 25134 14376
rect 25190 14320 32862 14376
rect 32918 14320 34610 14376
rect 34666 14320 34671 14376
rect 25129 14318 34671 14320
rect 25129 14315 25195 14318
rect 32857 14315 32923 14318
rect 34605 14315 34671 14318
rect 0 14152 800 14272
rect 29269 14242 29335 14245
rect 37089 14242 37155 14245
rect 29269 14240 37155 14242
rect 29269 14184 29274 14240
rect 29330 14184 37094 14240
rect 37150 14184 37155 14240
rect 29269 14182 37155 14184
rect 29269 14179 29335 14182
rect 37089 14179 37155 14182
rect 68093 14242 68159 14245
rect 69200 14242 70000 14272
rect 68093 14240 70000 14242
rect 68093 14184 68098 14240
rect 68154 14184 70000 14240
rect 68093 14182 70000 14184
rect 68093 14179 68159 14182
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 50290 14176 50606 14177
rect 50290 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50606 14176
rect 69200 14152 70000 14182
rect 50290 14111 50606 14112
rect 10409 14106 10475 14109
rect 17033 14106 17099 14109
rect 10409 14104 17099 14106
rect 10409 14048 10414 14104
rect 10470 14048 17038 14104
rect 17094 14048 17099 14104
rect 10409 14046 17099 14048
rect 10409 14043 10475 14046
rect 17033 14043 17099 14046
rect 35525 14108 35591 14109
rect 35525 14104 35572 14108
rect 35636 14106 35642 14108
rect 35525 14048 35530 14104
rect 35525 14044 35572 14048
rect 35636 14046 35682 14106
rect 35636 14044 35642 14046
rect 35525 14043 35591 14044
rect 7741 13970 7807 13973
rect 14733 13970 14799 13973
rect 20253 13970 20319 13973
rect 7741 13968 14799 13970
rect 7741 13912 7746 13968
rect 7802 13912 14738 13968
rect 14794 13912 14799 13968
rect 7741 13910 14799 13912
rect 7741 13907 7807 13910
rect 14733 13907 14799 13910
rect 18830 13968 20319 13970
rect 18830 13912 20258 13968
rect 20314 13912 20319 13968
rect 18830 13910 20319 13912
rect 8017 13834 8083 13837
rect 18830 13834 18890 13910
rect 20253 13907 20319 13910
rect 8017 13832 18890 13834
rect 8017 13776 8022 13832
rect 8078 13776 18890 13832
rect 8017 13774 18890 13776
rect 8017 13771 8083 13774
rect 19374 13772 19380 13836
rect 19444 13834 19450 13836
rect 19885 13834 19951 13837
rect 19444 13832 19951 13834
rect 19444 13776 19890 13832
rect 19946 13776 19951 13832
rect 19444 13774 19951 13776
rect 19444 13772 19450 13774
rect 19885 13771 19951 13774
rect 12893 13698 12959 13701
rect 16573 13698 16639 13701
rect 12893 13696 16639 13698
rect 12893 13640 12898 13696
rect 12954 13640 16578 13696
rect 16634 13640 16639 13696
rect 12893 13638 16639 13640
rect 12893 13635 12959 13638
rect 16573 13635 16639 13638
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 65650 13632 65966 13633
rect 65650 13568 65656 13632
rect 65720 13568 65736 13632
rect 65800 13568 65816 13632
rect 65880 13568 65896 13632
rect 65960 13568 65966 13632
rect 65650 13567 65966 13568
rect 19701 13562 19767 13565
rect 28717 13562 28783 13565
rect 19701 13560 28783 13562
rect 19701 13504 19706 13560
rect 19762 13504 28722 13560
rect 28778 13504 28783 13560
rect 19701 13502 28783 13504
rect 19701 13499 19767 13502
rect 28717 13499 28783 13502
rect 12893 13426 12959 13429
rect 16021 13426 16087 13429
rect 12893 13424 16087 13426
rect 12893 13368 12898 13424
rect 12954 13368 16026 13424
rect 16082 13368 16087 13424
rect 12893 13366 16087 13368
rect 12893 13363 12959 13366
rect 16021 13363 16087 13366
rect 16481 13426 16547 13429
rect 31385 13426 31451 13429
rect 16481 13424 31451 13426
rect 16481 13368 16486 13424
rect 16542 13368 31390 13424
rect 31446 13368 31451 13424
rect 16481 13366 31451 13368
rect 16481 13363 16547 13366
rect 31385 13363 31451 13366
rect 11237 13290 11303 13293
rect 14641 13290 14707 13293
rect 19057 13290 19123 13293
rect 11237 13288 19123 13290
rect 11237 13232 11242 13288
rect 11298 13232 14646 13288
rect 14702 13232 19062 13288
rect 19118 13232 19123 13288
rect 11237 13230 19123 13232
rect 11237 13227 11303 13230
rect 14641 13227 14707 13230
rect 19057 13227 19123 13230
rect 23749 13290 23815 13293
rect 24761 13290 24827 13293
rect 27061 13290 27127 13293
rect 23749 13288 27127 13290
rect 23749 13232 23754 13288
rect 23810 13232 24766 13288
rect 24822 13232 27066 13288
rect 27122 13232 27127 13288
rect 23749 13230 27127 13232
rect 23749 13227 23815 13230
rect 24761 13227 24827 13230
rect 27061 13227 27127 13230
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 50290 13088 50606 13089
rect 50290 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50606 13088
rect 50290 13023 50606 13024
rect 20805 13018 20871 13021
rect 23473 13018 23539 13021
rect 20805 13016 23539 13018
rect 20805 12960 20810 13016
rect 20866 12960 23478 13016
rect 23534 12960 23539 13016
rect 20805 12958 23539 12960
rect 20805 12955 20871 12958
rect 23473 12955 23539 12958
rect 25405 13018 25471 13021
rect 26141 13018 26207 13021
rect 25405 13016 26207 13018
rect 25405 12960 25410 13016
rect 25466 12960 26146 13016
rect 26202 12960 26207 13016
rect 25405 12958 26207 12960
rect 25405 12955 25471 12958
rect 26141 12955 26207 12958
rect 12525 12882 12591 12885
rect 24669 12882 24735 12885
rect 26325 12882 26391 12885
rect 12525 12880 26391 12882
rect 12525 12824 12530 12880
rect 12586 12824 24674 12880
rect 24730 12824 26330 12880
rect 26386 12824 26391 12880
rect 12525 12822 26391 12824
rect 12525 12819 12591 12822
rect 24669 12819 24735 12822
rect 26325 12819 26391 12822
rect 0 12656 800 12776
rect 4613 12746 4679 12749
rect 22369 12746 22435 12749
rect 4613 12744 22435 12746
rect 4613 12688 4618 12744
rect 4674 12688 22374 12744
rect 22430 12688 22435 12744
rect 4613 12686 22435 12688
rect 4613 12683 4679 12686
rect 22369 12683 22435 12686
rect 23473 12746 23539 12749
rect 26601 12746 26667 12749
rect 23473 12744 26667 12746
rect 23473 12688 23478 12744
rect 23534 12688 26606 12744
rect 26662 12688 26667 12744
rect 23473 12686 26667 12688
rect 23473 12683 23539 12686
rect 26601 12683 26667 12686
rect 67633 12746 67699 12749
rect 69200 12746 70000 12776
rect 67633 12744 70000 12746
rect 67633 12688 67638 12744
rect 67694 12688 70000 12744
rect 67633 12686 70000 12688
rect 67633 12683 67699 12686
rect 69200 12656 70000 12686
rect 17401 12610 17467 12613
rect 31293 12610 31359 12613
rect 17401 12608 31359 12610
rect 17401 12552 17406 12608
rect 17462 12552 31298 12608
rect 31354 12552 31359 12608
rect 17401 12550 31359 12552
rect 17401 12547 17467 12550
rect 31293 12547 31359 12550
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 65650 12544 65966 12545
rect 65650 12480 65656 12544
rect 65720 12480 65736 12544
rect 65800 12480 65816 12544
rect 65880 12480 65896 12544
rect 65960 12480 65966 12544
rect 65650 12479 65966 12480
rect 25313 12474 25379 12477
rect 29085 12474 29151 12477
rect 25313 12472 29151 12474
rect 25313 12416 25318 12472
rect 25374 12416 29090 12472
rect 29146 12416 29151 12472
rect 25313 12414 29151 12416
rect 25313 12411 25379 12414
rect 29085 12411 29151 12414
rect 16113 12338 16179 12341
rect 25405 12338 25471 12341
rect 16113 12336 25471 12338
rect 16113 12280 16118 12336
rect 16174 12280 25410 12336
rect 25466 12280 25471 12336
rect 16113 12278 25471 12280
rect 16113 12275 16179 12278
rect 25405 12275 25471 12278
rect 3417 12202 3483 12205
rect 12801 12202 12867 12205
rect 3417 12200 12867 12202
rect 3417 12144 3422 12200
rect 3478 12144 12806 12200
rect 12862 12144 12867 12200
rect 3417 12142 12867 12144
rect 3417 12139 3483 12142
rect 12801 12139 12867 12142
rect 14917 12202 14983 12205
rect 17861 12202 17927 12205
rect 19149 12202 19215 12205
rect 14917 12200 19215 12202
rect 14917 12144 14922 12200
rect 14978 12144 17866 12200
rect 17922 12144 19154 12200
rect 19210 12144 19215 12200
rect 14917 12142 19215 12144
rect 14917 12139 14983 12142
rect 17861 12139 17927 12142
rect 19149 12139 19215 12142
rect 21909 12202 21975 12205
rect 32397 12202 32463 12205
rect 21909 12200 32463 12202
rect 21909 12144 21914 12200
rect 21970 12144 32402 12200
rect 32458 12144 32463 12200
rect 21909 12142 32463 12144
rect 21909 12139 21975 12142
rect 32397 12139 32463 12142
rect 16757 12066 16823 12069
rect 17861 12068 17927 12069
rect 17861 12066 17908 12068
rect 16757 12064 17908 12066
rect 16757 12008 16762 12064
rect 16818 12008 17866 12064
rect 16757 12006 17908 12008
rect 16757 12003 16823 12006
rect 17861 12004 17908 12006
rect 17972 12004 17978 12068
rect 22921 12066 22987 12069
rect 25129 12066 25195 12069
rect 26233 12066 26299 12069
rect 22921 12064 26299 12066
rect 22921 12008 22926 12064
rect 22982 12008 25134 12064
rect 25190 12008 26238 12064
rect 26294 12008 26299 12064
rect 22921 12006 26299 12008
rect 17861 12003 17927 12004
rect 22921 12003 22987 12006
rect 25129 12003 25195 12006
rect 26233 12003 26299 12006
rect 29821 12066 29887 12069
rect 31109 12066 31175 12069
rect 29821 12064 31175 12066
rect 29821 12008 29826 12064
rect 29882 12008 31114 12064
rect 31170 12008 31175 12064
rect 29821 12006 31175 12008
rect 29821 12003 29887 12006
rect 31109 12003 31175 12006
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 50290 12000 50606 12001
rect 50290 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50606 12000
rect 50290 11935 50606 11936
rect 15101 11930 15167 11933
rect 18505 11930 18571 11933
rect 24761 11930 24827 11933
rect 35617 11932 35683 11933
rect 15101 11928 18571 11930
rect 15101 11872 15106 11928
rect 15162 11872 18510 11928
rect 18566 11872 18571 11928
rect 15101 11870 18571 11872
rect 15101 11867 15167 11870
rect 18505 11867 18571 11870
rect 24718 11928 24827 11930
rect 24718 11872 24766 11928
rect 24822 11872 24827 11928
rect 24718 11867 24827 11872
rect 35566 11868 35572 11932
rect 35636 11930 35683 11932
rect 35636 11928 35728 11930
rect 35678 11872 35728 11928
rect 35636 11870 35728 11872
rect 35636 11868 35683 11870
rect 35617 11867 35683 11868
rect 15469 11794 15535 11797
rect 23289 11794 23355 11797
rect 15469 11792 23355 11794
rect 15469 11736 15474 11792
rect 15530 11736 23294 11792
rect 23350 11736 23355 11792
rect 15469 11734 23355 11736
rect 15469 11731 15535 11734
rect 23289 11731 23355 11734
rect 21817 11658 21883 11661
rect 24117 11658 24183 11661
rect 24718 11658 24778 11867
rect 25129 11794 25195 11797
rect 26233 11794 26299 11797
rect 25129 11792 26299 11794
rect 25129 11736 25134 11792
rect 25190 11736 26238 11792
rect 26294 11736 26299 11792
rect 25129 11734 26299 11736
rect 25129 11731 25195 11734
rect 26233 11731 26299 11734
rect 21817 11656 22110 11658
rect 21817 11600 21822 11656
rect 21878 11600 22110 11656
rect 21817 11598 22110 11600
rect 21817 11595 21883 11598
rect 11053 11524 11119 11525
rect 11053 11522 11100 11524
rect 11008 11520 11100 11522
rect 11008 11464 11058 11520
rect 11008 11462 11100 11464
rect 11053 11460 11100 11462
rect 11164 11460 11170 11524
rect 22050 11522 22110 11598
rect 24117 11656 24778 11658
rect 24117 11600 24122 11656
rect 24178 11600 24778 11656
rect 24117 11598 24778 11600
rect 24117 11595 24183 11598
rect 28073 11522 28139 11525
rect 22050 11520 28139 11522
rect 22050 11464 28078 11520
rect 28134 11464 28139 11520
rect 22050 11462 28139 11464
rect 11053 11459 11119 11460
rect 28073 11459 28139 11462
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 65650 11456 65966 11457
rect 65650 11392 65656 11456
rect 65720 11392 65736 11456
rect 65800 11392 65816 11456
rect 65880 11392 65896 11456
rect 65960 11392 65966 11456
rect 65650 11391 65966 11392
rect 17309 11386 17375 11389
rect 23606 11386 23612 11388
rect 17309 11384 23612 11386
rect 17309 11328 17314 11384
rect 17370 11328 23612 11384
rect 17309 11326 23612 11328
rect 17309 11323 17375 11326
rect 23606 11324 23612 11326
rect 23676 11324 23682 11388
rect 29821 11386 29887 11389
rect 30281 11386 30347 11389
rect 32857 11386 32923 11389
rect 29821 11384 32923 11386
rect 29821 11328 29826 11384
rect 29882 11328 30286 11384
rect 30342 11328 32862 11384
rect 32918 11328 32923 11384
rect 29821 11326 32923 11328
rect 29821 11323 29887 11326
rect 30281 11323 30347 11326
rect 32857 11323 32923 11326
rect 0 11160 800 11280
rect 16481 11250 16547 11253
rect 32857 11250 32923 11253
rect 16481 11248 32923 11250
rect 16481 11192 16486 11248
rect 16542 11192 32862 11248
rect 32918 11192 32923 11248
rect 16481 11190 32923 11192
rect 16481 11187 16547 11190
rect 32857 11187 32923 11190
rect 34973 11250 35039 11253
rect 36997 11250 37063 11253
rect 34973 11248 37063 11250
rect 34973 11192 34978 11248
rect 35034 11192 37002 11248
rect 37058 11192 37063 11248
rect 34973 11190 37063 11192
rect 34973 11187 35039 11190
rect 36997 11187 37063 11190
rect 67633 11250 67699 11253
rect 69200 11250 70000 11280
rect 67633 11248 70000 11250
rect 67633 11192 67638 11248
rect 67694 11192 70000 11248
rect 67633 11190 70000 11192
rect 67633 11187 67699 11190
rect 69200 11160 70000 11190
rect 16757 11114 16823 11117
rect 29729 11114 29795 11117
rect 16757 11112 29795 11114
rect 16757 11056 16762 11112
rect 16818 11056 29734 11112
rect 29790 11056 29795 11112
rect 16757 11054 29795 11056
rect 16757 11051 16823 11054
rect 29729 11051 29795 11054
rect 28717 10978 28783 10981
rect 36077 10978 36143 10981
rect 28717 10976 36143 10978
rect 28717 10920 28722 10976
rect 28778 10920 36082 10976
rect 36138 10920 36143 10976
rect 28717 10918 36143 10920
rect 28717 10915 28783 10918
rect 36077 10915 36143 10918
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 19570 10847 19886 10848
rect 50290 10912 50606 10913
rect 50290 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50606 10912
rect 50290 10847 50606 10848
rect 9489 10706 9555 10709
rect 10777 10706 10843 10709
rect 21950 10706 21956 10708
rect 9489 10704 21956 10706
rect 9489 10648 9494 10704
rect 9550 10648 10782 10704
rect 10838 10648 21956 10704
rect 9489 10646 21956 10648
rect 9489 10643 9555 10646
rect 10777 10643 10843 10646
rect 21950 10644 21956 10646
rect 22020 10644 22026 10708
rect 4705 10570 4771 10573
rect 9121 10570 9187 10573
rect 4705 10568 9187 10570
rect 4705 10512 4710 10568
rect 4766 10512 9126 10568
rect 9182 10512 9187 10568
rect 4705 10510 9187 10512
rect 4705 10507 4771 10510
rect 9121 10507 9187 10510
rect 18965 10570 19031 10573
rect 30833 10570 30899 10573
rect 18965 10568 30899 10570
rect 18965 10512 18970 10568
rect 19026 10512 30838 10568
rect 30894 10512 30899 10568
rect 18965 10510 30899 10512
rect 18965 10507 19031 10510
rect 30833 10507 30899 10510
rect 28073 10434 28139 10437
rect 32305 10434 32371 10437
rect 28073 10432 32371 10434
rect 28073 10376 28078 10432
rect 28134 10376 32310 10432
rect 32366 10376 32371 10432
rect 28073 10374 32371 10376
rect 28073 10371 28139 10374
rect 32305 10371 32371 10374
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 65650 10368 65966 10369
rect 65650 10304 65656 10368
rect 65720 10304 65736 10368
rect 65800 10304 65816 10368
rect 65880 10304 65896 10368
rect 65960 10304 65966 10368
rect 65650 10303 65966 10304
rect 10726 10236 10732 10300
rect 10796 10298 10802 10300
rect 20621 10298 20687 10301
rect 10796 10296 20687 10298
rect 10796 10240 20626 10296
rect 20682 10240 20687 10296
rect 10796 10238 20687 10240
rect 10796 10236 10802 10238
rect 20621 10235 20687 10238
rect 27429 10162 27495 10165
rect 31201 10162 31267 10165
rect 33317 10162 33383 10165
rect 27429 10160 33383 10162
rect 27429 10104 27434 10160
rect 27490 10104 31206 10160
rect 31262 10104 33322 10160
rect 33378 10104 33383 10160
rect 27429 10102 33383 10104
rect 27429 10099 27495 10102
rect 31201 10099 31267 10102
rect 33317 10099 33383 10102
rect 18229 10026 18295 10029
rect 28809 10026 28875 10029
rect 18229 10024 28875 10026
rect 18229 9968 18234 10024
rect 18290 9968 28814 10024
rect 28870 9968 28875 10024
rect 18229 9966 28875 9968
rect 18229 9963 18295 9966
rect 28809 9963 28875 9966
rect 6085 9890 6151 9893
rect 10041 9890 10107 9893
rect 6085 9888 10107 9890
rect 6085 9832 6090 9888
rect 6146 9832 10046 9888
rect 10102 9832 10107 9888
rect 6085 9830 10107 9832
rect 6085 9827 6151 9830
rect 10041 9827 10107 9830
rect 19570 9824 19886 9825
rect 0 9664 800 9784
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 50290 9824 50606 9825
rect 50290 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50606 9824
rect 50290 9759 50606 9760
rect 6269 9754 6335 9757
rect 8109 9754 8175 9757
rect 6269 9752 8175 9754
rect 6269 9696 6274 9752
rect 6330 9696 8114 9752
rect 8170 9696 8175 9752
rect 6269 9694 8175 9696
rect 6269 9691 6335 9694
rect 8109 9691 8175 9694
rect 32305 9754 32371 9757
rect 68093 9754 68159 9757
rect 69200 9754 70000 9784
rect 32305 9752 32506 9754
rect 32305 9696 32310 9752
rect 32366 9696 32506 9752
rect 32305 9694 32506 9696
rect 32305 9691 32371 9694
rect 17125 9618 17191 9621
rect 24158 9618 24164 9620
rect 17125 9616 24164 9618
rect 17125 9560 17130 9616
rect 17186 9560 24164 9616
rect 17125 9558 24164 9560
rect 17125 9555 17191 9558
rect 24158 9556 24164 9558
rect 24228 9556 24234 9620
rect 32446 9618 32506 9694
rect 68093 9752 70000 9754
rect 68093 9696 68098 9752
rect 68154 9696 70000 9752
rect 68093 9694 70000 9696
rect 68093 9691 68159 9694
rect 69200 9664 70000 9694
rect 33317 9618 33383 9621
rect 38377 9618 38443 9621
rect 32446 9616 38443 9618
rect 32446 9560 33322 9616
rect 33378 9560 38382 9616
rect 38438 9560 38443 9616
rect 32446 9558 38443 9560
rect 33317 9555 33383 9558
rect 38377 9555 38443 9558
rect 26141 9482 26207 9485
rect 31477 9482 31543 9485
rect 26141 9480 31543 9482
rect 26141 9424 26146 9480
rect 26202 9424 31482 9480
rect 31538 9424 31543 9480
rect 26141 9422 31543 9424
rect 26141 9419 26207 9422
rect 31477 9419 31543 9422
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 65650 9280 65966 9281
rect 65650 9216 65656 9280
rect 65720 9216 65736 9280
rect 65800 9216 65816 9280
rect 65880 9216 65896 9280
rect 65960 9216 65966 9280
rect 65650 9215 65966 9216
rect 11053 8938 11119 8941
rect 21173 8938 21239 8941
rect 11053 8936 21239 8938
rect 11053 8880 11058 8936
rect 11114 8880 21178 8936
rect 21234 8880 21239 8936
rect 11053 8878 21239 8880
rect 11053 8875 11119 8878
rect 21173 8875 21239 8878
rect 7281 8802 7347 8805
rect 7833 8802 7899 8805
rect 11145 8802 11211 8805
rect 12014 8802 12020 8804
rect 7281 8800 12020 8802
rect 7281 8744 7286 8800
rect 7342 8744 7838 8800
rect 7894 8744 11150 8800
rect 11206 8744 12020 8800
rect 7281 8742 12020 8744
rect 7281 8739 7347 8742
rect 7833 8739 7899 8742
rect 11145 8739 11211 8742
rect 12014 8740 12020 8742
rect 12084 8740 12090 8804
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 50290 8736 50606 8737
rect 50290 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50606 8736
rect 50290 8671 50606 8672
rect 36537 8530 36603 8533
rect 38009 8530 38075 8533
rect 36537 8528 38075 8530
rect 36537 8472 36542 8528
rect 36598 8472 38014 8528
rect 38070 8472 38075 8528
rect 36537 8470 38075 8472
rect 36537 8467 36603 8470
rect 38009 8467 38075 8470
rect 7925 8394 7991 8397
rect 8385 8394 8451 8397
rect 7925 8392 8451 8394
rect 7925 8336 7930 8392
rect 7986 8336 8390 8392
rect 8446 8336 8451 8392
rect 7925 8334 8451 8336
rect 7925 8331 7991 8334
rect 8385 8331 8451 8334
rect 0 8168 800 8288
rect 67541 8258 67607 8261
rect 69200 8258 70000 8288
rect 67541 8256 70000 8258
rect 67541 8200 67546 8256
rect 67602 8200 70000 8256
rect 67541 8198 70000 8200
rect 67541 8195 67607 8198
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 65650 8192 65966 8193
rect 65650 8128 65656 8192
rect 65720 8128 65736 8192
rect 65800 8128 65816 8192
rect 65880 8128 65896 8192
rect 65960 8128 65966 8192
rect 69200 8168 70000 8198
rect 65650 8127 65966 8128
rect 5717 7850 5783 7853
rect 15837 7850 15903 7853
rect 5717 7848 15903 7850
rect 5717 7792 5722 7848
rect 5778 7792 15842 7848
rect 15898 7792 15903 7848
rect 5717 7790 15903 7792
rect 5717 7787 5783 7790
rect 15837 7787 15903 7790
rect 19570 7648 19886 7649
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 50290 7648 50606 7649
rect 50290 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50606 7648
rect 50290 7583 50606 7584
rect 11697 7442 11763 7445
rect 19374 7442 19380 7444
rect 11697 7440 19380 7442
rect 11697 7384 11702 7440
rect 11758 7384 19380 7440
rect 11697 7382 19380 7384
rect 11697 7379 11763 7382
rect 19374 7380 19380 7382
rect 19444 7380 19450 7444
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 65650 7104 65966 7105
rect 65650 7040 65656 7104
rect 65720 7040 65736 7104
rect 65800 7040 65816 7104
rect 65880 7040 65896 7104
rect 65960 7040 65966 7104
rect 65650 7039 65966 7040
rect 5901 7034 5967 7037
rect 11053 7034 11119 7037
rect 5901 7032 11119 7034
rect 5901 6976 5906 7032
rect 5962 6976 11058 7032
rect 11114 6976 11119 7032
rect 5901 6974 11119 6976
rect 5901 6971 5967 6974
rect 11053 6971 11119 6974
rect 11421 6898 11487 6901
rect 11973 6898 12039 6901
rect 16849 6898 16915 6901
rect 11421 6896 16915 6898
rect 11421 6840 11426 6896
rect 11482 6840 11978 6896
rect 12034 6840 16854 6896
rect 16910 6840 16915 6896
rect 11421 6838 16915 6840
rect 11421 6835 11487 6838
rect 11973 6835 12039 6838
rect 16849 6835 16915 6838
rect 0 6672 800 6792
rect 68093 6762 68159 6765
rect 69200 6762 70000 6792
rect 68093 6760 70000 6762
rect 68093 6704 68098 6760
rect 68154 6704 70000 6760
rect 68093 6702 70000 6704
rect 68093 6699 68159 6702
rect 69200 6672 70000 6702
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 50290 6560 50606 6561
rect 50290 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50606 6560
rect 50290 6495 50606 6496
rect 9213 6218 9279 6221
rect 12617 6218 12683 6221
rect 9213 6216 12683 6218
rect 9213 6160 9218 6216
rect 9274 6160 12622 6216
rect 12678 6160 12683 6216
rect 9213 6158 12683 6160
rect 9213 6155 9279 6158
rect 12617 6155 12683 6158
rect 10869 6082 10935 6085
rect 13445 6082 13511 6085
rect 10869 6080 13511 6082
rect 10869 6024 10874 6080
rect 10930 6024 13450 6080
rect 13506 6024 13511 6080
rect 10869 6022 13511 6024
rect 10869 6019 10935 6022
rect 13445 6019 13511 6022
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 65650 6016 65966 6017
rect 65650 5952 65656 6016
rect 65720 5952 65736 6016
rect 65800 5952 65816 6016
rect 65880 5952 65896 6016
rect 65960 5952 65966 6016
rect 65650 5951 65966 5952
rect 11053 5946 11119 5949
rect 12157 5946 12223 5949
rect 11053 5944 12223 5946
rect 11053 5888 11058 5944
rect 11114 5888 12162 5944
rect 12218 5888 12223 5944
rect 11053 5886 12223 5888
rect 11053 5883 11119 5886
rect 12157 5883 12223 5886
rect 5625 5810 5691 5813
rect 15377 5810 15443 5813
rect 5625 5808 15443 5810
rect 5625 5752 5630 5808
rect 5686 5752 15382 5808
rect 15438 5752 15443 5808
rect 5625 5750 15443 5752
rect 5625 5747 5691 5750
rect 15377 5747 15443 5750
rect 14917 5538 14983 5541
rect 17401 5538 17467 5541
rect 14917 5536 17467 5538
rect 14917 5480 14922 5536
rect 14978 5480 17406 5536
rect 17462 5480 17467 5536
rect 14917 5478 17467 5480
rect 14917 5475 14983 5478
rect 17401 5475 17467 5478
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 19570 5407 19886 5408
rect 50290 5472 50606 5473
rect 50290 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50606 5472
rect 50290 5407 50606 5408
rect 12157 5402 12223 5405
rect 16205 5402 16271 5405
rect 12157 5400 16271 5402
rect 12157 5344 12162 5400
rect 12218 5344 16210 5400
rect 16266 5344 16271 5400
rect 12157 5342 16271 5344
rect 12157 5339 12223 5342
rect 16205 5339 16271 5342
rect 0 5176 800 5296
rect 68093 5266 68159 5269
rect 69200 5266 70000 5296
rect 68093 5264 70000 5266
rect 68093 5208 68098 5264
rect 68154 5208 70000 5264
rect 68093 5206 70000 5208
rect 68093 5203 68159 5206
rect 69200 5176 70000 5206
rect 3969 5130 4035 5133
rect 7281 5130 7347 5133
rect 3969 5128 7347 5130
rect 3969 5072 3974 5128
rect 4030 5072 7286 5128
rect 7342 5072 7347 5128
rect 3969 5070 7347 5072
rect 3969 5067 4035 5070
rect 7281 5067 7347 5070
rect 11697 5130 11763 5133
rect 17309 5130 17375 5133
rect 11697 5128 17375 5130
rect 11697 5072 11702 5128
rect 11758 5072 17314 5128
rect 17370 5072 17375 5128
rect 11697 5070 17375 5072
rect 11697 5067 11763 5070
rect 17309 5067 17375 5070
rect 11973 4994 12039 4997
rect 15929 4994 15995 4997
rect 11973 4992 15995 4994
rect 11973 4936 11978 4992
rect 12034 4936 15934 4992
rect 15990 4936 15995 4992
rect 11973 4934 15995 4936
rect 11973 4931 12039 4934
rect 15929 4931 15995 4934
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 65650 4928 65966 4929
rect 65650 4864 65656 4928
rect 65720 4864 65736 4928
rect 65800 4864 65816 4928
rect 65880 4864 65896 4928
rect 65960 4864 65966 4928
rect 65650 4863 65966 4864
rect 8109 4722 8175 4725
rect 11329 4722 11395 4725
rect 22829 4722 22895 4725
rect 8109 4720 22895 4722
rect 8109 4664 8114 4720
rect 8170 4664 11334 4720
rect 11390 4664 22834 4720
rect 22890 4664 22895 4720
rect 8109 4662 22895 4664
rect 8109 4659 8175 4662
rect 11329 4659 11395 4662
rect 22829 4659 22895 4662
rect 9765 4586 9831 4589
rect 9949 4586 10015 4589
rect 26693 4586 26759 4589
rect 27797 4586 27863 4589
rect 9765 4584 27863 4586
rect 9765 4528 9770 4584
rect 9826 4528 9954 4584
rect 10010 4528 26698 4584
rect 26754 4528 27802 4584
rect 27858 4528 27863 4584
rect 9765 4526 27863 4528
rect 9765 4523 9831 4526
rect 9949 4523 10015 4526
rect 26693 4523 26759 4526
rect 27797 4523 27863 4526
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 50290 4384 50606 4385
rect 50290 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50606 4384
rect 50290 4319 50606 4320
rect 4981 4178 5047 4181
rect 8937 4178 9003 4181
rect 11421 4178 11487 4181
rect 4981 4176 11487 4178
rect 4981 4120 4986 4176
rect 5042 4120 8942 4176
rect 8998 4120 11426 4176
rect 11482 4120 11487 4176
rect 4981 4118 11487 4120
rect 4981 4115 5047 4118
rect 8937 4115 9003 4118
rect 11421 4115 11487 4118
rect 7649 4042 7715 4045
rect 10317 4042 10383 4045
rect 10593 4042 10659 4045
rect 10726 4042 10732 4044
rect 7649 4040 10426 4042
rect 7649 3984 7654 4040
rect 7710 3984 10322 4040
rect 10378 3984 10426 4040
rect 7649 3982 10426 3984
rect 7649 3979 7715 3982
rect 10317 3979 10426 3982
rect 10593 4040 10732 4042
rect 10593 3984 10598 4040
rect 10654 3984 10732 4040
rect 10593 3982 10732 3984
rect 10593 3979 10659 3982
rect 10726 3980 10732 3982
rect 10796 3980 10802 4044
rect 10961 4042 11027 4045
rect 19425 4042 19491 4045
rect 20805 4042 20871 4045
rect 10961 4040 20871 4042
rect 10961 3984 10966 4040
rect 11022 3984 19430 4040
rect 19486 3984 20810 4040
rect 20866 3984 20871 4040
rect 10961 3982 20871 3984
rect 10961 3979 11027 3982
rect 19425 3979 19491 3982
rect 20805 3979 20871 3982
rect 10366 3906 10426 3979
rect 10501 3906 10567 3909
rect 10366 3904 10567 3906
rect 10366 3848 10506 3904
rect 10562 3848 10567 3904
rect 10366 3846 10567 3848
rect 10501 3843 10567 3846
rect 11329 3904 11395 3909
rect 11329 3848 11334 3904
rect 11390 3848 11395 3904
rect 11329 3843 11395 3848
rect 16297 3906 16363 3909
rect 20437 3906 20503 3909
rect 16297 3904 20503 3906
rect 16297 3848 16302 3904
rect 16358 3848 20442 3904
rect 20498 3848 20503 3904
rect 16297 3846 20503 3848
rect 16297 3843 16363 3846
rect 20437 3843 20503 3846
rect 4210 3840 4526 3841
rect 0 3680 800 3800
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 4613 3770 4679 3773
rect 11332 3770 11392 3843
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 65650 3840 65966 3841
rect 65650 3776 65656 3840
rect 65720 3776 65736 3840
rect 65800 3776 65816 3840
rect 65880 3776 65896 3840
rect 65960 3776 65966 3840
rect 65650 3775 65966 3776
rect 4613 3768 11392 3770
rect 4613 3712 4618 3768
rect 4674 3712 11392 3768
rect 4613 3710 11392 3712
rect 14089 3770 14155 3773
rect 24485 3770 24551 3773
rect 14089 3768 24551 3770
rect 14089 3712 14094 3768
rect 14150 3712 24490 3768
rect 24546 3712 24551 3768
rect 14089 3710 24551 3712
rect 4613 3707 4679 3710
rect 14089 3707 14155 3710
rect 24485 3707 24551 3710
rect 67633 3770 67699 3773
rect 69200 3770 70000 3800
rect 67633 3768 70000 3770
rect 67633 3712 67638 3768
rect 67694 3712 70000 3768
rect 67633 3710 70000 3712
rect 67633 3707 67699 3710
rect 69200 3680 70000 3710
rect 10869 3634 10935 3637
rect 12157 3634 12223 3637
rect 15101 3634 15167 3637
rect 17902 3634 17908 3636
rect 10869 3632 12223 3634
rect 10869 3576 10874 3632
rect 10930 3576 12162 3632
rect 12218 3576 12223 3632
rect 10869 3574 12223 3576
rect 10869 3571 10935 3574
rect 12157 3571 12223 3574
rect 12390 3632 17908 3634
rect 12390 3576 15106 3632
rect 15162 3576 17908 3632
rect 12390 3574 17908 3576
rect 9305 3498 9371 3501
rect 12390 3498 12450 3574
rect 15101 3571 15167 3574
rect 17902 3572 17908 3574
rect 17972 3634 17978 3636
rect 26141 3634 26207 3637
rect 17972 3632 26207 3634
rect 17972 3576 26146 3632
rect 26202 3576 26207 3632
rect 17972 3574 26207 3576
rect 17972 3572 17978 3574
rect 26141 3571 26207 3574
rect 9305 3496 12450 3498
rect 9305 3440 9310 3496
rect 9366 3440 12450 3496
rect 9305 3438 12450 3440
rect 9305 3435 9371 3438
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 50290 3296 50606 3297
rect 50290 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50606 3296
rect 50290 3231 50606 3232
rect 6453 3226 6519 3229
rect 8661 3226 8727 3229
rect 6453 3224 8727 3226
rect 6453 3168 6458 3224
rect 6514 3168 8666 3224
rect 8722 3168 8727 3224
rect 6453 3166 8727 3168
rect 6453 3163 6519 3166
rect 8661 3163 8727 3166
rect 57881 3226 57947 3229
rect 60457 3226 60523 3229
rect 57881 3224 60523 3226
rect 57881 3168 57886 3224
rect 57942 3168 60462 3224
rect 60518 3168 60523 3224
rect 57881 3166 60523 3168
rect 57881 3163 57947 3166
rect 60457 3163 60523 3166
rect 11094 3028 11100 3092
rect 11164 3090 11170 3092
rect 15653 3090 15719 3093
rect 23749 3090 23815 3093
rect 11164 3088 23815 3090
rect 11164 3032 15658 3088
rect 15714 3032 23754 3088
rect 23810 3032 23815 3088
rect 11164 3030 23815 3032
rect 11164 3028 11170 3030
rect 15653 3027 15719 3030
rect 23749 3027 23815 3030
rect 11513 2954 11579 2957
rect 14089 2954 14155 2957
rect 15193 2954 15259 2957
rect 11513 2952 15259 2954
rect 11513 2896 11518 2952
rect 11574 2896 14094 2952
rect 14150 2896 15198 2952
rect 15254 2896 15259 2952
rect 11513 2894 15259 2896
rect 11513 2891 11579 2894
rect 14089 2891 14155 2894
rect 15193 2891 15259 2894
rect 9581 2818 9647 2821
rect 11881 2818 11947 2821
rect 12065 2820 12131 2821
rect 9581 2816 11947 2818
rect 9581 2760 9586 2816
rect 9642 2760 11886 2816
rect 11942 2760 11947 2816
rect 9581 2758 11947 2760
rect 9581 2755 9647 2758
rect 11881 2755 11947 2758
rect 12014 2756 12020 2820
rect 12084 2818 12131 2820
rect 23841 2818 23907 2821
rect 12084 2816 23907 2818
rect 12126 2760 23846 2816
rect 23902 2760 23907 2816
rect 12084 2758 23907 2760
rect 12084 2756 12131 2758
rect 12065 2755 12131 2756
rect 23841 2755 23907 2758
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 65650 2752 65966 2753
rect 65650 2688 65656 2752
rect 65720 2688 65736 2752
rect 65800 2688 65816 2752
rect 65880 2688 65896 2752
rect 65960 2688 65966 2752
rect 65650 2687 65966 2688
rect 7925 2682 7991 2685
rect 18229 2682 18295 2685
rect 7925 2680 18295 2682
rect 7925 2624 7930 2680
rect 7986 2624 18234 2680
rect 18290 2624 18295 2680
rect 7925 2622 18295 2624
rect 7925 2619 7991 2622
rect 18229 2619 18295 2622
rect 10041 2410 10107 2413
rect 25589 2410 25655 2413
rect 10041 2408 25655 2410
rect 10041 2352 10046 2408
rect 10102 2352 25594 2408
rect 25650 2352 25655 2408
rect 10041 2350 25655 2352
rect 10041 2347 10107 2350
rect 25589 2347 25655 2350
rect 0 2184 800 2304
rect 67633 2274 67699 2277
rect 69200 2274 70000 2304
rect 67633 2272 70000 2274
rect 67633 2216 67638 2272
rect 67694 2216 70000 2272
rect 67633 2214 70000 2216
rect 67633 2211 67699 2214
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
rect 50290 2208 50606 2209
rect 50290 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50606 2208
rect 69200 2184 70000 2214
rect 50290 2143 50606 2144
rect 6453 2138 6519 2141
rect 10869 2138 10935 2141
rect 15653 2138 15719 2141
rect 6453 2136 15719 2138
rect 6453 2080 6458 2136
rect 6514 2080 10874 2136
rect 10930 2080 15658 2136
rect 15714 2080 15719 2136
rect 6453 2078 15719 2080
rect 6453 2075 6519 2078
rect 10869 2075 10935 2078
rect 15653 2075 15719 2078
rect 6729 2002 6795 2005
rect 19057 2002 19123 2005
rect 6729 2000 19123 2002
rect 6729 1944 6734 2000
rect 6790 1944 19062 2000
rect 19118 1944 19123 2000
rect 6729 1942 19123 1944
rect 6729 1939 6795 1942
rect 19057 1939 19123 1942
rect 9029 1866 9095 1869
rect 15837 1866 15903 1869
rect 9029 1864 15903 1866
rect 9029 1808 9034 1864
rect 9090 1808 15842 1864
rect 15898 1808 15903 1864
rect 9029 1806 15903 1808
rect 9029 1803 9095 1806
rect 15837 1803 15903 1806
rect 12709 1322 12775 1325
rect 12893 1322 12959 1325
rect 12709 1320 12959 1322
rect 12709 1264 12714 1320
rect 12770 1264 12898 1320
rect 12954 1264 12959 1320
rect 12709 1262 12959 1264
rect 12709 1259 12775 1262
rect 12893 1259 12959 1262
<< via3 >>
rect 19576 57692 19640 57696
rect 19576 57636 19580 57692
rect 19580 57636 19636 57692
rect 19636 57636 19640 57692
rect 19576 57632 19640 57636
rect 19656 57692 19720 57696
rect 19656 57636 19660 57692
rect 19660 57636 19716 57692
rect 19716 57636 19720 57692
rect 19656 57632 19720 57636
rect 19736 57692 19800 57696
rect 19736 57636 19740 57692
rect 19740 57636 19796 57692
rect 19796 57636 19800 57692
rect 19736 57632 19800 57636
rect 19816 57692 19880 57696
rect 19816 57636 19820 57692
rect 19820 57636 19876 57692
rect 19876 57636 19880 57692
rect 19816 57632 19880 57636
rect 50296 57692 50360 57696
rect 50296 57636 50300 57692
rect 50300 57636 50356 57692
rect 50356 57636 50360 57692
rect 50296 57632 50360 57636
rect 50376 57692 50440 57696
rect 50376 57636 50380 57692
rect 50380 57636 50436 57692
rect 50436 57636 50440 57692
rect 50376 57632 50440 57636
rect 50456 57692 50520 57696
rect 50456 57636 50460 57692
rect 50460 57636 50516 57692
rect 50516 57636 50520 57692
rect 50456 57632 50520 57636
rect 50536 57692 50600 57696
rect 50536 57636 50540 57692
rect 50540 57636 50596 57692
rect 50596 57636 50600 57692
rect 50536 57632 50600 57636
rect 4216 57148 4280 57152
rect 4216 57092 4220 57148
rect 4220 57092 4276 57148
rect 4276 57092 4280 57148
rect 4216 57088 4280 57092
rect 4296 57148 4360 57152
rect 4296 57092 4300 57148
rect 4300 57092 4356 57148
rect 4356 57092 4360 57148
rect 4296 57088 4360 57092
rect 4376 57148 4440 57152
rect 4376 57092 4380 57148
rect 4380 57092 4436 57148
rect 4436 57092 4440 57148
rect 4376 57088 4440 57092
rect 4456 57148 4520 57152
rect 4456 57092 4460 57148
rect 4460 57092 4516 57148
rect 4516 57092 4520 57148
rect 4456 57088 4520 57092
rect 34936 57148 35000 57152
rect 34936 57092 34940 57148
rect 34940 57092 34996 57148
rect 34996 57092 35000 57148
rect 34936 57088 35000 57092
rect 35016 57148 35080 57152
rect 35016 57092 35020 57148
rect 35020 57092 35076 57148
rect 35076 57092 35080 57148
rect 35016 57088 35080 57092
rect 35096 57148 35160 57152
rect 35096 57092 35100 57148
rect 35100 57092 35156 57148
rect 35156 57092 35160 57148
rect 35096 57088 35160 57092
rect 35176 57148 35240 57152
rect 35176 57092 35180 57148
rect 35180 57092 35236 57148
rect 35236 57092 35240 57148
rect 35176 57088 35240 57092
rect 65656 57148 65720 57152
rect 65656 57092 65660 57148
rect 65660 57092 65716 57148
rect 65716 57092 65720 57148
rect 65656 57088 65720 57092
rect 65736 57148 65800 57152
rect 65736 57092 65740 57148
rect 65740 57092 65796 57148
rect 65796 57092 65800 57148
rect 65736 57088 65800 57092
rect 65816 57148 65880 57152
rect 65816 57092 65820 57148
rect 65820 57092 65876 57148
rect 65876 57092 65880 57148
rect 65816 57088 65880 57092
rect 65896 57148 65960 57152
rect 65896 57092 65900 57148
rect 65900 57092 65956 57148
rect 65956 57092 65960 57148
rect 65896 57088 65960 57092
rect 19576 56604 19640 56608
rect 19576 56548 19580 56604
rect 19580 56548 19636 56604
rect 19636 56548 19640 56604
rect 19576 56544 19640 56548
rect 19656 56604 19720 56608
rect 19656 56548 19660 56604
rect 19660 56548 19716 56604
rect 19716 56548 19720 56604
rect 19656 56544 19720 56548
rect 19736 56604 19800 56608
rect 19736 56548 19740 56604
rect 19740 56548 19796 56604
rect 19796 56548 19800 56604
rect 19736 56544 19800 56548
rect 19816 56604 19880 56608
rect 19816 56548 19820 56604
rect 19820 56548 19876 56604
rect 19876 56548 19880 56604
rect 19816 56544 19880 56548
rect 50296 56604 50360 56608
rect 50296 56548 50300 56604
rect 50300 56548 50356 56604
rect 50356 56548 50360 56604
rect 50296 56544 50360 56548
rect 50376 56604 50440 56608
rect 50376 56548 50380 56604
rect 50380 56548 50436 56604
rect 50436 56548 50440 56604
rect 50376 56544 50440 56548
rect 50456 56604 50520 56608
rect 50456 56548 50460 56604
rect 50460 56548 50516 56604
rect 50516 56548 50520 56604
rect 50456 56544 50520 56548
rect 50536 56604 50600 56608
rect 50536 56548 50540 56604
rect 50540 56548 50596 56604
rect 50596 56548 50600 56604
rect 50536 56544 50600 56548
rect 4216 56060 4280 56064
rect 4216 56004 4220 56060
rect 4220 56004 4276 56060
rect 4276 56004 4280 56060
rect 4216 56000 4280 56004
rect 4296 56060 4360 56064
rect 4296 56004 4300 56060
rect 4300 56004 4356 56060
rect 4356 56004 4360 56060
rect 4296 56000 4360 56004
rect 4376 56060 4440 56064
rect 4376 56004 4380 56060
rect 4380 56004 4436 56060
rect 4436 56004 4440 56060
rect 4376 56000 4440 56004
rect 4456 56060 4520 56064
rect 4456 56004 4460 56060
rect 4460 56004 4516 56060
rect 4516 56004 4520 56060
rect 4456 56000 4520 56004
rect 34936 56060 35000 56064
rect 34936 56004 34940 56060
rect 34940 56004 34996 56060
rect 34996 56004 35000 56060
rect 34936 56000 35000 56004
rect 35016 56060 35080 56064
rect 35016 56004 35020 56060
rect 35020 56004 35076 56060
rect 35076 56004 35080 56060
rect 35016 56000 35080 56004
rect 35096 56060 35160 56064
rect 35096 56004 35100 56060
rect 35100 56004 35156 56060
rect 35156 56004 35160 56060
rect 35096 56000 35160 56004
rect 35176 56060 35240 56064
rect 35176 56004 35180 56060
rect 35180 56004 35236 56060
rect 35236 56004 35240 56060
rect 35176 56000 35240 56004
rect 65656 56060 65720 56064
rect 65656 56004 65660 56060
rect 65660 56004 65716 56060
rect 65716 56004 65720 56060
rect 65656 56000 65720 56004
rect 65736 56060 65800 56064
rect 65736 56004 65740 56060
rect 65740 56004 65796 56060
rect 65796 56004 65800 56060
rect 65736 56000 65800 56004
rect 65816 56060 65880 56064
rect 65816 56004 65820 56060
rect 65820 56004 65876 56060
rect 65876 56004 65880 56060
rect 65816 56000 65880 56004
rect 65896 56060 65960 56064
rect 65896 56004 65900 56060
rect 65900 56004 65956 56060
rect 65956 56004 65960 56060
rect 65896 56000 65960 56004
rect 19576 55516 19640 55520
rect 19576 55460 19580 55516
rect 19580 55460 19636 55516
rect 19636 55460 19640 55516
rect 19576 55456 19640 55460
rect 19656 55516 19720 55520
rect 19656 55460 19660 55516
rect 19660 55460 19716 55516
rect 19716 55460 19720 55516
rect 19656 55456 19720 55460
rect 19736 55516 19800 55520
rect 19736 55460 19740 55516
rect 19740 55460 19796 55516
rect 19796 55460 19800 55516
rect 19736 55456 19800 55460
rect 19816 55516 19880 55520
rect 19816 55460 19820 55516
rect 19820 55460 19876 55516
rect 19876 55460 19880 55516
rect 19816 55456 19880 55460
rect 50296 55516 50360 55520
rect 50296 55460 50300 55516
rect 50300 55460 50356 55516
rect 50356 55460 50360 55516
rect 50296 55456 50360 55460
rect 50376 55516 50440 55520
rect 50376 55460 50380 55516
rect 50380 55460 50436 55516
rect 50436 55460 50440 55516
rect 50376 55456 50440 55460
rect 50456 55516 50520 55520
rect 50456 55460 50460 55516
rect 50460 55460 50516 55516
rect 50516 55460 50520 55516
rect 50456 55456 50520 55460
rect 50536 55516 50600 55520
rect 50536 55460 50540 55516
rect 50540 55460 50596 55516
rect 50596 55460 50600 55516
rect 50536 55456 50600 55460
rect 4216 54972 4280 54976
rect 4216 54916 4220 54972
rect 4220 54916 4276 54972
rect 4276 54916 4280 54972
rect 4216 54912 4280 54916
rect 4296 54972 4360 54976
rect 4296 54916 4300 54972
rect 4300 54916 4356 54972
rect 4356 54916 4360 54972
rect 4296 54912 4360 54916
rect 4376 54972 4440 54976
rect 4376 54916 4380 54972
rect 4380 54916 4436 54972
rect 4436 54916 4440 54972
rect 4376 54912 4440 54916
rect 4456 54972 4520 54976
rect 4456 54916 4460 54972
rect 4460 54916 4516 54972
rect 4516 54916 4520 54972
rect 4456 54912 4520 54916
rect 34936 54972 35000 54976
rect 34936 54916 34940 54972
rect 34940 54916 34996 54972
rect 34996 54916 35000 54972
rect 34936 54912 35000 54916
rect 35016 54972 35080 54976
rect 35016 54916 35020 54972
rect 35020 54916 35076 54972
rect 35076 54916 35080 54972
rect 35016 54912 35080 54916
rect 35096 54972 35160 54976
rect 35096 54916 35100 54972
rect 35100 54916 35156 54972
rect 35156 54916 35160 54972
rect 35096 54912 35160 54916
rect 35176 54972 35240 54976
rect 35176 54916 35180 54972
rect 35180 54916 35236 54972
rect 35236 54916 35240 54972
rect 35176 54912 35240 54916
rect 65656 54972 65720 54976
rect 65656 54916 65660 54972
rect 65660 54916 65716 54972
rect 65716 54916 65720 54972
rect 65656 54912 65720 54916
rect 65736 54972 65800 54976
rect 65736 54916 65740 54972
rect 65740 54916 65796 54972
rect 65796 54916 65800 54972
rect 65736 54912 65800 54916
rect 65816 54972 65880 54976
rect 65816 54916 65820 54972
rect 65820 54916 65876 54972
rect 65876 54916 65880 54972
rect 65816 54912 65880 54916
rect 65896 54972 65960 54976
rect 65896 54916 65900 54972
rect 65900 54916 65956 54972
rect 65956 54916 65960 54972
rect 65896 54912 65960 54916
rect 19576 54428 19640 54432
rect 19576 54372 19580 54428
rect 19580 54372 19636 54428
rect 19636 54372 19640 54428
rect 19576 54368 19640 54372
rect 19656 54428 19720 54432
rect 19656 54372 19660 54428
rect 19660 54372 19716 54428
rect 19716 54372 19720 54428
rect 19656 54368 19720 54372
rect 19736 54428 19800 54432
rect 19736 54372 19740 54428
rect 19740 54372 19796 54428
rect 19796 54372 19800 54428
rect 19736 54368 19800 54372
rect 19816 54428 19880 54432
rect 19816 54372 19820 54428
rect 19820 54372 19876 54428
rect 19876 54372 19880 54428
rect 19816 54368 19880 54372
rect 50296 54428 50360 54432
rect 50296 54372 50300 54428
rect 50300 54372 50356 54428
rect 50356 54372 50360 54428
rect 50296 54368 50360 54372
rect 50376 54428 50440 54432
rect 50376 54372 50380 54428
rect 50380 54372 50436 54428
rect 50436 54372 50440 54428
rect 50376 54368 50440 54372
rect 50456 54428 50520 54432
rect 50456 54372 50460 54428
rect 50460 54372 50516 54428
rect 50516 54372 50520 54428
rect 50456 54368 50520 54372
rect 50536 54428 50600 54432
rect 50536 54372 50540 54428
rect 50540 54372 50596 54428
rect 50596 54372 50600 54428
rect 50536 54368 50600 54372
rect 4216 53884 4280 53888
rect 4216 53828 4220 53884
rect 4220 53828 4276 53884
rect 4276 53828 4280 53884
rect 4216 53824 4280 53828
rect 4296 53884 4360 53888
rect 4296 53828 4300 53884
rect 4300 53828 4356 53884
rect 4356 53828 4360 53884
rect 4296 53824 4360 53828
rect 4376 53884 4440 53888
rect 4376 53828 4380 53884
rect 4380 53828 4436 53884
rect 4436 53828 4440 53884
rect 4376 53824 4440 53828
rect 4456 53884 4520 53888
rect 4456 53828 4460 53884
rect 4460 53828 4516 53884
rect 4516 53828 4520 53884
rect 4456 53824 4520 53828
rect 34936 53884 35000 53888
rect 34936 53828 34940 53884
rect 34940 53828 34996 53884
rect 34996 53828 35000 53884
rect 34936 53824 35000 53828
rect 35016 53884 35080 53888
rect 35016 53828 35020 53884
rect 35020 53828 35076 53884
rect 35076 53828 35080 53884
rect 35016 53824 35080 53828
rect 35096 53884 35160 53888
rect 35096 53828 35100 53884
rect 35100 53828 35156 53884
rect 35156 53828 35160 53884
rect 35096 53824 35160 53828
rect 35176 53884 35240 53888
rect 35176 53828 35180 53884
rect 35180 53828 35236 53884
rect 35236 53828 35240 53884
rect 35176 53824 35240 53828
rect 65656 53884 65720 53888
rect 65656 53828 65660 53884
rect 65660 53828 65716 53884
rect 65716 53828 65720 53884
rect 65656 53824 65720 53828
rect 65736 53884 65800 53888
rect 65736 53828 65740 53884
rect 65740 53828 65796 53884
rect 65796 53828 65800 53884
rect 65736 53824 65800 53828
rect 65816 53884 65880 53888
rect 65816 53828 65820 53884
rect 65820 53828 65876 53884
rect 65876 53828 65880 53884
rect 65816 53824 65880 53828
rect 65896 53884 65960 53888
rect 65896 53828 65900 53884
rect 65900 53828 65956 53884
rect 65956 53828 65960 53884
rect 65896 53824 65960 53828
rect 19576 53340 19640 53344
rect 19576 53284 19580 53340
rect 19580 53284 19636 53340
rect 19636 53284 19640 53340
rect 19576 53280 19640 53284
rect 19656 53340 19720 53344
rect 19656 53284 19660 53340
rect 19660 53284 19716 53340
rect 19716 53284 19720 53340
rect 19656 53280 19720 53284
rect 19736 53340 19800 53344
rect 19736 53284 19740 53340
rect 19740 53284 19796 53340
rect 19796 53284 19800 53340
rect 19736 53280 19800 53284
rect 19816 53340 19880 53344
rect 19816 53284 19820 53340
rect 19820 53284 19876 53340
rect 19876 53284 19880 53340
rect 19816 53280 19880 53284
rect 50296 53340 50360 53344
rect 50296 53284 50300 53340
rect 50300 53284 50356 53340
rect 50356 53284 50360 53340
rect 50296 53280 50360 53284
rect 50376 53340 50440 53344
rect 50376 53284 50380 53340
rect 50380 53284 50436 53340
rect 50436 53284 50440 53340
rect 50376 53280 50440 53284
rect 50456 53340 50520 53344
rect 50456 53284 50460 53340
rect 50460 53284 50516 53340
rect 50516 53284 50520 53340
rect 50456 53280 50520 53284
rect 50536 53340 50600 53344
rect 50536 53284 50540 53340
rect 50540 53284 50596 53340
rect 50596 53284 50600 53340
rect 50536 53280 50600 53284
rect 4216 52796 4280 52800
rect 4216 52740 4220 52796
rect 4220 52740 4276 52796
rect 4276 52740 4280 52796
rect 4216 52736 4280 52740
rect 4296 52796 4360 52800
rect 4296 52740 4300 52796
rect 4300 52740 4356 52796
rect 4356 52740 4360 52796
rect 4296 52736 4360 52740
rect 4376 52796 4440 52800
rect 4376 52740 4380 52796
rect 4380 52740 4436 52796
rect 4436 52740 4440 52796
rect 4376 52736 4440 52740
rect 4456 52796 4520 52800
rect 4456 52740 4460 52796
rect 4460 52740 4516 52796
rect 4516 52740 4520 52796
rect 4456 52736 4520 52740
rect 34936 52796 35000 52800
rect 34936 52740 34940 52796
rect 34940 52740 34996 52796
rect 34996 52740 35000 52796
rect 34936 52736 35000 52740
rect 35016 52796 35080 52800
rect 35016 52740 35020 52796
rect 35020 52740 35076 52796
rect 35076 52740 35080 52796
rect 35016 52736 35080 52740
rect 35096 52796 35160 52800
rect 35096 52740 35100 52796
rect 35100 52740 35156 52796
rect 35156 52740 35160 52796
rect 35096 52736 35160 52740
rect 35176 52796 35240 52800
rect 35176 52740 35180 52796
rect 35180 52740 35236 52796
rect 35236 52740 35240 52796
rect 35176 52736 35240 52740
rect 65656 52796 65720 52800
rect 65656 52740 65660 52796
rect 65660 52740 65716 52796
rect 65716 52740 65720 52796
rect 65656 52736 65720 52740
rect 65736 52796 65800 52800
rect 65736 52740 65740 52796
rect 65740 52740 65796 52796
rect 65796 52740 65800 52796
rect 65736 52736 65800 52740
rect 65816 52796 65880 52800
rect 65816 52740 65820 52796
rect 65820 52740 65876 52796
rect 65876 52740 65880 52796
rect 65816 52736 65880 52740
rect 65896 52796 65960 52800
rect 65896 52740 65900 52796
rect 65900 52740 65956 52796
rect 65956 52740 65960 52796
rect 65896 52736 65960 52740
rect 19576 52252 19640 52256
rect 19576 52196 19580 52252
rect 19580 52196 19636 52252
rect 19636 52196 19640 52252
rect 19576 52192 19640 52196
rect 19656 52252 19720 52256
rect 19656 52196 19660 52252
rect 19660 52196 19716 52252
rect 19716 52196 19720 52252
rect 19656 52192 19720 52196
rect 19736 52252 19800 52256
rect 19736 52196 19740 52252
rect 19740 52196 19796 52252
rect 19796 52196 19800 52252
rect 19736 52192 19800 52196
rect 19816 52252 19880 52256
rect 19816 52196 19820 52252
rect 19820 52196 19876 52252
rect 19876 52196 19880 52252
rect 19816 52192 19880 52196
rect 50296 52252 50360 52256
rect 50296 52196 50300 52252
rect 50300 52196 50356 52252
rect 50356 52196 50360 52252
rect 50296 52192 50360 52196
rect 50376 52252 50440 52256
rect 50376 52196 50380 52252
rect 50380 52196 50436 52252
rect 50436 52196 50440 52252
rect 50376 52192 50440 52196
rect 50456 52252 50520 52256
rect 50456 52196 50460 52252
rect 50460 52196 50516 52252
rect 50516 52196 50520 52252
rect 50456 52192 50520 52196
rect 50536 52252 50600 52256
rect 50536 52196 50540 52252
rect 50540 52196 50596 52252
rect 50596 52196 50600 52252
rect 50536 52192 50600 52196
rect 4216 51708 4280 51712
rect 4216 51652 4220 51708
rect 4220 51652 4276 51708
rect 4276 51652 4280 51708
rect 4216 51648 4280 51652
rect 4296 51708 4360 51712
rect 4296 51652 4300 51708
rect 4300 51652 4356 51708
rect 4356 51652 4360 51708
rect 4296 51648 4360 51652
rect 4376 51708 4440 51712
rect 4376 51652 4380 51708
rect 4380 51652 4436 51708
rect 4436 51652 4440 51708
rect 4376 51648 4440 51652
rect 4456 51708 4520 51712
rect 4456 51652 4460 51708
rect 4460 51652 4516 51708
rect 4516 51652 4520 51708
rect 4456 51648 4520 51652
rect 34936 51708 35000 51712
rect 34936 51652 34940 51708
rect 34940 51652 34996 51708
rect 34996 51652 35000 51708
rect 34936 51648 35000 51652
rect 35016 51708 35080 51712
rect 35016 51652 35020 51708
rect 35020 51652 35076 51708
rect 35076 51652 35080 51708
rect 35016 51648 35080 51652
rect 35096 51708 35160 51712
rect 35096 51652 35100 51708
rect 35100 51652 35156 51708
rect 35156 51652 35160 51708
rect 35096 51648 35160 51652
rect 35176 51708 35240 51712
rect 35176 51652 35180 51708
rect 35180 51652 35236 51708
rect 35236 51652 35240 51708
rect 35176 51648 35240 51652
rect 65656 51708 65720 51712
rect 65656 51652 65660 51708
rect 65660 51652 65716 51708
rect 65716 51652 65720 51708
rect 65656 51648 65720 51652
rect 65736 51708 65800 51712
rect 65736 51652 65740 51708
rect 65740 51652 65796 51708
rect 65796 51652 65800 51708
rect 65736 51648 65800 51652
rect 65816 51708 65880 51712
rect 65816 51652 65820 51708
rect 65820 51652 65876 51708
rect 65876 51652 65880 51708
rect 65816 51648 65880 51652
rect 65896 51708 65960 51712
rect 65896 51652 65900 51708
rect 65900 51652 65956 51708
rect 65956 51652 65960 51708
rect 65896 51648 65960 51652
rect 19576 51164 19640 51168
rect 19576 51108 19580 51164
rect 19580 51108 19636 51164
rect 19636 51108 19640 51164
rect 19576 51104 19640 51108
rect 19656 51164 19720 51168
rect 19656 51108 19660 51164
rect 19660 51108 19716 51164
rect 19716 51108 19720 51164
rect 19656 51104 19720 51108
rect 19736 51164 19800 51168
rect 19736 51108 19740 51164
rect 19740 51108 19796 51164
rect 19796 51108 19800 51164
rect 19736 51104 19800 51108
rect 19816 51164 19880 51168
rect 19816 51108 19820 51164
rect 19820 51108 19876 51164
rect 19876 51108 19880 51164
rect 19816 51104 19880 51108
rect 50296 51164 50360 51168
rect 50296 51108 50300 51164
rect 50300 51108 50356 51164
rect 50356 51108 50360 51164
rect 50296 51104 50360 51108
rect 50376 51164 50440 51168
rect 50376 51108 50380 51164
rect 50380 51108 50436 51164
rect 50436 51108 50440 51164
rect 50376 51104 50440 51108
rect 50456 51164 50520 51168
rect 50456 51108 50460 51164
rect 50460 51108 50516 51164
rect 50516 51108 50520 51164
rect 50456 51104 50520 51108
rect 50536 51164 50600 51168
rect 50536 51108 50540 51164
rect 50540 51108 50596 51164
rect 50596 51108 50600 51164
rect 50536 51104 50600 51108
rect 4216 50620 4280 50624
rect 4216 50564 4220 50620
rect 4220 50564 4276 50620
rect 4276 50564 4280 50620
rect 4216 50560 4280 50564
rect 4296 50620 4360 50624
rect 4296 50564 4300 50620
rect 4300 50564 4356 50620
rect 4356 50564 4360 50620
rect 4296 50560 4360 50564
rect 4376 50620 4440 50624
rect 4376 50564 4380 50620
rect 4380 50564 4436 50620
rect 4436 50564 4440 50620
rect 4376 50560 4440 50564
rect 4456 50620 4520 50624
rect 4456 50564 4460 50620
rect 4460 50564 4516 50620
rect 4516 50564 4520 50620
rect 4456 50560 4520 50564
rect 34936 50620 35000 50624
rect 34936 50564 34940 50620
rect 34940 50564 34996 50620
rect 34996 50564 35000 50620
rect 34936 50560 35000 50564
rect 35016 50620 35080 50624
rect 35016 50564 35020 50620
rect 35020 50564 35076 50620
rect 35076 50564 35080 50620
rect 35016 50560 35080 50564
rect 35096 50620 35160 50624
rect 35096 50564 35100 50620
rect 35100 50564 35156 50620
rect 35156 50564 35160 50620
rect 35096 50560 35160 50564
rect 35176 50620 35240 50624
rect 35176 50564 35180 50620
rect 35180 50564 35236 50620
rect 35236 50564 35240 50620
rect 35176 50560 35240 50564
rect 65656 50620 65720 50624
rect 65656 50564 65660 50620
rect 65660 50564 65716 50620
rect 65716 50564 65720 50620
rect 65656 50560 65720 50564
rect 65736 50620 65800 50624
rect 65736 50564 65740 50620
rect 65740 50564 65796 50620
rect 65796 50564 65800 50620
rect 65736 50560 65800 50564
rect 65816 50620 65880 50624
rect 65816 50564 65820 50620
rect 65820 50564 65876 50620
rect 65876 50564 65880 50620
rect 65816 50560 65880 50564
rect 65896 50620 65960 50624
rect 65896 50564 65900 50620
rect 65900 50564 65956 50620
rect 65956 50564 65960 50620
rect 65896 50560 65960 50564
rect 19576 50076 19640 50080
rect 19576 50020 19580 50076
rect 19580 50020 19636 50076
rect 19636 50020 19640 50076
rect 19576 50016 19640 50020
rect 19656 50076 19720 50080
rect 19656 50020 19660 50076
rect 19660 50020 19716 50076
rect 19716 50020 19720 50076
rect 19656 50016 19720 50020
rect 19736 50076 19800 50080
rect 19736 50020 19740 50076
rect 19740 50020 19796 50076
rect 19796 50020 19800 50076
rect 19736 50016 19800 50020
rect 19816 50076 19880 50080
rect 19816 50020 19820 50076
rect 19820 50020 19876 50076
rect 19876 50020 19880 50076
rect 19816 50016 19880 50020
rect 50296 50076 50360 50080
rect 50296 50020 50300 50076
rect 50300 50020 50356 50076
rect 50356 50020 50360 50076
rect 50296 50016 50360 50020
rect 50376 50076 50440 50080
rect 50376 50020 50380 50076
rect 50380 50020 50436 50076
rect 50436 50020 50440 50076
rect 50376 50016 50440 50020
rect 50456 50076 50520 50080
rect 50456 50020 50460 50076
rect 50460 50020 50516 50076
rect 50516 50020 50520 50076
rect 50456 50016 50520 50020
rect 50536 50076 50600 50080
rect 50536 50020 50540 50076
rect 50540 50020 50596 50076
rect 50596 50020 50600 50076
rect 50536 50016 50600 50020
rect 4216 49532 4280 49536
rect 4216 49476 4220 49532
rect 4220 49476 4276 49532
rect 4276 49476 4280 49532
rect 4216 49472 4280 49476
rect 4296 49532 4360 49536
rect 4296 49476 4300 49532
rect 4300 49476 4356 49532
rect 4356 49476 4360 49532
rect 4296 49472 4360 49476
rect 4376 49532 4440 49536
rect 4376 49476 4380 49532
rect 4380 49476 4436 49532
rect 4436 49476 4440 49532
rect 4376 49472 4440 49476
rect 4456 49532 4520 49536
rect 4456 49476 4460 49532
rect 4460 49476 4516 49532
rect 4516 49476 4520 49532
rect 4456 49472 4520 49476
rect 34936 49532 35000 49536
rect 34936 49476 34940 49532
rect 34940 49476 34996 49532
rect 34996 49476 35000 49532
rect 34936 49472 35000 49476
rect 35016 49532 35080 49536
rect 35016 49476 35020 49532
rect 35020 49476 35076 49532
rect 35076 49476 35080 49532
rect 35016 49472 35080 49476
rect 35096 49532 35160 49536
rect 35096 49476 35100 49532
rect 35100 49476 35156 49532
rect 35156 49476 35160 49532
rect 35096 49472 35160 49476
rect 35176 49532 35240 49536
rect 35176 49476 35180 49532
rect 35180 49476 35236 49532
rect 35236 49476 35240 49532
rect 35176 49472 35240 49476
rect 65656 49532 65720 49536
rect 65656 49476 65660 49532
rect 65660 49476 65716 49532
rect 65716 49476 65720 49532
rect 65656 49472 65720 49476
rect 65736 49532 65800 49536
rect 65736 49476 65740 49532
rect 65740 49476 65796 49532
rect 65796 49476 65800 49532
rect 65736 49472 65800 49476
rect 65816 49532 65880 49536
rect 65816 49476 65820 49532
rect 65820 49476 65876 49532
rect 65876 49476 65880 49532
rect 65816 49472 65880 49476
rect 65896 49532 65960 49536
rect 65896 49476 65900 49532
rect 65900 49476 65956 49532
rect 65956 49476 65960 49532
rect 65896 49472 65960 49476
rect 19576 48988 19640 48992
rect 19576 48932 19580 48988
rect 19580 48932 19636 48988
rect 19636 48932 19640 48988
rect 19576 48928 19640 48932
rect 19656 48988 19720 48992
rect 19656 48932 19660 48988
rect 19660 48932 19716 48988
rect 19716 48932 19720 48988
rect 19656 48928 19720 48932
rect 19736 48988 19800 48992
rect 19736 48932 19740 48988
rect 19740 48932 19796 48988
rect 19796 48932 19800 48988
rect 19736 48928 19800 48932
rect 19816 48988 19880 48992
rect 19816 48932 19820 48988
rect 19820 48932 19876 48988
rect 19876 48932 19880 48988
rect 19816 48928 19880 48932
rect 50296 48988 50360 48992
rect 50296 48932 50300 48988
rect 50300 48932 50356 48988
rect 50356 48932 50360 48988
rect 50296 48928 50360 48932
rect 50376 48988 50440 48992
rect 50376 48932 50380 48988
rect 50380 48932 50436 48988
rect 50436 48932 50440 48988
rect 50376 48928 50440 48932
rect 50456 48988 50520 48992
rect 50456 48932 50460 48988
rect 50460 48932 50516 48988
rect 50516 48932 50520 48988
rect 50456 48928 50520 48932
rect 50536 48988 50600 48992
rect 50536 48932 50540 48988
rect 50540 48932 50596 48988
rect 50596 48932 50600 48988
rect 50536 48928 50600 48932
rect 4216 48444 4280 48448
rect 4216 48388 4220 48444
rect 4220 48388 4276 48444
rect 4276 48388 4280 48444
rect 4216 48384 4280 48388
rect 4296 48444 4360 48448
rect 4296 48388 4300 48444
rect 4300 48388 4356 48444
rect 4356 48388 4360 48444
rect 4296 48384 4360 48388
rect 4376 48444 4440 48448
rect 4376 48388 4380 48444
rect 4380 48388 4436 48444
rect 4436 48388 4440 48444
rect 4376 48384 4440 48388
rect 4456 48444 4520 48448
rect 4456 48388 4460 48444
rect 4460 48388 4516 48444
rect 4516 48388 4520 48444
rect 4456 48384 4520 48388
rect 34936 48444 35000 48448
rect 34936 48388 34940 48444
rect 34940 48388 34996 48444
rect 34996 48388 35000 48444
rect 34936 48384 35000 48388
rect 35016 48444 35080 48448
rect 35016 48388 35020 48444
rect 35020 48388 35076 48444
rect 35076 48388 35080 48444
rect 35016 48384 35080 48388
rect 35096 48444 35160 48448
rect 35096 48388 35100 48444
rect 35100 48388 35156 48444
rect 35156 48388 35160 48444
rect 35096 48384 35160 48388
rect 35176 48444 35240 48448
rect 35176 48388 35180 48444
rect 35180 48388 35236 48444
rect 35236 48388 35240 48444
rect 35176 48384 35240 48388
rect 65656 48444 65720 48448
rect 65656 48388 65660 48444
rect 65660 48388 65716 48444
rect 65716 48388 65720 48444
rect 65656 48384 65720 48388
rect 65736 48444 65800 48448
rect 65736 48388 65740 48444
rect 65740 48388 65796 48444
rect 65796 48388 65800 48444
rect 65736 48384 65800 48388
rect 65816 48444 65880 48448
rect 65816 48388 65820 48444
rect 65820 48388 65876 48444
rect 65876 48388 65880 48444
rect 65816 48384 65880 48388
rect 65896 48444 65960 48448
rect 65896 48388 65900 48444
rect 65900 48388 65956 48444
rect 65956 48388 65960 48444
rect 65896 48384 65960 48388
rect 19576 47900 19640 47904
rect 19576 47844 19580 47900
rect 19580 47844 19636 47900
rect 19636 47844 19640 47900
rect 19576 47840 19640 47844
rect 19656 47900 19720 47904
rect 19656 47844 19660 47900
rect 19660 47844 19716 47900
rect 19716 47844 19720 47900
rect 19656 47840 19720 47844
rect 19736 47900 19800 47904
rect 19736 47844 19740 47900
rect 19740 47844 19796 47900
rect 19796 47844 19800 47900
rect 19736 47840 19800 47844
rect 19816 47900 19880 47904
rect 19816 47844 19820 47900
rect 19820 47844 19876 47900
rect 19876 47844 19880 47900
rect 19816 47840 19880 47844
rect 50296 47900 50360 47904
rect 50296 47844 50300 47900
rect 50300 47844 50356 47900
rect 50356 47844 50360 47900
rect 50296 47840 50360 47844
rect 50376 47900 50440 47904
rect 50376 47844 50380 47900
rect 50380 47844 50436 47900
rect 50436 47844 50440 47900
rect 50376 47840 50440 47844
rect 50456 47900 50520 47904
rect 50456 47844 50460 47900
rect 50460 47844 50516 47900
rect 50516 47844 50520 47900
rect 50456 47840 50520 47844
rect 50536 47900 50600 47904
rect 50536 47844 50540 47900
rect 50540 47844 50596 47900
rect 50596 47844 50600 47900
rect 50536 47840 50600 47844
rect 4216 47356 4280 47360
rect 4216 47300 4220 47356
rect 4220 47300 4276 47356
rect 4276 47300 4280 47356
rect 4216 47296 4280 47300
rect 4296 47356 4360 47360
rect 4296 47300 4300 47356
rect 4300 47300 4356 47356
rect 4356 47300 4360 47356
rect 4296 47296 4360 47300
rect 4376 47356 4440 47360
rect 4376 47300 4380 47356
rect 4380 47300 4436 47356
rect 4436 47300 4440 47356
rect 4376 47296 4440 47300
rect 4456 47356 4520 47360
rect 4456 47300 4460 47356
rect 4460 47300 4516 47356
rect 4516 47300 4520 47356
rect 4456 47296 4520 47300
rect 34936 47356 35000 47360
rect 34936 47300 34940 47356
rect 34940 47300 34996 47356
rect 34996 47300 35000 47356
rect 34936 47296 35000 47300
rect 35016 47356 35080 47360
rect 35016 47300 35020 47356
rect 35020 47300 35076 47356
rect 35076 47300 35080 47356
rect 35016 47296 35080 47300
rect 35096 47356 35160 47360
rect 35096 47300 35100 47356
rect 35100 47300 35156 47356
rect 35156 47300 35160 47356
rect 35096 47296 35160 47300
rect 35176 47356 35240 47360
rect 35176 47300 35180 47356
rect 35180 47300 35236 47356
rect 35236 47300 35240 47356
rect 35176 47296 35240 47300
rect 65656 47356 65720 47360
rect 65656 47300 65660 47356
rect 65660 47300 65716 47356
rect 65716 47300 65720 47356
rect 65656 47296 65720 47300
rect 65736 47356 65800 47360
rect 65736 47300 65740 47356
rect 65740 47300 65796 47356
rect 65796 47300 65800 47356
rect 65736 47296 65800 47300
rect 65816 47356 65880 47360
rect 65816 47300 65820 47356
rect 65820 47300 65876 47356
rect 65876 47300 65880 47356
rect 65816 47296 65880 47300
rect 65896 47356 65960 47360
rect 65896 47300 65900 47356
rect 65900 47300 65956 47356
rect 65956 47300 65960 47356
rect 65896 47296 65960 47300
rect 19576 46812 19640 46816
rect 19576 46756 19580 46812
rect 19580 46756 19636 46812
rect 19636 46756 19640 46812
rect 19576 46752 19640 46756
rect 19656 46812 19720 46816
rect 19656 46756 19660 46812
rect 19660 46756 19716 46812
rect 19716 46756 19720 46812
rect 19656 46752 19720 46756
rect 19736 46812 19800 46816
rect 19736 46756 19740 46812
rect 19740 46756 19796 46812
rect 19796 46756 19800 46812
rect 19736 46752 19800 46756
rect 19816 46812 19880 46816
rect 19816 46756 19820 46812
rect 19820 46756 19876 46812
rect 19876 46756 19880 46812
rect 19816 46752 19880 46756
rect 50296 46812 50360 46816
rect 50296 46756 50300 46812
rect 50300 46756 50356 46812
rect 50356 46756 50360 46812
rect 50296 46752 50360 46756
rect 50376 46812 50440 46816
rect 50376 46756 50380 46812
rect 50380 46756 50436 46812
rect 50436 46756 50440 46812
rect 50376 46752 50440 46756
rect 50456 46812 50520 46816
rect 50456 46756 50460 46812
rect 50460 46756 50516 46812
rect 50516 46756 50520 46812
rect 50456 46752 50520 46756
rect 50536 46812 50600 46816
rect 50536 46756 50540 46812
rect 50540 46756 50596 46812
rect 50596 46756 50600 46812
rect 50536 46752 50600 46756
rect 4216 46268 4280 46272
rect 4216 46212 4220 46268
rect 4220 46212 4276 46268
rect 4276 46212 4280 46268
rect 4216 46208 4280 46212
rect 4296 46268 4360 46272
rect 4296 46212 4300 46268
rect 4300 46212 4356 46268
rect 4356 46212 4360 46268
rect 4296 46208 4360 46212
rect 4376 46268 4440 46272
rect 4376 46212 4380 46268
rect 4380 46212 4436 46268
rect 4436 46212 4440 46268
rect 4376 46208 4440 46212
rect 4456 46268 4520 46272
rect 4456 46212 4460 46268
rect 4460 46212 4516 46268
rect 4516 46212 4520 46268
rect 4456 46208 4520 46212
rect 34936 46268 35000 46272
rect 34936 46212 34940 46268
rect 34940 46212 34996 46268
rect 34996 46212 35000 46268
rect 34936 46208 35000 46212
rect 35016 46268 35080 46272
rect 35016 46212 35020 46268
rect 35020 46212 35076 46268
rect 35076 46212 35080 46268
rect 35016 46208 35080 46212
rect 35096 46268 35160 46272
rect 35096 46212 35100 46268
rect 35100 46212 35156 46268
rect 35156 46212 35160 46268
rect 35096 46208 35160 46212
rect 35176 46268 35240 46272
rect 35176 46212 35180 46268
rect 35180 46212 35236 46268
rect 35236 46212 35240 46268
rect 35176 46208 35240 46212
rect 65656 46268 65720 46272
rect 65656 46212 65660 46268
rect 65660 46212 65716 46268
rect 65716 46212 65720 46268
rect 65656 46208 65720 46212
rect 65736 46268 65800 46272
rect 65736 46212 65740 46268
rect 65740 46212 65796 46268
rect 65796 46212 65800 46268
rect 65736 46208 65800 46212
rect 65816 46268 65880 46272
rect 65816 46212 65820 46268
rect 65820 46212 65876 46268
rect 65876 46212 65880 46268
rect 65816 46208 65880 46212
rect 65896 46268 65960 46272
rect 65896 46212 65900 46268
rect 65900 46212 65956 46268
rect 65956 46212 65960 46268
rect 65896 46208 65960 46212
rect 19576 45724 19640 45728
rect 19576 45668 19580 45724
rect 19580 45668 19636 45724
rect 19636 45668 19640 45724
rect 19576 45664 19640 45668
rect 19656 45724 19720 45728
rect 19656 45668 19660 45724
rect 19660 45668 19716 45724
rect 19716 45668 19720 45724
rect 19656 45664 19720 45668
rect 19736 45724 19800 45728
rect 19736 45668 19740 45724
rect 19740 45668 19796 45724
rect 19796 45668 19800 45724
rect 19736 45664 19800 45668
rect 19816 45724 19880 45728
rect 19816 45668 19820 45724
rect 19820 45668 19876 45724
rect 19876 45668 19880 45724
rect 19816 45664 19880 45668
rect 50296 45724 50360 45728
rect 50296 45668 50300 45724
rect 50300 45668 50356 45724
rect 50356 45668 50360 45724
rect 50296 45664 50360 45668
rect 50376 45724 50440 45728
rect 50376 45668 50380 45724
rect 50380 45668 50436 45724
rect 50436 45668 50440 45724
rect 50376 45664 50440 45668
rect 50456 45724 50520 45728
rect 50456 45668 50460 45724
rect 50460 45668 50516 45724
rect 50516 45668 50520 45724
rect 50456 45664 50520 45668
rect 50536 45724 50600 45728
rect 50536 45668 50540 45724
rect 50540 45668 50596 45724
rect 50596 45668 50600 45724
rect 50536 45664 50600 45668
rect 4216 45180 4280 45184
rect 4216 45124 4220 45180
rect 4220 45124 4276 45180
rect 4276 45124 4280 45180
rect 4216 45120 4280 45124
rect 4296 45180 4360 45184
rect 4296 45124 4300 45180
rect 4300 45124 4356 45180
rect 4356 45124 4360 45180
rect 4296 45120 4360 45124
rect 4376 45180 4440 45184
rect 4376 45124 4380 45180
rect 4380 45124 4436 45180
rect 4436 45124 4440 45180
rect 4376 45120 4440 45124
rect 4456 45180 4520 45184
rect 4456 45124 4460 45180
rect 4460 45124 4516 45180
rect 4516 45124 4520 45180
rect 4456 45120 4520 45124
rect 34936 45180 35000 45184
rect 34936 45124 34940 45180
rect 34940 45124 34996 45180
rect 34996 45124 35000 45180
rect 34936 45120 35000 45124
rect 35016 45180 35080 45184
rect 35016 45124 35020 45180
rect 35020 45124 35076 45180
rect 35076 45124 35080 45180
rect 35016 45120 35080 45124
rect 35096 45180 35160 45184
rect 35096 45124 35100 45180
rect 35100 45124 35156 45180
rect 35156 45124 35160 45180
rect 35096 45120 35160 45124
rect 35176 45180 35240 45184
rect 35176 45124 35180 45180
rect 35180 45124 35236 45180
rect 35236 45124 35240 45180
rect 35176 45120 35240 45124
rect 65656 45180 65720 45184
rect 65656 45124 65660 45180
rect 65660 45124 65716 45180
rect 65716 45124 65720 45180
rect 65656 45120 65720 45124
rect 65736 45180 65800 45184
rect 65736 45124 65740 45180
rect 65740 45124 65796 45180
rect 65796 45124 65800 45180
rect 65736 45120 65800 45124
rect 65816 45180 65880 45184
rect 65816 45124 65820 45180
rect 65820 45124 65876 45180
rect 65876 45124 65880 45180
rect 65816 45120 65880 45124
rect 65896 45180 65960 45184
rect 65896 45124 65900 45180
rect 65900 45124 65956 45180
rect 65956 45124 65960 45180
rect 65896 45120 65960 45124
rect 19576 44636 19640 44640
rect 19576 44580 19580 44636
rect 19580 44580 19636 44636
rect 19636 44580 19640 44636
rect 19576 44576 19640 44580
rect 19656 44636 19720 44640
rect 19656 44580 19660 44636
rect 19660 44580 19716 44636
rect 19716 44580 19720 44636
rect 19656 44576 19720 44580
rect 19736 44636 19800 44640
rect 19736 44580 19740 44636
rect 19740 44580 19796 44636
rect 19796 44580 19800 44636
rect 19736 44576 19800 44580
rect 19816 44636 19880 44640
rect 19816 44580 19820 44636
rect 19820 44580 19876 44636
rect 19876 44580 19880 44636
rect 19816 44576 19880 44580
rect 50296 44636 50360 44640
rect 50296 44580 50300 44636
rect 50300 44580 50356 44636
rect 50356 44580 50360 44636
rect 50296 44576 50360 44580
rect 50376 44636 50440 44640
rect 50376 44580 50380 44636
rect 50380 44580 50436 44636
rect 50436 44580 50440 44636
rect 50376 44576 50440 44580
rect 50456 44636 50520 44640
rect 50456 44580 50460 44636
rect 50460 44580 50516 44636
rect 50516 44580 50520 44636
rect 50456 44576 50520 44580
rect 50536 44636 50600 44640
rect 50536 44580 50540 44636
rect 50540 44580 50596 44636
rect 50596 44580 50600 44636
rect 50536 44576 50600 44580
rect 4216 44092 4280 44096
rect 4216 44036 4220 44092
rect 4220 44036 4276 44092
rect 4276 44036 4280 44092
rect 4216 44032 4280 44036
rect 4296 44092 4360 44096
rect 4296 44036 4300 44092
rect 4300 44036 4356 44092
rect 4356 44036 4360 44092
rect 4296 44032 4360 44036
rect 4376 44092 4440 44096
rect 4376 44036 4380 44092
rect 4380 44036 4436 44092
rect 4436 44036 4440 44092
rect 4376 44032 4440 44036
rect 4456 44092 4520 44096
rect 4456 44036 4460 44092
rect 4460 44036 4516 44092
rect 4516 44036 4520 44092
rect 4456 44032 4520 44036
rect 34936 44092 35000 44096
rect 34936 44036 34940 44092
rect 34940 44036 34996 44092
rect 34996 44036 35000 44092
rect 34936 44032 35000 44036
rect 35016 44092 35080 44096
rect 35016 44036 35020 44092
rect 35020 44036 35076 44092
rect 35076 44036 35080 44092
rect 35016 44032 35080 44036
rect 35096 44092 35160 44096
rect 35096 44036 35100 44092
rect 35100 44036 35156 44092
rect 35156 44036 35160 44092
rect 35096 44032 35160 44036
rect 35176 44092 35240 44096
rect 35176 44036 35180 44092
rect 35180 44036 35236 44092
rect 35236 44036 35240 44092
rect 35176 44032 35240 44036
rect 65656 44092 65720 44096
rect 65656 44036 65660 44092
rect 65660 44036 65716 44092
rect 65716 44036 65720 44092
rect 65656 44032 65720 44036
rect 65736 44092 65800 44096
rect 65736 44036 65740 44092
rect 65740 44036 65796 44092
rect 65796 44036 65800 44092
rect 65736 44032 65800 44036
rect 65816 44092 65880 44096
rect 65816 44036 65820 44092
rect 65820 44036 65876 44092
rect 65876 44036 65880 44092
rect 65816 44032 65880 44036
rect 65896 44092 65960 44096
rect 65896 44036 65900 44092
rect 65900 44036 65956 44092
rect 65956 44036 65960 44092
rect 65896 44032 65960 44036
rect 19576 43548 19640 43552
rect 19576 43492 19580 43548
rect 19580 43492 19636 43548
rect 19636 43492 19640 43548
rect 19576 43488 19640 43492
rect 19656 43548 19720 43552
rect 19656 43492 19660 43548
rect 19660 43492 19716 43548
rect 19716 43492 19720 43548
rect 19656 43488 19720 43492
rect 19736 43548 19800 43552
rect 19736 43492 19740 43548
rect 19740 43492 19796 43548
rect 19796 43492 19800 43548
rect 19736 43488 19800 43492
rect 19816 43548 19880 43552
rect 19816 43492 19820 43548
rect 19820 43492 19876 43548
rect 19876 43492 19880 43548
rect 19816 43488 19880 43492
rect 50296 43548 50360 43552
rect 50296 43492 50300 43548
rect 50300 43492 50356 43548
rect 50356 43492 50360 43548
rect 50296 43488 50360 43492
rect 50376 43548 50440 43552
rect 50376 43492 50380 43548
rect 50380 43492 50436 43548
rect 50436 43492 50440 43548
rect 50376 43488 50440 43492
rect 50456 43548 50520 43552
rect 50456 43492 50460 43548
rect 50460 43492 50516 43548
rect 50516 43492 50520 43548
rect 50456 43488 50520 43492
rect 50536 43548 50600 43552
rect 50536 43492 50540 43548
rect 50540 43492 50596 43548
rect 50596 43492 50600 43548
rect 50536 43488 50600 43492
rect 4216 43004 4280 43008
rect 4216 42948 4220 43004
rect 4220 42948 4276 43004
rect 4276 42948 4280 43004
rect 4216 42944 4280 42948
rect 4296 43004 4360 43008
rect 4296 42948 4300 43004
rect 4300 42948 4356 43004
rect 4356 42948 4360 43004
rect 4296 42944 4360 42948
rect 4376 43004 4440 43008
rect 4376 42948 4380 43004
rect 4380 42948 4436 43004
rect 4436 42948 4440 43004
rect 4376 42944 4440 42948
rect 4456 43004 4520 43008
rect 4456 42948 4460 43004
rect 4460 42948 4516 43004
rect 4516 42948 4520 43004
rect 4456 42944 4520 42948
rect 34936 43004 35000 43008
rect 34936 42948 34940 43004
rect 34940 42948 34996 43004
rect 34996 42948 35000 43004
rect 34936 42944 35000 42948
rect 35016 43004 35080 43008
rect 35016 42948 35020 43004
rect 35020 42948 35076 43004
rect 35076 42948 35080 43004
rect 35016 42944 35080 42948
rect 35096 43004 35160 43008
rect 35096 42948 35100 43004
rect 35100 42948 35156 43004
rect 35156 42948 35160 43004
rect 35096 42944 35160 42948
rect 35176 43004 35240 43008
rect 35176 42948 35180 43004
rect 35180 42948 35236 43004
rect 35236 42948 35240 43004
rect 35176 42944 35240 42948
rect 65656 43004 65720 43008
rect 65656 42948 65660 43004
rect 65660 42948 65716 43004
rect 65716 42948 65720 43004
rect 65656 42944 65720 42948
rect 65736 43004 65800 43008
rect 65736 42948 65740 43004
rect 65740 42948 65796 43004
rect 65796 42948 65800 43004
rect 65736 42944 65800 42948
rect 65816 43004 65880 43008
rect 65816 42948 65820 43004
rect 65820 42948 65876 43004
rect 65876 42948 65880 43004
rect 65816 42944 65880 42948
rect 65896 43004 65960 43008
rect 65896 42948 65900 43004
rect 65900 42948 65956 43004
rect 65956 42948 65960 43004
rect 65896 42944 65960 42948
rect 19576 42460 19640 42464
rect 19576 42404 19580 42460
rect 19580 42404 19636 42460
rect 19636 42404 19640 42460
rect 19576 42400 19640 42404
rect 19656 42460 19720 42464
rect 19656 42404 19660 42460
rect 19660 42404 19716 42460
rect 19716 42404 19720 42460
rect 19656 42400 19720 42404
rect 19736 42460 19800 42464
rect 19736 42404 19740 42460
rect 19740 42404 19796 42460
rect 19796 42404 19800 42460
rect 19736 42400 19800 42404
rect 19816 42460 19880 42464
rect 19816 42404 19820 42460
rect 19820 42404 19876 42460
rect 19876 42404 19880 42460
rect 19816 42400 19880 42404
rect 50296 42460 50360 42464
rect 50296 42404 50300 42460
rect 50300 42404 50356 42460
rect 50356 42404 50360 42460
rect 50296 42400 50360 42404
rect 50376 42460 50440 42464
rect 50376 42404 50380 42460
rect 50380 42404 50436 42460
rect 50436 42404 50440 42460
rect 50376 42400 50440 42404
rect 50456 42460 50520 42464
rect 50456 42404 50460 42460
rect 50460 42404 50516 42460
rect 50516 42404 50520 42460
rect 50456 42400 50520 42404
rect 50536 42460 50600 42464
rect 50536 42404 50540 42460
rect 50540 42404 50596 42460
rect 50596 42404 50600 42460
rect 50536 42400 50600 42404
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 34936 41916 35000 41920
rect 34936 41860 34940 41916
rect 34940 41860 34996 41916
rect 34996 41860 35000 41916
rect 34936 41856 35000 41860
rect 35016 41916 35080 41920
rect 35016 41860 35020 41916
rect 35020 41860 35076 41916
rect 35076 41860 35080 41916
rect 35016 41856 35080 41860
rect 35096 41916 35160 41920
rect 35096 41860 35100 41916
rect 35100 41860 35156 41916
rect 35156 41860 35160 41916
rect 35096 41856 35160 41860
rect 35176 41916 35240 41920
rect 35176 41860 35180 41916
rect 35180 41860 35236 41916
rect 35236 41860 35240 41916
rect 35176 41856 35240 41860
rect 65656 41916 65720 41920
rect 65656 41860 65660 41916
rect 65660 41860 65716 41916
rect 65716 41860 65720 41916
rect 65656 41856 65720 41860
rect 65736 41916 65800 41920
rect 65736 41860 65740 41916
rect 65740 41860 65796 41916
rect 65796 41860 65800 41916
rect 65736 41856 65800 41860
rect 65816 41916 65880 41920
rect 65816 41860 65820 41916
rect 65820 41860 65876 41916
rect 65876 41860 65880 41916
rect 65816 41856 65880 41860
rect 65896 41916 65960 41920
rect 65896 41860 65900 41916
rect 65900 41860 65956 41916
rect 65956 41860 65960 41916
rect 65896 41856 65960 41860
rect 19576 41372 19640 41376
rect 19576 41316 19580 41372
rect 19580 41316 19636 41372
rect 19636 41316 19640 41372
rect 19576 41312 19640 41316
rect 19656 41372 19720 41376
rect 19656 41316 19660 41372
rect 19660 41316 19716 41372
rect 19716 41316 19720 41372
rect 19656 41312 19720 41316
rect 19736 41372 19800 41376
rect 19736 41316 19740 41372
rect 19740 41316 19796 41372
rect 19796 41316 19800 41372
rect 19736 41312 19800 41316
rect 19816 41372 19880 41376
rect 19816 41316 19820 41372
rect 19820 41316 19876 41372
rect 19876 41316 19880 41372
rect 19816 41312 19880 41316
rect 50296 41372 50360 41376
rect 50296 41316 50300 41372
rect 50300 41316 50356 41372
rect 50356 41316 50360 41372
rect 50296 41312 50360 41316
rect 50376 41372 50440 41376
rect 50376 41316 50380 41372
rect 50380 41316 50436 41372
rect 50436 41316 50440 41372
rect 50376 41312 50440 41316
rect 50456 41372 50520 41376
rect 50456 41316 50460 41372
rect 50460 41316 50516 41372
rect 50516 41316 50520 41372
rect 50456 41312 50520 41316
rect 50536 41372 50600 41376
rect 50536 41316 50540 41372
rect 50540 41316 50596 41372
rect 50596 41316 50600 41372
rect 50536 41312 50600 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 34936 40828 35000 40832
rect 34936 40772 34940 40828
rect 34940 40772 34996 40828
rect 34996 40772 35000 40828
rect 34936 40768 35000 40772
rect 35016 40828 35080 40832
rect 35016 40772 35020 40828
rect 35020 40772 35076 40828
rect 35076 40772 35080 40828
rect 35016 40768 35080 40772
rect 35096 40828 35160 40832
rect 35096 40772 35100 40828
rect 35100 40772 35156 40828
rect 35156 40772 35160 40828
rect 35096 40768 35160 40772
rect 35176 40828 35240 40832
rect 35176 40772 35180 40828
rect 35180 40772 35236 40828
rect 35236 40772 35240 40828
rect 35176 40768 35240 40772
rect 65656 40828 65720 40832
rect 65656 40772 65660 40828
rect 65660 40772 65716 40828
rect 65716 40772 65720 40828
rect 65656 40768 65720 40772
rect 65736 40828 65800 40832
rect 65736 40772 65740 40828
rect 65740 40772 65796 40828
rect 65796 40772 65800 40828
rect 65736 40768 65800 40772
rect 65816 40828 65880 40832
rect 65816 40772 65820 40828
rect 65820 40772 65876 40828
rect 65876 40772 65880 40828
rect 65816 40768 65880 40772
rect 65896 40828 65960 40832
rect 65896 40772 65900 40828
rect 65900 40772 65956 40828
rect 65956 40772 65960 40828
rect 65896 40768 65960 40772
rect 19576 40284 19640 40288
rect 19576 40228 19580 40284
rect 19580 40228 19636 40284
rect 19636 40228 19640 40284
rect 19576 40224 19640 40228
rect 19656 40284 19720 40288
rect 19656 40228 19660 40284
rect 19660 40228 19716 40284
rect 19716 40228 19720 40284
rect 19656 40224 19720 40228
rect 19736 40284 19800 40288
rect 19736 40228 19740 40284
rect 19740 40228 19796 40284
rect 19796 40228 19800 40284
rect 19736 40224 19800 40228
rect 19816 40284 19880 40288
rect 19816 40228 19820 40284
rect 19820 40228 19876 40284
rect 19876 40228 19880 40284
rect 19816 40224 19880 40228
rect 50296 40284 50360 40288
rect 50296 40228 50300 40284
rect 50300 40228 50356 40284
rect 50356 40228 50360 40284
rect 50296 40224 50360 40228
rect 50376 40284 50440 40288
rect 50376 40228 50380 40284
rect 50380 40228 50436 40284
rect 50436 40228 50440 40284
rect 50376 40224 50440 40228
rect 50456 40284 50520 40288
rect 50456 40228 50460 40284
rect 50460 40228 50516 40284
rect 50516 40228 50520 40284
rect 50456 40224 50520 40228
rect 50536 40284 50600 40288
rect 50536 40228 50540 40284
rect 50540 40228 50596 40284
rect 50596 40228 50600 40284
rect 50536 40224 50600 40228
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 65656 39740 65720 39744
rect 65656 39684 65660 39740
rect 65660 39684 65716 39740
rect 65716 39684 65720 39740
rect 65656 39680 65720 39684
rect 65736 39740 65800 39744
rect 65736 39684 65740 39740
rect 65740 39684 65796 39740
rect 65796 39684 65800 39740
rect 65736 39680 65800 39684
rect 65816 39740 65880 39744
rect 65816 39684 65820 39740
rect 65820 39684 65876 39740
rect 65876 39684 65880 39740
rect 65816 39680 65880 39684
rect 65896 39740 65960 39744
rect 65896 39684 65900 39740
rect 65900 39684 65956 39740
rect 65956 39684 65960 39740
rect 65896 39680 65960 39684
rect 19576 39196 19640 39200
rect 19576 39140 19580 39196
rect 19580 39140 19636 39196
rect 19636 39140 19640 39196
rect 19576 39136 19640 39140
rect 19656 39196 19720 39200
rect 19656 39140 19660 39196
rect 19660 39140 19716 39196
rect 19716 39140 19720 39196
rect 19656 39136 19720 39140
rect 19736 39196 19800 39200
rect 19736 39140 19740 39196
rect 19740 39140 19796 39196
rect 19796 39140 19800 39196
rect 19736 39136 19800 39140
rect 19816 39196 19880 39200
rect 19816 39140 19820 39196
rect 19820 39140 19876 39196
rect 19876 39140 19880 39196
rect 19816 39136 19880 39140
rect 50296 39196 50360 39200
rect 50296 39140 50300 39196
rect 50300 39140 50356 39196
rect 50356 39140 50360 39196
rect 50296 39136 50360 39140
rect 50376 39196 50440 39200
rect 50376 39140 50380 39196
rect 50380 39140 50436 39196
rect 50436 39140 50440 39196
rect 50376 39136 50440 39140
rect 50456 39196 50520 39200
rect 50456 39140 50460 39196
rect 50460 39140 50516 39196
rect 50516 39140 50520 39196
rect 50456 39136 50520 39140
rect 50536 39196 50600 39200
rect 50536 39140 50540 39196
rect 50540 39140 50596 39196
rect 50596 39140 50600 39196
rect 50536 39136 50600 39140
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 65656 38652 65720 38656
rect 65656 38596 65660 38652
rect 65660 38596 65716 38652
rect 65716 38596 65720 38652
rect 65656 38592 65720 38596
rect 65736 38652 65800 38656
rect 65736 38596 65740 38652
rect 65740 38596 65796 38652
rect 65796 38596 65800 38652
rect 65736 38592 65800 38596
rect 65816 38652 65880 38656
rect 65816 38596 65820 38652
rect 65820 38596 65876 38652
rect 65876 38596 65880 38652
rect 65816 38592 65880 38596
rect 65896 38652 65960 38656
rect 65896 38596 65900 38652
rect 65900 38596 65956 38652
rect 65956 38596 65960 38652
rect 65896 38592 65960 38596
rect 19576 38108 19640 38112
rect 19576 38052 19580 38108
rect 19580 38052 19636 38108
rect 19636 38052 19640 38108
rect 19576 38048 19640 38052
rect 19656 38108 19720 38112
rect 19656 38052 19660 38108
rect 19660 38052 19716 38108
rect 19716 38052 19720 38108
rect 19656 38048 19720 38052
rect 19736 38108 19800 38112
rect 19736 38052 19740 38108
rect 19740 38052 19796 38108
rect 19796 38052 19800 38108
rect 19736 38048 19800 38052
rect 19816 38108 19880 38112
rect 19816 38052 19820 38108
rect 19820 38052 19876 38108
rect 19876 38052 19880 38108
rect 19816 38048 19880 38052
rect 50296 38108 50360 38112
rect 50296 38052 50300 38108
rect 50300 38052 50356 38108
rect 50356 38052 50360 38108
rect 50296 38048 50360 38052
rect 50376 38108 50440 38112
rect 50376 38052 50380 38108
rect 50380 38052 50436 38108
rect 50436 38052 50440 38108
rect 50376 38048 50440 38052
rect 50456 38108 50520 38112
rect 50456 38052 50460 38108
rect 50460 38052 50516 38108
rect 50516 38052 50520 38108
rect 50456 38048 50520 38052
rect 50536 38108 50600 38112
rect 50536 38052 50540 38108
rect 50540 38052 50596 38108
rect 50596 38052 50600 38108
rect 50536 38048 50600 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 65656 37564 65720 37568
rect 65656 37508 65660 37564
rect 65660 37508 65716 37564
rect 65716 37508 65720 37564
rect 65656 37504 65720 37508
rect 65736 37564 65800 37568
rect 65736 37508 65740 37564
rect 65740 37508 65796 37564
rect 65796 37508 65800 37564
rect 65736 37504 65800 37508
rect 65816 37564 65880 37568
rect 65816 37508 65820 37564
rect 65820 37508 65876 37564
rect 65876 37508 65880 37564
rect 65816 37504 65880 37508
rect 65896 37564 65960 37568
rect 65896 37508 65900 37564
rect 65900 37508 65956 37564
rect 65956 37508 65960 37564
rect 65896 37504 65960 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 50296 37020 50360 37024
rect 50296 36964 50300 37020
rect 50300 36964 50356 37020
rect 50356 36964 50360 37020
rect 50296 36960 50360 36964
rect 50376 37020 50440 37024
rect 50376 36964 50380 37020
rect 50380 36964 50436 37020
rect 50436 36964 50440 37020
rect 50376 36960 50440 36964
rect 50456 37020 50520 37024
rect 50456 36964 50460 37020
rect 50460 36964 50516 37020
rect 50516 36964 50520 37020
rect 50456 36960 50520 36964
rect 50536 37020 50600 37024
rect 50536 36964 50540 37020
rect 50540 36964 50596 37020
rect 50596 36964 50600 37020
rect 50536 36960 50600 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 65656 36476 65720 36480
rect 65656 36420 65660 36476
rect 65660 36420 65716 36476
rect 65716 36420 65720 36476
rect 65656 36416 65720 36420
rect 65736 36476 65800 36480
rect 65736 36420 65740 36476
rect 65740 36420 65796 36476
rect 65796 36420 65800 36476
rect 65736 36416 65800 36420
rect 65816 36476 65880 36480
rect 65816 36420 65820 36476
rect 65820 36420 65876 36476
rect 65876 36420 65880 36476
rect 65816 36416 65880 36420
rect 65896 36476 65960 36480
rect 65896 36420 65900 36476
rect 65900 36420 65956 36476
rect 65956 36420 65960 36476
rect 65896 36416 65960 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 50296 35932 50360 35936
rect 50296 35876 50300 35932
rect 50300 35876 50356 35932
rect 50356 35876 50360 35932
rect 50296 35872 50360 35876
rect 50376 35932 50440 35936
rect 50376 35876 50380 35932
rect 50380 35876 50436 35932
rect 50436 35876 50440 35932
rect 50376 35872 50440 35876
rect 50456 35932 50520 35936
rect 50456 35876 50460 35932
rect 50460 35876 50516 35932
rect 50516 35876 50520 35932
rect 50456 35872 50520 35876
rect 50536 35932 50600 35936
rect 50536 35876 50540 35932
rect 50540 35876 50596 35932
rect 50596 35876 50600 35932
rect 50536 35872 50600 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 65656 35388 65720 35392
rect 65656 35332 65660 35388
rect 65660 35332 65716 35388
rect 65716 35332 65720 35388
rect 65656 35328 65720 35332
rect 65736 35388 65800 35392
rect 65736 35332 65740 35388
rect 65740 35332 65796 35388
rect 65796 35332 65800 35388
rect 65736 35328 65800 35332
rect 65816 35388 65880 35392
rect 65816 35332 65820 35388
rect 65820 35332 65876 35388
rect 65876 35332 65880 35388
rect 65816 35328 65880 35332
rect 65896 35388 65960 35392
rect 65896 35332 65900 35388
rect 65900 35332 65956 35388
rect 65956 35332 65960 35388
rect 65896 35328 65960 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 50296 34844 50360 34848
rect 50296 34788 50300 34844
rect 50300 34788 50356 34844
rect 50356 34788 50360 34844
rect 50296 34784 50360 34788
rect 50376 34844 50440 34848
rect 50376 34788 50380 34844
rect 50380 34788 50436 34844
rect 50436 34788 50440 34844
rect 50376 34784 50440 34788
rect 50456 34844 50520 34848
rect 50456 34788 50460 34844
rect 50460 34788 50516 34844
rect 50516 34788 50520 34844
rect 50456 34784 50520 34788
rect 50536 34844 50600 34848
rect 50536 34788 50540 34844
rect 50540 34788 50596 34844
rect 50596 34788 50600 34844
rect 50536 34784 50600 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 65656 34300 65720 34304
rect 65656 34244 65660 34300
rect 65660 34244 65716 34300
rect 65716 34244 65720 34300
rect 65656 34240 65720 34244
rect 65736 34300 65800 34304
rect 65736 34244 65740 34300
rect 65740 34244 65796 34300
rect 65796 34244 65800 34300
rect 65736 34240 65800 34244
rect 65816 34300 65880 34304
rect 65816 34244 65820 34300
rect 65820 34244 65876 34300
rect 65876 34244 65880 34300
rect 65816 34240 65880 34244
rect 65896 34300 65960 34304
rect 65896 34244 65900 34300
rect 65900 34244 65956 34300
rect 65956 34244 65960 34300
rect 65896 34240 65960 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 50296 33756 50360 33760
rect 50296 33700 50300 33756
rect 50300 33700 50356 33756
rect 50356 33700 50360 33756
rect 50296 33696 50360 33700
rect 50376 33756 50440 33760
rect 50376 33700 50380 33756
rect 50380 33700 50436 33756
rect 50436 33700 50440 33756
rect 50376 33696 50440 33700
rect 50456 33756 50520 33760
rect 50456 33700 50460 33756
rect 50460 33700 50516 33756
rect 50516 33700 50520 33756
rect 50456 33696 50520 33700
rect 50536 33756 50600 33760
rect 50536 33700 50540 33756
rect 50540 33700 50596 33756
rect 50596 33700 50600 33756
rect 50536 33696 50600 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 65656 33212 65720 33216
rect 65656 33156 65660 33212
rect 65660 33156 65716 33212
rect 65716 33156 65720 33212
rect 65656 33152 65720 33156
rect 65736 33212 65800 33216
rect 65736 33156 65740 33212
rect 65740 33156 65796 33212
rect 65796 33156 65800 33212
rect 65736 33152 65800 33156
rect 65816 33212 65880 33216
rect 65816 33156 65820 33212
rect 65820 33156 65876 33212
rect 65876 33156 65880 33212
rect 65816 33152 65880 33156
rect 65896 33212 65960 33216
rect 65896 33156 65900 33212
rect 65900 33156 65956 33212
rect 65956 33156 65960 33212
rect 65896 33152 65960 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 50296 32668 50360 32672
rect 50296 32612 50300 32668
rect 50300 32612 50356 32668
rect 50356 32612 50360 32668
rect 50296 32608 50360 32612
rect 50376 32668 50440 32672
rect 50376 32612 50380 32668
rect 50380 32612 50436 32668
rect 50436 32612 50440 32668
rect 50376 32608 50440 32612
rect 50456 32668 50520 32672
rect 50456 32612 50460 32668
rect 50460 32612 50516 32668
rect 50516 32612 50520 32668
rect 50456 32608 50520 32612
rect 50536 32668 50600 32672
rect 50536 32612 50540 32668
rect 50540 32612 50596 32668
rect 50596 32612 50600 32668
rect 50536 32608 50600 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 65656 32124 65720 32128
rect 65656 32068 65660 32124
rect 65660 32068 65716 32124
rect 65716 32068 65720 32124
rect 65656 32064 65720 32068
rect 65736 32124 65800 32128
rect 65736 32068 65740 32124
rect 65740 32068 65796 32124
rect 65796 32068 65800 32124
rect 65736 32064 65800 32068
rect 65816 32124 65880 32128
rect 65816 32068 65820 32124
rect 65820 32068 65876 32124
rect 65876 32068 65880 32124
rect 65816 32064 65880 32068
rect 65896 32124 65960 32128
rect 65896 32068 65900 32124
rect 65900 32068 65956 32124
rect 65956 32068 65960 32124
rect 65896 32064 65960 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 50296 31580 50360 31584
rect 50296 31524 50300 31580
rect 50300 31524 50356 31580
rect 50356 31524 50360 31580
rect 50296 31520 50360 31524
rect 50376 31580 50440 31584
rect 50376 31524 50380 31580
rect 50380 31524 50436 31580
rect 50436 31524 50440 31580
rect 50376 31520 50440 31524
rect 50456 31580 50520 31584
rect 50456 31524 50460 31580
rect 50460 31524 50516 31580
rect 50516 31524 50520 31580
rect 50456 31520 50520 31524
rect 50536 31580 50600 31584
rect 50536 31524 50540 31580
rect 50540 31524 50596 31580
rect 50596 31524 50600 31580
rect 50536 31520 50600 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 65656 31036 65720 31040
rect 65656 30980 65660 31036
rect 65660 30980 65716 31036
rect 65716 30980 65720 31036
rect 65656 30976 65720 30980
rect 65736 31036 65800 31040
rect 65736 30980 65740 31036
rect 65740 30980 65796 31036
rect 65796 30980 65800 31036
rect 65736 30976 65800 30980
rect 65816 31036 65880 31040
rect 65816 30980 65820 31036
rect 65820 30980 65876 31036
rect 65876 30980 65880 31036
rect 65816 30976 65880 30980
rect 65896 31036 65960 31040
rect 65896 30980 65900 31036
rect 65900 30980 65956 31036
rect 65956 30980 65960 31036
rect 65896 30976 65960 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 50296 30492 50360 30496
rect 50296 30436 50300 30492
rect 50300 30436 50356 30492
rect 50356 30436 50360 30492
rect 50296 30432 50360 30436
rect 50376 30492 50440 30496
rect 50376 30436 50380 30492
rect 50380 30436 50436 30492
rect 50436 30436 50440 30492
rect 50376 30432 50440 30436
rect 50456 30492 50520 30496
rect 50456 30436 50460 30492
rect 50460 30436 50516 30492
rect 50516 30436 50520 30492
rect 50456 30432 50520 30436
rect 50536 30492 50600 30496
rect 50536 30436 50540 30492
rect 50540 30436 50596 30492
rect 50596 30436 50600 30492
rect 50536 30432 50600 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 65656 29948 65720 29952
rect 65656 29892 65660 29948
rect 65660 29892 65716 29948
rect 65716 29892 65720 29948
rect 65656 29888 65720 29892
rect 65736 29948 65800 29952
rect 65736 29892 65740 29948
rect 65740 29892 65796 29948
rect 65796 29892 65800 29948
rect 65736 29888 65800 29892
rect 65816 29948 65880 29952
rect 65816 29892 65820 29948
rect 65820 29892 65876 29948
rect 65876 29892 65880 29948
rect 65816 29888 65880 29892
rect 65896 29948 65960 29952
rect 65896 29892 65900 29948
rect 65900 29892 65956 29948
rect 65956 29892 65960 29948
rect 65896 29888 65960 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 50296 29404 50360 29408
rect 50296 29348 50300 29404
rect 50300 29348 50356 29404
rect 50356 29348 50360 29404
rect 50296 29344 50360 29348
rect 50376 29404 50440 29408
rect 50376 29348 50380 29404
rect 50380 29348 50436 29404
rect 50436 29348 50440 29404
rect 50376 29344 50440 29348
rect 50456 29404 50520 29408
rect 50456 29348 50460 29404
rect 50460 29348 50516 29404
rect 50516 29348 50520 29404
rect 50456 29344 50520 29348
rect 50536 29404 50600 29408
rect 50536 29348 50540 29404
rect 50540 29348 50596 29404
rect 50596 29348 50600 29404
rect 50536 29344 50600 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 65656 28860 65720 28864
rect 65656 28804 65660 28860
rect 65660 28804 65716 28860
rect 65716 28804 65720 28860
rect 65656 28800 65720 28804
rect 65736 28860 65800 28864
rect 65736 28804 65740 28860
rect 65740 28804 65796 28860
rect 65796 28804 65800 28860
rect 65736 28800 65800 28804
rect 65816 28860 65880 28864
rect 65816 28804 65820 28860
rect 65820 28804 65876 28860
rect 65876 28804 65880 28860
rect 65816 28800 65880 28804
rect 65896 28860 65960 28864
rect 65896 28804 65900 28860
rect 65900 28804 65956 28860
rect 65956 28804 65960 28860
rect 65896 28800 65960 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 50296 28316 50360 28320
rect 50296 28260 50300 28316
rect 50300 28260 50356 28316
rect 50356 28260 50360 28316
rect 50296 28256 50360 28260
rect 50376 28316 50440 28320
rect 50376 28260 50380 28316
rect 50380 28260 50436 28316
rect 50436 28260 50440 28316
rect 50376 28256 50440 28260
rect 50456 28316 50520 28320
rect 50456 28260 50460 28316
rect 50460 28260 50516 28316
rect 50516 28260 50520 28316
rect 50456 28256 50520 28260
rect 50536 28316 50600 28320
rect 50536 28260 50540 28316
rect 50540 28260 50596 28316
rect 50596 28260 50600 28316
rect 50536 28256 50600 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 65656 27772 65720 27776
rect 65656 27716 65660 27772
rect 65660 27716 65716 27772
rect 65716 27716 65720 27772
rect 65656 27712 65720 27716
rect 65736 27772 65800 27776
rect 65736 27716 65740 27772
rect 65740 27716 65796 27772
rect 65796 27716 65800 27772
rect 65736 27712 65800 27716
rect 65816 27772 65880 27776
rect 65816 27716 65820 27772
rect 65820 27716 65876 27772
rect 65876 27716 65880 27772
rect 65816 27712 65880 27716
rect 65896 27772 65960 27776
rect 65896 27716 65900 27772
rect 65900 27716 65956 27772
rect 65956 27716 65960 27772
rect 65896 27712 65960 27716
rect 23428 27704 23492 27708
rect 23428 27648 23478 27704
rect 23478 27648 23492 27704
rect 23428 27644 23492 27648
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 50296 27228 50360 27232
rect 50296 27172 50300 27228
rect 50300 27172 50356 27228
rect 50356 27172 50360 27228
rect 50296 27168 50360 27172
rect 50376 27228 50440 27232
rect 50376 27172 50380 27228
rect 50380 27172 50436 27228
rect 50436 27172 50440 27228
rect 50376 27168 50440 27172
rect 50456 27228 50520 27232
rect 50456 27172 50460 27228
rect 50460 27172 50516 27228
rect 50516 27172 50520 27228
rect 50456 27168 50520 27172
rect 50536 27228 50600 27232
rect 50536 27172 50540 27228
rect 50540 27172 50596 27228
rect 50596 27172 50600 27228
rect 50536 27168 50600 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 65656 26684 65720 26688
rect 65656 26628 65660 26684
rect 65660 26628 65716 26684
rect 65716 26628 65720 26684
rect 65656 26624 65720 26628
rect 65736 26684 65800 26688
rect 65736 26628 65740 26684
rect 65740 26628 65796 26684
rect 65796 26628 65800 26684
rect 65736 26624 65800 26628
rect 65816 26684 65880 26688
rect 65816 26628 65820 26684
rect 65820 26628 65876 26684
rect 65876 26628 65880 26684
rect 65816 26624 65880 26628
rect 65896 26684 65960 26688
rect 65896 26628 65900 26684
rect 65900 26628 65956 26684
rect 65956 26628 65960 26684
rect 65896 26624 65960 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 50296 26140 50360 26144
rect 50296 26084 50300 26140
rect 50300 26084 50356 26140
rect 50356 26084 50360 26140
rect 50296 26080 50360 26084
rect 50376 26140 50440 26144
rect 50376 26084 50380 26140
rect 50380 26084 50436 26140
rect 50436 26084 50440 26140
rect 50376 26080 50440 26084
rect 50456 26140 50520 26144
rect 50456 26084 50460 26140
rect 50460 26084 50516 26140
rect 50516 26084 50520 26140
rect 50456 26080 50520 26084
rect 50536 26140 50600 26144
rect 50536 26084 50540 26140
rect 50540 26084 50596 26140
rect 50596 26084 50600 26140
rect 50536 26080 50600 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 65656 25596 65720 25600
rect 65656 25540 65660 25596
rect 65660 25540 65716 25596
rect 65716 25540 65720 25596
rect 65656 25536 65720 25540
rect 65736 25596 65800 25600
rect 65736 25540 65740 25596
rect 65740 25540 65796 25596
rect 65796 25540 65800 25596
rect 65736 25536 65800 25540
rect 65816 25596 65880 25600
rect 65816 25540 65820 25596
rect 65820 25540 65876 25596
rect 65876 25540 65880 25596
rect 65816 25536 65880 25540
rect 65896 25596 65960 25600
rect 65896 25540 65900 25596
rect 65900 25540 65956 25596
rect 65956 25540 65960 25596
rect 65896 25536 65960 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 50296 25052 50360 25056
rect 50296 24996 50300 25052
rect 50300 24996 50356 25052
rect 50356 24996 50360 25052
rect 50296 24992 50360 24996
rect 50376 25052 50440 25056
rect 50376 24996 50380 25052
rect 50380 24996 50436 25052
rect 50436 24996 50440 25052
rect 50376 24992 50440 24996
rect 50456 25052 50520 25056
rect 50456 24996 50460 25052
rect 50460 24996 50516 25052
rect 50516 24996 50520 25052
rect 50456 24992 50520 24996
rect 50536 25052 50600 25056
rect 50536 24996 50540 25052
rect 50540 24996 50596 25052
rect 50596 24996 50600 25052
rect 50536 24992 50600 24996
rect 23428 24712 23492 24716
rect 23428 24656 23442 24712
rect 23442 24656 23492 24712
rect 23428 24652 23492 24656
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 65656 24508 65720 24512
rect 65656 24452 65660 24508
rect 65660 24452 65716 24508
rect 65716 24452 65720 24508
rect 65656 24448 65720 24452
rect 65736 24508 65800 24512
rect 65736 24452 65740 24508
rect 65740 24452 65796 24508
rect 65796 24452 65800 24508
rect 65736 24448 65800 24452
rect 65816 24508 65880 24512
rect 65816 24452 65820 24508
rect 65820 24452 65876 24508
rect 65876 24452 65880 24508
rect 65816 24448 65880 24452
rect 65896 24508 65960 24512
rect 65896 24452 65900 24508
rect 65900 24452 65956 24508
rect 65956 24452 65960 24508
rect 65896 24448 65960 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 50296 23964 50360 23968
rect 50296 23908 50300 23964
rect 50300 23908 50356 23964
rect 50356 23908 50360 23964
rect 50296 23904 50360 23908
rect 50376 23964 50440 23968
rect 50376 23908 50380 23964
rect 50380 23908 50436 23964
rect 50436 23908 50440 23964
rect 50376 23904 50440 23908
rect 50456 23964 50520 23968
rect 50456 23908 50460 23964
rect 50460 23908 50516 23964
rect 50516 23908 50520 23964
rect 50456 23904 50520 23908
rect 50536 23964 50600 23968
rect 50536 23908 50540 23964
rect 50540 23908 50596 23964
rect 50596 23908 50600 23964
rect 50536 23904 50600 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 65656 23420 65720 23424
rect 65656 23364 65660 23420
rect 65660 23364 65716 23420
rect 65716 23364 65720 23420
rect 65656 23360 65720 23364
rect 65736 23420 65800 23424
rect 65736 23364 65740 23420
rect 65740 23364 65796 23420
rect 65796 23364 65800 23420
rect 65736 23360 65800 23364
rect 65816 23420 65880 23424
rect 65816 23364 65820 23420
rect 65820 23364 65876 23420
rect 65876 23364 65880 23420
rect 65816 23360 65880 23364
rect 65896 23420 65960 23424
rect 65896 23364 65900 23420
rect 65900 23364 65956 23420
rect 65956 23364 65960 23420
rect 65896 23360 65960 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 50296 22876 50360 22880
rect 50296 22820 50300 22876
rect 50300 22820 50356 22876
rect 50356 22820 50360 22876
rect 50296 22816 50360 22820
rect 50376 22876 50440 22880
rect 50376 22820 50380 22876
rect 50380 22820 50436 22876
rect 50436 22820 50440 22876
rect 50376 22816 50440 22820
rect 50456 22876 50520 22880
rect 50456 22820 50460 22876
rect 50460 22820 50516 22876
rect 50516 22820 50520 22876
rect 50456 22816 50520 22820
rect 50536 22876 50600 22880
rect 50536 22820 50540 22876
rect 50540 22820 50596 22876
rect 50596 22820 50600 22876
rect 50536 22816 50600 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 65656 22332 65720 22336
rect 65656 22276 65660 22332
rect 65660 22276 65716 22332
rect 65716 22276 65720 22332
rect 65656 22272 65720 22276
rect 65736 22332 65800 22336
rect 65736 22276 65740 22332
rect 65740 22276 65796 22332
rect 65796 22276 65800 22332
rect 65736 22272 65800 22276
rect 65816 22332 65880 22336
rect 65816 22276 65820 22332
rect 65820 22276 65876 22332
rect 65876 22276 65880 22332
rect 65816 22272 65880 22276
rect 65896 22332 65960 22336
rect 65896 22276 65900 22332
rect 65900 22276 65956 22332
rect 65956 22276 65960 22332
rect 65896 22272 65960 22276
rect 23612 22264 23676 22268
rect 23612 22208 23626 22264
rect 23626 22208 23676 22264
rect 23612 22204 23676 22208
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 50296 21788 50360 21792
rect 50296 21732 50300 21788
rect 50300 21732 50356 21788
rect 50356 21732 50360 21788
rect 50296 21728 50360 21732
rect 50376 21788 50440 21792
rect 50376 21732 50380 21788
rect 50380 21732 50436 21788
rect 50436 21732 50440 21788
rect 50376 21728 50440 21732
rect 50456 21788 50520 21792
rect 50456 21732 50460 21788
rect 50460 21732 50516 21788
rect 50516 21732 50520 21788
rect 50456 21728 50520 21732
rect 50536 21788 50600 21792
rect 50536 21732 50540 21788
rect 50540 21732 50596 21788
rect 50596 21732 50600 21788
rect 50536 21728 50600 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 65656 21244 65720 21248
rect 65656 21188 65660 21244
rect 65660 21188 65716 21244
rect 65716 21188 65720 21244
rect 65656 21184 65720 21188
rect 65736 21244 65800 21248
rect 65736 21188 65740 21244
rect 65740 21188 65796 21244
rect 65796 21188 65800 21244
rect 65736 21184 65800 21188
rect 65816 21244 65880 21248
rect 65816 21188 65820 21244
rect 65820 21188 65876 21244
rect 65876 21188 65880 21244
rect 65816 21184 65880 21188
rect 65896 21244 65960 21248
rect 65896 21188 65900 21244
rect 65900 21188 65956 21244
rect 65956 21188 65960 21244
rect 65896 21184 65960 21188
rect 24164 20708 24228 20772
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 50296 20700 50360 20704
rect 50296 20644 50300 20700
rect 50300 20644 50356 20700
rect 50356 20644 50360 20700
rect 50296 20640 50360 20644
rect 50376 20700 50440 20704
rect 50376 20644 50380 20700
rect 50380 20644 50436 20700
rect 50436 20644 50440 20700
rect 50376 20640 50440 20644
rect 50456 20700 50520 20704
rect 50456 20644 50460 20700
rect 50460 20644 50516 20700
rect 50516 20644 50520 20700
rect 50456 20640 50520 20644
rect 50536 20700 50600 20704
rect 50536 20644 50540 20700
rect 50540 20644 50596 20700
rect 50596 20644 50600 20700
rect 50536 20640 50600 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 65656 20156 65720 20160
rect 65656 20100 65660 20156
rect 65660 20100 65716 20156
rect 65716 20100 65720 20156
rect 65656 20096 65720 20100
rect 65736 20156 65800 20160
rect 65736 20100 65740 20156
rect 65740 20100 65796 20156
rect 65796 20100 65800 20156
rect 65736 20096 65800 20100
rect 65816 20156 65880 20160
rect 65816 20100 65820 20156
rect 65820 20100 65876 20156
rect 65876 20100 65880 20156
rect 65816 20096 65880 20100
rect 65896 20156 65960 20160
rect 65896 20100 65900 20156
rect 65900 20100 65956 20156
rect 65956 20100 65960 20156
rect 65896 20096 65960 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 50296 19612 50360 19616
rect 50296 19556 50300 19612
rect 50300 19556 50356 19612
rect 50356 19556 50360 19612
rect 50296 19552 50360 19556
rect 50376 19612 50440 19616
rect 50376 19556 50380 19612
rect 50380 19556 50436 19612
rect 50436 19556 50440 19612
rect 50376 19552 50440 19556
rect 50456 19612 50520 19616
rect 50456 19556 50460 19612
rect 50460 19556 50516 19612
rect 50516 19556 50520 19612
rect 50456 19552 50520 19556
rect 50536 19612 50600 19616
rect 50536 19556 50540 19612
rect 50540 19556 50596 19612
rect 50596 19556 50600 19612
rect 50536 19552 50600 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 65656 19068 65720 19072
rect 65656 19012 65660 19068
rect 65660 19012 65716 19068
rect 65716 19012 65720 19068
rect 65656 19008 65720 19012
rect 65736 19068 65800 19072
rect 65736 19012 65740 19068
rect 65740 19012 65796 19068
rect 65796 19012 65800 19068
rect 65736 19008 65800 19012
rect 65816 19068 65880 19072
rect 65816 19012 65820 19068
rect 65820 19012 65876 19068
rect 65876 19012 65880 19068
rect 65816 19008 65880 19012
rect 65896 19068 65960 19072
rect 65896 19012 65900 19068
rect 65900 19012 65956 19068
rect 65956 19012 65960 19068
rect 65896 19008 65960 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 50296 18524 50360 18528
rect 50296 18468 50300 18524
rect 50300 18468 50356 18524
rect 50356 18468 50360 18524
rect 50296 18464 50360 18468
rect 50376 18524 50440 18528
rect 50376 18468 50380 18524
rect 50380 18468 50436 18524
rect 50436 18468 50440 18524
rect 50376 18464 50440 18468
rect 50456 18524 50520 18528
rect 50456 18468 50460 18524
rect 50460 18468 50516 18524
rect 50516 18468 50520 18524
rect 50456 18464 50520 18468
rect 50536 18524 50600 18528
rect 50536 18468 50540 18524
rect 50540 18468 50596 18524
rect 50596 18468 50600 18524
rect 50536 18464 50600 18468
rect 21956 18184 22020 18188
rect 21956 18128 22006 18184
rect 22006 18128 22020 18184
rect 21956 18124 22020 18128
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 65656 17980 65720 17984
rect 65656 17924 65660 17980
rect 65660 17924 65716 17980
rect 65716 17924 65720 17980
rect 65656 17920 65720 17924
rect 65736 17980 65800 17984
rect 65736 17924 65740 17980
rect 65740 17924 65796 17980
rect 65796 17924 65800 17980
rect 65736 17920 65800 17924
rect 65816 17980 65880 17984
rect 65816 17924 65820 17980
rect 65820 17924 65876 17980
rect 65876 17924 65880 17980
rect 65816 17920 65880 17924
rect 65896 17980 65960 17984
rect 65896 17924 65900 17980
rect 65900 17924 65956 17980
rect 65956 17924 65960 17980
rect 65896 17920 65960 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 50296 17436 50360 17440
rect 50296 17380 50300 17436
rect 50300 17380 50356 17436
rect 50356 17380 50360 17436
rect 50296 17376 50360 17380
rect 50376 17436 50440 17440
rect 50376 17380 50380 17436
rect 50380 17380 50436 17436
rect 50436 17380 50440 17436
rect 50376 17376 50440 17380
rect 50456 17436 50520 17440
rect 50456 17380 50460 17436
rect 50460 17380 50516 17436
rect 50516 17380 50520 17436
rect 50456 17376 50520 17380
rect 50536 17436 50600 17440
rect 50536 17380 50540 17436
rect 50540 17380 50596 17436
rect 50596 17380 50600 17436
rect 50536 17376 50600 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 65656 16892 65720 16896
rect 65656 16836 65660 16892
rect 65660 16836 65716 16892
rect 65716 16836 65720 16892
rect 65656 16832 65720 16836
rect 65736 16892 65800 16896
rect 65736 16836 65740 16892
rect 65740 16836 65796 16892
rect 65796 16836 65800 16892
rect 65736 16832 65800 16836
rect 65816 16892 65880 16896
rect 65816 16836 65820 16892
rect 65820 16836 65876 16892
rect 65876 16836 65880 16892
rect 65816 16832 65880 16836
rect 65896 16892 65960 16896
rect 65896 16836 65900 16892
rect 65900 16836 65956 16892
rect 65956 16836 65960 16892
rect 65896 16832 65960 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 50296 16348 50360 16352
rect 50296 16292 50300 16348
rect 50300 16292 50356 16348
rect 50356 16292 50360 16348
rect 50296 16288 50360 16292
rect 50376 16348 50440 16352
rect 50376 16292 50380 16348
rect 50380 16292 50436 16348
rect 50436 16292 50440 16348
rect 50376 16288 50440 16292
rect 50456 16348 50520 16352
rect 50456 16292 50460 16348
rect 50460 16292 50516 16348
rect 50516 16292 50520 16348
rect 50456 16288 50520 16292
rect 50536 16348 50600 16352
rect 50536 16292 50540 16348
rect 50540 16292 50596 16348
rect 50596 16292 50600 16348
rect 50536 16288 50600 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 65656 15804 65720 15808
rect 65656 15748 65660 15804
rect 65660 15748 65716 15804
rect 65716 15748 65720 15804
rect 65656 15744 65720 15748
rect 65736 15804 65800 15808
rect 65736 15748 65740 15804
rect 65740 15748 65796 15804
rect 65796 15748 65800 15804
rect 65736 15744 65800 15748
rect 65816 15804 65880 15808
rect 65816 15748 65820 15804
rect 65820 15748 65876 15804
rect 65876 15748 65880 15804
rect 65816 15744 65880 15748
rect 65896 15804 65960 15808
rect 65896 15748 65900 15804
rect 65900 15748 65956 15804
rect 65956 15748 65960 15804
rect 65896 15744 65960 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 50296 15260 50360 15264
rect 50296 15204 50300 15260
rect 50300 15204 50356 15260
rect 50356 15204 50360 15260
rect 50296 15200 50360 15204
rect 50376 15260 50440 15264
rect 50376 15204 50380 15260
rect 50380 15204 50436 15260
rect 50436 15204 50440 15260
rect 50376 15200 50440 15204
rect 50456 15260 50520 15264
rect 50456 15204 50460 15260
rect 50460 15204 50516 15260
rect 50516 15204 50520 15260
rect 50456 15200 50520 15204
rect 50536 15260 50600 15264
rect 50536 15204 50540 15260
rect 50540 15204 50596 15260
rect 50596 15204 50600 15260
rect 50536 15200 50600 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 65656 14716 65720 14720
rect 65656 14660 65660 14716
rect 65660 14660 65716 14716
rect 65716 14660 65720 14716
rect 65656 14656 65720 14660
rect 65736 14716 65800 14720
rect 65736 14660 65740 14716
rect 65740 14660 65796 14716
rect 65796 14660 65800 14716
rect 65736 14656 65800 14660
rect 65816 14716 65880 14720
rect 65816 14660 65820 14716
rect 65820 14660 65876 14716
rect 65876 14660 65880 14716
rect 65816 14656 65880 14660
rect 65896 14716 65960 14720
rect 65896 14660 65900 14716
rect 65900 14660 65956 14716
rect 65956 14660 65960 14716
rect 65896 14656 65960 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 50296 14172 50360 14176
rect 50296 14116 50300 14172
rect 50300 14116 50356 14172
rect 50356 14116 50360 14172
rect 50296 14112 50360 14116
rect 50376 14172 50440 14176
rect 50376 14116 50380 14172
rect 50380 14116 50436 14172
rect 50436 14116 50440 14172
rect 50376 14112 50440 14116
rect 50456 14172 50520 14176
rect 50456 14116 50460 14172
rect 50460 14116 50516 14172
rect 50516 14116 50520 14172
rect 50456 14112 50520 14116
rect 50536 14172 50600 14176
rect 50536 14116 50540 14172
rect 50540 14116 50596 14172
rect 50596 14116 50600 14172
rect 50536 14112 50600 14116
rect 35572 14104 35636 14108
rect 35572 14048 35586 14104
rect 35586 14048 35636 14104
rect 35572 14044 35636 14048
rect 19380 13772 19444 13836
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 65656 13628 65720 13632
rect 65656 13572 65660 13628
rect 65660 13572 65716 13628
rect 65716 13572 65720 13628
rect 65656 13568 65720 13572
rect 65736 13628 65800 13632
rect 65736 13572 65740 13628
rect 65740 13572 65796 13628
rect 65796 13572 65800 13628
rect 65736 13568 65800 13572
rect 65816 13628 65880 13632
rect 65816 13572 65820 13628
rect 65820 13572 65876 13628
rect 65876 13572 65880 13628
rect 65816 13568 65880 13572
rect 65896 13628 65960 13632
rect 65896 13572 65900 13628
rect 65900 13572 65956 13628
rect 65956 13572 65960 13628
rect 65896 13568 65960 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 50296 13084 50360 13088
rect 50296 13028 50300 13084
rect 50300 13028 50356 13084
rect 50356 13028 50360 13084
rect 50296 13024 50360 13028
rect 50376 13084 50440 13088
rect 50376 13028 50380 13084
rect 50380 13028 50436 13084
rect 50436 13028 50440 13084
rect 50376 13024 50440 13028
rect 50456 13084 50520 13088
rect 50456 13028 50460 13084
rect 50460 13028 50516 13084
rect 50516 13028 50520 13084
rect 50456 13024 50520 13028
rect 50536 13084 50600 13088
rect 50536 13028 50540 13084
rect 50540 13028 50596 13084
rect 50596 13028 50600 13084
rect 50536 13024 50600 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 65656 12540 65720 12544
rect 65656 12484 65660 12540
rect 65660 12484 65716 12540
rect 65716 12484 65720 12540
rect 65656 12480 65720 12484
rect 65736 12540 65800 12544
rect 65736 12484 65740 12540
rect 65740 12484 65796 12540
rect 65796 12484 65800 12540
rect 65736 12480 65800 12484
rect 65816 12540 65880 12544
rect 65816 12484 65820 12540
rect 65820 12484 65876 12540
rect 65876 12484 65880 12540
rect 65816 12480 65880 12484
rect 65896 12540 65960 12544
rect 65896 12484 65900 12540
rect 65900 12484 65956 12540
rect 65956 12484 65960 12540
rect 65896 12480 65960 12484
rect 17908 12064 17972 12068
rect 17908 12008 17922 12064
rect 17922 12008 17972 12064
rect 17908 12004 17972 12008
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 50296 11996 50360 12000
rect 50296 11940 50300 11996
rect 50300 11940 50356 11996
rect 50356 11940 50360 11996
rect 50296 11936 50360 11940
rect 50376 11996 50440 12000
rect 50376 11940 50380 11996
rect 50380 11940 50436 11996
rect 50436 11940 50440 11996
rect 50376 11936 50440 11940
rect 50456 11996 50520 12000
rect 50456 11940 50460 11996
rect 50460 11940 50516 11996
rect 50516 11940 50520 11996
rect 50456 11936 50520 11940
rect 50536 11996 50600 12000
rect 50536 11940 50540 11996
rect 50540 11940 50596 11996
rect 50596 11940 50600 11996
rect 50536 11936 50600 11940
rect 35572 11928 35636 11932
rect 35572 11872 35622 11928
rect 35622 11872 35636 11928
rect 35572 11868 35636 11872
rect 11100 11520 11164 11524
rect 11100 11464 11114 11520
rect 11114 11464 11164 11520
rect 11100 11460 11164 11464
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 65656 11452 65720 11456
rect 65656 11396 65660 11452
rect 65660 11396 65716 11452
rect 65716 11396 65720 11452
rect 65656 11392 65720 11396
rect 65736 11452 65800 11456
rect 65736 11396 65740 11452
rect 65740 11396 65796 11452
rect 65796 11396 65800 11452
rect 65736 11392 65800 11396
rect 65816 11452 65880 11456
rect 65816 11396 65820 11452
rect 65820 11396 65876 11452
rect 65876 11396 65880 11452
rect 65816 11392 65880 11396
rect 65896 11452 65960 11456
rect 65896 11396 65900 11452
rect 65900 11396 65956 11452
rect 65956 11396 65960 11452
rect 65896 11392 65960 11396
rect 23612 11324 23676 11388
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 50296 10908 50360 10912
rect 50296 10852 50300 10908
rect 50300 10852 50356 10908
rect 50356 10852 50360 10908
rect 50296 10848 50360 10852
rect 50376 10908 50440 10912
rect 50376 10852 50380 10908
rect 50380 10852 50436 10908
rect 50436 10852 50440 10908
rect 50376 10848 50440 10852
rect 50456 10908 50520 10912
rect 50456 10852 50460 10908
rect 50460 10852 50516 10908
rect 50516 10852 50520 10908
rect 50456 10848 50520 10852
rect 50536 10908 50600 10912
rect 50536 10852 50540 10908
rect 50540 10852 50596 10908
rect 50596 10852 50600 10908
rect 50536 10848 50600 10852
rect 21956 10644 22020 10708
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 65656 10364 65720 10368
rect 65656 10308 65660 10364
rect 65660 10308 65716 10364
rect 65716 10308 65720 10364
rect 65656 10304 65720 10308
rect 65736 10364 65800 10368
rect 65736 10308 65740 10364
rect 65740 10308 65796 10364
rect 65796 10308 65800 10364
rect 65736 10304 65800 10308
rect 65816 10364 65880 10368
rect 65816 10308 65820 10364
rect 65820 10308 65876 10364
rect 65876 10308 65880 10364
rect 65816 10304 65880 10308
rect 65896 10364 65960 10368
rect 65896 10308 65900 10364
rect 65900 10308 65956 10364
rect 65956 10308 65960 10364
rect 65896 10304 65960 10308
rect 10732 10236 10796 10300
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 50296 9820 50360 9824
rect 50296 9764 50300 9820
rect 50300 9764 50356 9820
rect 50356 9764 50360 9820
rect 50296 9760 50360 9764
rect 50376 9820 50440 9824
rect 50376 9764 50380 9820
rect 50380 9764 50436 9820
rect 50436 9764 50440 9820
rect 50376 9760 50440 9764
rect 50456 9820 50520 9824
rect 50456 9764 50460 9820
rect 50460 9764 50516 9820
rect 50516 9764 50520 9820
rect 50456 9760 50520 9764
rect 50536 9820 50600 9824
rect 50536 9764 50540 9820
rect 50540 9764 50596 9820
rect 50596 9764 50600 9820
rect 50536 9760 50600 9764
rect 24164 9556 24228 9620
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 65656 9276 65720 9280
rect 65656 9220 65660 9276
rect 65660 9220 65716 9276
rect 65716 9220 65720 9276
rect 65656 9216 65720 9220
rect 65736 9276 65800 9280
rect 65736 9220 65740 9276
rect 65740 9220 65796 9276
rect 65796 9220 65800 9276
rect 65736 9216 65800 9220
rect 65816 9276 65880 9280
rect 65816 9220 65820 9276
rect 65820 9220 65876 9276
rect 65876 9220 65880 9276
rect 65816 9216 65880 9220
rect 65896 9276 65960 9280
rect 65896 9220 65900 9276
rect 65900 9220 65956 9276
rect 65956 9220 65960 9276
rect 65896 9216 65960 9220
rect 12020 8740 12084 8804
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 50296 8732 50360 8736
rect 50296 8676 50300 8732
rect 50300 8676 50356 8732
rect 50356 8676 50360 8732
rect 50296 8672 50360 8676
rect 50376 8732 50440 8736
rect 50376 8676 50380 8732
rect 50380 8676 50436 8732
rect 50436 8676 50440 8732
rect 50376 8672 50440 8676
rect 50456 8732 50520 8736
rect 50456 8676 50460 8732
rect 50460 8676 50516 8732
rect 50516 8676 50520 8732
rect 50456 8672 50520 8676
rect 50536 8732 50600 8736
rect 50536 8676 50540 8732
rect 50540 8676 50596 8732
rect 50596 8676 50600 8732
rect 50536 8672 50600 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 65656 8188 65720 8192
rect 65656 8132 65660 8188
rect 65660 8132 65716 8188
rect 65716 8132 65720 8188
rect 65656 8128 65720 8132
rect 65736 8188 65800 8192
rect 65736 8132 65740 8188
rect 65740 8132 65796 8188
rect 65796 8132 65800 8188
rect 65736 8128 65800 8132
rect 65816 8188 65880 8192
rect 65816 8132 65820 8188
rect 65820 8132 65876 8188
rect 65876 8132 65880 8188
rect 65816 8128 65880 8132
rect 65896 8188 65960 8192
rect 65896 8132 65900 8188
rect 65900 8132 65956 8188
rect 65956 8132 65960 8188
rect 65896 8128 65960 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 50296 7644 50360 7648
rect 50296 7588 50300 7644
rect 50300 7588 50356 7644
rect 50356 7588 50360 7644
rect 50296 7584 50360 7588
rect 50376 7644 50440 7648
rect 50376 7588 50380 7644
rect 50380 7588 50436 7644
rect 50436 7588 50440 7644
rect 50376 7584 50440 7588
rect 50456 7644 50520 7648
rect 50456 7588 50460 7644
rect 50460 7588 50516 7644
rect 50516 7588 50520 7644
rect 50456 7584 50520 7588
rect 50536 7644 50600 7648
rect 50536 7588 50540 7644
rect 50540 7588 50596 7644
rect 50596 7588 50600 7644
rect 50536 7584 50600 7588
rect 19380 7380 19444 7444
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 65656 7100 65720 7104
rect 65656 7044 65660 7100
rect 65660 7044 65716 7100
rect 65716 7044 65720 7100
rect 65656 7040 65720 7044
rect 65736 7100 65800 7104
rect 65736 7044 65740 7100
rect 65740 7044 65796 7100
rect 65796 7044 65800 7100
rect 65736 7040 65800 7044
rect 65816 7100 65880 7104
rect 65816 7044 65820 7100
rect 65820 7044 65876 7100
rect 65876 7044 65880 7100
rect 65816 7040 65880 7044
rect 65896 7100 65960 7104
rect 65896 7044 65900 7100
rect 65900 7044 65956 7100
rect 65956 7044 65960 7100
rect 65896 7040 65960 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 50296 6556 50360 6560
rect 50296 6500 50300 6556
rect 50300 6500 50356 6556
rect 50356 6500 50360 6556
rect 50296 6496 50360 6500
rect 50376 6556 50440 6560
rect 50376 6500 50380 6556
rect 50380 6500 50436 6556
rect 50436 6500 50440 6556
rect 50376 6496 50440 6500
rect 50456 6556 50520 6560
rect 50456 6500 50460 6556
rect 50460 6500 50516 6556
rect 50516 6500 50520 6556
rect 50456 6496 50520 6500
rect 50536 6556 50600 6560
rect 50536 6500 50540 6556
rect 50540 6500 50596 6556
rect 50596 6500 50600 6556
rect 50536 6496 50600 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 65656 6012 65720 6016
rect 65656 5956 65660 6012
rect 65660 5956 65716 6012
rect 65716 5956 65720 6012
rect 65656 5952 65720 5956
rect 65736 6012 65800 6016
rect 65736 5956 65740 6012
rect 65740 5956 65796 6012
rect 65796 5956 65800 6012
rect 65736 5952 65800 5956
rect 65816 6012 65880 6016
rect 65816 5956 65820 6012
rect 65820 5956 65876 6012
rect 65876 5956 65880 6012
rect 65816 5952 65880 5956
rect 65896 6012 65960 6016
rect 65896 5956 65900 6012
rect 65900 5956 65956 6012
rect 65956 5956 65960 6012
rect 65896 5952 65960 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 50296 5468 50360 5472
rect 50296 5412 50300 5468
rect 50300 5412 50356 5468
rect 50356 5412 50360 5468
rect 50296 5408 50360 5412
rect 50376 5468 50440 5472
rect 50376 5412 50380 5468
rect 50380 5412 50436 5468
rect 50436 5412 50440 5468
rect 50376 5408 50440 5412
rect 50456 5468 50520 5472
rect 50456 5412 50460 5468
rect 50460 5412 50516 5468
rect 50516 5412 50520 5468
rect 50456 5408 50520 5412
rect 50536 5468 50600 5472
rect 50536 5412 50540 5468
rect 50540 5412 50596 5468
rect 50596 5412 50600 5468
rect 50536 5408 50600 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 65656 4924 65720 4928
rect 65656 4868 65660 4924
rect 65660 4868 65716 4924
rect 65716 4868 65720 4924
rect 65656 4864 65720 4868
rect 65736 4924 65800 4928
rect 65736 4868 65740 4924
rect 65740 4868 65796 4924
rect 65796 4868 65800 4924
rect 65736 4864 65800 4868
rect 65816 4924 65880 4928
rect 65816 4868 65820 4924
rect 65820 4868 65876 4924
rect 65876 4868 65880 4924
rect 65816 4864 65880 4868
rect 65896 4924 65960 4928
rect 65896 4868 65900 4924
rect 65900 4868 65956 4924
rect 65956 4868 65960 4924
rect 65896 4864 65960 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 50296 4380 50360 4384
rect 50296 4324 50300 4380
rect 50300 4324 50356 4380
rect 50356 4324 50360 4380
rect 50296 4320 50360 4324
rect 50376 4380 50440 4384
rect 50376 4324 50380 4380
rect 50380 4324 50436 4380
rect 50436 4324 50440 4380
rect 50376 4320 50440 4324
rect 50456 4380 50520 4384
rect 50456 4324 50460 4380
rect 50460 4324 50516 4380
rect 50516 4324 50520 4380
rect 50456 4320 50520 4324
rect 50536 4380 50600 4384
rect 50536 4324 50540 4380
rect 50540 4324 50596 4380
rect 50596 4324 50600 4380
rect 50536 4320 50600 4324
rect 10732 3980 10796 4044
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 65656 3836 65720 3840
rect 65656 3780 65660 3836
rect 65660 3780 65716 3836
rect 65716 3780 65720 3836
rect 65656 3776 65720 3780
rect 65736 3836 65800 3840
rect 65736 3780 65740 3836
rect 65740 3780 65796 3836
rect 65796 3780 65800 3836
rect 65736 3776 65800 3780
rect 65816 3836 65880 3840
rect 65816 3780 65820 3836
rect 65820 3780 65876 3836
rect 65876 3780 65880 3836
rect 65816 3776 65880 3780
rect 65896 3836 65960 3840
rect 65896 3780 65900 3836
rect 65900 3780 65956 3836
rect 65956 3780 65960 3836
rect 65896 3776 65960 3780
rect 17908 3572 17972 3636
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 50296 3292 50360 3296
rect 50296 3236 50300 3292
rect 50300 3236 50356 3292
rect 50356 3236 50360 3292
rect 50296 3232 50360 3236
rect 50376 3292 50440 3296
rect 50376 3236 50380 3292
rect 50380 3236 50436 3292
rect 50436 3236 50440 3292
rect 50376 3232 50440 3236
rect 50456 3292 50520 3296
rect 50456 3236 50460 3292
rect 50460 3236 50516 3292
rect 50516 3236 50520 3292
rect 50456 3232 50520 3236
rect 50536 3292 50600 3296
rect 50536 3236 50540 3292
rect 50540 3236 50596 3292
rect 50596 3236 50600 3292
rect 50536 3232 50600 3236
rect 11100 3028 11164 3092
rect 12020 2816 12084 2820
rect 12020 2760 12070 2816
rect 12070 2760 12084 2816
rect 12020 2756 12084 2760
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 65656 2748 65720 2752
rect 65656 2692 65660 2748
rect 65660 2692 65716 2748
rect 65716 2692 65720 2748
rect 65656 2688 65720 2692
rect 65736 2748 65800 2752
rect 65736 2692 65740 2748
rect 65740 2692 65796 2748
rect 65796 2692 65800 2748
rect 65736 2688 65800 2692
rect 65816 2748 65880 2752
rect 65816 2692 65820 2748
rect 65820 2692 65876 2748
rect 65876 2692 65880 2748
rect 65816 2688 65880 2692
rect 65896 2748 65960 2752
rect 65896 2692 65900 2748
rect 65900 2692 65956 2748
rect 65956 2692 65960 2748
rect 65896 2688 65960 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
rect 50296 2204 50360 2208
rect 50296 2148 50300 2204
rect 50300 2148 50356 2204
rect 50356 2148 50360 2204
rect 50296 2144 50360 2148
rect 50376 2204 50440 2208
rect 50376 2148 50380 2204
rect 50380 2148 50436 2204
rect 50436 2148 50440 2204
rect 50376 2144 50440 2148
rect 50456 2204 50520 2208
rect 50456 2148 50460 2204
rect 50460 2148 50516 2204
rect 50516 2148 50520 2204
rect 50456 2144 50520 2148
rect 50536 2204 50600 2208
rect 50536 2148 50540 2204
rect 50540 2148 50596 2204
rect 50596 2148 50600 2204
rect 50536 2144 50600 2148
<< metal4 >>
rect 4208 57152 4528 57712
rect 4208 57088 4216 57152
rect 4280 57088 4296 57152
rect 4360 57088 4376 57152
rect 4440 57088 4456 57152
rect 4520 57088 4528 57152
rect 4208 56064 4528 57088
rect 4208 56000 4216 56064
rect 4280 56000 4296 56064
rect 4360 56000 4376 56064
rect 4440 56000 4456 56064
rect 4520 56000 4528 56064
rect 4208 54976 4528 56000
rect 4208 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4528 54976
rect 4208 53888 4528 54912
rect 4208 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4528 53888
rect 4208 52800 4528 53824
rect 4208 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4528 52800
rect 4208 51712 4528 52736
rect 4208 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4528 51712
rect 4208 50624 4528 51648
rect 4208 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4528 50624
rect 4208 49536 4528 50560
rect 4208 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4528 49536
rect 4208 48448 4528 49472
rect 4208 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4528 48448
rect 4208 47360 4528 48384
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 46272 4528 47296
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 45184 4528 46208
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 44096 4528 45120
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 43008 4528 44032
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 41920 4528 42944
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 19568 57696 19888 57712
rect 19568 57632 19576 57696
rect 19640 57632 19656 57696
rect 19720 57632 19736 57696
rect 19800 57632 19816 57696
rect 19880 57632 19888 57696
rect 19568 56608 19888 57632
rect 19568 56544 19576 56608
rect 19640 56544 19656 56608
rect 19720 56544 19736 56608
rect 19800 56544 19816 56608
rect 19880 56544 19888 56608
rect 19568 55520 19888 56544
rect 19568 55456 19576 55520
rect 19640 55456 19656 55520
rect 19720 55456 19736 55520
rect 19800 55456 19816 55520
rect 19880 55456 19888 55520
rect 19568 54432 19888 55456
rect 19568 54368 19576 54432
rect 19640 54368 19656 54432
rect 19720 54368 19736 54432
rect 19800 54368 19816 54432
rect 19880 54368 19888 54432
rect 19568 53344 19888 54368
rect 19568 53280 19576 53344
rect 19640 53280 19656 53344
rect 19720 53280 19736 53344
rect 19800 53280 19816 53344
rect 19880 53280 19888 53344
rect 19568 52256 19888 53280
rect 19568 52192 19576 52256
rect 19640 52192 19656 52256
rect 19720 52192 19736 52256
rect 19800 52192 19816 52256
rect 19880 52192 19888 52256
rect 19568 51168 19888 52192
rect 19568 51104 19576 51168
rect 19640 51104 19656 51168
rect 19720 51104 19736 51168
rect 19800 51104 19816 51168
rect 19880 51104 19888 51168
rect 19568 50080 19888 51104
rect 19568 50016 19576 50080
rect 19640 50016 19656 50080
rect 19720 50016 19736 50080
rect 19800 50016 19816 50080
rect 19880 50016 19888 50080
rect 19568 48992 19888 50016
rect 19568 48928 19576 48992
rect 19640 48928 19656 48992
rect 19720 48928 19736 48992
rect 19800 48928 19816 48992
rect 19880 48928 19888 48992
rect 19568 47904 19888 48928
rect 19568 47840 19576 47904
rect 19640 47840 19656 47904
rect 19720 47840 19736 47904
rect 19800 47840 19816 47904
rect 19880 47840 19888 47904
rect 19568 46816 19888 47840
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 45728 19888 46752
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 44640 19888 45664
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 43552 19888 44576
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 42464 19888 43488
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 41376 19888 42400
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 40288 19888 41312
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 39200 19888 40224
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 38112 19888 39136
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 37024 19888 38048
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 34928 57152 35248 57712
rect 34928 57088 34936 57152
rect 35000 57088 35016 57152
rect 35080 57088 35096 57152
rect 35160 57088 35176 57152
rect 35240 57088 35248 57152
rect 34928 56064 35248 57088
rect 34928 56000 34936 56064
rect 35000 56000 35016 56064
rect 35080 56000 35096 56064
rect 35160 56000 35176 56064
rect 35240 56000 35248 56064
rect 34928 54976 35248 56000
rect 34928 54912 34936 54976
rect 35000 54912 35016 54976
rect 35080 54912 35096 54976
rect 35160 54912 35176 54976
rect 35240 54912 35248 54976
rect 34928 53888 35248 54912
rect 34928 53824 34936 53888
rect 35000 53824 35016 53888
rect 35080 53824 35096 53888
rect 35160 53824 35176 53888
rect 35240 53824 35248 53888
rect 34928 52800 35248 53824
rect 34928 52736 34936 52800
rect 35000 52736 35016 52800
rect 35080 52736 35096 52800
rect 35160 52736 35176 52800
rect 35240 52736 35248 52800
rect 34928 51712 35248 52736
rect 34928 51648 34936 51712
rect 35000 51648 35016 51712
rect 35080 51648 35096 51712
rect 35160 51648 35176 51712
rect 35240 51648 35248 51712
rect 34928 50624 35248 51648
rect 34928 50560 34936 50624
rect 35000 50560 35016 50624
rect 35080 50560 35096 50624
rect 35160 50560 35176 50624
rect 35240 50560 35248 50624
rect 34928 49536 35248 50560
rect 34928 49472 34936 49536
rect 35000 49472 35016 49536
rect 35080 49472 35096 49536
rect 35160 49472 35176 49536
rect 35240 49472 35248 49536
rect 34928 48448 35248 49472
rect 34928 48384 34936 48448
rect 35000 48384 35016 48448
rect 35080 48384 35096 48448
rect 35160 48384 35176 48448
rect 35240 48384 35248 48448
rect 34928 47360 35248 48384
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 46272 35248 47296
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 45184 35248 46208
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 44096 35248 45120
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 43008 35248 44032
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 41920 35248 42944
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 40832 35248 41856
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 39744 35248 40768
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 38656 35248 39680
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 23427 27708 23493 27709
rect 23427 27644 23428 27708
rect 23492 27644 23493 27708
rect 23427 27643 23493 27644
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 23430 24717 23490 27643
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 23427 24716 23493 24717
rect 23427 24652 23428 24716
rect 23492 24652 23493 24716
rect 23427 24651 23493 24652
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 23611 22268 23677 22269
rect 23611 22204 23612 22268
rect 23676 22204 23677 22268
rect 23611 22203 23677 22204
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 21955 18188 22021 18189
rect 21955 18124 21956 18188
rect 22020 18124 22021 18188
rect 21955 18123 22021 18124
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19379 13836 19445 13837
rect 19379 13772 19380 13836
rect 19444 13772 19445 13836
rect 19379 13771 19445 13772
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 17907 12068 17973 12069
rect 17907 12004 17908 12068
rect 17972 12004 17973 12068
rect 17907 12003 17973 12004
rect 11099 11524 11165 11525
rect 11099 11460 11100 11524
rect 11164 11460 11165 11524
rect 11099 11459 11165 11460
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 10731 10300 10797 10301
rect 10731 10236 10732 10300
rect 10796 10236 10797 10300
rect 10731 10235 10797 10236
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 10734 4045 10794 10235
rect 10731 4044 10797 4045
rect 10731 3980 10732 4044
rect 10796 3980 10797 4044
rect 10731 3979 10797 3980
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 11102 3093 11162 11459
rect 12019 8804 12085 8805
rect 12019 8740 12020 8804
rect 12084 8740 12085 8804
rect 12019 8739 12085 8740
rect 11099 3092 11165 3093
rect 11099 3028 11100 3092
rect 11164 3028 11165 3092
rect 11099 3027 11165 3028
rect 12022 2821 12082 8739
rect 17910 3637 17970 12003
rect 19382 7445 19442 13771
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 21958 10709 22018 18123
rect 23614 11389 23674 22203
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 24163 20772 24229 20773
rect 24163 20708 24164 20772
rect 24228 20708 24229 20772
rect 24163 20707 24229 20708
rect 23611 11388 23677 11389
rect 23611 11324 23612 11388
rect 23676 11324 23677 11388
rect 23611 11323 23677 11324
rect 21955 10708 22021 10709
rect 21955 10644 21956 10708
rect 22020 10644 22021 10708
rect 21955 10643 22021 10644
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 24166 9621 24226 20707
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 50288 57696 50608 57712
rect 50288 57632 50296 57696
rect 50360 57632 50376 57696
rect 50440 57632 50456 57696
rect 50520 57632 50536 57696
rect 50600 57632 50608 57696
rect 50288 56608 50608 57632
rect 50288 56544 50296 56608
rect 50360 56544 50376 56608
rect 50440 56544 50456 56608
rect 50520 56544 50536 56608
rect 50600 56544 50608 56608
rect 50288 55520 50608 56544
rect 50288 55456 50296 55520
rect 50360 55456 50376 55520
rect 50440 55456 50456 55520
rect 50520 55456 50536 55520
rect 50600 55456 50608 55520
rect 50288 54432 50608 55456
rect 50288 54368 50296 54432
rect 50360 54368 50376 54432
rect 50440 54368 50456 54432
rect 50520 54368 50536 54432
rect 50600 54368 50608 54432
rect 50288 53344 50608 54368
rect 50288 53280 50296 53344
rect 50360 53280 50376 53344
rect 50440 53280 50456 53344
rect 50520 53280 50536 53344
rect 50600 53280 50608 53344
rect 50288 52256 50608 53280
rect 50288 52192 50296 52256
rect 50360 52192 50376 52256
rect 50440 52192 50456 52256
rect 50520 52192 50536 52256
rect 50600 52192 50608 52256
rect 50288 51168 50608 52192
rect 50288 51104 50296 51168
rect 50360 51104 50376 51168
rect 50440 51104 50456 51168
rect 50520 51104 50536 51168
rect 50600 51104 50608 51168
rect 50288 50080 50608 51104
rect 50288 50016 50296 50080
rect 50360 50016 50376 50080
rect 50440 50016 50456 50080
rect 50520 50016 50536 50080
rect 50600 50016 50608 50080
rect 50288 48992 50608 50016
rect 50288 48928 50296 48992
rect 50360 48928 50376 48992
rect 50440 48928 50456 48992
rect 50520 48928 50536 48992
rect 50600 48928 50608 48992
rect 50288 47904 50608 48928
rect 50288 47840 50296 47904
rect 50360 47840 50376 47904
rect 50440 47840 50456 47904
rect 50520 47840 50536 47904
rect 50600 47840 50608 47904
rect 50288 46816 50608 47840
rect 50288 46752 50296 46816
rect 50360 46752 50376 46816
rect 50440 46752 50456 46816
rect 50520 46752 50536 46816
rect 50600 46752 50608 46816
rect 50288 45728 50608 46752
rect 50288 45664 50296 45728
rect 50360 45664 50376 45728
rect 50440 45664 50456 45728
rect 50520 45664 50536 45728
rect 50600 45664 50608 45728
rect 50288 44640 50608 45664
rect 50288 44576 50296 44640
rect 50360 44576 50376 44640
rect 50440 44576 50456 44640
rect 50520 44576 50536 44640
rect 50600 44576 50608 44640
rect 50288 43552 50608 44576
rect 50288 43488 50296 43552
rect 50360 43488 50376 43552
rect 50440 43488 50456 43552
rect 50520 43488 50536 43552
rect 50600 43488 50608 43552
rect 50288 42464 50608 43488
rect 50288 42400 50296 42464
rect 50360 42400 50376 42464
rect 50440 42400 50456 42464
rect 50520 42400 50536 42464
rect 50600 42400 50608 42464
rect 50288 41376 50608 42400
rect 50288 41312 50296 41376
rect 50360 41312 50376 41376
rect 50440 41312 50456 41376
rect 50520 41312 50536 41376
rect 50600 41312 50608 41376
rect 50288 40288 50608 41312
rect 50288 40224 50296 40288
rect 50360 40224 50376 40288
rect 50440 40224 50456 40288
rect 50520 40224 50536 40288
rect 50600 40224 50608 40288
rect 50288 39200 50608 40224
rect 50288 39136 50296 39200
rect 50360 39136 50376 39200
rect 50440 39136 50456 39200
rect 50520 39136 50536 39200
rect 50600 39136 50608 39200
rect 50288 38112 50608 39136
rect 50288 38048 50296 38112
rect 50360 38048 50376 38112
rect 50440 38048 50456 38112
rect 50520 38048 50536 38112
rect 50600 38048 50608 38112
rect 50288 37024 50608 38048
rect 50288 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50608 37024
rect 50288 35936 50608 36960
rect 50288 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50608 35936
rect 50288 34848 50608 35872
rect 50288 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50608 34848
rect 50288 33760 50608 34784
rect 50288 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50608 33760
rect 50288 32672 50608 33696
rect 50288 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50608 32672
rect 50288 31584 50608 32608
rect 50288 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50608 31584
rect 50288 30496 50608 31520
rect 50288 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50608 30496
rect 50288 29408 50608 30432
rect 50288 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50608 29408
rect 50288 28320 50608 29344
rect 50288 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50608 28320
rect 50288 27232 50608 28256
rect 50288 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50608 27232
rect 50288 26144 50608 27168
rect 50288 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50608 26144
rect 50288 25056 50608 26080
rect 50288 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50608 25056
rect 50288 23968 50608 24992
rect 50288 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50608 23968
rect 50288 22880 50608 23904
rect 50288 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50608 22880
rect 50288 21792 50608 22816
rect 50288 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50608 21792
rect 50288 20704 50608 21728
rect 50288 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50608 20704
rect 50288 19616 50608 20640
rect 50288 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50608 19616
rect 50288 18528 50608 19552
rect 50288 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50608 18528
rect 50288 17440 50608 18464
rect 50288 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50608 17440
rect 50288 16352 50608 17376
rect 50288 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50608 16352
rect 50288 15264 50608 16288
rect 50288 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50608 15264
rect 50288 14176 50608 15200
rect 50288 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50608 14176
rect 35571 14108 35637 14109
rect 35571 14044 35572 14108
rect 35636 14044 35637 14108
rect 35571 14043 35637 14044
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 35574 11933 35634 14043
rect 50288 13088 50608 14112
rect 50288 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50608 13088
rect 50288 12000 50608 13024
rect 50288 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50608 12000
rect 35571 11932 35637 11933
rect 35571 11868 35572 11932
rect 35636 11868 35637 11932
rect 35571 11867 35637 11868
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 24163 9620 24229 9621
rect 24163 9556 24164 9620
rect 24228 9556 24229 9620
rect 24163 9555 24229 9556
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19379 7444 19445 7445
rect 19379 7380 19380 7444
rect 19444 7380 19445 7444
rect 19379 7379 19445 7380
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 17907 3636 17973 3637
rect 17907 3572 17908 3636
rect 17972 3572 17973 3636
rect 17907 3571 17973 3572
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 12019 2820 12085 2821
rect 12019 2756 12020 2820
rect 12084 2756 12085 2820
rect 12019 2755 12085 2756
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
rect 50288 10912 50608 11936
rect 50288 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50608 10912
rect 50288 9824 50608 10848
rect 50288 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50608 9824
rect 50288 8736 50608 9760
rect 50288 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50608 8736
rect 50288 7648 50608 8672
rect 50288 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50608 7648
rect 50288 6560 50608 7584
rect 50288 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50608 6560
rect 50288 5472 50608 6496
rect 50288 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50608 5472
rect 50288 4384 50608 5408
rect 50288 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50608 4384
rect 50288 3296 50608 4320
rect 50288 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50608 3296
rect 50288 2208 50608 3232
rect 50288 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50608 2208
rect 50288 2128 50608 2144
rect 65648 57152 65968 57712
rect 65648 57088 65656 57152
rect 65720 57088 65736 57152
rect 65800 57088 65816 57152
rect 65880 57088 65896 57152
rect 65960 57088 65968 57152
rect 65648 56064 65968 57088
rect 65648 56000 65656 56064
rect 65720 56000 65736 56064
rect 65800 56000 65816 56064
rect 65880 56000 65896 56064
rect 65960 56000 65968 56064
rect 65648 54976 65968 56000
rect 65648 54912 65656 54976
rect 65720 54912 65736 54976
rect 65800 54912 65816 54976
rect 65880 54912 65896 54976
rect 65960 54912 65968 54976
rect 65648 53888 65968 54912
rect 65648 53824 65656 53888
rect 65720 53824 65736 53888
rect 65800 53824 65816 53888
rect 65880 53824 65896 53888
rect 65960 53824 65968 53888
rect 65648 52800 65968 53824
rect 65648 52736 65656 52800
rect 65720 52736 65736 52800
rect 65800 52736 65816 52800
rect 65880 52736 65896 52800
rect 65960 52736 65968 52800
rect 65648 51712 65968 52736
rect 65648 51648 65656 51712
rect 65720 51648 65736 51712
rect 65800 51648 65816 51712
rect 65880 51648 65896 51712
rect 65960 51648 65968 51712
rect 65648 50624 65968 51648
rect 65648 50560 65656 50624
rect 65720 50560 65736 50624
rect 65800 50560 65816 50624
rect 65880 50560 65896 50624
rect 65960 50560 65968 50624
rect 65648 49536 65968 50560
rect 65648 49472 65656 49536
rect 65720 49472 65736 49536
rect 65800 49472 65816 49536
rect 65880 49472 65896 49536
rect 65960 49472 65968 49536
rect 65648 48448 65968 49472
rect 65648 48384 65656 48448
rect 65720 48384 65736 48448
rect 65800 48384 65816 48448
rect 65880 48384 65896 48448
rect 65960 48384 65968 48448
rect 65648 47360 65968 48384
rect 65648 47296 65656 47360
rect 65720 47296 65736 47360
rect 65800 47296 65816 47360
rect 65880 47296 65896 47360
rect 65960 47296 65968 47360
rect 65648 46272 65968 47296
rect 65648 46208 65656 46272
rect 65720 46208 65736 46272
rect 65800 46208 65816 46272
rect 65880 46208 65896 46272
rect 65960 46208 65968 46272
rect 65648 45184 65968 46208
rect 65648 45120 65656 45184
rect 65720 45120 65736 45184
rect 65800 45120 65816 45184
rect 65880 45120 65896 45184
rect 65960 45120 65968 45184
rect 65648 44096 65968 45120
rect 65648 44032 65656 44096
rect 65720 44032 65736 44096
rect 65800 44032 65816 44096
rect 65880 44032 65896 44096
rect 65960 44032 65968 44096
rect 65648 43008 65968 44032
rect 65648 42944 65656 43008
rect 65720 42944 65736 43008
rect 65800 42944 65816 43008
rect 65880 42944 65896 43008
rect 65960 42944 65968 43008
rect 65648 41920 65968 42944
rect 65648 41856 65656 41920
rect 65720 41856 65736 41920
rect 65800 41856 65816 41920
rect 65880 41856 65896 41920
rect 65960 41856 65968 41920
rect 65648 40832 65968 41856
rect 65648 40768 65656 40832
rect 65720 40768 65736 40832
rect 65800 40768 65816 40832
rect 65880 40768 65896 40832
rect 65960 40768 65968 40832
rect 65648 39744 65968 40768
rect 65648 39680 65656 39744
rect 65720 39680 65736 39744
rect 65800 39680 65816 39744
rect 65880 39680 65896 39744
rect 65960 39680 65968 39744
rect 65648 38656 65968 39680
rect 65648 38592 65656 38656
rect 65720 38592 65736 38656
rect 65800 38592 65816 38656
rect 65880 38592 65896 38656
rect 65960 38592 65968 38656
rect 65648 37568 65968 38592
rect 65648 37504 65656 37568
rect 65720 37504 65736 37568
rect 65800 37504 65816 37568
rect 65880 37504 65896 37568
rect 65960 37504 65968 37568
rect 65648 36480 65968 37504
rect 65648 36416 65656 36480
rect 65720 36416 65736 36480
rect 65800 36416 65816 36480
rect 65880 36416 65896 36480
rect 65960 36416 65968 36480
rect 65648 35392 65968 36416
rect 65648 35328 65656 35392
rect 65720 35328 65736 35392
rect 65800 35328 65816 35392
rect 65880 35328 65896 35392
rect 65960 35328 65968 35392
rect 65648 34304 65968 35328
rect 65648 34240 65656 34304
rect 65720 34240 65736 34304
rect 65800 34240 65816 34304
rect 65880 34240 65896 34304
rect 65960 34240 65968 34304
rect 65648 33216 65968 34240
rect 65648 33152 65656 33216
rect 65720 33152 65736 33216
rect 65800 33152 65816 33216
rect 65880 33152 65896 33216
rect 65960 33152 65968 33216
rect 65648 32128 65968 33152
rect 65648 32064 65656 32128
rect 65720 32064 65736 32128
rect 65800 32064 65816 32128
rect 65880 32064 65896 32128
rect 65960 32064 65968 32128
rect 65648 31040 65968 32064
rect 65648 30976 65656 31040
rect 65720 30976 65736 31040
rect 65800 30976 65816 31040
rect 65880 30976 65896 31040
rect 65960 30976 65968 31040
rect 65648 29952 65968 30976
rect 65648 29888 65656 29952
rect 65720 29888 65736 29952
rect 65800 29888 65816 29952
rect 65880 29888 65896 29952
rect 65960 29888 65968 29952
rect 65648 28864 65968 29888
rect 65648 28800 65656 28864
rect 65720 28800 65736 28864
rect 65800 28800 65816 28864
rect 65880 28800 65896 28864
rect 65960 28800 65968 28864
rect 65648 27776 65968 28800
rect 65648 27712 65656 27776
rect 65720 27712 65736 27776
rect 65800 27712 65816 27776
rect 65880 27712 65896 27776
rect 65960 27712 65968 27776
rect 65648 26688 65968 27712
rect 65648 26624 65656 26688
rect 65720 26624 65736 26688
rect 65800 26624 65816 26688
rect 65880 26624 65896 26688
rect 65960 26624 65968 26688
rect 65648 25600 65968 26624
rect 65648 25536 65656 25600
rect 65720 25536 65736 25600
rect 65800 25536 65816 25600
rect 65880 25536 65896 25600
rect 65960 25536 65968 25600
rect 65648 24512 65968 25536
rect 65648 24448 65656 24512
rect 65720 24448 65736 24512
rect 65800 24448 65816 24512
rect 65880 24448 65896 24512
rect 65960 24448 65968 24512
rect 65648 23424 65968 24448
rect 65648 23360 65656 23424
rect 65720 23360 65736 23424
rect 65800 23360 65816 23424
rect 65880 23360 65896 23424
rect 65960 23360 65968 23424
rect 65648 22336 65968 23360
rect 65648 22272 65656 22336
rect 65720 22272 65736 22336
rect 65800 22272 65816 22336
rect 65880 22272 65896 22336
rect 65960 22272 65968 22336
rect 65648 21248 65968 22272
rect 65648 21184 65656 21248
rect 65720 21184 65736 21248
rect 65800 21184 65816 21248
rect 65880 21184 65896 21248
rect 65960 21184 65968 21248
rect 65648 20160 65968 21184
rect 65648 20096 65656 20160
rect 65720 20096 65736 20160
rect 65800 20096 65816 20160
rect 65880 20096 65896 20160
rect 65960 20096 65968 20160
rect 65648 19072 65968 20096
rect 65648 19008 65656 19072
rect 65720 19008 65736 19072
rect 65800 19008 65816 19072
rect 65880 19008 65896 19072
rect 65960 19008 65968 19072
rect 65648 17984 65968 19008
rect 65648 17920 65656 17984
rect 65720 17920 65736 17984
rect 65800 17920 65816 17984
rect 65880 17920 65896 17984
rect 65960 17920 65968 17984
rect 65648 16896 65968 17920
rect 65648 16832 65656 16896
rect 65720 16832 65736 16896
rect 65800 16832 65816 16896
rect 65880 16832 65896 16896
rect 65960 16832 65968 16896
rect 65648 15808 65968 16832
rect 65648 15744 65656 15808
rect 65720 15744 65736 15808
rect 65800 15744 65816 15808
rect 65880 15744 65896 15808
rect 65960 15744 65968 15808
rect 65648 14720 65968 15744
rect 65648 14656 65656 14720
rect 65720 14656 65736 14720
rect 65800 14656 65816 14720
rect 65880 14656 65896 14720
rect 65960 14656 65968 14720
rect 65648 13632 65968 14656
rect 65648 13568 65656 13632
rect 65720 13568 65736 13632
rect 65800 13568 65816 13632
rect 65880 13568 65896 13632
rect 65960 13568 65968 13632
rect 65648 12544 65968 13568
rect 65648 12480 65656 12544
rect 65720 12480 65736 12544
rect 65800 12480 65816 12544
rect 65880 12480 65896 12544
rect 65960 12480 65968 12544
rect 65648 11456 65968 12480
rect 65648 11392 65656 11456
rect 65720 11392 65736 11456
rect 65800 11392 65816 11456
rect 65880 11392 65896 11456
rect 65960 11392 65968 11456
rect 65648 10368 65968 11392
rect 65648 10304 65656 10368
rect 65720 10304 65736 10368
rect 65800 10304 65816 10368
rect 65880 10304 65896 10368
rect 65960 10304 65968 10368
rect 65648 9280 65968 10304
rect 65648 9216 65656 9280
rect 65720 9216 65736 9280
rect 65800 9216 65816 9280
rect 65880 9216 65896 9280
rect 65960 9216 65968 9280
rect 65648 8192 65968 9216
rect 65648 8128 65656 8192
rect 65720 8128 65736 8192
rect 65800 8128 65816 8192
rect 65880 8128 65896 8192
rect 65960 8128 65968 8192
rect 65648 7104 65968 8128
rect 65648 7040 65656 7104
rect 65720 7040 65736 7104
rect 65800 7040 65816 7104
rect 65880 7040 65896 7104
rect 65960 7040 65968 7104
rect 65648 6016 65968 7040
rect 65648 5952 65656 6016
rect 65720 5952 65736 6016
rect 65800 5952 65816 6016
rect 65880 5952 65896 6016
rect 65960 5952 65968 6016
rect 65648 4928 65968 5952
rect 65648 4864 65656 4928
rect 65720 4864 65736 4928
rect 65800 4864 65816 4928
rect 65880 4864 65896 4928
rect 65960 4864 65968 4928
rect 65648 3840 65968 4864
rect 65648 3776 65656 3840
rect 65720 3776 65736 3840
rect 65800 3776 65816 3840
rect 65880 3776 65896 3840
rect 65960 3776 65968 3840
rect 65648 2752 65968 3776
rect 65648 2688 65656 2752
rect 65720 2688 65736 2752
rect 65800 2688 65816 2752
rect 65880 2688 65896 2752
rect 65960 2688 65968 2752
rect 65648 2128 65968 2688
use sky130_fd_sc_hd__diode_2  ANTENNA__0775__B dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2760 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0776__B
timestamp 1649977179
transform 1 0 3496 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0781__A
timestamp 1649977179
transform -1 0 4232 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0781__C
timestamp 1649977179
transform 1 0 2668 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0782__A
timestamp 1649977179
transform 1 0 2392 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0784__C
timestamp 1649977179
transform -1 0 6440 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0787__B1
timestamp 1649977179
transform 1 0 6808 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0789__A2
timestamp 1649977179
transform -1 0 7084 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0793__A
timestamp 1649977179
transform 1 0 10028 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0793__B
timestamp 1649977179
transform 1 0 8648 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0796__A
timestamp 1649977179
transform -1 0 8464 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0800__A1
timestamp 1649977179
transform 1 0 10304 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0800__A2
timestamp 1649977179
transform 1 0 10856 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0800__B1
timestamp 1649977179
transform 1 0 12236 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0803__A
timestamp 1649977179
transform -1 0 7544 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0804__A1
timestamp 1649977179
transform 1 0 7176 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0805__D
timestamp 1649977179
transform 1 0 7728 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0806__A1
timestamp 1649977179
transform 1 0 8924 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0808__A
timestamp 1649977179
transform 1 0 2484 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0809__A
timestamp 1649977179
transform -1 0 3036 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0810__B2
timestamp 1649977179
transform -1 0 10672 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0812__A1
timestamp 1649977179
transform -1 0 9292 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0837__A
timestamp 1649977179
transform -1 0 33396 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0847__D1
timestamp 1649977179
transform 1 0 30912 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0867__D
timestamp 1649977179
transform -1 0 36800 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0868__D
timestamp 1649977179
transform -1 0 36800 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0869__A
timestamp 1649977179
transform -1 0 41768 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0869__B
timestamp 1649977179
transform 1 0 40664 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0869__C
timestamp 1649977179
transform 1 0 41032 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0874__A
timestamp 1649977179
transform -1 0 39100 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0874__B
timestamp 1649977179
transform -1 0 38824 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0874__C
timestamp 1649977179
transform 1 0 38916 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0876__A
timestamp 1649977179
transform 1 0 40204 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0876__B
timestamp 1649977179
transform -1 0 41768 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0879__A1
timestamp 1649977179
transform 1 0 40756 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0880__A1
timestamp 1649977179
transform -1 0 42320 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0881__D
timestamp 1649977179
transform 1 0 40664 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0896__B
timestamp 1649977179
transform -1 0 18768 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0908__A
timestamp 1649977179
transform 1 0 2944 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0909__A
timestamp 1649977179
transform 1 0 21160 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0911__A
timestamp 1649977179
transform -1 0 20608 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0912__A1
timestamp 1649977179
transform 1 0 2852 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0912__C1
timestamp 1649977179
transform 1 0 3772 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0913__A
timestamp 1649977179
transform 1 0 3772 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0914__C1
timestamp 1649977179
transform -1 0 2944 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0915__A
timestamp 1649977179
transform 1 0 2944 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0916__A1
timestamp 1649977179
transform -1 0 2852 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0916__C1
timestamp 1649977179
transform 1 0 2392 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0917__A
timestamp 1649977179
transform -1 0 2392 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0918__C1
timestamp 1649977179
transform 1 0 3496 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0919__A
timestamp 1649977179
transform -1 0 4508 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0920__A
timestamp 1649977179
transform 1 0 14996 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0925__A
timestamp 1649977179
transform 1 0 12880 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0927__A
timestamp 1649977179
transform 1 0 11040 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0929__A
timestamp 1649977179
transform 1 0 8188 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0931__A
timestamp 1649977179
transform 1 0 13248 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0933__A
timestamp 1649977179
transform 1 0 10856 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0936__A
timestamp 1649977179
transform 1 0 10580 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0938__A
timestamp 1649977179
transform 1 0 12328 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0939__B
timestamp 1649977179
transform -1 0 21988 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0946__A1
timestamp 1649977179
transform 1 0 6532 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0947__A
timestamp 1649977179
transform 1 0 2116 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0950__A
timestamp 1649977179
transform -1 0 1748 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0951__A1
timestamp 1649977179
transform 1 0 3772 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0952__A
timestamp 1649977179
transform -1 0 2116 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0954__A1
timestamp 1649977179
transform -1 0 3956 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0955__A
timestamp 1649977179
transform 1 0 18860 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0956__A
timestamp 1649977179
transform 1 0 3772 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0958__A1
timestamp 1649977179
transform 1 0 4048 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0959__A
timestamp 1649977179
transform -1 0 18768 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0961__A1
timestamp 1649977179
transform 1 0 3772 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0962__A
timestamp 1649977179
transform 1 0 20792 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0965__A1
timestamp 1649977179
transform 1 0 7176 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0966__A
timestamp 1649977179
transform 1 0 21436 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0968__A1
timestamp 1649977179
transform -1 0 12880 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0969__A
timestamp 1649977179
transform 1 0 18308 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0971__A1
timestamp 1649977179
transform 1 0 9200 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0972__A
timestamp 1649977179
transform -1 0 23460 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0975__A1
timestamp 1649977179
transform 1 0 8096 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0976__A
timestamp 1649977179
transform 1 0 20424 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0978__A1
timestamp 1649977179
transform 1 0 10764 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0979__A
timestamp 1649977179
transform 1 0 18308 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0982__B
timestamp 1649977179
transform 1 0 21252 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0988__A1
timestamp 1649977179
transform 1 0 9844 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0991__A
timestamp 1649977179
transform 1 0 5612 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0992__A1
timestamp 1649977179
transform 1 0 4692 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0993__A
timestamp 1649977179
transform 1 0 3036 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0994__A
timestamp 1649977179
transform -1 0 17296 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0996__A1
timestamp 1649977179
transform 1 0 2944 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0997__A
timestamp 1649977179
transform 1 0 3588 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0998__A1
timestamp 1649977179
transform 1 0 3128 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1000__A1
timestamp 1649977179
transform 1 0 6348 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1003__A1
timestamp 1649977179
transform 1 0 7176 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1005__A1
timestamp 1649977179
transform 1 0 9660 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1008__A1
timestamp 1649977179
transform 1 0 8280 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1010__A1
timestamp 1649977179
transform -1 0 6440 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1012__A1
timestamp 1649977179
transform 1 0 10120 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1016__B_N
timestamp 1649977179
transform 1 0 16008 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1020__A
timestamp 1649977179
transform 1 0 18492 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1023__A
timestamp 1649977179
transform 1 0 16652 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1025__A
timestamp 1649977179
transform -1 0 5888 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1026__A1
timestamp 1649977179
transform 1 0 6440 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1027__A
timestamp 1649977179
transform 1 0 4324 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1029__A1
timestamp 1649977179
transform 1 0 3036 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1030__A
timestamp 1649977179
transform 1 0 9016 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1031__A1
timestamp 1649977179
transform 1 0 5980 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1033__A1
timestamp 1649977179
transform 1 0 11868 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1034__A
timestamp 1649977179
transform 1 0 2760 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1035__A1
timestamp 1649977179
transform 1 0 4232 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1039__A1
timestamp 1649977179
transform -1 0 16192 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1042__A1
timestamp 1649977179
transform -1 0 18400 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1044__A1
timestamp 1649977179
transform 1 0 15916 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1046__A1
timestamp 1649977179
transform 1 0 17756 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1048__A1
timestamp 1649977179
transform 1 0 18400 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1054__A
timestamp 1649977179
transform 1 0 20700 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1057__A
timestamp 1649977179
transform 1 0 18584 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1061__A1
timestamp 1649977179
transform 1 0 14536 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1063__A1
timestamp 1649977179
transform 1 0 12880 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1065__A1
timestamp 1649977179
transform -1 0 19504 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1067__A1
timestamp 1649977179
transform -1 0 17480 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1069__A1
timestamp 1649977179
transform 1 0 19596 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1073__A
timestamp 1649977179
transform 1 0 20424 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1075__A1
timestamp 1649977179
transform -1 0 24656 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1077__A1
timestamp 1649977179
transform 1 0 24380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1079__A1
timestamp 1649977179
transform -1 0 20608 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1081__A1
timestamp 1649977179
transform -1 0 25484 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1083__A1
timestamp 1649977179
transform -1 0 22724 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1089__A
timestamp 1649977179
transform -1 0 14352 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1092__A
timestamp 1649977179
transform 1 0 14076 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1095__A1
timestamp 1649977179
transform 1 0 11960 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1097__A1
timestamp 1649977179
transform 1 0 12696 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1099__A1
timestamp 1649977179
transform 1 0 11224 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1101__A1
timestamp 1649977179
transform 1 0 12604 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1104__A1
timestamp 1649977179
transform 1 0 13432 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1108__A1
timestamp 1649977179
transform 1 0 17756 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1110__A1
timestamp 1649977179
transform 1 0 18216 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1112__A1
timestamp 1649977179
transform 1 0 17204 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1114__A1
timestamp 1649977179
transform 1 0 16468 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1117__A1
timestamp 1649977179
transform 1 0 18676 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1120__A
timestamp 1649977179
transform -1 0 24840 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1121__A
timestamp 1649977179
transform 1 0 20332 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1125__A
timestamp 1649977179
transform 1 0 23736 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1127__A
timestamp 1649977179
transform 1 0 22264 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1130__A1
timestamp 1649977179
transform 1 0 26404 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1131__A
timestamp 1649977179
transform 1 0 25024 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1133__A1
timestamp 1649977179
transform 1 0 26220 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1134__A
timestamp 1649977179
transform 1 0 27968 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1136__A1
timestamp 1649977179
transform 1 0 26956 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1137__A
timestamp 1649977179
transform 1 0 23092 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1141__A
timestamp 1649977179
transform 1 0 23092 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1143__A1
timestamp 1649977179
transform 1 0 24656 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1144__A
timestamp 1649977179
transform 1 0 28428 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1148__A1
timestamp 1649977179
transform -1 0 27968 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1149__A
timestamp 1649977179
transform -1 0 27140 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1151__A1
timestamp 1649977179
transform -1 0 26588 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1152__A
timestamp 1649977179
transform 1 0 27692 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1154__A1
timestamp 1649977179
transform -1 0 27324 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1155__A
timestamp 1649977179
transform 1 0 26312 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1159__A1
timestamp 1649977179
transform 1 0 29072 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1160__A
timestamp 1649977179
transform -1 0 26036 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1162__A1
timestamp 1649977179
transform 1 0 30360 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1163__A
timestamp 1649977179
transform -1 0 24564 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1165__A1
timestamp 1649977179
transform 1 0 27508 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1169__A
timestamp 1649977179
transform 1 0 31648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1171__A
timestamp 1649977179
transform 1 0 27232 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1174__A1
timestamp 1649977179
transform 1 0 27784 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1176__A1
timestamp 1649977179
transform 1 0 27692 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1179__A1
timestamp 1649977179
transform 1 0 29624 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1183__A1
timestamp 1649977179
transform 1 0 28888 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1187__A1
timestamp 1649977179
transform 1 0 36616 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1188__A
timestamp 1649977179
transform 1 0 34040 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1189__A1
timestamp 1649977179
transform 1 0 34684 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1192__A1
timestamp 1649977179
transform 1 0 32108 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1194__A1
timestamp 1649977179
transform 1 0 36616 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1196__A1
timestamp 1649977179
transform 1 0 36708 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1198__A1
timestamp 1649977179
transform 1 0 30912 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1203__A
timestamp 1649977179
transform 1 0 32844 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1205__A
timestamp 1649977179
transform 1 0 30544 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1208__A1
timestamp 1649977179
transform 1 0 35788 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1211__A1
timestamp 1649977179
transform -1 0 39008 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1213__A1
timestamp 1649977179
transform -1 0 38364 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1217__A1
timestamp 1649977179
transform 1 0 34040 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1221__A1
timestamp 1649977179
transform 1 0 36432 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1222__A
timestamp 1649977179
transform 1 0 39100 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1224__A1
timestamp 1649977179
transform -1 0 37444 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1226__A1
timestamp 1649977179
transform -1 0 38548 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1228__A1
timestamp 1649977179
transform 1 0 36616 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1230__A1
timestamp 1649977179
transform 1 0 38180 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1232__A1
timestamp 1649977179
transform 1 0 36524 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1236__A
timestamp 1649977179
transform 1 0 32384 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1238__A
timestamp 1649977179
transform -1 0 31740 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1240__A
timestamp 1649977179
transform 1 0 40020 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1243__A1
timestamp 1649977179
transform 1 0 36248 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1244__A
timestamp 1649977179
transform 1 0 36616 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1245__A1
timestamp 1649977179
transform 1 0 38456 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1246__A
timestamp 1649977179
transform -1 0 39652 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1247__A1
timestamp 1649977179
transform -1 0 38548 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1248__A
timestamp 1649977179
transform 1 0 34224 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1251__A1
timestamp 1649977179
transform 1 0 33396 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1256__A1
timestamp 1649977179
transform -1 0 33488 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1258__A1
timestamp 1649977179
transform 1 0 33948 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1259__A
timestamp 1649977179
transform 1 0 39100 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1260__A1
timestamp 1649977179
transform 1 0 36616 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1262__A1
timestamp 1649977179
transform -1 0 37720 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1264__A1
timestamp 1649977179
transform -1 0 38456 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1267__A1
timestamp 1649977179
transform 1 0 31464 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1271__A
timestamp 1649977179
transform 1 0 29716 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1273__A
timestamp 1649977179
transform 1 0 26312 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1276__A1
timestamp 1649977179
transform -1 0 26588 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1278__A1
timestamp 1649977179
transform -1 0 25760 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1280__A1
timestamp 1649977179
transform 1 0 26036 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1285__A1
timestamp 1649977179
transform 1 0 25576 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1289__A1
timestamp 1649977179
transform 1 0 34040 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1291__A1
timestamp 1649977179
transform 1 0 33120 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1293__A1
timestamp 1649977179
transform -1 0 32936 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1295__A1
timestamp 1649977179
transform 1 0 35512 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1298__A1
timestamp 1649977179
transform -1 0 31648 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1300__A1
timestamp 1649977179
transform -1 0 28704 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1303__A
timestamp 1649977179
transform 1 0 23736 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1306__A
timestamp 1649977179
transform -1 0 23368 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1309__A1
timestamp 1649977179
transform 1 0 29348 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1311__A1
timestamp 1649977179
transform 1 0 27784 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1313__A1
timestamp 1649977179
transform 1 0 27508 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1317__A1
timestamp 1649977179
transform 1 0 22080 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1319__A1
timestamp 1649977179
transform 1 0 23092 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1323__A1
timestamp 1649977179
transform 1 0 26772 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1325__A1
timestamp 1649977179
transform 1 0 23736 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1327__A1
timestamp 1649977179
transform 1 0 26956 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1330__A1
timestamp 1649977179
transform 1 0 24472 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1330__C1
timestamp 1649977179
transform 1 0 26128 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1332__A1
timestamp 1649977179
transform 1 0 23828 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1332__C1
timestamp 1649977179
transform 1 0 23736 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1334__A1
timestamp 1649977179
transform 1 0 23184 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1334__C1
timestamp 1649977179
transform -1 0 23920 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1339__A
timestamp 1649977179
transform -1 0 10856 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1345__A1
timestamp 1649977179
transform 1 0 8280 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1345__C1
timestamp 1649977179
transform -1 0 9200 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1347__A1
timestamp 1649977179
transform 1 0 7176 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1347__C1
timestamp 1649977179
transform 1 0 9108 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1350__A1
timestamp 1649977179
transform 1 0 8924 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1352__A1
timestamp 1649977179
transform 1 0 5704 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1354__A1
timestamp 1649977179
transform 1 0 4784 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1358__A1
timestamp 1649977179
transform -1 0 5060 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1360__A1
timestamp 1649977179
transform -1 0 7360 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1363__A1
timestamp 1649977179
transform -1 0 8372 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1365__A1
timestamp 1649977179
transform 1 0 7176 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1367__A1
timestamp 1649977179
transform -1 0 4784 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1369__A1
timestamp 1649977179
transform -1 0 4968 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1374__B
timestamp 1649977179
transform 1 0 20424 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1386__A1
timestamp 1649977179
transform -1 0 18308 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1387__B2
timestamp 1649977179
transform -1 0 21068 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1393__A1
timestamp 1649977179
transform 1 0 10856 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1394__A
timestamp 1649977179
transform -1 0 20056 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1399__A1
timestamp 1649977179
transform 1 0 13432 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1402__A1
timestamp 1649977179
transform -1 0 22540 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1404__A1
timestamp 1649977179
transform -1 0 18492 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1405__A1
timestamp 1649977179
transform -1 0 23276 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1418__B2
timestamp 1649977179
transform -1 0 24564 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1419__A1
timestamp 1649977179
transform -1 0 21344 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1420__A1
timestamp 1649977179
transform 1 0 8280 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1422__A1
timestamp 1649977179
transform -1 0 18032 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1431__A
timestamp 1649977179
transform 1 0 22264 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1432__A1
timestamp 1649977179
transform 1 0 20332 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1433__A1
timestamp 1649977179
transform -1 0 20608 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1440__A1
timestamp 1649977179
transform -1 0 25300 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1446__B1
timestamp 1649977179
transform -1 0 17388 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1455__C1
timestamp 1649977179
transform -1 0 17296 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1462__A1
timestamp 1649977179
transform 1 0 25024 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1463__A1
timestamp 1649977179
transform -1 0 29164 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1465__B1
timestamp 1649977179
transform 1 0 17020 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1471__B2
timestamp 1649977179
transform 1 0 21988 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1505__A
timestamp 1649977179
transform 1 0 22816 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1506__B1
timestamp 1649977179
transform 1 0 10856 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1508__A
timestamp 1649977179
transform 1 0 32108 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1514__A
timestamp 1649977179
transform 1 0 9660 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1515__A
timestamp 1649977179
transform 1 0 23736 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1516__A
timestamp 1649977179
transform -1 0 27784 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1517__A
timestamp 1649977179
transform 1 0 25760 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1518__A
timestamp 1649977179
transform 1 0 7636 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1519__A
timestamp 1649977179
transform 1 0 5428 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1520__A
timestamp 1649977179
transform 1 0 5612 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1521__A
timestamp 1649977179
transform 1 0 5520 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1678__RESET_B
timestamp 1649977179
transform 1 0 33672 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_wb_clk_i_A
timestamp 1649977179
transform 1 0 21804 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_0_0_wb_clk_i_A
timestamp 1649977179
transform 1 0 7636 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_1_0_wb_clk_i_A
timestamp 1649977179
transform 1 0 8924 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_2_0_wb_clk_i_A
timestamp 1649977179
transform 1 0 15088 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_3_0_wb_clk_i_A
timestamp 1649977179
transform 1 0 15180 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_4_0_wb_clk_i_A
timestamp 1649977179
transform 1 0 8924 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_5_0_wb_clk_i_A
timestamp 1649977179
transform 1 0 7544 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_6_0_wb_clk_i_A
timestamp 1649977179
transform 1 0 13432 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_7_0_wb_clk_i_A
timestamp 1649977179
transform -1 0 14444 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_8_0_wb_clk_i_A
timestamp 1649977179
transform -1 0 30084 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_9_0_wb_clk_i_A
timestamp 1649977179
transform 1 0 26956 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_10_0_wb_clk_i_A
timestamp 1649977179
transform 1 0 34040 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_11_0_wb_clk_i_A
timestamp 1649977179
transform 1 0 34500 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_12_0_wb_clk_i_A
timestamp 1649977179
transform 1 0 28796 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_13_0_wb_clk_i_A
timestamp 1649977179
transform -1 0 28060 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_14_0_wb_clk_i_A
timestamp 1649977179
transform 1 0 34868 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_15_0_wb_clk_i_A
timestamp 1649977179
transform 1 0 35144 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1649977179
transform -1 0 4232 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1649977179
transform -1 0 3312 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1649977179
transform -1 0 5060 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1649977179
transform -1 0 15916 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1649977179
transform -1 0 21160 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1649977179
transform -1 0 3956 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1649977179
transform -1 0 19412 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1649977179
transform -1 0 21988 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1649977179
transform -1 0 10396 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1649977179
transform -1 0 4508 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1649977179
transform -1 0 11040 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1649977179
transform -1 0 10488 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1649977179
transform -1 0 9752 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1649977179
transform -1 0 3496 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1649977179
transform -1 0 4048 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1649977179
transform -1 0 16192 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1649977179
transform -1 0 12328 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1649977179
transform -1 0 6624 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1649977179
transform -1 0 24564 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1649977179
transform -1 0 9936 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1649977179
transform -1 0 11684 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1649977179
transform -1 0 4600 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1649977179
transform -1 0 5152 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1649977179
transform -1 0 16192 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1649977179
transform -1 0 13616 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1649977179
transform -1 0 8464 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1649977179
transform -1 0 6072 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1649977179
transform -1 0 5520 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1649977179
transform -1 0 4784 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output30_A
timestamp 1649977179
transform 1 0 21712 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output31_A
timestamp 1649977179
transform 1 0 30084 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output32_A
timestamp 1649977179
transform 1 0 39192 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output33_A
timestamp 1649977179
transform 1 0 47564 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output34_A
timestamp 1649977179
transform 1 0 56304 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output35_A
timestamp 1649977179
transform 1 0 64952 0 -1 57664
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2484 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3036 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31
timestamp 1649977179
transform 1 0 3956 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37
timestamp 1649977179
transform 1 0 4508 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44
timestamp 1649977179
transform 1 0 5152 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52
timestamp 1649977179
transform 1 0 5888 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57
timestamp 1649977179
transform 1 0 6348 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_62
timestamp 1649977179
transform 1 0 6808 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_74
timestamp 1649977179
transform 1 0 7912 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_80
timestamp 1649977179
transform 1 0 8464 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_85 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 8924 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_92
timestamp 1649977179
transform 1 0 9568 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_100
timestamp 1649977179
transform 1 0 10304 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_108
timestamp 1649977179
transform 1 0 11040 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_113
timestamp 1649977179
transform 1 0 11500 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_122
timestamp 1649977179
transform 1 0 12328 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_136
timestamp 1649977179
transform 1 0 13616 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_145
timestamp 1649977179
transform 1 0 14444 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_153
timestamp 1649977179
transform 1 0 15180 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_161
timestamp 1649977179
transform 1 0 15916 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_167
timestamp 1649977179
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_173
timestamp 1649977179
transform 1 0 17020 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_181
timestamp 1649977179
transform 1 0 17756 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_189
timestamp 1649977179
transform 1 0 18492 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_195
timestamp 1649977179
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_199
timestamp 1649977179
transform 1 0 19412 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_206
timestamp 1649977179
transform 1 0 20056 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_213
timestamp 1649977179
transform 1 0 20700 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_220
timestamp 1649977179
transform 1 0 21344 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_227
timestamp 1649977179
transform 1 0 21988 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_234
timestamp 1649977179
transform 1 0 22632 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_241
timestamp 1649977179
transform 1 0 23276 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_248
timestamp 1649977179
transform 1 0 23920 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_255
timestamp 1649977179
transform 1 0 24564 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_262
timestamp 1649977179
transform 1 0 25208 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_269
timestamp 1649977179
transform 1 0 25852 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_276
timestamp 1649977179
transform 1 0 26496 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_281
timestamp 1649977179
transform 1 0 26956 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_290
timestamp 1649977179
transform 1 0 27784 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_297
timestamp 1649977179
transform 1 0 28428 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_304
timestamp 1649977179
transform 1 0 29072 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_309
timestamp 1649977179
transform 1 0 29532 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_318
timestamp 1649977179
transform 1 0 30360 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_325
timestamp 1649977179
transform 1 0 31004 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_332
timestamp 1649977179
transform 1 0 31648 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_337
timestamp 1649977179
transform 1 0 32108 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_346
timestamp 1649977179
transform 1 0 32936 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_353
timestamp 1649977179
transform 1 0 33580 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_360
timestamp 1649977179
transform 1 0 34224 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_368
timestamp 1649977179
transform 1 0 34960 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_375
timestamp 1649977179
transform 1 0 35604 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_382 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 36248 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_390 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 36984 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_396
timestamp 1649977179
transform 1 0 37536 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_403
timestamp 1649977179
transform 1 0 38180 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_410
timestamp 1649977179
transform 1 0 38824 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_418
timestamp 1649977179
transform 1 0 39560 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_424
timestamp 1649977179
transform 1 0 40112 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_431
timestamp 1649977179
transform 1 0 40756 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_438
timestamp 1649977179
transform 1 0 41400 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_446
timestamp 1649977179
transform 1 0 42136 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_452
timestamp 1649977179
transform 1 0 42688 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_459
timestamp 1649977179
transform 1 0 43332 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_466
timestamp 1649977179
transform 1 0 43976 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_474
timestamp 1649977179
transform 1 0 44712 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_480
timestamp 1649977179
transform 1 0 45264 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_487
timestamp 1649977179
transform 1 0 45908 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_494
timestamp 1649977179
transform 1 0 46552 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_502
timestamp 1649977179
transform 1 0 47288 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_508
timestamp 1649977179
transform 1 0 47840 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_515
timestamp 1649977179
transform 1 0 48484 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_522
timestamp 1649977179
transform 1 0 49128 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_530
timestamp 1649977179
transform 1 0 49864 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_536
timestamp 1649977179
transform 1 0 50416 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_543
timestamp 1649977179
transform 1 0 51060 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_550
timestamp 1649977179
transform 1 0 51704 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_558
timestamp 1649977179
transform 1 0 52440 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_564
timestamp 1649977179
transform 1 0 52992 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_571
timestamp 1649977179
transform 1 0 53636 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_578
timestamp 1649977179
transform 1 0 54280 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_586
timestamp 1649977179
transform 1 0 55016 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_592
timestamp 1649977179
transform 1 0 55568 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_599
timestamp 1649977179
transform 1 0 56212 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_606
timestamp 1649977179
transform 1 0 56856 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_614
timestamp 1649977179
transform 1 0 57592 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_620
timestamp 1649977179
transform 1 0 58144 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_627
timestamp 1649977179
transform 1 0 58788 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_634
timestamp 1649977179
transform 1 0 59432 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_642
timestamp 1649977179
transform 1 0 60168 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_648
timestamp 1649977179
transform 1 0 60720 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_655
timestamp 1649977179
transform 1 0 61364 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_662
timestamp 1649977179
transform 1 0 62008 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_670
timestamp 1649977179
transform 1 0 62744 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_676
timestamp 1649977179
transform 1 0 63296 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_683
timestamp 1649977179
transform 1 0 63940 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_695
timestamp 1649977179
transform 1 0 65044 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_699
timestamp 1649977179
transform 1 0 65412 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_701
timestamp 1649977179
transform 1 0 65596 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_713
timestamp 1649977179
transform 1 0 66700 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_724
timestamp 1649977179
transform 1 0 67712 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_729
timestamp 1649977179
transform 1 0 68172 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1649977179
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_15
timestamp 1649977179
transform 1 0 2484 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_23
timestamp 1649977179
transform 1 0 3220 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_26
timestamp 1649977179
transform 1 0 3496 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_32
timestamp 1649977179
transform 1 0 4048 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_38
timestamp 1649977179
transform 1 0 4600 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_44
timestamp 1649977179
transform 1 0 5152 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_52
timestamp 1649977179
transform 1 0 5888 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_61
timestamp 1649977179
transform 1 0 6716 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_81
timestamp 1649977179
transform 1 0 8556 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_85
timestamp 1649977179
transform 1 0 8924 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_102
timestamp 1649977179
transform 1 0 10488 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_108
timestamp 1649977179
transform 1 0 11040 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_117
timestamp 1649977179
transform 1 0 11868 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_131
timestamp 1649977179
transform 1 0 13156 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_151
timestamp 1649977179
transform 1 0 14996 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_159
timestamp 1649977179
transform 1 0 15732 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1649977179
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_173
timestamp 1649977179
transform 1 0 17020 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_181
timestamp 1649977179
transform 1 0 17756 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_192
timestamp 1649977179
transform 1 0 18768 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_199
timestamp 1649977179
transform 1 0 19412 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_206
timestamp 1649977179
transform 1 0 20056 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_213
timestamp 1649977179
transform 1 0 20700 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_220
timestamp 1649977179
transform 1 0 21344 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_227
timestamp 1649977179
transform 1 0 21988 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_234
timestamp 1649977179
transform 1 0 22632 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_241
timestamp 1649977179
transform 1 0 23276 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_248
timestamp 1649977179
transform 1 0 23920 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_255
timestamp 1649977179
transform 1 0 24564 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_262
timestamp 1649977179
transform 1 0 25208 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_269
timestamp 1649977179
transform 1 0 25852 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_276
timestamp 1649977179
transform 1 0 26496 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_281
timestamp 1649977179
transform 1 0 26956 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_290
timestamp 1649977179
transform 1 0 27784 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_297
timestamp 1649977179
transform 1 0 28428 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_304
timestamp 1649977179
transform 1 0 29072 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_311
timestamp 1649977179
transform 1 0 29716 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_318
timestamp 1649977179
transform 1 0 30360 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_325
timestamp 1649977179
transform 1 0 31004 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_332
timestamp 1649977179
transform 1 0 31648 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_337
timestamp 1649977179
transform 1 0 32108 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_346
timestamp 1649977179
transform 1 0 32936 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_353
timestamp 1649977179
transform 1 0 33580 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_360
timestamp 1649977179
transform 1 0 34224 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_367
timestamp 1649977179
transform 1 0 34868 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_1_376
timestamp 1649977179
transform 1 0 35696 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_1_385
timestamp 1649977179
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 1649977179
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_396
timestamp 1649977179
transform 1 0 37536 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_403
timestamp 1649977179
transform 1 0 38180 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_410
timestamp 1649977179
transform 1 0 38824 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_417
timestamp 1649977179
transform 1 0 39468 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_424
timestamp 1649977179
transform 1 0 40112 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_431
timestamp 1649977179
transform 1 0 40756 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_438
timestamp 1649977179
transform 1 0 41400 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_446
timestamp 1649977179
transform 1 0 42136 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_452
timestamp 1649977179
transform 1 0 42688 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_459
timestamp 1649977179
transform 1 0 43332 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_466
timestamp 1649977179
transform 1 0 43976 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_473
timestamp 1649977179
transform 1 0 44620 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_480
timestamp 1649977179
transform 1 0 45264 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_487
timestamp 1649977179
transform 1 0 45908 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_494
timestamp 1649977179
transform 1 0 46552 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_502
timestamp 1649977179
transform 1 0 47288 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_508
timestamp 1649977179
transform 1 0 47840 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_515
timestamp 1649977179
transform 1 0 48484 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_522
timestamp 1649977179
transform 1 0 49128 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_529
timestamp 1649977179
transform 1 0 49772 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_536
timestamp 1649977179
transform 1 0 50416 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_543
timestamp 1649977179
transform 1 0 51060 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_550
timestamp 1649977179
transform 1 0 51704 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_558
timestamp 1649977179
transform 1 0 52440 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_564
timestamp 1649977179
transform 1 0 52992 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_571
timestamp 1649977179
transform 1 0 53636 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_578
timestamp 1649977179
transform 1 0 54280 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_585
timestamp 1649977179
transform 1 0 54924 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_592
timestamp 1649977179
transform 1 0 55568 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_599
timestamp 1649977179
transform 1 0 56212 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_606
timestamp 1649977179
transform 1 0 56856 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_614
timestamp 1649977179
transform 1 0 57592 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_620
timestamp 1649977179
transform 1 0 58144 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_627
timestamp 1649977179
transform 1 0 58788 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_634
timestamp 1649977179
transform 1 0 59432 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_641
timestamp 1649977179
transform 1 0 60076 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_648
timestamp 1649977179
transform 1 0 60720 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_655
timestamp 1649977179
transform 1 0 61364 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_662
timestamp 1649977179
transform 1 0 62008 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_670
timestamp 1649977179
transform 1 0 62744 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_676
timestamp 1649977179
transform 1 0 63296 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_688
timestamp 1649977179
transform 1 0 64400 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_700
timestamp 1649977179
transform 1 0 65504 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_712
timestamp 1649977179
transform 1 0 66608 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_724
timestamp 1649977179
transform 1 0 67712 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_729
timestamp 1649977179
transform 1 0 68172 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_3
timestamp 1649977179
transform 1 0 1380 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_11
timestamp 1649977179
transform 1 0 2116 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_14
timestamp 1649977179
transform 1 0 2392 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_20
timestamp 1649977179
transform 1 0 2944 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_29
timestamp 1649977179
transform 1 0 3772 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_34
timestamp 1649977179
transform 1 0 4232 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_40
timestamp 1649977179
transform 1 0 4784 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_60
timestamp 1649977179
transform 1 0 6624 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_67
timestamp 1649977179
transform 1 0 7268 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_76
timestamp 1649977179
transform 1 0 8096 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_88
timestamp 1649977179
transform 1 0 9200 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_108
timestamp 1649977179
transform 1 0 11040 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_117
timestamp 1649977179
transform 1 0 11868 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_123
timestamp 1649977179
transform 1 0 12420 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_128
timestamp 1649977179
transform 1 0 12880 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_136
timestamp 1649977179
transform 1 0 13616 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_141
timestamp 1649977179
transform 1 0 14076 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_147
timestamp 1649977179
transform 1 0 14628 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_155
timestamp 1649977179
transform 1 0 15364 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_161
timestamp 1649977179
transform 1 0 15916 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_175
timestamp 1649977179
transform 1 0 17204 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_181
timestamp 1649977179
transform 1 0 17756 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_185
timestamp 1649977179
transform 1 0 18124 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_192
timestamp 1649977179
transform 1 0 18768 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_207
timestamp 1649977179
transform 1 0 20148 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_214
timestamp 1649977179
transform 1 0 20792 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_222
timestamp 1649977179
transform 1 0 21528 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_226
timestamp 1649977179
transform 1 0 21896 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_2_235
timestamp 1649977179
transform 1 0 22724 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_243
timestamp 1649977179
transform 1 0 23460 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_247
timestamp 1649977179
transform 1 0 23828 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1649977179
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_256
timestamp 1649977179
transform 1 0 24656 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_2_265
timestamp 1649977179
transform 1 0 25484 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_2_274
timestamp 1649977179
transform 1 0 26312 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_2_283
timestamp 1649977179
transform 1 0 27140 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_2_292
timestamp 1649977179
transform 1 0 27968 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_300
timestamp 1649977179
transform 1 0 28704 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_304
timestamp 1649977179
transform 1 0 29072 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_309
timestamp 1649977179
transform 1 0 29532 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_316
timestamp 1649977179
transform 1 0 30176 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_2_325
timestamp 1649977179
transform 1 0 31004 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_2_334
timestamp 1649977179
transform 1 0 31832 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_2_343
timestamp 1649977179
transform 1 0 32660 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_2_352
timestamp 1649977179
transform 1 0 33488 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1649977179
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_377
timestamp 1649977179
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_389
timestamp 1649977179
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_401
timestamp 1649977179
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_413
timestamp 1649977179
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp 1649977179
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_424
timestamp 1649977179
transform 1 0 40112 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_431
timestamp 1649977179
transform 1 0 40756 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_438
timestamp 1649977179
transform 1 0 41400 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_445
timestamp 1649977179
transform 1 0 42044 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_454
timestamp 1649977179
transform 1 0 42872 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_461
timestamp 1649977179
transform 1 0 43516 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_473
timestamp 1649977179
transform 1 0 44620 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_477
timestamp 1649977179
transform 1 0 44988 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_481
timestamp 1649977179
transform 1 0 45356 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_488
timestamp 1649977179
transform 1 0 46000 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_495
timestamp 1649977179
transform 1 0 46644 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_502
timestamp 1649977179
transform 1 0 47288 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_2_511
timestamp 1649977179
transform 1 0 48116 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_519
timestamp 1649977179
transform 1 0 48852 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_523
timestamp 1649977179
transform 1 0 49220 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_531
timestamp 1649977179
transform 1 0 49956 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_533
timestamp 1649977179
transform 1 0 50140 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_538
timestamp 1649977179
transform 1 0 50600 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_545
timestamp 1649977179
transform 1 0 51244 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_552
timestamp 1649977179
transform 1 0 51888 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_560
timestamp 1649977179
transform 1 0 52624 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_565
timestamp 1649977179
transform 1 0 53084 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_572
timestamp 1649977179
transform 1 0 53728 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_584
timestamp 1649977179
transform 1 0 54832 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_592
timestamp 1649977179
transform 1 0 55568 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_599
timestamp 1649977179
transform 1 0 56212 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_606
timestamp 1649977179
transform 1 0 56856 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_613
timestamp 1649977179
transform 1 0 57500 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_620
timestamp 1649977179
transform 1 0 58144 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_627
timestamp 1649977179
transform 1 0 58788 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_634
timestamp 1649977179
transform 1 0 59432 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_642
timestamp 1649977179
transform 1 0 60168 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_648
timestamp 1649977179
transform 1 0 60720 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_655
timestamp 1649977179
transform 1 0 61364 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_662
timestamp 1649977179
transform 1 0 62008 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_674
timestamp 1649977179
transform 1 0 63112 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_686
timestamp 1649977179
transform 1 0 64216 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_698
timestamp 1649977179
transform 1 0 65320 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_701
timestamp 1649977179
transform 1 0 65596 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_713
timestamp 1649977179
transform 1 0 66700 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_725
timestamp 1649977179
transform 1 0 67804 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_3
timestamp 1649977179
transform 1 0 1380 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_7
timestamp 1649977179
transform 1 0 1748 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_16
timestamp 1649977179
transform 1 0 2576 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_36
timestamp 1649977179
transform 1 0 4416 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_40
timestamp 1649977179
transform 1 0 4784 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_43
timestamp 1649977179
transform 1 0 5060 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_52
timestamp 1649977179
transform 1 0 5888 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_65
timestamp 1649977179
transform 1 0 7084 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_72
timestamp 1649977179
transform 1 0 7728 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_80
timestamp 1649977179
transform 1 0 8464 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_88
timestamp 1649977179
transform 1 0 9200 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_96
timestamp 1649977179
transform 1 0 9936 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_108
timestamp 1649977179
transform 1 0 11040 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_115
timestamp 1649977179
transform 1 0 11684 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_135
timestamp 1649977179
transform 1 0 13524 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_143
timestamp 1649977179
transform 1 0 14260 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_151
timestamp 1649977179
transform 1 0 14996 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_159
timestamp 1649977179
transform 1 0 15732 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1649977179
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_181
timestamp 1649977179
transform 1 0 17756 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_190
timestamp 1649977179
transform 1 0 18584 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_197
timestamp 1649977179
transform 1 0 19228 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_204
timestamp 1649977179
transform 1 0 19872 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_220
timestamp 1649977179
transform 1 0 21344 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_225
timestamp 1649977179
transform 1 0 21804 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_234
timestamp 1649977179
transform 1 0 22632 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_3_258
timestamp 1649977179
transform 1 0 24840 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_266
timestamp 1649977179
transform 1 0 25576 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1649977179
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1649977179
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_297
timestamp 1649977179
transform 1 0 28428 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_306
timestamp 1649977179
transform 1 0 29256 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_3_330
timestamp 1649977179
transform 1 0 31464 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1649977179
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_349
timestamp 1649977179
transform 1 0 33212 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_353
timestamp 1649977179
transform 1 0 33580 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_356
timestamp 1649977179
transform 1 0 33856 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_380
timestamp 1649977179
transform 1 0 36064 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1649977179
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_405
timestamp 1649977179
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_417
timestamp 1649977179
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_429
timestamp 1649977179
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_441
timestamp 1649977179
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 1649977179
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_449
timestamp 1649977179
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_461
timestamp 1649977179
transform 1 0 43516 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_473
timestamp 1649977179
transform 1 0 44620 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_485
timestamp 1649977179
transform 1 0 45724 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_497
timestamp 1649977179
transform 1 0 46828 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_503
timestamp 1649977179
transform 1 0 47380 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_505
timestamp 1649977179
transform 1 0 47564 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_517
timestamp 1649977179
transform 1 0 48668 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_529
timestamp 1649977179
transform 1 0 49772 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_541
timestamp 1649977179
transform 1 0 50876 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_553
timestamp 1649977179
transform 1 0 51980 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_559
timestamp 1649977179
transform 1 0 52532 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_561
timestamp 1649977179
transform 1 0 52716 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_573
timestamp 1649977179
transform 1 0 53820 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_585
timestamp 1649977179
transform 1 0 54924 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_597
timestamp 1649977179
transform 1 0 56028 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_602
timestamp 1649977179
transform 1 0 56488 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_609
timestamp 1649977179
transform 1 0 57132 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_615
timestamp 1649977179
transform 1 0 57684 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_620
timestamp 1649977179
transform 1 0 58144 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_627
timestamp 1649977179
transform 1 0 58788 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_634
timestamp 1649977179
transform 1 0 59432 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_641
timestamp 1649977179
transform 1 0 60076 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_648
timestamp 1649977179
transform 1 0 60720 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_655
timestamp 1649977179
transform 1 0 61364 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_667
timestamp 1649977179
transform 1 0 62468 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_671
timestamp 1649977179
transform 1 0 62836 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_673
timestamp 1649977179
transform 1 0 63020 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_685
timestamp 1649977179
transform 1 0 64124 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_697
timestamp 1649977179
transform 1 0 65228 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_709
timestamp 1649977179
transform 1 0 66332 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_724
timestamp 1649977179
transform 1 0 67712 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_729
timestamp 1649977179
transform 1 0 68172 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_3
timestamp 1649977179
transform 1 0 1380 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_12
timestamp 1649977179
transform 1 0 2208 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_21
timestamp 1649977179
transform 1 0 3036 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1649977179
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_31
timestamp 1649977179
transform 1 0 3956 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_39
timestamp 1649977179
transform 1 0 4692 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_42
timestamp 1649977179
transform 1 0 4968 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_48
timestamp 1649977179
transform 1 0 5520 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_54
timestamp 1649977179
transform 1 0 6072 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_60
timestamp 1649977179
transform 1 0 6624 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_80
timestamp 1649977179
transform 1 0 8464 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_88
timestamp 1649977179
transform 1 0 9200 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_96
timestamp 1649977179
transform 1 0 9936 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_104
timestamp 1649977179
transform 1 0 10672 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_112
timestamp 1649977179
transform 1 0 11408 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_125
timestamp 1649977179
transform 1 0 12604 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_131
timestamp 1649977179
transform 1 0 13156 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_136
timestamp 1649977179
transform 1 0 13616 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_157
timestamp 1649977179
transform 1 0 15548 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_165
timestamp 1649977179
transform 1 0 16284 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_169
timestamp 1649977179
transform 1 0 16652 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_192
timestamp 1649977179
transform 1 0 18768 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_207
timestamp 1649977179
transform 1 0 20148 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_214
timestamp 1649977179
transform 1 0 20792 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_221
timestamp 1649977179
transform 1 0 21436 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_229
timestamp 1649977179
transform 1 0 22172 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_238
timestamp 1649977179
transform 1 0 23000 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_248
timestamp 1649977179
transform 1 0 23920 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_261
timestamp 1649977179
transform 1 0 25116 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_275
timestamp 1649977179
transform 1 0 26404 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_281
timestamp 1649977179
transform 1 0 26956 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_289
timestamp 1649977179
transform 1 0 27692 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_292
timestamp 1649977179
transform 1 0 27968 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_304
timestamp 1649977179
transform 1 0 29072 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_317
timestamp 1649977179
transform 1 0 30268 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_329
timestamp 1649977179
transform 1 0 31372 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_349
timestamp 1649977179
transform 1 0 33212 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_361
timestamp 1649977179
transform 1 0 34316 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1649977179
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_377
timestamp 1649977179
transform 1 0 35788 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_381
timestamp 1649977179
transform 1 0 36156 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_385
timestamp 1649977179
transform 1 0 36524 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_392
timestamp 1649977179
transform 1 0 37168 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_404
timestamp 1649977179
transform 1 0 38272 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_416
timestamp 1649977179
transform 1 0 39376 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_421
timestamp 1649977179
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_433
timestamp 1649977179
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_445
timestamp 1649977179
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_457
timestamp 1649977179
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_469
timestamp 1649977179
transform 1 0 44252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 1649977179
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_477
timestamp 1649977179
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_489
timestamp 1649977179
transform 1 0 46092 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_501
timestamp 1649977179
transform 1 0 47196 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_513
timestamp 1649977179
transform 1 0 48300 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_525
timestamp 1649977179
transform 1 0 49404 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_531
timestamp 1649977179
transform 1 0 49956 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_533
timestamp 1649977179
transform 1 0 50140 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_545
timestamp 1649977179
transform 1 0 51244 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_557
timestamp 1649977179
transform 1 0 52348 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_569
timestamp 1649977179
transform 1 0 53452 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_581
timestamp 1649977179
transform 1 0 54556 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_587
timestamp 1649977179
transform 1 0 55108 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_589
timestamp 1649977179
transform 1 0 55292 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_601
timestamp 1649977179
transform 1 0 56396 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_609
timestamp 1649977179
transform 1 0 57132 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_613
timestamp 1649977179
transform 1 0 57500 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_620
timestamp 1649977179
transform 1 0 58144 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_627
timestamp 1649977179
transform 1 0 58788 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_634
timestamp 1649977179
transform 1 0 59432 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_642
timestamp 1649977179
transform 1 0 60168 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_648
timestamp 1649977179
transform 1 0 60720 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_660
timestamp 1649977179
transform 1 0 61824 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_672
timestamp 1649977179
transform 1 0 62928 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_684
timestamp 1649977179
transform 1 0 64032 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_696
timestamp 1649977179
transform 1 0 65136 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_701
timestamp 1649977179
transform 1 0 65596 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_713
timestamp 1649977179
transform 1 0 66700 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_725
timestamp 1649977179
transform 1 0 67804 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_3
timestamp 1649977179
transform 1 0 1380 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_7
timestamp 1649977179
transform 1 0 1748 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_16
timestamp 1649977179
transform 1 0 2576 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_22
timestamp 1649977179
transform 1 0 3128 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_28
timestamp 1649977179
transform 1 0 3680 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_48
timestamp 1649977179
transform 1 0 5520 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_62
timestamp 1649977179
transform 1 0 6808 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_66
timestamp 1649977179
transform 1 0 7176 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_72
timestamp 1649977179
transform 1 0 7728 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_81
timestamp 1649977179
transform 1 0 8556 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_88
timestamp 1649977179
transform 1 0 9200 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_108
timestamp 1649977179
transform 1 0 11040 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_122
timestamp 1649977179
transform 1 0 12328 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_128
timestamp 1649977179
transform 1 0 12880 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_136
timestamp 1649977179
transform 1 0 13616 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_148
timestamp 1649977179
transform 1 0 14720 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_158
timestamp 1649977179
transform 1 0 15640 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_164
timestamp 1649977179
transform 1 0 16192 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_179
timestamp 1649977179
transform 1 0 17572 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_190
timestamp 1649977179
transform 1 0 18584 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_204
timestamp 1649977179
transform 1 0 19872 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_220
timestamp 1649977179
transform 1 0 21344 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_5_225
timestamp 1649977179
transform 1 0 21804 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_230
timestamp 1649977179
transform 1 0 22264 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_250
timestamp 1649977179
transform 1 0 24104 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_254
timestamp 1649977179
transform 1 0 24472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_260
timestamp 1649977179
transform 1 0 25024 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_276
timestamp 1649977179
transform 1 0 26496 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_283
timestamp 1649977179
transform 1 0 27140 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_295
timestamp 1649977179
transform 1 0 28244 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_303
timestamp 1649977179
transform 1 0 28980 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_309
timestamp 1649977179
transform 1 0 29532 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_317
timestamp 1649977179
transform 1 0 30268 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_326
timestamp 1649977179
transform 1 0 31096 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_334
timestamp 1649977179
transform 1 0 31832 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1649977179
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_361
timestamp 1649977179
transform 1 0 34316 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_368
timestamp 1649977179
transform 1 0 34960 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_380
timestamp 1649977179
transform 1 0 36064 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_384
timestamp 1649977179
transform 1 0 36432 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_5_393
timestamp 1649977179
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_405
timestamp 1649977179
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_417
timestamp 1649977179
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_429
timestamp 1649977179
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_441
timestamp 1649977179
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1649977179
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_449
timestamp 1649977179
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_461
timestamp 1649977179
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_473
timestamp 1649977179
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_485
timestamp 1649977179
transform 1 0 45724 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_497
timestamp 1649977179
transform 1 0 46828 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_503
timestamp 1649977179
transform 1 0 47380 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_505
timestamp 1649977179
transform 1 0 47564 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_517
timestamp 1649977179
transform 1 0 48668 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_529
timestamp 1649977179
transform 1 0 49772 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_541
timestamp 1649977179
transform 1 0 50876 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_553
timestamp 1649977179
transform 1 0 51980 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_559
timestamp 1649977179
transform 1 0 52532 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_561
timestamp 1649977179
transform 1 0 52716 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_573
timestamp 1649977179
transform 1 0 53820 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_585
timestamp 1649977179
transform 1 0 54924 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_597
timestamp 1649977179
transform 1 0 56028 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_609
timestamp 1649977179
transform 1 0 57132 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_615
timestamp 1649977179
transform 1 0 57684 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_617
timestamp 1649977179
transform 1 0 57868 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_625
timestamp 1649977179
transform 1 0 58604 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_630
timestamp 1649977179
transform 1 0 59064 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_637
timestamp 1649977179
transform 1 0 59708 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_644
timestamp 1649977179
transform 1 0 60352 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_656
timestamp 1649977179
transform 1 0 61456 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_668
timestamp 1649977179
transform 1 0 62560 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_673
timestamp 1649977179
transform 1 0 63020 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_685
timestamp 1649977179
transform 1 0 64124 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_697
timestamp 1649977179
transform 1 0 65228 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_709
timestamp 1649977179
transform 1 0 66332 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_721
timestamp 1649977179
transform 1 0 67436 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_727
timestamp 1649977179
transform 1 0 67988 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_729
timestamp 1649977179
transform 1 0 68172 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_3
timestamp 1649977179
transform 1 0 1380 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_7
timestamp 1649977179
transform 1 0 1748 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_24
timestamp 1649977179
transform 1 0 3312 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_29
timestamp 1649977179
transform 1 0 3772 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_37
timestamp 1649977179
transform 1 0 4508 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_42
timestamp 1649977179
transform 1 0 4968 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_54
timestamp 1649977179
transform 1 0 6072 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_68
timestamp 1649977179
transform 1 0 7360 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_80
timestamp 1649977179
transform 1 0 8464 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_85
timestamp 1649977179
transform 1 0 8924 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_88
timestamp 1649977179
transform 1 0 9200 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_94
timestamp 1649977179
transform 1 0 9752 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_102
timestamp 1649977179
transform 1 0 10488 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_110
timestamp 1649977179
transform 1 0 11224 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_121
timestamp 1649977179
transform 1 0 12236 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_6_132
timestamp 1649977179
transform 1 0 13248 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_141
timestamp 1649977179
transform 1 0 14076 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_145
timestamp 1649977179
transform 1 0 14444 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_156
timestamp 1649977179
transform 1 0 15456 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_162
timestamp 1649977179
transform 1 0 16008 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_169
timestamp 1649977179
transform 1 0 16652 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_173
timestamp 1649977179
transform 1 0 17020 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_177
timestamp 1649977179
transform 1 0 17388 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_184
timestamp 1649977179
transform 1 0 18032 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_191
timestamp 1649977179
transform 1 0 18676 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1649977179
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_203
timestamp 1649977179
transform 1 0 19780 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_215
timestamp 1649977179
transform 1 0 20884 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1649977179
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1649977179
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1649977179
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1649977179
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_253
timestamp 1649977179
transform 1 0 24380 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_257
timestamp 1649977179
transform 1 0 24748 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_263
timestamp 1649977179
transform 1 0 25300 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_269
timestamp 1649977179
transform 1 0 25852 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_289
timestamp 1649977179
transform 1 0 27692 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_298
timestamp 1649977179
transform 1 0 28520 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_306
timestamp 1649977179
transform 1 0 29256 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1649977179
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_321
timestamp 1649977179
transform 1 0 30636 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_329
timestamp 1649977179
transform 1 0 31372 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_338
timestamp 1649977179
transform 1 0 32200 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_349
timestamp 1649977179
transform 1 0 33212 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_360
timestamp 1649977179
transform 1 0 34224 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1649977179
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_377
timestamp 1649977179
transform 1 0 35788 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_381
timestamp 1649977179
transform 1 0 36156 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_385
timestamp 1649977179
transform 1 0 36524 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_393
timestamp 1649977179
transform 1 0 37260 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_400
timestamp 1649977179
transform 1 0 37904 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_412
timestamp 1649977179
transform 1 0 39008 0 1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_6_421
timestamp 1649977179
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_433
timestamp 1649977179
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_445
timestamp 1649977179
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_457
timestamp 1649977179
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_469
timestamp 1649977179
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 1649977179
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_477
timestamp 1649977179
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_489
timestamp 1649977179
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_501
timestamp 1649977179
transform 1 0 47196 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_513
timestamp 1649977179
transform 1 0 48300 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_525
timestamp 1649977179
transform 1 0 49404 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_531
timestamp 1649977179
transform 1 0 49956 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_533
timestamp 1649977179
transform 1 0 50140 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_545
timestamp 1649977179
transform 1 0 51244 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_557
timestamp 1649977179
transform 1 0 52348 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_569
timestamp 1649977179
transform 1 0 53452 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_581
timestamp 1649977179
transform 1 0 54556 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_587
timestamp 1649977179
transform 1 0 55108 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_589
timestamp 1649977179
transform 1 0 55292 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_601
timestamp 1649977179
transform 1 0 56396 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_613
timestamp 1649977179
transform 1 0 57500 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_625
timestamp 1649977179
transform 1 0 58604 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_637
timestamp 1649977179
transform 1 0 59708 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_643
timestamp 1649977179
transform 1 0 60260 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_645
timestamp 1649977179
transform 1 0 60444 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_657
timestamp 1649977179
transform 1 0 61548 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_669
timestamp 1649977179
transform 1 0 62652 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_681
timestamp 1649977179
transform 1 0 63756 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_693
timestamp 1649977179
transform 1 0 64860 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_699
timestamp 1649977179
transform 1 0 65412 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_701
timestamp 1649977179
transform 1 0 65596 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_713
timestamp 1649977179
transform 1 0 66700 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_725
timestamp 1649977179
transform 1 0 67804 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_729
timestamp 1649977179
transform 1 0 68172 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_3
timestamp 1649977179
transform 1 0 1380 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_12
timestamp 1649977179
transform 1 0 2208 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_16
timestamp 1649977179
transform 1 0 2576 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_33
timestamp 1649977179
transform 1 0 4140 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_45
timestamp 1649977179
transform 1 0 5244 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_49
timestamp 1649977179
transform 1 0 5612 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_52
timestamp 1649977179
transform 1 0 5888 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_57
timestamp 1649977179
transform 1 0 6348 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_61
timestamp 1649977179
transform 1 0 6716 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_65
timestamp 1649977179
transform 1 0 7084 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_68
timestamp 1649977179
transform 1 0 7360 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_77
timestamp 1649977179
transform 1 0 8188 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_89
timestamp 1649977179
transform 1 0 9292 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_93
timestamp 1649977179
transform 1 0 9660 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_96
timestamp 1649977179
transform 1 0 9936 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_102
timestamp 1649977179
transform 1 0 10488 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_108
timestamp 1649977179
transform 1 0 11040 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_120
timestamp 1649977179
transform 1 0 12144 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_134
timestamp 1649977179
transform 1 0 13432 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_138
timestamp 1649977179
transform 1 0 13800 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_147
timestamp 1649977179
transform 1 0 14628 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_159
timestamp 1649977179
transform 1 0 15732 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1649977179
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_169
timestamp 1649977179
transform 1 0 16652 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_186
timestamp 1649977179
transform 1 0 18216 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_190
timestamp 1649977179
transform 1 0 18584 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_199
timestamp 1649977179
transform 1 0 19412 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_206
timestamp 1649977179
transform 1 0 20056 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_212
timestamp 1649977179
transform 1 0 20608 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_218
timestamp 1649977179
transform 1 0 21160 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_235
timestamp 1649977179
transform 1 0 22724 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_244
timestamp 1649977179
transform 1 0 23552 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_252
timestamp 1649977179
transform 1 0 24288 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_260
timestamp 1649977179
transform 1 0 25024 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_267
timestamp 1649977179
transform 1 0 25668 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1649977179
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_281
timestamp 1649977179
transform 1 0 26956 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_289
timestamp 1649977179
transform 1 0 27692 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_301
timestamp 1649977179
transform 1 0 28796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_321
timestamp 1649977179
transform 1 0 30636 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_332
timestamp 1649977179
transform 1 0 31648 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_7_337
timestamp 1649977179
transform 1 0 32108 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_348
timestamp 1649977179
transform 1 0 33120 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_364
timestamp 1649977179
transform 1 0 34592 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_388
timestamp 1649977179
transform 1 0 36800 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_393
timestamp 1649977179
transform 1 0 37260 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_401
timestamp 1649977179
transform 1 0 37996 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_415
timestamp 1649977179
transform 1 0 39284 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_427
timestamp 1649977179
transform 1 0 40388 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_439
timestamp 1649977179
transform 1 0 41492 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1649977179
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_449
timestamp 1649977179
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_461
timestamp 1649977179
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_473
timestamp 1649977179
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_485
timestamp 1649977179
transform 1 0 45724 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_497
timestamp 1649977179
transform 1 0 46828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_503
timestamp 1649977179
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_505
timestamp 1649977179
transform 1 0 47564 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_517
timestamp 1649977179
transform 1 0 48668 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_529
timestamp 1649977179
transform 1 0 49772 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_541
timestamp 1649977179
transform 1 0 50876 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_553
timestamp 1649977179
transform 1 0 51980 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_559
timestamp 1649977179
transform 1 0 52532 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_561
timestamp 1649977179
transform 1 0 52716 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_573
timestamp 1649977179
transform 1 0 53820 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_585
timestamp 1649977179
transform 1 0 54924 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_597
timestamp 1649977179
transform 1 0 56028 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_609
timestamp 1649977179
transform 1 0 57132 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_615
timestamp 1649977179
transform 1 0 57684 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_617
timestamp 1649977179
transform 1 0 57868 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_629
timestamp 1649977179
transform 1 0 58972 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_641
timestamp 1649977179
transform 1 0 60076 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_653
timestamp 1649977179
transform 1 0 61180 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_665
timestamp 1649977179
transform 1 0 62284 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_671
timestamp 1649977179
transform 1 0 62836 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_673
timestamp 1649977179
transform 1 0 63020 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_685
timestamp 1649977179
transform 1 0 64124 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_697
timestamp 1649977179
transform 1 0 65228 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_709
timestamp 1649977179
transform 1 0 66332 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_721
timestamp 1649977179
transform 1 0 67436 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_727
timestamp 1649977179
transform 1 0 67988 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_729
timestamp 1649977179
transform 1 0 68172 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_3
timestamp 1649977179
transform 1 0 1380 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_15
timestamp 1649977179
transform 1 0 2484 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_21
timestamp 1649977179
transform 1 0 3036 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1649977179
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_31
timestamp 1649977179
transform 1 0 3956 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_43
timestamp 1649977179
transform 1 0 5060 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_47
timestamp 1649977179
transform 1 0 5428 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_56
timestamp 1649977179
transform 1 0 6256 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_62
timestamp 1649977179
transform 1 0 6808 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_71
timestamp 1649977179
transform 1 0 7636 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_77
timestamp 1649977179
transform 1 0 8188 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_80
timestamp 1649977179
transform 1 0 8464 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_85
timestamp 1649977179
transform 1 0 8924 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_103
timestamp 1649977179
transform 1 0 10580 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_107
timestamp 1649977179
transform 1 0 10948 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_115
timestamp 1649977179
transform 1 0 11684 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_119
timestamp 1649977179
transform 1 0 12052 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_122
timestamp 1649977179
transform 1 0 12328 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_129
timestamp 1649977179
transform 1 0 12972 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_136
timestamp 1649977179
transform 1 0 13616 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_8_141
timestamp 1649977179
transform 1 0 14076 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_154
timestamp 1649977179
transform 1 0 15272 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_162
timestamp 1649977179
transform 1 0 16008 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_171
timestamp 1649977179
transform 1 0 16836 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_175
timestamp 1649977179
transform 1 0 17204 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_179
timestamp 1649977179
transform 1 0 17572 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_186
timestamp 1649977179
transform 1 0 18216 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_192
timestamp 1649977179
transform 1 0 18768 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_200
timestamp 1649977179
transform 1 0 19504 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_204
timestamp 1649977179
transform 1 0 19872 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_221
timestamp 1649977179
transform 1 0 21436 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_227
timestamp 1649977179
transform 1 0 21988 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_244
timestamp 1649977179
transform 1 0 23552 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_253
timestamp 1649977179
transform 1 0 24380 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_264
timestamp 1649977179
transform 1 0 25392 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_272
timestamp 1649977179
transform 1 0 26128 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_278
timestamp 1649977179
transform 1 0 26680 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_290
timestamp 1649977179
transform 1 0 27784 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_302
timestamp 1649977179
transform 1 0 28888 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_8_309
timestamp 1649977179
transform 1 0 29532 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_315
timestamp 1649977179
transform 1 0 30084 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_322
timestamp 1649977179
transform 1 0 30728 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_340
timestamp 1649977179
transform 1 0 32384 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_352
timestamp 1649977179
transform 1 0 33488 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_373
timestamp 1649977179
transform 1 0 35420 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_385
timestamp 1649977179
transform 1 0 36524 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_397
timestamp 1649977179
transform 1 0 37628 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_409
timestamp 1649977179
transform 1 0 38732 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_417
timestamp 1649977179
transform 1 0 39468 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_421
timestamp 1649977179
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_433
timestamp 1649977179
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_445
timestamp 1649977179
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_457
timestamp 1649977179
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 1649977179
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1649977179
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_477
timestamp 1649977179
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_489
timestamp 1649977179
transform 1 0 46092 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_501
timestamp 1649977179
transform 1 0 47196 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_513
timestamp 1649977179
transform 1 0 48300 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_525
timestamp 1649977179
transform 1 0 49404 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_531
timestamp 1649977179
transform 1 0 49956 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_533
timestamp 1649977179
transform 1 0 50140 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_545
timestamp 1649977179
transform 1 0 51244 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_557
timestamp 1649977179
transform 1 0 52348 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_569
timestamp 1649977179
transform 1 0 53452 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_581
timestamp 1649977179
transform 1 0 54556 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_587
timestamp 1649977179
transform 1 0 55108 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_589
timestamp 1649977179
transform 1 0 55292 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_601
timestamp 1649977179
transform 1 0 56396 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_613
timestamp 1649977179
transform 1 0 57500 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_625
timestamp 1649977179
transform 1 0 58604 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_637
timestamp 1649977179
transform 1 0 59708 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_643
timestamp 1649977179
transform 1 0 60260 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_645
timestamp 1649977179
transform 1 0 60444 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_657
timestamp 1649977179
transform 1 0 61548 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_669
timestamp 1649977179
transform 1 0 62652 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_681
timestamp 1649977179
transform 1 0 63756 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_693
timestamp 1649977179
transform 1 0 64860 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_699
timestamp 1649977179
transform 1 0 65412 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_701
timestamp 1649977179
transform 1 0 65596 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_713
timestamp 1649977179
transform 1 0 66700 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_725
timestamp 1649977179
transform 1 0 67804 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_729
timestamp 1649977179
transform 1 0 68172 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_3
timestamp 1649977179
transform 1 0 1380 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_11
timestamp 1649977179
transform 1 0 2116 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_16
timestamp 1649977179
transform 1 0 2576 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_22
timestamp 1649977179
transform 1 0 3128 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_30
timestamp 1649977179
transform 1 0 3864 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_9_49
timestamp 1649977179
transform 1 0 5612 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1649977179
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_57
timestamp 1649977179
transform 1 0 6348 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_63
timestamp 1649977179
transform 1 0 6900 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_83
timestamp 1649977179
transform 1 0 8740 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_89
timestamp 1649977179
transform 1 0 9292 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_95
timestamp 1649977179
transform 1 0 9844 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_101
timestamp 1649977179
transform 1 0 10396 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_105
timestamp 1649977179
transform 1 0 10764 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_108
timestamp 1649977179
transform 1 0 11040 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_122
timestamp 1649977179
transform 1 0 12328 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_142
timestamp 1649977179
transform 1 0 14168 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_158
timestamp 1649977179
transform 1 0 15640 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_164
timestamp 1649977179
transform 1 0 16192 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_169
timestamp 1649977179
transform 1 0 16652 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_176
timestamp 1649977179
transform 1 0 17296 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_183
timestamp 1649977179
transform 1 0 17940 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_187
timestamp 1649977179
transform 1 0 18308 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_198
timestamp 1649977179
transform 1 0 19320 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_206
timestamp 1649977179
transform 1 0 20056 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_212
timestamp 1649977179
transform 1 0 20608 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_220
timestamp 1649977179
transform 1 0 21344 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_225
timestamp 1649977179
transform 1 0 21804 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_235
timestamp 1649977179
transform 1 0 22724 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_241
timestamp 1649977179
transform 1 0 23276 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_249
timestamp 1649977179
transform 1 0 24012 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_263
timestamp 1649977179
transform 1 0 25300 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_267
timestamp 1649977179
transform 1 0 25668 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_276
timestamp 1649977179
transform 1 0 26496 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_297
timestamp 1649977179
transform 1 0 28428 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_307
timestamp 1649977179
transform 1 0 29348 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_316
timestamp 1649977179
transform 1 0 30176 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_328
timestamp 1649977179
transform 1 0 31280 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_9_337
timestamp 1649977179
transform 1 0 32108 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_343
timestamp 1649977179
transform 1 0 32660 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_346
timestamp 1649977179
transform 1 0 32936 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_358
timestamp 1649977179
transform 1 0 34040 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_364
timestamp 1649977179
transform 1 0 34592 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_381
timestamp 1649977179
transform 1 0 36156 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_389
timestamp 1649977179
transform 1 0 36892 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_395
timestamp 1649977179
transform 1 0 37444 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_407
timestamp 1649977179
transform 1 0 38548 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_419
timestamp 1649977179
transform 1 0 39652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_431
timestamp 1649977179
transform 1 0 40756 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_443
timestamp 1649977179
transform 1 0 41860 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 1649977179
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_449
timestamp 1649977179
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_461
timestamp 1649977179
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_473
timestamp 1649977179
transform 1 0 44620 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_485
timestamp 1649977179
transform 1 0 45724 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_497
timestamp 1649977179
transform 1 0 46828 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_503
timestamp 1649977179
transform 1 0 47380 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_505
timestamp 1649977179
transform 1 0 47564 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_517
timestamp 1649977179
transform 1 0 48668 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_529
timestamp 1649977179
transform 1 0 49772 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_541
timestamp 1649977179
transform 1 0 50876 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_553
timestamp 1649977179
transform 1 0 51980 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_559
timestamp 1649977179
transform 1 0 52532 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_561
timestamp 1649977179
transform 1 0 52716 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_573
timestamp 1649977179
transform 1 0 53820 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_585
timestamp 1649977179
transform 1 0 54924 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_597
timestamp 1649977179
transform 1 0 56028 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_609
timestamp 1649977179
transform 1 0 57132 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_615
timestamp 1649977179
transform 1 0 57684 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_617
timestamp 1649977179
transform 1 0 57868 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_629
timestamp 1649977179
transform 1 0 58972 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_641
timestamp 1649977179
transform 1 0 60076 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_653
timestamp 1649977179
transform 1 0 61180 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_665
timestamp 1649977179
transform 1 0 62284 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_671
timestamp 1649977179
transform 1 0 62836 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_673
timestamp 1649977179
transform 1 0 63020 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_685
timestamp 1649977179
transform 1 0 64124 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_697
timestamp 1649977179
transform 1 0 65228 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_709
timestamp 1649977179
transform 1 0 66332 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_721
timestamp 1649977179
transform 1 0 67436 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_727
timestamp 1649977179
transform 1 0 67988 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_729
timestamp 1649977179
transform 1 0 68172 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_3
timestamp 1649977179
transform 1 0 1380 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_7
timestamp 1649977179
transform 1 0 1748 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_13
timestamp 1649977179
transform 1 0 2300 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_19
timestamp 1649977179
transform 1 0 2852 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1649977179
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1649977179
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_41
timestamp 1649977179
transform 1 0 4876 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_47
timestamp 1649977179
transform 1 0 5428 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_53
timestamp 1649977179
transform 1 0 5980 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_10_69
timestamp 1649977179
transform 1 0 7452 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_79
timestamp 1649977179
transform 1 0 8372 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1649977179
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_87
timestamp 1649977179
transform 1 0 9108 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_99
timestamp 1649977179
transform 1 0 10212 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_107
timestamp 1649977179
transform 1 0 10948 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_125
timestamp 1649977179
transform 1 0 12604 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_133
timestamp 1649977179
transform 1 0 13340 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_136
timestamp 1649977179
transform 1 0 13616 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_141
timestamp 1649977179
transform 1 0 14076 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_151
timestamp 1649977179
transform 1 0 14996 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_158
timestamp 1649977179
transform 1 0 15640 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_170
timestamp 1649977179
transform 1 0 16744 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_180
timestamp 1649977179
transform 1 0 17664 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_192
timestamp 1649977179
transform 1 0 18768 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_197
timestamp 1649977179
transform 1 0 19228 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_219
timestamp 1649977179
transform 1 0 21252 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_233
timestamp 1649977179
transform 1 0 22540 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_239
timestamp 1649977179
transform 1 0 23092 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_242
timestamp 1649977179
transform 1 0 23368 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_248
timestamp 1649977179
transform 1 0 23920 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_253
timestamp 1649977179
transform 1 0 24380 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_256
timestamp 1649977179
transform 1 0 24656 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_268
timestamp 1649977179
transform 1 0 25760 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_274
timestamp 1649977179
transform 1 0 26312 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_286
timestamp 1649977179
transform 1 0 27416 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_294
timestamp 1649977179
transform 1 0 28152 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_302
timestamp 1649977179
transform 1 0 28888 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_309
timestamp 1649977179
transform 1 0 29532 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_326
timestamp 1649977179
transform 1 0 31096 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_336
timestamp 1649977179
transform 1 0 32016 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_360
timestamp 1649977179
transform 1 0 34224 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_365
timestamp 1649977179
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_377
timestamp 1649977179
transform 1 0 35788 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_395
timestamp 1649977179
transform 1 0 37444 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_399
timestamp 1649977179
transform 1 0 37812 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_416
timestamp 1649977179
transform 1 0 39376 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_421
timestamp 1649977179
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_433
timestamp 1649977179
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_445
timestamp 1649977179
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_457
timestamp 1649977179
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_469
timestamp 1649977179
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp 1649977179
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_477
timestamp 1649977179
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_489
timestamp 1649977179
transform 1 0 46092 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_501
timestamp 1649977179
transform 1 0 47196 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_513
timestamp 1649977179
transform 1 0 48300 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_525
timestamp 1649977179
transform 1 0 49404 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_531
timestamp 1649977179
transform 1 0 49956 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_533
timestamp 1649977179
transform 1 0 50140 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_545
timestamp 1649977179
transform 1 0 51244 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_557
timestamp 1649977179
transform 1 0 52348 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_569
timestamp 1649977179
transform 1 0 53452 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_581
timestamp 1649977179
transform 1 0 54556 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_587
timestamp 1649977179
transform 1 0 55108 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_589
timestamp 1649977179
transform 1 0 55292 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_601
timestamp 1649977179
transform 1 0 56396 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_613
timestamp 1649977179
transform 1 0 57500 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_625
timestamp 1649977179
transform 1 0 58604 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_637
timestamp 1649977179
transform 1 0 59708 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_643
timestamp 1649977179
transform 1 0 60260 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_645
timestamp 1649977179
transform 1 0 60444 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_657
timestamp 1649977179
transform 1 0 61548 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_669
timestamp 1649977179
transform 1 0 62652 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_681
timestamp 1649977179
transform 1 0 63756 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_693
timestamp 1649977179
transform 1 0 64860 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_699
timestamp 1649977179
transform 1 0 65412 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_701
timestamp 1649977179
transform 1 0 65596 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_713
timestamp 1649977179
transform 1 0 66700 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_725
timestamp 1649977179
transform 1 0 67804 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_3
timestamp 1649977179
transform 1 0 1380 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_14
timestamp 1649977179
transform 1 0 2392 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_34
timestamp 1649977179
transform 1 0 4232 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_42
timestamp 1649977179
transform 1 0 4968 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_52
timestamp 1649977179
transform 1 0 5888 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_57
timestamp 1649977179
transform 1 0 6348 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_68
timestamp 1649977179
transform 1 0 7360 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_77
timestamp 1649977179
transform 1 0 8188 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_99
timestamp 1649977179
transform 1 0 10212 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1649977179
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1649977179
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1649977179
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1649977179
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_137
timestamp 1649977179
transform 1 0 13708 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_11_149
timestamp 1649977179
transform 1 0 14812 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_158
timestamp 1649977179
transform 1 0 15640 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_164
timestamp 1649977179
transform 1 0 16192 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_185
timestamp 1649977179
transform 1 0 18124 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_191
timestamp 1649977179
transform 1 0 18676 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_200
timestamp 1649977179
transform 1 0 19504 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_208
timestamp 1649977179
transform 1 0 20240 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_220
timestamp 1649977179
transform 1 0 21344 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_225
timestamp 1649977179
transform 1 0 21804 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_243
timestamp 1649977179
transform 1 0 23460 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_255
timestamp 1649977179
transform 1 0 24564 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_11_266
timestamp 1649977179
transform 1 0 25576 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_278
timestamp 1649977179
transform 1 0 26680 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_281
timestamp 1649977179
transform 1 0 26956 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_11_291
timestamp 1649977179
transform 1 0 27876 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_297
timestamp 1649977179
transform 1 0 28428 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_309
timestamp 1649977179
transform 1 0 29532 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_315
timestamp 1649977179
transform 1 0 30084 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_327
timestamp 1649977179
transform 1 0 31188 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_332
timestamp 1649977179
transform 1 0 31648 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_353
timestamp 1649977179
transform 1 0 33580 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_360
timestamp 1649977179
transform 1 0 34224 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_364
timestamp 1649977179
transform 1 0 34592 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_370
timestamp 1649977179
transform 1 0 35144 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_382
timestamp 1649977179
transform 1 0 36248 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_388
timestamp 1649977179
transform 1 0 36800 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_393
timestamp 1649977179
transform 1 0 37260 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_402
timestamp 1649977179
transform 1 0 38088 0 -1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_11_426
timestamp 1649977179
transform 1 0 40296 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_438
timestamp 1649977179
transform 1 0 41400 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_446
timestamp 1649977179
transform 1 0 42136 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_449
timestamp 1649977179
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_461
timestamp 1649977179
transform 1 0 43516 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_473
timestamp 1649977179
transform 1 0 44620 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_485
timestamp 1649977179
transform 1 0 45724 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_497
timestamp 1649977179
transform 1 0 46828 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_503
timestamp 1649977179
transform 1 0 47380 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_505
timestamp 1649977179
transform 1 0 47564 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_517
timestamp 1649977179
transform 1 0 48668 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_529
timestamp 1649977179
transform 1 0 49772 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_541
timestamp 1649977179
transform 1 0 50876 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_553
timestamp 1649977179
transform 1 0 51980 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_559
timestamp 1649977179
transform 1 0 52532 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_561
timestamp 1649977179
transform 1 0 52716 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_573
timestamp 1649977179
transform 1 0 53820 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_585
timestamp 1649977179
transform 1 0 54924 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_597
timestamp 1649977179
transform 1 0 56028 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_609
timestamp 1649977179
transform 1 0 57132 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_615
timestamp 1649977179
transform 1 0 57684 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_617
timestamp 1649977179
transform 1 0 57868 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_629
timestamp 1649977179
transform 1 0 58972 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_641
timestamp 1649977179
transform 1 0 60076 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_653
timestamp 1649977179
transform 1 0 61180 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_665
timestamp 1649977179
transform 1 0 62284 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_671
timestamp 1649977179
transform 1 0 62836 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_673
timestamp 1649977179
transform 1 0 63020 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_685
timestamp 1649977179
transform 1 0 64124 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_697
timestamp 1649977179
transform 1 0 65228 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_709
timestamp 1649977179
transform 1 0 66332 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_724
timestamp 1649977179
transform 1 0 67712 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_729
timestamp 1649977179
transform 1 0 68172 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_3
timestamp 1649977179
transform 1 0 1380 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_14
timestamp 1649977179
transform 1 0 2392 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_20
timestamp 1649977179
transform 1 0 2944 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_12_45
timestamp 1649977179
transform 1 0 5244 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_51
timestamp 1649977179
transform 1 0 5796 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_62
timestamp 1649977179
transform 1 0 6808 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_68
timestamp 1649977179
transform 1 0 7360 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_80
timestamp 1649977179
transform 1 0 8464 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_95
timestamp 1649977179
transform 1 0 9844 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_102
timestamp 1649977179
transform 1 0 10488 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_12_110
timestamp 1649977179
transform 1 0 11224 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_116
timestamp 1649977179
transform 1 0 11776 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1649977179
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1649977179
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_141
timestamp 1649977179
transform 1 0 14076 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_145
timestamp 1649977179
transform 1 0 14444 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_162
timestamp 1649977179
transform 1 0 16008 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_174
timestamp 1649977179
transform 1 0 17112 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_177
timestamp 1649977179
transform 1 0 17388 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1649977179
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1649977179
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_202
timestamp 1649977179
transform 1 0 19688 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_212
timestamp 1649977179
transform 1 0 20608 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_220
timestamp 1649977179
transform 1 0 21344 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_228
timestamp 1649977179
transform 1 0 22080 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_232
timestamp 1649977179
transform 1 0 22448 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_236
timestamp 1649977179
transform 1 0 22816 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_242
timestamp 1649977179
transform 1 0 23368 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_248
timestamp 1649977179
transform 1 0 23920 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_258
timestamp 1649977179
transform 1 0 24840 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_266
timestamp 1649977179
transform 1 0 25576 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_283
timestamp 1649977179
transform 1 0 27140 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_303
timestamp 1649977179
transform 1 0 28980 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1649977179
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_314
timestamp 1649977179
transform 1 0 29992 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_318
timestamp 1649977179
transform 1 0 30360 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_329
timestamp 1649977179
transform 1 0 31372 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_341
timestamp 1649977179
transform 1 0 32476 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_345
timestamp 1649977179
transform 1 0 32844 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_354
timestamp 1649977179
transform 1 0 33672 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_360
timestamp 1649977179
transform 1 0 34224 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_365
timestamp 1649977179
transform 1 0 34684 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_369
timestamp 1649977179
transform 1 0 35052 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_381
timestamp 1649977179
transform 1 0 36156 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_385
timestamp 1649977179
transform 1 0 36524 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_388
timestamp 1649977179
transform 1 0 36800 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_400
timestamp 1649977179
transform 1 0 37904 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_409
timestamp 1649977179
transform 1 0 38732 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_415
timestamp 1649977179
transform 1 0 39284 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_419
timestamp 1649977179
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_421
timestamp 1649977179
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_433
timestamp 1649977179
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_445
timestamp 1649977179
transform 1 0 42044 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_457
timestamp 1649977179
transform 1 0 43148 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_469
timestamp 1649977179
transform 1 0 44252 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 1649977179
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_477
timestamp 1649977179
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_489
timestamp 1649977179
transform 1 0 46092 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_501
timestamp 1649977179
transform 1 0 47196 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_513
timestamp 1649977179
transform 1 0 48300 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_525
timestamp 1649977179
transform 1 0 49404 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_531
timestamp 1649977179
transform 1 0 49956 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_533
timestamp 1649977179
transform 1 0 50140 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_545
timestamp 1649977179
transform 1 0 51244 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_557
timestamp 1649977179
transform 1 0 52348 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_569
timestamp 1649977179
transform 1 0 53452 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_581
timestamp 1649977179
transform 1 0 54556 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_587
timestamp 1649977179
transform 1 0 55108 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_589
timestamp 1649977179
transform 1 0 55292 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_601
timestamp 1649977179
transform 1 0 56396 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_613
timestamp 1649977179
transform 1 0 57500 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_625
timestamp 1649977179
transform 1 0 58604 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_637
timestamp 1649977179
transform 1 0 59708 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_643
timestamp 1649977179
transform 1 0 60260 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_645
timestamp 1649977179
transform 1 0 60444 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_657
timestamp 1649977179
transform 1 0 61548 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_669
timestamp 1649977179
transform 1 0 62652 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_681
timestamp 1649977179
transform 1 0 63756 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_693
timestamp 1649977179
transform 1 0 64860 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_699
timestamp 1649977179
transform 1 0 65412 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_701
timestamp 1649977179
transform 1 0 65596 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_713
timestamp 1649977179
transform 1 0 66700 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_725
timestamp 1649977179
transform 1 0 67804 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1649977179
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1649977179
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_27
timestamp 1649977179
transform 1 0 3588 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_37
timestamp 1649977179
transform 1 0 4508 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_43
timestamp 1649977179
transform 1 0 5060 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_52
timestamp 1649977179
transform 1 0 5888 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_67
timestamp 1649977179
transform 1 0 7268 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_73
timestamp 1649977179
transform 1 0 7820 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_88
timestamp 1649977179
transform 1 0 9200 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_97
timestamp 1649977179
transform 1 0 10028 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_108
timestamp 1649977179
transform 1 0 11040 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_121
timestamp 1649977179
transform 1 0 12236 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_144
timestamp 1649977179
transform 1 0 14352 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_157
timestamp 1649977179
transform 1 0 15548 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_165
timestamp 1649977179
transform 1 0 16284 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_176
timestamp 1649977179
transform 1 0 17296 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_184
timestamp 1649977179
transform 1 0 18032 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_194
timestamp 1649977179
transform 1 0 18952 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_203
timestamp 1649977179
transform 1 0 19780 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_13_216
timestamp 1649977179
transform 1 0 20976 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_225
timestamp 1649977179
transform 1 0 21804 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_234
timestamp 1649977179
transform 1 0 22632 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_247
timestamp 1649977179
transform 1 0 23828 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_267
timestamp 1649977179
transform 1 0 25668 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_273
timestamp 1649977179
transform 1 0 26220 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_276
timestamp 1649977179
transform 1 0 26496 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_281
timestamp 1649977179
transform 1 0 26956 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_292
timestamp 1649977179
transform 1 0 27968 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_300
timestamp 1649977179
transform 1 0 28704 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_312
timestamp 1649977179
transform 1 0 29808 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_320
timestamp 1649977179
transform 1 0 30544 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_332
timestamp 1649977179
transform 1 0 31648 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_337
timestamp 1649977179
transform 1 0 32108 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_351
timestamp 1649977179
transform 1 0 33396 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_355
timestamp 1649977179
transform 1 0 33764 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_364
timestamp 1649977179
transform 1 0 34592 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_376
timestamp 1649977179
transform 1 0 35696 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_382
timestamp 1649977179
transform 1 0 36248 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_388
timestamp 1649977179
transform 1 0 36800 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_393
timestamp 1649977179
transform 1 0 37260 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_405
timestamp 1649977179
transform 1 0 38364 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_13_427
timestamp 1649977179
transform 1 0 40388 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_439
timestamp 1649977179
transform 1 0 41492 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_447
timestamp 1649977179
transform 1 0 42228 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_449
timestamp 1649977179
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_461
timestamp 1649977179
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_473
timestamp 1649977179
transform 1 0 44620 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_485
timestamp 1649977179
transform 1 0 45724 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_497
timestamp 1649977179
transform 1 0 46828 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_503
timestamp 1649977179
transform 1 0 47380 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_505
timestamp 1649977179
transform 1 0 47564 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_517
timestamp 1649977179
transform 1 0 48668 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_529
timestamp 1649977179
transform 1 0 49772 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_541
timestamp 1649977179
transform 1 0 50876 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_553
timestamp 1649977179
transform 1 0 51980 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_559
timestamp 1649977179
transform 1 0 52532 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_561
timestamp 1649977179
transform 1 0 52716 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_573
timestamp 1649977179
transform 1 0 53820 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_585
timestamp 1649977179
transform 1 0 54924 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_597
timestamp 1649977179
transform 1 0 56028 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_609
timestamp 1649977179
transform 1 0 57132 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_615
timestamp 1649977179
transform 1 0 57684 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_617
timestamp 1649977179
transform 1 0 57868 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_629
timestamp 1649977179
transform 1 0 58972 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_641
timestamp 1649977179
transform 1 0 60076 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_653
timestamp 1649977179
transform 1 0 61180 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_665
timestamp 1649977179
transform 1 0 62284 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_671
timestamp 1649977179
transform 1 0 62836 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_673
timestamp 1649977179
transform 1 0 63020 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_685
timestamp 1649977179
transform 1 0 64124 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_697
timestamp 1649977179
transform 1 0 65228 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_709
timestamp 1649977179
transform 1 0 66332 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_721
timestamp 1649977179
transform 1 0 67436 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_727
timestamp 1649977179
transform 1 0 67988 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_729
timestamp 1649977179
transform 1 0 68172 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1649977179
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1649977179
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1649977179
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_45
timestamp 1649977179
transform 1 0 5244 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_57
timestamp 1649977179
transform 1 0 6348 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_61
timestamp 1649977179
transform 1 0 6716 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_65
timestamp 1649977179
transform 1 0 7084 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1649977179
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1649977179
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_90
timestamp 1649977179
transform 1 0 9384 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_99
timestamp 1649977179
transform 1 0 10212 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_113
timestamp 1649977179
transform 1 0 11500 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_122
timestamp 1649977179
transform 1 0 12328 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_134
timestamp 1649977179
transform 1 0 13432 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_148
timestamp 1649977179
transform 1 0 14720 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_154
timestamp 1649977179
transform 1 0 15272 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_169
timestamp 1649977179
transform 1 0 16652 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_175
timestamp 1649977179
transform 1 0 17204 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1649977179
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1649977179
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_197
timestamp 1649977179
transform 1 0 19228 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_215
timestamp 1649977179
transform 1 0 20884 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_224
timestamp 1649977179
transform 1 0 21712 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_230
timestamp 1649977179
transform 1 0 22264 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_236
timestamp 1649977179
transform 1 0 22816 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_240
timestamp 1649977179
transform 1 0 23184 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1649977179
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1649977179
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_253
timestamp 1649977179
transform 1 0 24380 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_259
timestamp 1649977179
transform 1 0 24932 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_262
timestamp 1649977179
transform 1 0 25208 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_268
timestamp 1649977179
transform 1 0 25760 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_277
timestamp 1649977179
transform 1 0 26588 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_286
timestamp 1649977179
transform 1 0 27416 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_293
timestamp 1649977179
transform 1 0 28060 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_304
timestamp 1649977179
transform 1 0 29072 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_316
timestamp 1649977179
transform 1 0 30176 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_322
timestamp 1649977179
transform 1 0 30728 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_331
timestamp 1649977179
transform 1 0 31556 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_335
timestamp 1649977179
transform 1 0 31924 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_346
timestamp 1649977179
transform 1 0 32936 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_355
timestamp 1649977179
transform 1 0 33764 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1649977179
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_370
timestamp 1649977179
transform 1 0 35144 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_376
timestamp 1649977179
transform 1 0 35696 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_384
timestamp 1649977179
transform 1 0 36432 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_387
timestamp 1649977179
transform 1 0 36708 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_399
timestamp 1649977179
transform 1 0 37812 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_405
timestamp 1649977179
transform 1 0 38364 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_417
timestamp 1649977179
transform 1 0 39468 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_421
timestamp 1649977179
transform 1 0 39836 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_429
timestamp 1649977179
transform 1 0 40572 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_432
timestamp 1649977179
transform 1 0 40848 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_444
timestamp 1649977179
transform 1 0 41952 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_456
timestamp 1649977179
transform 1 0 43056 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_468
timestamp 1649977179
transform 1 0 44160 0 1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_14_477
timestamp 1649977179
transform 1 0 44988 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_489
timestamp 1649977179
transform 1 0 46092 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_501
timestamp 1649977179
transform 1 0 47196 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_513
timestamp 1649977179
transform 1 0 48300 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_525
timestamp 1649977179
transform 1 0 49404 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_531
timestamp 1649977179
transform 1 0 49956 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_533
timestamp 1649977179
transform 1 0 50140 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_545
timestamp 1649977179
transform 1 0 51244 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_557
timestamp 1649977179
transform 1 0 52348 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_569
timestamp 1649977179
transform 1 0 53452 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_581
timestamp 1649977179
transform 1 0 54556 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_587
timestamp 1649977179
transform 1 0 55108 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_589
timestamp 1649977179
transform 1 0 55292 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_601
timestamp 1649977179
transform 1 0 56396 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_613
timestamp 1649977179
transform 1 0 57500 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_625
timestamp 1649977179
transform 1 0 58604 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_637
timestamp 1649977179
transform 1 0 59708 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_643
timestamp 1649977179
transform 1 0 60260 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_645
timestamp 1649977179
transform 1 0 60444 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_657
timestamp 1649977179
transform 1 0 61548 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_669
timestamp 1649977179
transform 1 0 62652 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_681
timestamp 1649977179
transform 1 0 63756 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_693
timestamp 1649977179
transform 1 0 64860 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_699
timestamp 1649977179
transform 1 0 65412 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_701
timestamp 1649977179
transform 1 0 65596 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_713
timestamp 1649977179
transform 1 0 66700 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_725
timestamp 1649977179
transform 1 0 67804 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_729
timestamp 1649977179
transform 1 0 68172 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_10
timestamp 1649977179
transform 1 0 2024 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_16
timestamp 1649977179
transform 1 0 2576 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_28
timestamp 1649977179
transform 1 0 3680 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_36
timestamp 1649977179
transform 1 0 4416 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_40
timestamp 1649977179
transform 1 0 4784 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_52
timestamp 1649977179
transform 1 0 5888 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_57
timestamp 1649977179
transform 1 0 6348 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_61
timestamp 1649977179
transform 1 0 6716 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_81
timestamp 1649977179
transform 1 0 8556 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_88
timestamp 1649977179
transform 1 0 9200 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_100
timestamp 1649977179
transform 1 0 10304 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_106
timestamp 1649977179
transform 1 0 10856 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_113
timestamp 1649977179
transform 1 0 11500 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_125
timestamp 1649977179
transform 1 0 12604 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_15_147
timestamp 1649977179
transform 1 0 14628 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_155
timestamp 1649977179
transform 1 0 15364 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1649977179
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_169
timestamp 1649977179
transform 1 0 16652 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_173
timestamp 1649977179
transform 1 0 17020 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_176
timestamp 1649977179
transform 1 0 17296 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_184
timestamp 1649977179
transform 1 0 18032 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_195
timestamp 1649977179
transform 1 0 19044 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_207
timestamp 1649977179
transform 1 0 20148 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_220
timestamp 1649977179
transform 1 0 21344 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_225
timestamp 1649977179
transform 1 0 21804 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_232
timestamp 1649977179
transform 1 0 22448 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_238
timestamp 1649977179
transform 1 0 23000 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_241
timestamp 1649977179
transform 1 0 23276 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_247
timestamp 1649977179
transform 1 0 23828 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_264
timestamp 1649977179
transform 1 0 25392 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_276
timestamp 1649977179
transform 1 0 26496 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_281
timestamp 1649977179
transform 1 0 26956 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_287
timestamp 1649977179
transform 1 0 27508 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_295
timestamp 1649977179
transform 1 0 28244 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_15_309
timestamp 1649977179
transform 1 0 29532 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_315
timestamp 1649977179
transform 1 0 30084 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_319
timestamp 1649977179
transform 1 0 30452 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_331
timestamp 1649977179
transform 1 0 31556 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1649977179
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_344
timestamp 1649977179
transform 1 0 32752 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_350
timestamp 1649977179
transform 1 0 33304 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_359
timestamp 1649977179
transform 1 0 34132 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_363
timestamp 1649977179
transform 1 0 34500 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_380
timestamp 1649977179
transform 1 0 36064 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_387
timestamp 1649977179
transform 1 0 36708 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1649977179
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_393
timestamp 1649977179
transform 1 0 37260 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_397
timestamp 1649977179
transform 1 0 37628 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_408
timestamp 1649977179
transform 1 0 38640 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_428
timestamp 1649977179
transform 1 0 40480 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_438
timestamp 1649977179
transform 1 0 41400 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_446
timestamp 1649977179
transform 1 0 42136 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_449
timestamp 1649977179
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_461
timestamp 1649977179
transform 1 0 43516 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_473
timestamp 1649977179
transform 1 0 44620 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_485
timestamp 1649977179
transform 1 0 45724 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_497
timestamp 1649977179
transform 1 0 46828 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_503
timestamp 1649977179
transform 1 0 47380 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_505
timestamp 1649977179
transform 1 0 47564 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_517
timestamp 1649977179
transform 1 0 48668 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_529
timestamp 1649977179
transform 1 0 49772 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_541
timestamp 1649977179
transform 1 0 50876 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_553
timestamp 1649977179
transform 1 0 51980 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_559
timestamp 1649977179
transform 1 0 52532 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_561
timestamp 1649977179
transform 1 0 52716 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_573
timestamp 1649977179
transform 1 0 53820 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_585
timestamp 1649977179
transform 1 0 54924 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_597
timestamp 1649977179
transform 1 0 56028 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_609
timestamp 1649977179
transform 1 0 57132 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_615
timestamp 1649977179
transform 1 0 57684 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_617
timestamp 1649977179
transform 1 0 57868 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_629
timestamp 1649977179
transform 1 0 58972 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_641
timestamp 1649977179
transform 1 0 60076 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_653
timestamp 1649977179
transform 1 0 61180 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_665
timestamp 1649977179
transform 1 0 62284 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_671
timestamp 1649977179
transform 1 0 62836 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_673
timestamp 1649977179
transform 1 0 63020 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_685
timestamp 1649977179
transform 1 0 64124 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_697
timestamp 1649977179
transform 1 0 65228 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_709
timestamp 1649977179
transform 1 0 66332 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_721
timestamp 1649977179
transform 1 0 67436 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_727
timestamp 1649977179
transform 1 0 67988 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_729
timestamp 1649977179
transform 1 0 68172 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_3
timestamp 1649977179
transform 1 0 1380 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_13
timestamp 1649977179
transform 1 0 2300 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_19
timestamp 1649977179
transform 1 0 2852 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1649977179
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_45
timestamp 1649977179
transform 1 0 5244 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_54
timestamp 1649977179
transform 1 0 6072 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_63
timestamp 1649977179
transform 1 0 6900 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_67
timestamp 1649977179
transform 1 0 7268 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_79
timestamp 1649977179
transform 1 0 8372 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1649977179
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_85
timestamp 1649977179
transform 1 0 8924 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_16_104
timestamp 1649977179
transform 1 0 10672 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_110
timestamp 1649977179
transform 1 0 11224 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_116
timestamp 1649977179
transform 1 0 11776 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_128
timestamp 1649977179
transform 1 0 12880 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_134
timestamp 1649977179
transform 1 0 13432 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_16_141
timestamp 1649977179
transform 1 0 14076 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_147
timestamp 1649977179
transform 1 0 14628 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_157
timestamp 1649977179
transform 1 0 15548 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_16_174
timestamp 1649977179
transform 1 0 17112 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_182
timestamp 1649977179
transform 1 0 17848 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_192
timestamp 1649977179
transform 1 0 18768 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_197
timestamp 1649977179
transform 1 0 19228 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_201
timestamp 1649977179
transform 1 0 19596 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_207
timestamp 1649977179
transform 1 0 20148 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_16_218
timestamp 1649977179
transform 1 0 21160 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_226
timestamp 1649977179
transform 1 0 21896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_232
timestamp 1649977179
transform 1 0 22448 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_240
timestamp 1649977179
transform 1 0 23184 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_248
timestamp 1649977179
transform 1 0 23920 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_260
timestamp 1649977179
transform 1 0 25024 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_16_273
timestamp 1649977179
transform 1 0 26220 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_289
timestamp 1649977179
transform 1 0 27692 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_304
timestamp 1649977179
transform 1 0 29072 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_309
timestamp 1649977179
transform 1 0 29532 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_313
timestamp 1649977179
transform 1 0 29900 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_327
timestamp 1649977179
transform 1 0 31188 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_335
timestamp 1649977179
transform 1 0 31924 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_346
timestamp 1649977179
transform 1 0 32936 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_353
timestamp 1649977179
transform 1 0 33580 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_357
timestamp 1649977179
transform 1 0 33948 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_360
timestamp 1649977179
transform 1 0 34224 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_373
timestamp 1649977179
transform 1 0 35420 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_377
timestamp 1649977179
transform 1 0 35788 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_383
timestamp 1649977179
transform 1 0 36340 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_392
timestamp 1649977179
transform 1 0 37168 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_412
timestamp 1649977179
transform 1 0 39008 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_16_421
timestamp 1649977179
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_433
timestamp 1649977179
transform 1 0 40940 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_445
timestamp 1649977179
transform 1 0 42044 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_457
timestamp 1649977179
transform 1 0 43148 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_469
timestamp 1649977179
transform 1 0 44252 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_475
timestamp 1649977179
transform 1 0 44804 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_477
timestamp 1649977179
transform 1 0 44988 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_489
timestamp 1649977179
transform 1 0 46092 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_501
timestamp 1649977179
transform 1 0 47196 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_513
timestamp 1649977179
transform 1 0 48300 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_525
timestamp 1649977179
transform 1 0 49404 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_531
timestamp 1649977179
transform 1 0 49956 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_533
timestamp 1649977179
transform 1 0 50140 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_545
timestamp 1649977179
transform 1 0 51244 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_557
timestamp 1649977179
transform 1 0 52348 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_569
timestamp 1649977179
transform 1 0 53452 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_581
timestamp 1649977179
transform 1 0 54556 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_587
timestamp 1649977179
transform 1 0 55108 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_589
timestamp 1649977179
transform 1 0 55292 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_601
timestamp 1649977179
transform 1 0 56396 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_613
timestamp 1649977179
transform 1 0 57500 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_625
timestamp 1649977179
transform 1 0 58604 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_637
timestamp 1649977179
transform 1 0 59708 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_643
timestamp 1649977179
transform 1 0 60260 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_645
timestamp 1649977179
transform 1 0 60444 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_657
timestamp 1649977179
transform 1 0 61548 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_669
timestamp 1649977179
transform 1 0 62652 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_681
timestamp 1649977179
transform 1 0 63756 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_693
timestamp 1649977179
transform 1 0 64860 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_699
timestamp 1649977179
transform 1 0 65412 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_701
timestamp 1649977179
transform 1 0 65596 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_713
timestamp 1649977179
transform 1 0 66700 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_725
timestamp 1649977179
transform 1 0 67804 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_3
timestamp 1649977179
transform 1 0 1380 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_13
timestamp 1649977179
transform 1 0 2300 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_22
timestamp 1649977179
transform 1 0 3128 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_28
timestamp 1649977179
transform 1 0 3680 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_34
timestamp 1649977179
transform 1 0 4232 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_46
timestamp 1649977179
transform 1 0 5336 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_52
timestamp 1649977179
transform 1 0 5888 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_62
timestamp 1649977179
transform 1 0 6808 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_68
timestamp 1649977179
transform 1 0 7360 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_88
timestamp 1649977179
transform 1 0 9200 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_100
timestamp 1649977179
transform 1 0 10304 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_108
timestamp 1649977179
transform 1 0 11040 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_118
timestamp 1649977179
transform 1 0 11960 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_124
timestamp 1649977179
transform 1 0 12512 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_130
timestamp 1649977179
transform 1 0 13064 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_153
timestamp 1649977179
transform 1 0 15180 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_162
timestamp 1649977179
transform 1 0 16008 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_178
timestamp 1649977179
transform 1 0 17480 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_184
timestamp 1649977179
transform 1 0 18032 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_190
timestamp 1649977179
transform 1 0 18584 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_200
timestamp 1649977179
transform 1 0 19504 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_208
timestamp 1649977179
transform 1 0 20240 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_216
timestamp 1649977179
transform 1 0 20976 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_225
timestamp 1649977179
transform 1 0 21804 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_237
timestamp 1649977179
transform 1 0 22908 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_248
timestamp 1649977179
transform 1 0 23920 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_256
timestamp 1649977179
transform 1 0 24656 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_262
timestamp 1649977179
transform 1 0 25208 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_268
timestamp 1649977179
transform 1 0 25760 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_276
timestamp 1649977179
transform 1 0 26496 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_281
timestamp 1649977179
transform 1 0 26956 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_293
timestamp 1649977179
transform 1 0 28060 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_299
timestamp 1649977179
transform 1 0 28612 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_305
timestamp 1649977179
transform 1 0 29164 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_17_319
timestamp 1649977179
transform 1 0 30452 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_331
timestamp 1649977179
transform 1 0 31556 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1649977179
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_337
timestamp 1649977179
transform 1 0 32108 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_347
timestamp 1649977179
transform 1 0 33028 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_354
timestamp 1649977179
transform 1 0 33672 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_362
timestamp 1649977179
transform 1 0 34408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_365
timestamp 1649977179
transform 1 0 34684 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_372
timestamp 1649977179
transform 1 0 35328 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_387
timestamp 1649977179
transform 1 0 36708 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1649977179
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_403
timestamp 1649977179
transform 1 0 38180 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_415
timestamp 1649977179
transform 1 0 39284 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_427
timestamp 1649977179
transform 1 0 40388 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_439
timestamp 1649977179
transform 1 0 41492 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_447
timestamp 1649977179
transform 1 0 42228 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_449
timestamp 1649977179
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_461
timestamp 1649977179
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_473
timestamp 1649977179
transform 1 0 44620 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_485
timestamp 1649977179
transform 1 0 45724 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_497
timestamp 1649977179
transform 1 0 46828 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_503
timestamp 1649977179
transform 1 0 47380 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_505
timestamp 1649977179
transform 1 0 47564 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_517
timestamp 1649977179
transform 1 0 48668 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_529
timestamp 1649977179
transform 1 0 49772 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_541
timestamp 1649977179
transform 1 0 50876 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_553
timestamp 1649977179
transform 1 0 51980 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_559
timestamp 1649977179
transform 1 0 52532 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_561
timestamp 1649977179
transform 1 0 52716 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_573
timestamp 1649977179
transform 1 0 53820 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_585
timestamp 1649977179
transform 1 0 54924 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_597
timestamp 1649977179
transform 1 0 56028 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_609
timestamp 1649977179
transform 1 0 57132 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_615
timestamp 1649977179
transform 1 0 57684 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_617
timestamp 1649977179
transform 1 0 57868 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_629
timestamp 1649977179
transform 1 0 58972 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_641
timestamp 1649977179
transform 1 0 60076 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_653
timestamp 1649977179
transform 1 0 61180 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_665
timestamp 1649977179
transform 1 0 62284 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_671
timestamp 1649977179
transform 1 0 62836 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_673
timestamp 1649977179
transform 1 0 63020 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_685
timestamp 1649977179
transform 1 0 64124 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_697
timestamp 1649977179
transform 1 0 65228 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_709
timestamp 1649977179
transform 1 0 66332 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_724
timestamp 1649977179
transform 1 0 67712 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_729
timestamp 1649977179
transform 1 0 68172 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_3
timestamp 1649977179
transform 1 0 1380 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_11
timestamp 1649977179
transform 1 0 2116 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_23
timestamp 1649977179
transform 1 0 3220 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1649977179
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_31
timestamp 1649977179
transform 1 0 3956 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_51
timestamp 1649977179
transform 1 0 5796 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_63
timestamp 1649977179
transform 1 0 6900 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_75
timestamp 1649977179
transform 1 0 8004 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1649977179
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_87
timestamp 1649977179
transform 1 0 9108 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_102
timestamp 1649977179
transform 1 0 10488 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_111
timestamp 1649977179
transform 1 0 11316 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_123
timestamp 1649977179
transform 1 0 12420 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1649977179
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1649977179
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_151
timestamp 1649977179
transform 1 0 14996 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_162
timestamp 1649977179
transform 1 0 16008 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_170
timestamp 1649977179
transform 1 0 16744 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_176
timestamp 1649977179
transform 1 0 17296 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_183
timestamp 1649977179
transform 1 0 17940 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1649977179
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1649977179
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_197
timestamp 1649977179
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_209
timestamp 1649977179
transform 1 0 20332 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_216
timestamp 1649977179
transform 1 0 20976 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_224
timestamp 1649977179
transform 1 0 21712 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_231
timestamp 1649977179
transform 1 0 22356 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_239
timestamp 1649977179
transform 1 0 23092 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_245
timestamp 1649977179
transform 1 0 23644 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_248
timestamp 1649977179
transform 1 0 23920 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_256
timestamp 1649977179
transform 1 0 24656 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_271
timestamp 1649977179
transform 1 0 26036 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_277
timestamp 1649977179
transform 1 0 26588 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_283
timestamp 1649977179
transform 1 0 27140 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_294
timestamp 1649977179
transform 1 0 28152 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_302
timestamp 1649977179
transform 1 0 28888 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_309
timestamp 1649977179
transform 1 0 29532 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_317
timestamp 1649977179
transform 1 0 30268 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_325
timestamp 1649977179
transform 1 0 31004 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_335
timestamp 1649977179
transform 1 0 31924 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_351
timestamp 1649977179
transform 1 0 33396 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_359
timestamp 1649977179
transform 1 0 34132 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1649977179
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_381
timestamp 1649977179
transform 1 0 36156 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_385
timestamp 1649977179
transform 1 0 36524 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_394
timestamp 1649977179
transform 1 0 37352 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_398
timestamp 1649977179
transform 1 0 37720 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_407
timestamp 1649977179
transform 1 0 38548 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_419
timestamp 1649977179
transform 1 0 39652 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_437
timestamp 1649977179
transform 1 0 41308 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_449
timestamp 1649977179
transform 1 0 42412 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_461
timestamp 1649977179
transform 1 0 43516 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_473
timestamp 1649977179
transform 1 0 44620 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_477
timestamp 1649977179
transform 1 0 44988 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_489
timestamp 1649977179
transform 1 0 46092 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_501
timestamp 1649977179
transform 1 0 47196 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_513
timestamp 1649977179
transform 1 0 48300 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_525
timestamp 1649977179
transform 1 0 49404 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_531
timestamp 1649977179
transform 1 0 49956 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_533
timestamp 1649977179
transform 1 0 50140 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_545
timestamp 1649977179
transform 1 0 51244 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_557
timestamp 1649977179
transform 1 0 52348 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_569
timestamp 1649977179
transform 1 0 53452 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_581
timestamp 1649977179
transform 1 0 54556 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_587
timestamp 1649977179
transform 1 0 55108 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_589
timestamp 1649977179
transform 1 0 55292 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_601
timestamp 1649977179
transform 1 0 56396 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_613
timestamp 1649977179
transform 1 0 57500 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_625
timestamp 1649977179
transform 1 0 58604 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_637
timestamp 1649977179
transform 1 0 59708 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_643
timestamp 1649977179
transform 1 0 60260 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_645
timestamp 1649977179
transform 1 0 60444 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_657
timestamp 1649977179
transform 1 0 61548 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_669
timestamp 1649977179
transform 1 0 62652 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_681
timestamp 1649977179
transform 1 0 63756 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_693
timestamp 1649977179
transform 1 0 64860 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_699
timestamp 1649977179
transform 1 0 65412 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_701
timestamp 1649977179
transform 1 0 65596 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_713
timestamp 1649977179
transform 1 0 66700 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_725
timestamp 1649977179
transform 1 0 67804 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3
timestamp 1649977179
transform 1 0 1380 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_7
timestamp 1649977179
transform 1 0 1748 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_16
timestamp 1649977179
transform 1 0 2576 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_20
timestamp 1649977179
transform 1 0 2944 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_37
timestamp 1649977179
transform 1 0 4508 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_49
timestamp 1649977179
transform 1 0 5612 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1649977179
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_57
timestamp 1649977179
transform 1 0 6348 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_65
timestamp 1649977179
transform 1 0 7084 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_73
timestamp 1649977179
transform 1 0 7820 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_79
timestamp 1649977179
transform 1 0 8372 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_91
timestamp 1649977179
transform 1 0 9476 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_100
timestamp 1649977179
transform 1 0 10304 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_108
timestamp 1649977179
transform 1 0 11040 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_117
timestamp 1649977179
transform 1 0 11868 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_125
timestamp 1649977179
transform 1 0 12604 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_129
timestamp 1649977179
transform 1 0 12972 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_146
timestamp 1649977179
transform 1 0 14536 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_150
timestamp 1649977179
transform 1 0 14904 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_153
timestamp 1649977179
transform 1 0 15180 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_157
timestamp 1649977179
transform 1 0 15548 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_164
timestamp 1649977179
transform 1 0 16192 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_169
timestamp 1649977179
transform 1 0 16652 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_189
timestamp 1649977179
transform 1 0 18492 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_195
timestamp 1649977179
transform 1 0 19044 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_212
timestamp 1649977179
transform 1 0 20608 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_230
timestamp 1649977179
transform 1 0 22264 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_238
timestamp 1649977179
transform 1 0 23000 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_246
timestamp 1649977179
transform 1 0 23736 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_260
timestamp 1649977179
transform 1 0 25024 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_272
timestamp 1649977179
transform 1 0 26128 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_287
timestamp 1649977179
transform 1 0 27508 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_291
timestamp 1649977179
transform 1 0 27876 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_302
timestamp 1649977179
transform 1 0 28888 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_316
timestamp 1649977179
transform 1 0 30176 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_320
timestamp 1649977179
transform 1 0 30544 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 1649977179
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1649977179
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_337
timestamp 1649977179
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_349
timestamp 1649977179
transform 1 0 33212 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_355
timestamp 1649977179
transform 1 0 33764 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_367
timestamp 1649977179
transform 1 0 34868 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_375
timestamp 1649977179
transform 1 0 35604 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_388
timestamp 1649977179
transform 1 0 36800 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_393
timestamp 1649977179
transform 1 0 37260 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_401
timestamp 1649977179
transform 1 0 37996 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_407
timestamp 1649977179
transform 1 0 38548 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_419
timestamp 1649977179
transform 1 0 39652 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_427
timestamp 1649977179
transform 1 0 40388 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_432
timestamp 1649977179
transform 1 0 40848 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_439
timestamp 1649977179
transform 1 0 41492 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_447
timestamp 1649977179
transform 1 0 42228 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_449
timestamp 1649977179
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_461
timestamp 1649977179
transform 1 0 43516 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_473
timestamp 1649977179
transform 1 0 44620 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_485
timestamp 1649977179
transform 1 0 45724 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_497
timestamp 1649977179
transform 1 0 46828 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_503
timestamp 1649977179
transform 1 0 47380 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_505
timestamp 1649977179
transform 1 0 47564 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_517
timestamp 1649977179
transform 1 0 48668 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_529
timestamp 1649977179
transform 1 0 49772 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_541
timestamp 1649977179
transform 1 0 50876 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_553
timestamp 1649977179
transform 1 0 51980 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_559
timestamp 1649977179
transform 1 0 52532 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_561
timestamp 1649977179
transform 1 0 52716 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_573
timestamp 1649977179
transform 1 0 53820 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_585
timestamp 1649977179
transform 1 0 54924 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_597
timestamp 1649977179
transform 1 0 56028 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_609
timestamp 1649977179
transform 1 0 57132 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_615
timestamp 1649977179
transform 1 0 57684 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_617
timestamp 1649977179
transform 1 0 57868 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_629
timestamp 1649977179
transform 1 0 58972 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_641
timestamp 1649977179
transform 1 0 60076 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_653
timestamp 1649977179
transform 1 0 61180 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_665
timestamp 1649977179
transform 1 0 62284 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_671
timestamp 1649977179
transform 1 0 62836 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_673
timestamp 1649977179
transform 1 0 63020 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_685
timestamp 1649977179
transform 1 0 64124 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_697
timestamp 1649977179
transform 1 0 65228 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_709
timestamp 1649977179
transform 1 0 66332 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_724
timestamp 1649977179
transform 1 0 67712 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_729
timestamp 1649977179
transform 1 0 68172 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1649977179
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_20
timestamp 1649977179
transform 1 0 2944 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_20_31
timestamp 1649977179
transform 1 0 3956 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_43
timestamp 1649977179
transform 1 0 5060 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_55
timestamp 1649977179
transform 1 0 6164 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_61
timestamp 1649977179
transform 1 0 6716 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_78
timestamp 1649977179
transform 1 0 8280 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_20_92
timestamp 1649977179
transform 1 0 9568 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_104
timestamp 1649977179
transform 1 0 10672 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_116
timestamp 1649977179
transform 1 0 11776 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_124
timestamp 1649977179
transform 1 0 12512 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_135
timestamp 1649977179
transform 1 0 13524 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1649977179
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_141
timestamp 1649977179
transform 1 0 14076 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_149
timestamp 1649977179
transform 1 0 14812 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_153
timestamp 1649977179
transform 1 0 15180 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_161
timestamp 1649977179
transform 1 0 15916 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_169
timestamp 1649977179
transform 1 0 16652 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_175
timestamp 1649977179
transform 1 0 17204 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_180
timestamp 1649977179
transform 1 0 17664 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_186
timestamp 1649977179
transform 1 0 18216 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_192
timestamp 1649977179
transform 1 0 18768 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_202
timestamp 1649977179
transform 1 0 19688 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_217
timestamp 1649977179
transform 1 0 21068 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_227
timestamp 1649977179
transform 1 0 21988 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_236
timestamp 1649977179
transform 1 0 22816 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_247
timestamp 1649977179
transform 1 0 23828 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1649977179
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_253
timestamp 1649977179
transform 1 0 24380 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_258
timestamp 1649977179
transform 1 0 24840 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_267
timestamp 1649977179
transform 1 0 25668 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_277
timestamp 1649977179
transform 1 0 26588 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_281
timestamp 1649977179
transform 1 0 26956 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_289
timestamp 1649977179
transform 1 0 27692 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_301
timestamp 1649977179
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1649977179
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_309
timestamp 1649977179
transform 1 0 29532 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_313
timestamp 1649977179
transform 1 0 29900 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_321
timestamp 1649977179
transform 1 0 30636 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_20_336
timestamp 1649977179
transform 1 0 32016 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_348
timestamp 1649977179
transform 1 0 33120 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_356
timestamp 1649977179
transform 1 0 33856 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_360
timestamp 1649977179
transform 1 0 34224 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_365
timestamp 1649977179
transform 1 0 34684 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_376
timestamp 1649977179
transform 1 0 35696 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_386
timestamp 1649977179
transform 1 0 36616 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_399
timestamp 1649977179
transform 1 0 37812 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_405
timestamp 1649977179
transform 1 0 38364 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_417
timestamp 1649977179
transform 1 0 39468 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_437
timestamp 1649977179
transform 1 0 41308 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_449
timestamp 1649977179
transform 1 0 42412 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_461
timestamp 1649977179
transform 1 0 43516 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_473
timestamp 1649977179
transform 1 0 44620 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_477
timestamp 1649977179
transform 1 0 44988 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_489
timestamp 1649977179
transform 1 0 46092 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_501
timestamp 1649977179
transform 1 0 47196 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_513
timestamp 1649977179
transform 1 0 48300 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_525
timestamp 1649977179
transform 1 0 49404 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_531
timestamp 1649977179
transform 1 0 49956 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_533
timestamp 1649977179
transform 1 0 50140 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_545
timestamp 1649977179
transform 1 0 51244 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_557
timestamp 1649977179
transform 1 0 52348 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_569
timestamp 1649977179
transform 1 0 53452 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_581
timestamp 1649977179
transform 1 0 54556 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_587
timestamp 1649977179
transform 1 0 55108 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_589
timestamp 1649977179
transform 1 0 55292 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_601
timestamp 1649977179
transform 1 0 56396 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_613
timestamp 1649977179
transform 1 0 57500 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_625
timestamp 1649977179
transform 1 0 58604 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_637
timestamp 1649977179
transform 1 0 59708 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_643
timestamp 1649977179
transform 1 0 60260 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_645
timestamp 1649977179
transform 1 0 60444 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_657
timestamp 1649977179
transform 1 0 61548 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_669
timestamp 1649977179
transform 1 0 62652 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_681
timestamp 1649977179
transform 1 0 63756 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_693
timestamp 1649977179
transform 1 0 64860 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_699
timestamp 1649977179
transform 1 0 65412 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_701
timestamp 1649977179
transform 1 0 65596 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_713
timestamp 1649977179
transform 1 0 66700 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_725
timestamp 1649977179
transform 1 0 67804 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_10
timestamp 1649977179
transform 1 0 2024 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_14
timestamp 1649977179
transform 1 0 2392 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_23
timestamp 1649977179
transform 1 0 3220 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_43
timestamp 1649977179
transform 1 0 5060 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1649977179
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_73
timestamp 1649977179
transform 1 0 7820 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_79
timestamp 1649977179
transform 1 0 8372 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_87
timestamp 1649977179
transform 1 0 9108 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_101
timestamp 1649977179
transform 1 0 10396 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_109
timestamp 1649977179
transform 1 0 11132 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_123
timestamp 1649977179
transform 1 0 12420 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_137
timestamp 1649977179
transform 1 0 13708 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_145
timestamp 1649977179
transform 1 0 14444 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_153
timestamp 1649977179
transform 1 0 15180 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_159
timestamp 1649977179
transform 1 0 15732 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1649977179
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_169
timestamp 1649977179
transform 1 0 16652 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_181
timestamp 1649977179
transform 1 0 17756 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_190
timestamp 1649977179
transform 1 0 18584 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_198
timestamp 1649977179
transform 1 0 19320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_205
timestamp 1649977179
transform 1 0 19964 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_211
timestamp 1649977179
transform 1 0 20516 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1649977179
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_225
timestamp 1649977179
transform 1 0 21804 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_229
timestamp 1649977179
transform 1 0 22172 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_232
timestamp 1649977179
transform 1 0 22448 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_238
timestamp 1649977179
transform 1 0 23000 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_241
timestamp 1649977179
transform 1 0 23276 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_249
timestamp 1649977179
transform 1 0 24012 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_257
timestamp 1649977179
transform 1 0 24748 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_267
timestamp 1649977179
transform 1 0 25668 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_273
timestamp 1649977179
transform 1 0 26220 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1649977179
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_281
timestamp 1649977179
transform 1 0 26956 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_287
timestamp 1649977179
transform 1 0 27508 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_291
timestamp 1649977179
transform 1 0 27876 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_294
timestamp 1649977179
transform 1 0 28152 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_302
timestamp 1649977179
transform 1 0 28888 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_310
timestamp 1649977179
transform 1 0 29624 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_322
timestamp 1649977179
transform 1 0 30728 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_334
timestamp 1649977179
transform 1 0 31832 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_353
timestamp 1649977179
transform 1 0 33580 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_361
timestamp 1649977179
transform 1 0 34316 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_368
timestamp 1649977179
transform 1 0 34960 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_388
timestamp 1649977179
transform 1 0 36800 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_393
timestamp 1649977179
transform 1 0 37260 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_405
timestamp 1649977179
transform 1 0 38364 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_417
timestamp 1649977179
transform 1 0 39468 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_429
timestamp 1649977179
transform 1 0 40572 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_441
timestamp 1649977179
transform 1 0 41676 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_447
timestamp 1649977179
transform 1 0 42228 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_449
timestamp 1649977179
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_461
timestamp 1649977179
transform 1 0 43516 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_473
timestamp 1649977179
transform 1 0 44620 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_485
timestamp 1649977179
transform 1 0 45724 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_497
timestamp 1649977179
transform 1 0 46828 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_503
timestamp 1649977179
transform 1 0 47380 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_505
timestamp 1649977179
transform 1 0 47564 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_517
timestamp 1649977179
transform 1 0 48668 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_529
timestamp 1649977179
transform 1 0 49772 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_541
timestamp 1649977179
transform 1 0 50876 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_553
timestamp 1649977179
transform 1 0 51980 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_559
timestamp 1649977179
transform 1 0 52532 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_561
timestamp 1649977179
transform 1 0 52716 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_573
timestamp 1649977179
transform 1 0 53820 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_585
timestamp 1649977179
transform 1 0 54924 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_597
timestamp 1649977179
transform 1 0 56028 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_609
timestamp 1649977179
transform 1 0 57132 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_615
timestamp 1649977179
transform 1 0 57684 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_617
timestamp 1649977179
transform 1 0 57868 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_629
timestamp 1649977179
transform 1 0 58972 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_641
timestamp 1649977179
transform 1 0 60076 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_653
timestamp 1649977179
transform 1 0 61180 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_665
timestamp 1649977179
transform 1 0 62284 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_671
timestamp 1649977179
transform 1 0 62836 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_673
timestamp 1649977179
transform 1 0 63020 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_685
timestamp 1649977179
transform 1 0 64124 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_697
timestamp 1649977179
transform 1 0 65228 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_709
timestamp 1649977179
transform 1 0 66332 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_721
timestamp 1649977179
transform 1 0 67436 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_727
timestamp 1649977179
transform 1 0 67988 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_729
timestamp 1649977179
transform 1 0 68172 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_3
timestamp 1649977179
transform 1 0 1380 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_11
timestamp 1649977179
transform 1 0 2116 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_19
timestamp 1649977179
transform 1 0 2852 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1649977179
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1649977179
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_41
timestamp 1649977179
transform 1 0 4876 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_52
timestamp 1649977179
transform 1 0 5888 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_58
timestamp 1649977179
transform 1 0 6440 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_64
timestamp 1649977179
transform 1 0 6992 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_68
timestamp 1649977179
transform 1 0 7360 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_76
timestamp 1649977179
transform 1 0 8096 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_80
timestamp 1649977179
transform 1 0 8464 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_85
timestamp 1649977179
transform 1 0 8924 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_93
timestamp 1649977179
transform 1 0 9660 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_102
timestamp 1649977179
transform 1 0 10488 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_113
timestamp 1649977179
transform 1 0 11500 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_117
timestamp 1649977179
transform 1 0 11868 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_122
timestamp 1649977179
transform 1 0 12328 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_136
timestamp 1649977179
transform 1 0 13616 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_22_141
timestamp 1649977179
transform 1 0 14076 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_152
timestamp 1649977179
transform 1 0 15088 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_166
timestamp 1649977179
transform 1 0 16376 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_180
timestamp 1649977179
transform 1 0 17664 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_188
timestamp 1649977179
transform 1 0 18400 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_192
timestamp 1649977179
transform 1 0 18768 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_201
timestamp 1649977179
transform 1 0 19596 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_209
timestamp 1649977179
transform 1 0 20332 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_212
timestamp 1649977179
transform 1 0 20608 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_220
timestamp 1649977179
transform 1 0 21344 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_224
timestamp 1649977179
transform 1 0 21712 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_227
timestamp 1649977179
transform 1 0 21988 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_233
timestamp 1649977179
transform 1 0 22540 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_22_241
timestamp 1649977179
transform 1 0 23276 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_249
timestamp 1649977179
transform 1 0 24012 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_22_255
timestamp 1649977179
transform 1 0 24564 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_269
timestamp 1649977179
transform 1 0 25852 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_289
timestamp 1649977179
transform 1 0 27692 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_293
timestamp 1649977179
transform 1 0 28060 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_298
timestamp 1649977179
transform 1 0 28520 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_304
timestamp 1649977179
transform 1 0 29072 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_309
timestamp 1649977179
transform 1 0 29532 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_319
timestamp 1649977179
transform 1 0 30452 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_328
timestamp 1649977179
transform 1 0 31280 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_334
timestamp 1649977179
transform 1 0 31832 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_349
timestamp 1649977179
transform 1 0 33212 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_361
timestamp 1649977179
transform 1 0 34316 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_375
timestamp 1649977179
transform 1 0 35604 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_387
timestamp 1649977179
transform 1 0 36708 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_394
timestamp 1649977179
transform 1 0 37352 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_406
timestamp 1649977179
transform 1 0 38456 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_412
timestamp 1649977179
transform 1 0 39008 0 1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_22_421
timestamp 1649977179
transform 1 0 39836 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_433
timestamp 1649977179
transform 1 0 40940 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_445
timestamp 1649977179
transform 1 0 42044 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_457
timestamp 1649977179
transform 1 0 43148 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_469
timestamp 1649977179
transform 1 0 44252 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_475
timestamp 1649977179
transform 1 0 44804 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_477
timestamp 1649977179
transform 1 0 44988 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_489
timestamp 1649977179
transform 1 0 46092 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_501
timestamp 1649977179
transform 1 0 47196 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_513
timestamp 1649977179
transform 1 0 48300 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_525
timestamp 1649977179
transform 1 0 49404 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_531
timestamp 1649977179
transform 1 0 49956 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_533
timestamp 1649977179
transform 1 0 50140 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_545
timestamp 1649977179
transform 1 0 51244 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_557
timestamp 1649977179
transform 1 0 52348 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_569
timestamp 1649977179
transform 1 0 53452 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_581
timestamp 1649977179
transform 1 0 54556 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_587
timestamp 1649977179
transform 1 0 55108 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_589
timestamp 1649977179
transform 1 0 55292 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_601
timestamp 1649977179
transform 1 0 56396 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_613
timestamp 1649977179
transform 1 0 57500 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_625
timestamp 1649977179
transform 1 0 58604 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_637
timestamp 1649977179
transform 1 0 59708 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_643
timestamp 1649977179
transform 1 0 60260 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_645
timestamp 1649977179
transform 1 0 60444 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_657
timestamp 1649977179
transform 1 0 61548 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_669
timestamp 1649977179
transform 1 0 62652 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_681
timestamp 1649977179
transform 1 0 63756 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_693
timestamp 1649977179
transform 1 0 64860 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_699
timestamp 1649977179
transform 1 0 65412 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_701
timestamp 1649977179
transform 1 0 65596 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_713
timestamp 1649977179
transform 1 0 66700 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_725
timestamp 1649977179
transform 1 0 67804 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_729
timestamp 1649977179
transform 1 0 68172 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1649977179
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_15
timestamp 1649977179
transform 1 0 2484 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_19
timestamp 1649977179
transform 1 0 2852 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_25
timestamp 1649977179
transform 1 0 3404 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_31
timestamp 1649977179
transform 1 0 3956 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_39
timestamp 1649977179
transform 1 0 4692 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_47
timestamp 1649977179
transform 1 0 5428 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1649977179
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_57
timestamp 1649977179
transform 1 0 6348 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_61
timestamp 1649977179
transform 1 0 6716 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_64
timestamp 1649977179
transform 1 0 6992 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_76
timestamp 1649977179
transform 1 0 8096 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_82
timestamp 1649977179
transform 1 0 8648 0 -1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_23_93
timestamp 1649977179
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1649977179
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1649977179
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_113
timestamp 1649977179
transform 1 0 11500 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_119
timestamp 1649977179
transform 1 0 12052 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_123
timestamp 1649977179
transform 1 0 12420 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_132
timestamp 1649977179
transform 1 0 13248 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_23_147
timestamp 1649977179
transform 1 0 14628 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_155
timestamp 1649977179
transform 1 0 15364 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_164
timestamp 1649977179
transform 1 0 16192 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_169
timestamp 1649977179
transform 1 0 16652 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_175
timestamp 1649977179
transform 1 0 17204 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_183
timestamp 1649977179
transform 1 0 17940 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_189
timestamp 1649977179
transform 1 0 18492 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_209
timestamp 1649977179
transform 1 0 20332 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_220
timestamp 1649977179
transform 1 0 21344 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_232
timestamp 1649977179
transform 1 0 22448 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_252
timestamp 1649977179
transform 1 0 24288 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_265
timestamp 1649977179
transform 1 0 25484 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_271
timestamp 1649977179
transform 1 0 26036 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 1649977179
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_281
timestamp 1649977179
transform 1 0 26956 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_286
timestamp 1649977179
transform 1 0 27416 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_293
timestamp 1649977179
transform 1 0 28060 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_302
timestamp 1649977179
transform 1 0 28888 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_311
timestamp 1649977179
transform 1 0 29716 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_322
timestamp 1649977179
transform 1 0 30728 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_326
timestamp 1649977179
transform 1 0 31096 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_330
timestamp 1649977179
transform 1 0 31464 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_23_345
timestamp 1649977179
transform 1 0 32844 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_351
timestamp 1649977179
transform 1 0 33396 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_357
timestamp 1649977179
transform 1 0 33948 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_371
timestamp 1649977179
transform 1 0 35236 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_383
timestamp 1649977179
transform 1 0 36340 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_388
timestamp 1649977179
transform 1 0 36800 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_401
timestamp 1649977179
transform 1 0 37996 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_429
timestamp 1649977179
transform 1 0 40572 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_441
timestamp 1649977179
transform 1 0 41676 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_447
timestamp 1649977179
transform 1 0 42228 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_449
timestamp 1649977179
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_461
timestamp 1649977179
transform 1 0 43516 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_473
timestamp 1649977179
transform 1 0 44620 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_485
timestamp 1649977179
transform 1 0 45724 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_497
timestamp 1649977179
transform 1 0 46828 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_503
timestamp 1649977179
transform 1 0 47380 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_505
timestamp 1649977179
transform 1 0 47564 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_517
timestamp 1649977179
transform 1 0 48668 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_529
timestamp 1649977179
transform 1 0 49772 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_541
timestamp 1649977179
transform 1 0 50876 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_553
timestamp 1649977179
transform 1 0 51980 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_559
timestamp 1649977179
transform 1 0 52532 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_561
timestamp 1649977179
transform 1 0 52716 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_573
timestamp 1649977179
transform 1 0 53820 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_585
timestamp 1649977179
transform 1 0 54924 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_597
timestamp 1649977179
transform 1 0 56028 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_609
timestamp 1649977179
transform 1 0 57132 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_615
timestamp 1649977179
transform 1 0 57684 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_617
timestamp 1649977179
transform 1 0 57868 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_629
timestamp 1649977179
transform 1 0 58972 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_641
timestamp 1649977179
transform 1 0 60076 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_653
timestamp 1649977179
transform 1 0 61180 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_665
timestamp 1649977179
transform 1 0 62284 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_671
timestamp 1649977179
transform 1 0 62836 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_673
timestamp 1649977179
transform 1 0 63020 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_685
timestamp 1649977179
transform 1 0 64124 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_697
timestamp 1649977179
transform 1 0 65228 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_709
timestamp 1649977179
transform 1 0 66332 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_721
timestamp 1649977179
transform 1 0 67436 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_727
timestamp 1649977179
transform 1 0 67988 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_729
timestamp 1649977179
transform 1 0 68172 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_3
timestamp 1649977179
transform 1 0 1380 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_12
timestamp 1649977179
transform 1 0 2208 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_22
timestamp 1649977179
transform 1 0 3128 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_24_45
timestamp 1649977179
transform 1 0 5244 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_60
timestamp 1649977179
transform 1 0 6624 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_69
timestamp 1649977179
transform 1 0 7452 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_80
timestamp 1649977179
transform 1 0 8464 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_92
timestamp 1649977179
transform 1 0 9568 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_96
timestamp 1649977179
transform 1 0 9936 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_104
timestamp 1649977179
transform 1 0 10672 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_114
timestamp 1649977179
transform 1 0 11592 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_123
timestamp 1649977179
transform 1 0 12420 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_127
timestamp 1649977179
transform 1 0 12788 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_136
timestamp 1649977179
transform 1 0 13616 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_141
timestamp 1649977179
transform 1 0 14076 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_144
timestamp 1649977179
transform 1 0 14352 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_151
timestamp 1649977179
transform 1 0 14996 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_167
timestamp 1649977179
transform 1 0 16468 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_179
timestamp 1649977179
transform 1 0 17572 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_187
timestamp 1649977179
transform 1 0 18308 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_192
timestamp 1649977179
transform 1 0 18768 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_202
timestamp 1649977179
transform 1 0 19688 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_216
timestamp 1649977179
transform 1 0 20976 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_220
timestamp 1649977179
transform 1 0 21344 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_223
timestamp 1649977179
transform 1 0 21620 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_247
timestamp 1649977179
transform 1 0 23828 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1649977179
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_257
timestamp 1649977179
transform 1 0 24748 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_261
timestamp 1649977179
transform 1 0 25116 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_266
timestamp 1649977179
transform 1 0 25576 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_270
timestamp 1649977179
transform 1 0 25944 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_287
timestamp 1649977179
transform 1 0 27508 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_24_300
timestamp 1649977179
transform 1 0 28704 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_24_317
timestamp 1649977179
transform 1 0 30268 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_323
timestamp 1649977179
transform 1 0 30820 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_326
timestamp 1649977179
transform 1 0 31096 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_340
timestamp 1649977179
transform 1 0 32384 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_344
timestamp 1649977179
transform 1 0 32752 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_353
timestamp 1649977179
transform 1 0 33580 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_357
timestamp 1649977179
transform 1 0 33948 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_360
timestamp 1649977179
transform 1 0 34224 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_370
timestamp 1649977179
transform 1 0 35144 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_390
timestamp 1649977179
transform 1 0 36984 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_398
timestamp 1649977179
transform 1 0 37720 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_416
timestamp 1649977179
transform 1 0 39376 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_421
timestamp 1649977179
transform 1 0 39836 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_433
timestamp 1649977179
transform 1 0 40940 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_445
timestamp 1649977179
transform 1 0 42044 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_457
timestamp 1649977179
transform 1 0 43148 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_469
timestamp 1649977179
transform 1 0 44252 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_475
timestamp 1649977179
transform 1 0 44804 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_477
timestamp 1649977179
transform 1 0 44988 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_489
timestamp 1649977179
transform 1 0 46092 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_501
timestamp 1649977179
transform 1 0 47196 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_513
timestamp 1649977179
transform 1 0 48300 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_525
timestamp 1649977179
transform 1 0 49404 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_531
timestamp 1649977179
transform 1 0 49956 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_533
timestamp 1649977179
transform 1 0 50140 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_545
timestamp 1649977179
transform 1 0 51244 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_557
timestamp 1649977179
transform 1 0 52348 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_569
timestamp 1649977179
transform 1 0 53452 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_581
timestamp 1649977179
transform 1 0 54556 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_587
timestamp 1649977179
transform 1 0 55108 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_589
timestamp 1649977179
transform 1 0 55292 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_601
timestamp 1649977179
transform 1 0 56396 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_613
timestamp 1649977179
transform 1 0 57500 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_625
timestamp 1649977179
transform 1 0 58604 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_637
timestamp 1649977179
transform 1 0 59708 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_643
timestamp 1649977179
transform 1 0 60260 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_645
timestamp 1649977179
transform 1 0 60444 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_657
timestamp 1649977179
transform 1 0 61548 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_669
timestamp 1649977179
transform 1 0 62652 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_681
timestamp 1649977179
transform 1 0 63756 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_693
timestamp 1649977179
transform 1 0 64860 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_699
timestamp 1649977179
transform 1 0 65412 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_701
timestamp 1649977179
transform 1 0 65596 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_713
timestamp 1649977179
transform 1 0 66700 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_725
timestamp 1649977179
transform 1 0 67804 0 1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1649977179
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_15
timestamp 1649977179
transform 1 0 2484 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_19
timestamp 1649977179
transform 1 0 2852 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_28
timestamp 1649977179
transform 1 0 3680 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_34
timestamp 1649977179
transform 1 0 4232 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_46
timestamp 1649977179
transform 1 0 5336 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_52
timestamp 1649977179
transform 1 0 5888 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_57
timestamp 1649977179
transform 1 0 6348 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_66
timestamp 1649977179
transform 1 0 7176 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_78
timestamp 1649977179
transform 1 0 8280 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_86
timestamp 1649977179
transform 1 0 9016 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_92
timestamp 1649977179
transform 1 0 9568 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_100
timestamp 1649977179
transform 1 0 10304 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_108
timestamp 1649977179
transform 1 0 11040 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_123
timestamp 1649977179
transform 1 0 12420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_135
timestamp 1649977179
transform 1 0 13524 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_143
timestamp 1649977179
transform 1 0 14260 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_154
timestamp 1649977179
transform 1 0 15272 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_166
timestamp 1649977179
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1649977179
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_187
timestamp 1649977179
transform 1 0 18308 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_193
timestamp 1649977179
transform 1 0 18860 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_199
timestamp 1649977179
transform 1 0 19412 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_207
timestamp 1649977179
transform 1 0 20148 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_212
timestamp 1649977179
transform 1 0 20608 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_220
timestamp 1649977179
transform 1 0 21344 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_225
timestamp 1649977179
transform 1 0 21804 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_229
timestamp 1649977179
transform 1 0 22172 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_239
timestamp 1649977179
transform 1 0 23092 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_247
timestamp 1649977179
transform 1 0 23828 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_251
timestamp 1649977179
transform 1 0 24196 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_268
timestamp 1649977179
transform 1 0 25760 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_276
timestamp 1649977179
transform 1 0 26496 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_285
timestamp 1649977179
transform 1 0 27324 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_293
timestamp 1649977179
transform 1 0 28060 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_302
timestamp 1649977179
transform 1 0 28888 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_312
timestamp 1649977179
transform 1 0 29808 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_326
timestamp 1649977179
transform 1 0 31096 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_334
timestamp 1649977179
transform 1 0 31832 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_353
timestamp 1649977179
transform 1 0 33580 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_359
timestamp 1649977179
transform 1 0 34132 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_370
timestamp 1649977179
transform 1 0 35144 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_382
timestamp 1649977179
transform 1 0 36248 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_390
timestamp 1649977179
transform 1 0 36984 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_398
timestamp 1649977179
transform 1 0 37720 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_406
timestamp 1649977179
transform 1 0 38456 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_424
timestamp 1649977179
transform 1 0 40112 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_436
timestamp 1649977179
transform 1 0 41216 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_449
timestamp 1649977179
transform 1 0 42412 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_461
timestamp 1649977179
transform 1 0 43516 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_473
timestamp 1649977179
transform 1 0 44620 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_485
timestamp 1649977179
transform 1 0 45724 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_497
timestamp 1649977179
transform 1 0 46828 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_503
timestamp 1649977179
transform 1 0 47380 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_505
timestamp 1649977179
transform 1 0 47564 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_517
timestamp 1649977179
transform 1 0 48668 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_529
timestamp 1649977179
transform 1 0 49772 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_541
timestamp 1649977179
transform 1 0 50876 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_553
timestamp 1649977179
transform 1 0 51980 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_559
timestamp 1649977179
transform 1 0 52532 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_561
timestamp 1649977179
transform 1 0 52716 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_573
timestamp 1649977179
transform 1 0 53820 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_585
timestamp 1649977179
transform 1 0 54924 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_597
timestamp 1649977179
transform 1 0 56028 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_609
timestamp 1649977179
transform 1 0 57132 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_615
timestamp 1649977179
transform 1 0 57684 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_617
timestamp 1649977179
transform 1 0 57868 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_629
timestamp 1649977179
transform 1 0 58972 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_641
timestamp 1649977179
transform 1 0 60076 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_653
timestamp 1649977179
transform 1 0 61180 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_665
timestamp 1649977179
transform 1 0 62284 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_671
timestamp 1649977179
transform 1 0 62836 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_673
timestamp 1649977179
transform 1 0 63020 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_685
timestamp 1649977179
transform 1 0 64124 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_697
timestamp 1649977179
transform 1 0 65228 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_709
timestamp 1649977179
transform 1 0 66332 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_724
timestamp 1649977179
transform 1 0 67712 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_729
timestamp 1649977179
transform 1 0 68172 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_3
timestamp 1649977179
transform 1 0 1380 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_9
timestamp 1649977179
transform 1 0 1932 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_16
timestamp 1649977179
transform 1 0 2576 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_31
timestamp 1649977179
transform 1 0 3956 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_40
timestamp 1649977179
transform 1 0 4784 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_48
timestamp 1649977179
transform 1 0 5520 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_59
timestamp 1649977179
transform 1 0 6532 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_65
timestamp 1649977179
transform 1 0 7084 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_72
timestamp 1649977179
transform 1 0 7728 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_78
timestamp 1649977179
transform 1 0 8280 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_26_101
timestamp 1649977179
transform 1 0 10396 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_107
timestamp 1649977179
transform 1 0 10948 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_116
timestamp 1649977179
transform 1 0 11776 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_136
timestamp 1649977179
transform 1 0 13616 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1649977179
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_153
timestamp 1649977179
transform 1 0 15180 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_157
timestamp 1649977179
transform 1 0 15548 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_163
timestamp 1649977179
transform 1 0 16100 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_169
timestamp 1649977179
transform 1 0 16652 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_181
timestamp 1649977179
transform 1 0 17756 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_193
timestamp 1649977179
transform 1 0 18860 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_205
timestamp 1649977179
transform 1 0 19964 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_225
timestamp 1649977179
transform 1 0 21804 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_233
timestamp 1649977179
transform 1 0 22540 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_26_243
timestamp 1649977179
transform 1 0 23460 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1649977179
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_253
timestamp 1649977179
transform 1 0 24380 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_257
timestamp 1649977179
transform 1 0 24748 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_263
timestamp 1649977179
transform 1 0 25300 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_271
timestamp 1649977179
transform 1 0 26036 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_277
timestamp 1649977179
transform 1 0 26588 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_283
timestamp 1649977179
transform 1 0 27140 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_291
timestamp 1649977179
transform 1 0 27876 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_300
timestamp 1649977179
transform 1 0 28704 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_309
timestamp 1649977179
transform 1 0 29532 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_321
timestamp 1649977179
transform 1 0 30636 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_330
timestamp 1649977179
transform 1 0 31464 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_342
timestamp 1649977179
transform 1 0 32568 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_349
timestamp 1649977179
transform 1 0 33212 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_360
timestamp 1649977179
transform 1 0 34224 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_373
timestamp 1649977179
transform 1 0 35420 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_379
timestamp 1649977179
transform 1 0 35972 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_389
timestamp 1649977179
transform 1 0 36892 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_401
timestamp 1649977179
transform 1 0 37996 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_413
timestamp 1649977179
transform 1 0 39100 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_419
timestamp 1649977179
transform 1 0 39652 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_421
timestamp 1649977179
transform 1 0 39836 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_433
timestamp 1649977179
transform 1 0 40940 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_445
timestamp 1649977179
transform 1 0 42044 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_457
timestamp 1649977179
transform 1 0 43148 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_469
timestamp 1649977179
transform 1 0 44252 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_475
timestamp 1649977179
transform 1 0 44804 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_477
timestamp 1649977179
transform 1 0 44988 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_489
timestamp 1649977179
transform 1 0 46092 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_501
timestamp 1649977179
transform 1 0 47196 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_513
timestamp 1649977179
transform 1 0 48300 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_525
timestamp 1649977179
transform 1 0 49404 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_531
timestamp 1649977179
transform 1 0 49956 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_533
timestamp 1649977179
transform 1 0 50140 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_545
timestamp 1649977179
transform 1 0 51244 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_557
timestamp 1649977179
transform 1 0 52348 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_569
timestamp 1649977179
transform 1 0 53452 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_581
timestamp 1649977179
transform 1 0 54556 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_587
timestamp 1649977179
transform 1 0 55108 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_589
timestamp 1649977179
transform 1 0 55292 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_601
timestamp 1649977179
transform 1 0 56396 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_613
timestamp 1649977179
transform 1 0 57500 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_625
timestamp 1649977179
transform 1 0 58604 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_637
timestamp 1649977179
transform 1 0 59708 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_643
timestamp 1649977179
transform 1 0 60260 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_645
timestamp 1649977179
transform 1 0 60444 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_657
timestamp 1649977179
transform 1 0 61548 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_669
timestamp 1649977179
transform 1 0 62652 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_681
timestamp 1649977179
transform 1 0 63756 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_693
timestamp 1649977179
transform 1 0 64860 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_699
timestamp 1649977179
transform 1 0 65412 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_701
timestamp 1649977179
transform 1 0 65596 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_713
timestamp 1649977179
transform 1 0 66700 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_725
timestamp 1649977179
transform 1 0 67804 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_11
timestamp 1649977179
transform 1 0 2116 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_23
timestamp 1649977179
transform 1 0 3220 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_43
timestamp 1649977179
transform 1 0 5060 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_52
timestamp 1649977179
transform 1 0 5888 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_57
timestamp 1649977179
transform 1 0 6348 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_61
timestamp 1649977179
transform 1 0 6716 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_72
timestamp 1649977179
transform 1 0 7728 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_84
timestamp 1649977179
transform 1 0 8832 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_90
timestamp 1649977179
transform 1 0 9384 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_102
timestamp 1649977179
transform 1 0 10488 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_108
timestamp 1649977179
transform 1 0 11040 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_113
timestamp 1649977179
transform 1 0 11500 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_122
timestamp 1649977179
transform 1 0 12328 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_128
timestamp 1649977179
transform 1 0 12880 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_140
timestamp 1649977179
transform 1 0 13984 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_152
timestamp 1649977179
transform 1 0 15088 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_164
timestamp 1649977179
transform 1 0 16192 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_185
timestamp 1649977179
transform 1 0 18124 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_193
timestamp 1649977179
transform 1 0 18860 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_205
timestamp 1649977179
transform 1 0 19964 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_209
timestamp 1649977179
transform 1 0 20332 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_212
timestamp 1649977179
transform 1 0 20608 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_220
timestamp 1649977179
transform 1 0 21344 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_229
timestamp 1649977179
transform 1 0 22172 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_249
timestamp 1649977179
transform 1 0 24012 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_257
timestamp 1649977179
transform 1 0 24748 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_266
timestamp 1649977179
transform 1 0 25576 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_272
timestamp 1649977179
transform 1 0 26128 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_275
timestamp 1649977179
transform 1 0 26404 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1649977179
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_281
timestamp 1649977179
transform 1 0 26956 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_289
timestamp 1649977179
transform 1 0 27692 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_292
timestamp 1649977179
transform 1 0 27968 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_304
timestamp 1649977179
transform 1 0 29072 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_332
timestamp 1649977179
transform 1 0 31648 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_337
timestamp 1649977179
transform 1 0 32108 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_345
timestamp 1649977179
transform 1 0 32844 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_356
timestamp 1649977179
transform 1 0 33856 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_364
timestamp 1649977179
transform 1 0 34592 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_381
timestamp 1649977179
transform 1 0 36156 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_385
timestamp 1649977179
transform 1 0 36524 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_388
timestamp 1649977179
transform 1 0 36800 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_401
timestamp 1649977179
transform 1 0 37996 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_409
timestamp 1649977179
transform 1 0 38732 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_428
timestamp 1649977179
transform 1 0 40480 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_440
timestamp 1649977179
transform 1 0 41584 0 -1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_27_449
timestamp 1649977179
transform 1 0 42412 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_461
timestamp 1649977179
transform 1 0 43516 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_473
timestamp 1649977179
transform 1 0 44620 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_485
timestamp 1649977179
transform 1 0 45724 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_497
timestamp 1649977179
transform 1 0 46828 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_503
timestamp 1649977179
transform 1 0 47380 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_505
timestamp 1649977179
transform 1 0 47564 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_517
timestamp 1649977179
transform 1 0 48668 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_529
timestamp 1649977179
transform 1 0 49772 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_541
timestamp 1649977179
transform 1 0 50876 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_553
timestamp 1649977179
transform 1 0 51980 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_559
timestamp 1649977179
transform 1 0 52532 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_561
timestamp 1649977179
transform 1 0 52716 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_573
timestamp 1649977179
transform 1 0 53820 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_585
timestamp 1649977179
transform 1 0 54924 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_597
timestamp 1649977179
transform 1 0 56028 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_609
timestamp 1649977179
transform 1 0 57132 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_615
timestamp 1649977179
transform 1 0 57684 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_617
timestamp 1649977179
transform 1 0 57868 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_629
timestamp 1649977179
transform 1 0 58972 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_641
timestamp 1649977179
transform 1 0 60076 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_653
timestamp 1649977179
transform 1 0 61180 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_665
timestamp 1649977179
transform 1 0 62284 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_671
timestamp 1649977179
transform 1 0 62836 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_673
timestamp 1649977179
transform 1 0 63020 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_685
timestamp 1649977179
transform 1 0 64124 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_697
timestamp 1649977179
transform 1 0 65228 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_709
timestamp 1649977179
transform 1 0 66332 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_721
timestamp 1649977179
transform 1 0 67436 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_727
timestamp 1649977179
transform 1 0 67988 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_729
timestamp 1649977179
transform 1 0 68172 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_3
timestamp 1649977179
transform 1 0 1380 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_28_12
timestamp 1649977179
transform 1 0 2208 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_24
timestamp 1649977179
transform 1 0 3312 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1649977179
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_41
timestamp 1649977179
transform 1 0 4876 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_61
timestamp 1649977179
transform 1 0 6716 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_67
timestamp 1649977179
transform 1 0 7268 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_76
timestamp 1649977179
transform 1 0 8096 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_28_90
timestamp 1649977179
transform 1 0 9384 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_28_101
timestamp 1649977179
transform 1 0 10396 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_109
timestamp 1649977179
transform 1 0 11132 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_116
timestamp 1649977179
transform 1 0 11776 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_136
timestamp 1649977179
transform 1 0 13616 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_157
timestamp 1649977179
transform 1 0 15548 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_171
timestamp 1649977179
transform 1 0 16836 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_177
timestamp 1649977179
transform 1 0 17388 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_183
timestamp 1649977179
transform 1 0 17940 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_189
timestamp 1649977179
transform 1 0 18492 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_192
timestamp 1649977179
transform 1 0 18768 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_202
timestamp 1649977179
transform 1 0 19688 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_208
timestamp 1649977179
transform 1 0 20240 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_211
timestamp 1649977179
transform 1 0 20516 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_217
timestamp 1649977179
transform 1 0 21068 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_226
timestamp 1649977179
transform 1 0 21896 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_232
timestamp 1649977179
transform 1 0 22448 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_238
timestamp 1649977179
transform 1 0 23000 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_248
timestamp 1649977179
transform 1 0 23920 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_258
timestamp 1649977179
transform 1 0 24840 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_264
timestamp 1649977179
transform 1 0 25392 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_273
timestamp 1649977179
transform 1 0 26220 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_293
timestamp 1649977179
transform 1 0 28060 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_305
timestamp 1649977179
transform 1 0 29164 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_309
timestamp 1649977179
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_321
timestamp 1649977179
transform 1 0 30636 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_327
timestamp 1649977179
transform 1 0 31188 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_331
timestamp 1649977179
transform 1 0 31556 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_339
timestamp 1649977179
transform 1 0 32292 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_351
timestamp 1649977179
transform 1 0 33396 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1649977179
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_367
timestamp 1649977179
transform 1 0 34868 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_379
timestamp 1649977179
transform 1 0 35972 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_384
timestamp 1649977179
transform 1 0 36432 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_393
timestamp 1649977179
transform 1 0 37260 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_402
timestamp 1649977179
transform 1 0 38088 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_408
timestamp 1649977179
transform 1 0 38640 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_421
timestamp 1649977179
transform 1 0 39836 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_433
timestamp 1649977179
transform 1 0 40940 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_445
timestamp 1649977179
transform 1 0 42044 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_457
timestamp 1649977179
transform 1 0 43148 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_469
timestamp 1649977179
transform 1 0 44252 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_475
timestamp 1649977179
transform 1 0 44804 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_477
timestamp 1649977179
transform 1 0 44988 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_489
timestamp 1649977179
transform 1 0 46092 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_501
timestamp 1649977179
transform 1 0 47196 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_513
timestamp 1649977179
transform 1 0 48300 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_525
timestamp 1649977179
transform 1 0 49404 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_531
timestamp 1649977179
transform 1 0 49956 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_533
timestamp 1649977179
transform 1 0 50140 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_545
timestamp 1649977179
transform 1 0 51244 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_557
timestamp 1649977179
transform 1 0 52348 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_569
timestamp 1649977179
transform 1 0 53452 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_581
timestamp 1649977179
transform 1 0 54556 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_587
timestamp 1649977179
transform 1 0 55108 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_589
timestamp 1649977179
transform 1 0 55292 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_601
timestamp 1649977179
transform 1 0 56396 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_613
timestamp 1649977179
transform 1 0 57500 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_625
timestamp 1649977179
transform 1 0 58604 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_637
timestamp 1649977179
transform 1 0 59708 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_643
timestamp 1649977179
transform 1 0 60260 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_645
timestamp 1649977179
transform 1 0 60444 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_657
timestamp 1649977179
transform 1 0 61548 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_669
timestamp 1649977179
transform 1 0 62652 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_681
timestamp 1649977179
transform 1 0 63756 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_693
timestamp 1649977179
transform 1 0 64860 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_699
timestamp 1649977179
transform 1 0 65412 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_701
timestamp 1649977179
transform 1 0 65596 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_713
timestamp 1649977179
transform 1 0 66700 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_725
timestamp 1649977179
transform 1 0 67804 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_729
timestamp 1649977179
transform 1 0 68172 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_3
timestamp 1649977179
transform 1 0 1380 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_11
timestamp 1649977179
transform 1 0 2116 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_15
timestamp 1649977179
transform 1 0 2484 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_39
timestamp 1649977179
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1649977179
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1649977179
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_57
timestamp 1649977179
transform 1 0 6348 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_66
timestamp 1649977179
transform 1 0 7176 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_88
timestamp 1649977179
transform 1 0 9200 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_92
timestamp 1649977179
transform 1 0 9568 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_101
timestamp 1649977179
transform 1 0 10396 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_107
timestamp 1649977179
transform 1 0 10948 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1649977179
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1649977179
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_125
timestamp 1649977179
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_137
timestamp 1649977179
transform 1 0 13708 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_143
timestamp 1649977179
transform 1 0 14260 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_152
timestamp 1649977179
transform 1 0 15088 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_164
timestamp 1649977179
transform 1 0 16192 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_29_169
timestamp 1649977179
transform 1 0 16652 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_29_180
timestamp 1649977179
transform 1 0 17664 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_188
timestamp 1649977179
transform 1 0 18400 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_200
timestamp 1649977179
transform 1 0 19504 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_220
timestamp 1649977179
transform 1 0 21344 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_229
timestamp 1649977179
transform 1 0 22172 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_249
timestamp 1649977179
transform 1 0 24012 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_261
timestamp 1649977179
transform 1 0 25116 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_265
timestamp 1649977179
transform 1 0 25484 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_271
timestamp 1649977179
transform 1 0 26036 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 1649977179
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_281
timestamp 1649977179
transform 1 0 26956 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_287
timestamp 1649977179
transform 1 0 27508 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_294
timestamp 1649977179
transform 1 0 28152 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_314
timestamp 1649977179
transform 1 0 29992 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_326
timestamp 1649977179
transform 1 0 31096 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_334
timestamp 1649977179
transform 1 0 31832 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_339
timestamp 1649977179
transform 1 0 32292 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_347
timestamp 1649977179
transform 1 0 33028 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_353
timestamp 1649977179
transform 1 0 33580 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_359
timestamp 1649977179
transform 1 0 34132 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_362
timestamp 1649977179
transform 1 0 34408 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_382
timestamp 1649977179
transform 1 0 36248 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_388
timestamp 1649977179
transform 1 0 36800 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_393
timestamp 1649977179
transform 1 0 37260 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_403
timestamp 1649977179
transform 1 0 38180 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_411
timestamp 1649977179
transform 1 0 38916 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_429
timestamp 1649977179
transform 1 0 40572 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_441
timestamp 1649977179
transform 1 0 41676 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_447
timestamp 1649977179
transform 1 0 42228 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_449
timestamp 1649977179
transform 1 0 42412 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_461
timestamp 1649977179
transform 1 0 43516 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_473
timestamp 1649977179
transform 1 0 44620 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_485
timestamp 1649977179
transform 1 0 45724 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_497
timestamp 1649977179
transform 1 0 46828 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_503
timestamp 1649977179
transform 1 0 47380 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_505
timestamp 1649977179
transform 1 0 47564 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_517
timestamp 1649977179
transform 1 0 48668 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_529
timestamp 1649977179
transform 1 0 49772 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_541
timestamp 1649977179
transform 1 0 50876 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_553
timestamp 1649977179
transform 1 0 51980 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_559
timestamp 1649977179
transform 1 0 52532 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_561
timestamp 1649977179
transform 1 0 52716 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_573
timestamp 1649977179
transform 1 0 53820 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_585
timestamp 1649977179
transform 1 0 54924 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_597
timestamp 1649977179
transform 1 0 56028 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_609
timestamp 1649977179
transform 1 0 57132 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_615
timestamp 1649977179
transform 1 0 57684 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_617
timestamp 1649977179
transform 1 0 57868 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_629
timestamp 1649977179
transform 1 0 58972 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_641
timestamp 1649977179
transform 1 0 60076 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_653
timestamp 1649977179
transform 1 0 61180 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_665
timestamp 1649977179
transform 1 0 62284 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_671
timestamp 1649977179
transform 1 0 62836 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_673
timestamp 1649977179
transform 1 0 63020 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_685
timestamp 1649977179
transform 1 0 64124 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_697
timestamp 1649977179
transform 1 0 65228 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_709
timestamp 1649977179
transform 1 0 66332 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_721
timestamp 1649977179
transform 1 0 67436 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_727
timestamp 1649977179
transform 1 0 67988 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_729
timestamp 1649977179
transform 1 0 68172 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_3
timestamp 1649977179
transform 1 0 1380 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_16
timestamp 1649977179
transform 1 0 2576 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1649977179
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_44
timestamp 1649977179
transform 1 0 5152 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_50
timestamp 1649977179
transform 1 0 5704 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_62
timestamp 1649977179
transform 1 0 6808 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_68
timestamp 1649977179
transform 1 0 7360 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_80
timestamp 1649977179
transform 1 0 8464 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1649977179
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_97
timestamp 1649977179
transform 1 0 10028 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_30_116
timestamp 1649977179
transform 1 0 11776 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_128
timestamp 1649977179
transform 1 0 12880 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_136
timestamp 1649977179
transform 1 0 13616 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_149
timestamp 1649977179
transform 1 0 14812 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_158
timestamp 1649977179
transform 1 0 15640 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_165
timestamp 1649977179
transform 1 0 16284 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_171
timestamp 1649977179
transform 1 0 16836 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_191
timestamp 1649977179
transform 1 0 18676 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1649977179
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_197
timestamp 1649977179
transform 1 0 19228 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_201
timestamp 1649977179
transform 1 0 19596 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_215
timestamp 1649977179
transform 1 0 20884 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_219
timestamp 1649977179
transform 1 0 21252 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_227
timestamp 1649977179
transform 1 0 21988 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_237
timestamp 1649977179
transform 1 0 22908 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_245
timestamp 1649977179
transform 1 0 23644 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_248
timestamp 1649977179
transform 1 0 23920 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_30_253
timestamp 1649977179
transform 1 0 24380 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_258
timestamp 1649977179
transform 1 0 24840 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_267
timestamp 1649977179
transform 1 0 25668 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_273
timestamp 1649977179
transform 1 0 26220 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_290
timestamp 1649977179
transform 1 0 27784 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_302
timestamp 1649977179
transform 1 0 28888 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_30_309
timestamp 1649977179
transform 1 0 29532 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_318
timestamp 1649977179
transform 1 0 30360 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_330
timestamp 1649977179
transform 1 0 31464 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_30_349
timestamp 1649977179
transform 1 0 33212 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_360
timestamp 1649977179
transform 1 0 34224 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_373
timestamp 1649977179
transform 1 0 35420 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_384
timestamp 1649977179
transform 1 0 36432 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_396
timestamp 1649977179
transform 1 0 37536 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_416
timestamp 1649977179
transform 1 0 39376 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_421
timestamp 1649977179
transform 1 0 39836 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_427
timestamp 1649977179
transform 1 0 40388 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_435
timestamp 1649977179
transform 1 0 41124 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_443
timestamp 1649977179
transform 1 0 41860 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_455
timestamp 1649977179
transform 1 0 42964 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_467
timestamp 1649977179
transform 1 0 44068 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_475
timestamp 1649977179
transform 1 0 44804 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_477
timestamp 1649977179
transform 1 0 44988 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_489
timestamp 1649977179
transform 1 0 46092 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_501
timestamp 1649977179
transform 1 0 47196 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_513
timestamp 1649977179
transform 1 0 48300 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_525
timestamp 1649977179
transform 1 0 49404 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_531
timestamp 1649977179
transform 1 0 49956 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_533
timestamp 1649977179
transform 1 0 50140 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_545
timestamp 1649977179
transform 1 0 51244 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_557
timestamp 1649977179
transform 1 0 52348 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_569
timestamp 1649977179
transform 1 0 53452 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_581
timestamp 1649977179
transform 1 0 54556 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_587
timestamp 1649977179
transform 1 0 55108 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_589
timestamp 1649977179
transform 1 0 55292 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_601
timestamp 1649977179
transform 1 0 56396 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_613
timestamp 1649977179
transform 1 0 57500 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_625
timestamp 1649977179
transform 1 0 58604 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_637
timestamp 1649977179
transform 1 0 59708 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_643
timestamp 1649977179
transform 1 0 60260 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_645
timestamp 1649977179
transform 1 0 60444 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_657
timestamp 1649977179
transform 1 0 61548 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_669
timestamp 1649977179
transform 1 0 62652 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_681
timestamp 1649977179
transform 1 0 63756 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_693
timestamp 1649977179
transform 1 0 64860 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_699
timestamp 1649977179
transform 1 0 65412 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_701
timestamp 1649977179
transform 1 0 65596 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_713
timestamp 1649977179
transform 1 0 66700 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_725
timestamp 1649977179
transform 1 0 67804 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_729
timestamp 1649977179
transform 1 0 68172 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_3
timestamp 1649977179
transform 1 0 1380 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_11
timestamp 1649977179
transform 1 0 2116 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_17
timestamp 1649977179
transform 1 0 2668 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_29
timestamp 1649977179
transform 1 0 3772 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_41
timestamp 1649977179
transform 1 0 4876 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_53
timestamp 1649977179
transform 1 0 5980 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_62
timestamp 1649977179
transform 1 0 6808 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_68
timestamp 1649977179
transform 1 0 7360 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_74
timestamp 1649977179
transform 1 0 7912 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_78
timestamp 1649977179
transform 1 0 8280 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_84
timestamp 1649977179
transform 1 0 8832 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_92
timestamp 1649977179
transform 1 0 9568 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_95
timestamp 1649977179
transform 1 0 9844 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_107
timestamp 1649977179
transform 1 0 10948 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1649977179
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_113
timestamp 1649977179
transform 1 0 11500 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_119
timestamp 1649977179
transform 1 0 12052 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_136
timestamp 1649977179
transform 1 0 13616 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_152
timestamp 1649977179
transform 1 0 15088 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_159
timestamp 1649977179
transform 1 0 15732 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1649977179
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_174
timestamp 1649977179
transform 1 0 17112 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_181
timestamp 1649977179
transform 1 0 17756 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_187
timestamp 1649977179
transform 1 0 18308 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_203
timestamp 1649977179
transform 1 0 19780 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_217
timestamp 1649977179
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1649977179
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_235
timestamp 1649977179
transform 1 0 22724 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_239
timestamp 1649977179
transform 1 0 23092 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_250
timestamp 1649977179
transform 1 0 24104 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_254
timestamp 1649977179
transform 1 0 24472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_258
timestamp 1649977179
transform 1 0 24840 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_264
timestamp 1649977179
transform 1 0 25392 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_273
timestamp 1649977179
transform 1 0 26220 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 1649977179
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_283
timestamp 1649977179
transform 1 0 27140 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_289
timestamp 1649977179
transform 1 0 27692 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_295
timestamp 1649977179
transform 1 0 28244 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_312
timestamp 1649977179
transform 1 0 29808 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_324
timestamp 1649977179
transform 1 0 30912 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_328
timestamp 1649977179
transform 1 0 31280 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_337
timestamp 1649977179
transform 1 0 32108 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_345
timestamp 1649977179
transform 1 0 32844 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_361
timestamp 1649977179
transform 1 0 34316 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_375
timestamp 1649977179
transform 1 0 35604 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_379
timestamp 1649977179
transform 1 0 35972 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_383
timestamp 1649977179
transform 1 0 36340 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1649977179
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_398
timestamp 1649977179
transform 1 0 37720 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_407
timestamp 1649977179
transform 1 0 38548 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_413
timestamp 1649977179
transform 1 0 39100 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_419
timestamp 1649977179
transform 1 0 39652 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_425
timestamp 1649977179
transform 1 0 40204 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_436
timestamp 1649977179
transform 1 0 41216 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_442
timestamp 1649977179
transform 1 0 41768 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_31_449
timestamp 1649977179
transform 1 0 42412 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_461
timestamp 1649977179
transform 1 0 43516 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_473
timestamp 1649977179
transform 1 0 44620 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_485
timestamp 1649977179
transform 1 0 45724 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_497
timestamp 1649977179
transform 1 0 46828 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_503
timestamp 1649977179
transform 1 0 47380 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_505
timestamp 1649977179
transform 1 0 47564 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_517
timestamp 1649977179
transform 1 0 48668 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_529
timestamp 1649977179
transform 1 0 49772 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_541
timestamp 1649977179
transform 1 0 50876 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_553
timestamp 1649977179
transform 1 0 51980 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_559
timestamp 1649977179
transform 1 0 52532 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_561
timestamp 1649977179
transform 1 0 52716 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_573
timestamp 1649977179
transform 1 0 53820 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_585
timestamp 1649977179
transform 1 0 54924 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_597
timestamp 1649977179
transform 1 0 56028 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_609
timestamp 1649977179
transform 1 0 57132 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_615
timestamp 1649977179
transform 1 0 57684 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_617
timestamp 1649977179
transform 1 0 57868 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_629
timestamp 1649977179
transform 1 0 58972 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_641
timestamp 1649977179
transform 1 0 60076 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_653
timestamp 1649977179
transform 1 0 61180 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_665
timestamp 1649977179
transform 1 0 62284 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_671
timestamp 1649977179
transform 1 0 62836 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_673
timestamp 1649977179
transform 1 0 63020 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_685
timestamp 1649977179
transform 1 0 64124 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_697
timestamp 1649977179
transform 1 0 65228 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_709
timestamp 1649977179
transform 1 0 66332 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_721
timestamp 1649977179
transform 1 0 67436 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_727
timestamp 1649977179
transform 1 0 67988 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_729
timestamp 1649977179
transform 1 0 68172 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_3
timestamp 1649977179
transform 1 0 1380 0 1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_32_14
timestamp 1649977179
transform 1 0 2392 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_26
timestamp 1649977179
transform 1 0 3496 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1649977179
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_41
timestamp 1649977179
transform 1 0 4876 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_58
timestamp 1649977179
transform 1 0 6440 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_70
timestamp 1649977179
transform 1 0 7544 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_80
timestamp 1649977179
transform 1 0 8464 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_93
timestamp 1649977179
transform 1 0 9660 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_113
timestamp 1649977179
transform 1 0 11500 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_125
timestamp 1649977179
transform 1 0 12604 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_133
timestamp 1649977179
transform 1 0 13340 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_136
timestamp 1649977179
transform 1 0 13616 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_141
timestamp 1649977179
transform 1 0 14076 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_156
timestamp 1649977179
transform 1 0 15456 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_167
timestamp 1649977179
transform 1 0 16468 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_173
timestamp 1649977179
transform 1 0 17020 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_181
timestamp 1649977179
transform 1 0 17756 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_192
timestamp 1649977179
transform 1 0 18768 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_207
timestamp 1649977179
transform 1 0 20148 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_221
timestamp 1649977179
transform 1 0 21436 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_234
timestamp 1649977179
transform 1 0 22632 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_248
timestamp 1649977179
transform 1 0 23920 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_253
timestamp 1649977179
transform 1 0 24380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_261
timestamp 1649977179
transform 1 0 25116 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_273
timestamp 1649977179
transform 1 0 26220 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_280
timestamp 1649977179
transform 1 0 26864 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_288
timestamp 1649977179
transform 1 0 27600 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_297
timestamp 1649977179
transform 1 0 28428 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_303
timestamp 1649977179
transform 1 0 28980 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 1649977179
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_309
timestamp 1649977179
transform 1 0 29532 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_315
timestamp 1649977179
transform 1 0 30084 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_325
timestamp 1649977179
transform 1 0 31004 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_338
timestamp 1649977179
transform 1 0 32200 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_345
timestamp 1649977179
transform 1 0 32844 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_351
timestamp 1649977179
transform 1 0 33396 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_360
timestamp 1649977179
transform 1 0 34224 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_365
timestamp 1649977179
transform 1 0 34684 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_369
timestamp 1649977179
transform 1 0 35052 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_384
timestamp 1649977179
transform 1 0 36432 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_392
timestamp 1649977179
transform 1 0 37168 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_401
timestamp 1649977179
transform 1 0 37996 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_407
timestamp 1649977179
transform 1 0 38548 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_413
timestamp 1649977179
transform 1 0 39100 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_419
timestamp 1649977179
transform 1 0 39652 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_421
timestamp 1649977179
transform 1 0 39836 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_430
timestamp 1649977179
transform 1 0 40664 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_436
timestamp 1649977179
transform 1 0 41216 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_442
timestamp 1649977179
transform 1 0 41768 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_448
timestamp 1649977179
transform 1 0 42320 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_460
timestamp 1649977179
transform 1 0 43424 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_472
timestamp 1649977179
transform 1 0 44528 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_477
timestamp 1649977179
transform 1 0 44988 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_489
timestamp 1649977179
transform 1 0 46092 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_501
timestamp 1649977179
transform 1 0 47196 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_513
timestamp 1649977179
transform 1 0 48300 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_525
timestamp 1649977179
transform 1 0 49404 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_531
timestamp 1649977179
transform 1 0 49956 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_533
timestamp 1649977179
transform 1 0 50140 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_545
timestamp 1649977179
transform 1 0 51244 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_557
timestamp 1649977179
transform 1 0 52348 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_569
timestamp 1649977179
transform 1 0 53452 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_581
timestamp 1649977179
transform 1 0 54556 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_587
timestamp 1649977179
transform 1 0 55108 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_589
timestamp 1649977179
transform 1 0 55292 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_601
timestamp 1649977179
transform 1 0 56396 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_613
timestamp 1649977179
transform 1 0 57500 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_625
timestamp 1649977179
transform 1 0 58604 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_637
timestamp 1649977179
transform 1 0 59708 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_643
timestamp 1649977179
transform 1 0 60260 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_645
timestamp 1649977179
transform 1 0 60444 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_657
timestamp 1649977179
transform 1 0 61548 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_669
timestamp 1649977179
transform 1 0 62652 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_681
timestamp 1649977179
transform 1 0 63756 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_693
timestamp 1649977179
transform 1 0 64860 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_699
timestamp 1649977179
transform 1 0 65412 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_701
timestamp 1649977179
transform 1 0 65596 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_713
timestamp 1649977179
transform 1 0 66700 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_725
timestamp 1649977179
transform 1 0 67804 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_3
timestamp 1649977179
transform 1 0 1380 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_18
timestamp 1649977179
transform 1 0 2760 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_42
timestamp 1649977179
transform 1 0 4968 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_49
timestamp 1649977179
transform 1 0 5612 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1649977179
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_60
timestamp 1649977179
transform 1 0 6624 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_70
timestamp 1649977179
transform 1 0 7544 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_85
timestamp 1649977179
transform 1 0 8924 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_99
timestamp 1649977179
transform 1 0 10212 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1649977179
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_113
timestamp 1649977179
transform 1 0 11500 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_119
timestamp 1649977179
transform 1 0 12052 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_125
timestamp 1649977179
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_137
timestamp 1649977179
transform 1 0 13708 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_146
timestamp 1649977179
transform 1 0 14536 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_33_160
timestamp 1649977179
transform 1 0 15824 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_33_173
timestamp 1649977179
transform 1 0 17020 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_179
timestamp 1649977179
transform 1 0 17572 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_183
timestamp 1649977179
transform 1 0 17940 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_189
timestamp 1649977179
transform 1 0 18492 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_201
timestamp 1649977179
transform 1 0 19596 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_212
timestamp 1649977179
transform 1 0 20608 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_220
timestamp 1649977179
transform 1 0 21344 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_232
timestamp 1649977179
transform 1 0 22448 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_33_246
timestamp 1649977179
transform 1 0 23736 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_252
timestamp 1649977179
transform 1 0 24288 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_256
timestamp 1649977179
transform 1 0 24656 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_262
timestamp 1649977179
transform 1 0 25208 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_273
timestamp 1649977179
transform 1 0 26220 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1649977179
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_281
timestamp 1649977179
transform 1 0 26956 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_33_289
timestamp 1649977179
transform 1 0 27692 0 -1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_33_306
timestamp 1649977179
transform 1 0 29256 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_318
timestamp 1649977179
transform 1 0 30360 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_326
timestamp 1649977179
transform 1 0 31096 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_332
timestamp 1649977179
transform 1 0 31648 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_337
timestamp 1649977179
transform 1 0 32108 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_347
timestamp 1649977179
transform 1 0 33028 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_351
timestamp 1649977179
transform 1 0 33396 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_355
timestamp 1649977179
transform 1 0 33764 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_364
timestamp 1649977179
transform 1 0 34592 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_368
timestamp 1649977179
transform 1 0 34960 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_385
timestamp 1649977179
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 1649977179
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_393
timestamp 1649977179
transform 1 0 37260 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_33_402
timestamp 1649977179
transform 1 0 38088 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_426
timestamp 1649977179
transform 1 0 40296 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_432
timestamp 1649977179
transform 1 0 40848 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_444
timestamp 1649977179
transform 1 0 41952 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_455
timestamp 1649977179
transform 1 0 42964 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_467
timestamp 1649977179
transform 1 0 44068 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_479
timestamp 1649977179
transform 1 0 45172 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_491
timestamp 1649977179
transform 1 0 46276 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_503
timestamp 1649977179
transform 1 0 47380 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_505
timestamp 1649977179
transform 1 0 47564 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_517
timestamp 1649977179
transform 1 0 48668 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_529
timestamp 1649977179
transform 1 0 49772 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_541
timestamp 1649977179
transform 1 0 50876 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_553
timestamp 1649977179
transform 1 0 51980 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_559
timestamp 1649977179
transform 1 0 52532 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_561
timestamp 1649977179
transform 1 0 52716 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_573
timestamp 1649977179
transform 1 0 53820 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_585
timestamp 1649977179
transform 1 0 54924 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_597
timestamp 1649977179
transform 1 0 56028 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_609
timestamp 1649977179
transform 1 0 57132 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_615
timestamp 1649977179
transform 1 0 57684 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_617
timestamp 1649977179
transform 1 0 57868 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_629
timestamp 1649977179
transform 1 0 58972 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_641
timestamp 1649977179
transform 1 0 60076 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_653
timestamp 1649977179
transform 1 0 61180 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_665
timestamp 1649977179
transform 1 0 62284 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_671
timestamp 1649977179
transform 1 0 62836 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_673
timestamp 1649977179
transform 1 0 63020 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_685
timestamp 1649977179
transform 1 0 64124 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_697
timestamp 1649977179
transform 1 0 65228 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_709
timestamp 1649977179
transform 1 0 66332 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_724
timestamp 1649977179
transform 1 0 67712 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_729
timestamp 1649977179
transform 1 0 68172 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_3
timestamp 1649977179
transform 1 0 1380 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_18
timestamp 1649977179
transform 1 0 2760 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_24
timestamp 1649977179
transform 1 0 3312 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1649977179
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_41
timestamp 1649977179
transform 1 0 4876 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_51
timestamp 1649977179
transform 1 0 5796 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_55
timestamp 1649977179
transform 1 0 6164 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_58
timestamp 1649977179
transform 1 0 6440 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_70
timestamp 1649977179
transform 1 0 7544 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_80
timestamp 1649977179
transform 1 0 8464 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_87
timestamp 1649977179
transform 1 0 9108 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_91
timestamp 1649977179
transform 1 0 9476 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_108
timestamp 1649977179
transform 1 0 11040 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_130
timestamp 1649977179
transform 1 0 13064 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_136
timestamp 1649977179
transform 1 0 13616 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_148
timestamp 1649977179
transform 1 0 14720 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_170
timestamp 1649977179
transform 1 0 16744 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_176
timestamp 1649977179
transform 1 0 17296 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_187
timestamp 1649977179
transform 1 0 18308 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1649977179
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_205
timestamp 1649977179
transform 1 0 19964 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_34_215
timestamp 1649977179
transform 1 0 20884 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_34_228
timestamp 1649977179
transform 1 0 22080 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_34_244
timestamp 1649977179
transform 1 0 23552 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_260
timestamp 1649977179
transform 1 0 25024 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_269
timestamp 1649977179
transform 1 0 25852 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_273
timestamp 1649977179
transform 1 0 26220 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_290
timestamp 1649977179
transform 1 0 27784 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_297
timestamp 1649977179
transform 1 0 28428 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_304
timestamp 1649977179
transform 1 0 29072 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_316
timestamp 1649977179
transform 1 0 30176 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_326
timestamp 1649977179
transform 1 0 31096 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_330
timestamp 1649977179
transform 1 0 31464 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_333
timestamp 1649977179
transform 1 0 31740 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_337
timestamp 1649977179
transform 1 0 32108 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_343
timestamp 1649977179
transform 1 0 32660 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_349
timestamp 1649977179
transform 1 0 33212 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_360
timestamp 1649977179
transform 1 0 34224 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_368
timestamp 1649977179
transform 1 0 34960 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_382
timestamp 1649977179
transform 1 0 36248 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_388
timestamp 1649977179
transform 1 0 36800 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_397
timestamp 1649977179
transform 1 0 37628 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_403
timestamp 1649977179
transform 1 0 38180 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_409
timestamp 1649977179
transform 1 0 38732 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_415
timestamp 1649977179
transform 1 0 39284 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_419
timestamp 1649977179
transform 1 0 39652 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_421
timestamp 1649977179
transform 1 0 39836 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_429
timestamp 1649977179
transform 1 0 40572 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_433
timestamp 1649977179
transform 1 0 40940 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_444
timestamp 1649977179
transform 1 0 41952 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_456
timestamp 1649977179
transform 1 0 43056 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_468
timestamp 1649977179
transform 1 0 44160 0 1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_34_477
timestamp 1649977179
transform 1 0 44988 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_489
timestamp 1649977179
transform 1 0 46092 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_501
timestamp 1649977179
transform 1 0 47196 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_513
timestamp 1649977179
transform 1 0 48300 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_525
timestamp 1649977179
transform 1 0 49404 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_531
timestamp 1649977179
transform 1 0 49956 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_533
timestamp 1649977179
transform 1 0 50140 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_545
timestamp 1649977179
transform 1 0 51244 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_557
timestamp 1649977179
transform 1 0 52348 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_569
timestamp 1649977179
transform 1 0 53452 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_581
timestamp 1649977179
transform 1 0 54556 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_587
timestamp 1649977179
transform 1 0 55108 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_589
timestamp 1649977179
transform 1 0 55292 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_601
timestamp 1649977179
transform 1 0 56396 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_613
timestamp 1649977179
transform 1 0 57500 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_625
timestamp 1649977179
transform 1 0 58604 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_637
timestamp 1649977179
transform 1 0 59708 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_643
timestamp 1649977179
transform 1 0 60260 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_645
timestamp 1649977179
transform 1 0 60444 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_657
timestamp 1649977179
transform 1 0 61548 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_669
timestamp 1649977179
transform 1 0 62652 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_681
timestamp 1649977179
transform 1 0 63756 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_693
timestamp 1649977179
transform 1 0 64860 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_699
timestamp 1649977179
transform 1 0 65412 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_701
timestamp 1649977179
transform 1 0 65596 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_713
timestamp 1649977179
transform 1 0 66700 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_725
timestamp 1649977179
transform 1 0 67804 0 1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 1649977179
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_15
timestamp 1649977179
transform 1 0 2484 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_35
timestamp 1649977179
transform 1 0 4324 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_47
timestamp 1649977179
transform 1 0 5428 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1649977179
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_73
timestamp 1649977179
transform 1 0 7820 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_82
timestamp 1649977179
transform 1 0 8648 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_94
timestamp 1649977179
transform 1 0 9752 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_100
timestamp 1649977179
transform 1 0 10304 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_121
timestamp 1649977179
transform 1 0 12236 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_127
timestamp 1649977179
transform 1 0 12788 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_139
timestamp 1649977179
transform 1 0 13892 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_151
timestamp 1649977179
transform 1 0 14996 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_35_160
timestamp 1649977179
transform 1 0 15824 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_35_174
timestamp 1649977179
transform 1 0 17112 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_185
timestamp 1649977179
transform 1 0 18124 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_191
timestamp 1649977179
transform 1 0 18676 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_211
timestamp 1649977179
transform 1 0 20516 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_218
timestamp 1649977179
transform 1 0 21160 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_35_225
timestamp 1649977179
transform 1 0 21804 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_229
timestamp 1649977179
transform 1 0 22172 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_243
timestamp 1649977179
transform 1 0 23460 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_257
timestamp 1649977179
transform 1 0 24748 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_263
timestamp 1649977179
transform 1 0 25300 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_275
timestamp 1649977179
transform 1 0 26404 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1649977179
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_281
timestamp 1649977179
transform 1 0 26956 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_285
timestamp 1649977179
transform 1 0 27324 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_295
timestamp 1649977179
transform 1 0 28244 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_307
timestamp 1649977179
transform 1 0 29348 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_315
timestamp 1649977179
transform 1 0 30084 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_332
timestamp 1649977179
transform 1 0 31648 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_35_337
timestamp 1649977179
transform 1 0 32108 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_35_342
timestamp 1649977179
transform 1 0 32568 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_366
timestamp 1649977179
transform 1 0 34776 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_380
timestamp 1649977179
transform 1 0 36064 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_388
timestamp 1649977179
transform 1 0 36800 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_35_393
timestamp 1649977179
transform 1 0 37260 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_404
timestamp 1649977179
transform 1 0 38272 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_410
timestamp 1649977179
transform 1 0 38824 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_422
timestamp 1649977179
transform 1 0 39928 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_434
timestamp 1649977179
transform 1 0 41032 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_442
timestamp 1649977179
transform 1 0 41768 0 -1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_35_457
timestamp 1649977179
transform 1 0 43148 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_469
timestamp 1649977179
transform 1 0 44252 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_481
timestamp 1649977179
transform 1 0 45356 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_493
timestamp 1649977179
transform 1 0 46460 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_501
timestamp 1649977179
transform 1 0 47196 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_505
timestamp 1649977179
transform 1 0 47564 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_517
timestamp 1649977179
transform 1 0 48668 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_529
timestamp 1649977179
transform 1 0 49772 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_541
timestamp 1649977179
transform 1 0 50876 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_553
timestamp 1649977179
transform 1 0 51980 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_559
timestamp 1649977179
transform 1 0 52532 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_561
timestamp 1649977179
transform 1 0 52716 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_573
timestamp 1649977179
transform 1 0 53820 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_585
timestamp 1649977179
transform 1 0 54924 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_597
timestamp 1649977179
transform 1 0 56028 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_609
timestamp 1649977179
transform 1 0 57132 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_615
timestamp 1649977179
transform 1 0 57684 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_617
timestamp 1649977179
transform 1 0 57868 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_629
timestamp 1649977179
transform 1 0 58972 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_641
timestamp 1649977179
transform 1 0 60076 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_653
timestamp 1649977179
transform 1 0 61180 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_665
timestamp 1649977179
transform 1 0 62284 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_671
timestamp 1649977179
transform 1 0 62836 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_673
timestamp 1649977179
transform 1 0 63020 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_685
timestamp 1649977179
transform 1 0 64124 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_697
timestamp 1649977179
transform 1 0 65228 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_709
timestamp 1649977179
transform 1 0 66332 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_721
timestamp 1649977179
transform 1 0 67436 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_727
timestamp 1649977179
transform 1 0 67988 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_729
timestamp 1649977179
transform 1 0 68172 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_3
timestamp 1649977179
transform 1 0 1380 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_11
timestamp 1649977179
transform 1 0 2116 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_36_22
timestamp 1649977179
transform 1 0 3128 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_29
timestamp 1649977179
transform 1 0 3772 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_49
timestamp 1649977179
transform 1 0 5612 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_58
timestamp 1649977179
transform 1 0 6440 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_71
timestamp 1649977179
transform 1 0 7636 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_80
timestamp 1649977179
transform 1 0 8464 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_95
timestamp 1649977179
transform 1 0 9844 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_107
timestamp 1649977179
transform 1 0 10948 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_115
timestamp 1649977179
transform 1 0 11684 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_120
timestamp 1649977179
transform 1 0 12144 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_132
timestamp 1649977179
transform 1 0 13248 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_157
timestamp 1649977179
transform 1 0 15548 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_169
timestamp 1649977179
transform 1 0 16652 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_177
timestamp 1649977179
transform 1 0 17388 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_185
timestamp 1649977179
transform 1 0 18124 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_193
timestamp 1649977179
transform 1 0 18860 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_36_205
timestamp 1649977179
transform 1 0 19964 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_217
timestamp 1649977179
transform 1 0 21068 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_36_230
timestamp 1649977179
transform 1 0 22264 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_36_243
timestamp 1649977179
transform 1 0 23460 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1649977179
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_255
timestamp 1649977179
transform 1 0 24564 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_274
timestamp 1649977179
transform 1 0 26312 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_36_286
timestamp 1649977179
transform 1 0 27416 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_36_299
timestamp 1649977179
transform 1 0 28612 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1649977179
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_314
timestamp 1649977179
transform 1 0 29992 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_320
timestamp 1649977179
transform 1 0 30544 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_324
timestamp 1649977179
transform 1 0 30912 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_341
timestamp 1649977179
transform 1 0 32476 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_353
timestamp 1649977179
transform 1 0 33580 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_359
timestamp 1649977179
transform 1 0 34132 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1649977179
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_365
timestamp 1649977179
transform 1 0 34684 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_369
timestamp 1649977179
transform 1 0 35052 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_372
timestamp 1649977179
transform 1 0 35328 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_382
timestamp 1649977179
transform 1 0 36248 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_388
timestamp 1649977179
transform 1 0 36800 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_400
timestamp 1649977179
transform 1 0 37904 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_406
timestamp 1649977179
transform 1 0 38456 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_418
timestamp 1649977179
transform 1 0 39560 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_437
timestamp 1649977179
transform 1 0 41308 0 1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_36_448
timestamp 1649977179
transform 1 0 42320 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_460
timestamp 1649977179
transform 1 0 43424 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_472
timestamp 1649977179
transform 1 0 44528 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_477
timestamp 1649977179
transform 1 0 44988 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_489
timestamp 1649977179
transform 1 0 46092 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_501
timestamp 1649977179
transform 1 0 47196 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_513
timestamp 1649977179
transform 1 0 48300 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_525
timestamp 1649977179
transform 1 0 49404 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_531
timestamp 1649977179
transform 1 0 49956 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_533
timestamp 1649977179
transform 1 0 50140 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_545
timestamp 1649977179
transform 1 0 51244 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_557
timestamp 1649977179
transform 1 0 52348 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_569
timestamp 1649977179
transform 1 0 53452 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_581
timestamp 1649977179
transform 1 0 54556 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_587
timestamp 1649977179
transform 1 0 55108 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_589
timestamp 1649977179
transform 1 0 55292 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_601
timestamp 1649977179
transform 1 0 56396 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_613
timestamp 1649977179
transform 1 0 57500 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_625
timestamp 1649977179
transform 1 0 58604 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_637
timestamp 1649977179
transform 1 0 59708 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_643
timestamp 1649977179
transform 1 0 60260 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_645
timestamp 1649977179
transform 1 0 60444 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_657
timestamp 1649977179
transform 1 0 61548 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_669
timestamp 1649977179
transform 1 0 62652 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_681
timestamp 1649977179
transform 1 0 63756 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_693
timestamp 1649977179
transform 1 0 64860 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_699
timestamp 1649977179
transform 1 0 65412 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_701
timestamp 1649977179
transform 1 0 65596 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_713
timestamp 1649977179
transform 1 0 66700 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_725
timestamp 1649977179
transform 1 0 67804 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_729
timestamp 1649977179
transform 1 0 68172 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_3
timestamp 1649977179
transform 1 0 1380 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_11
timestamp 1649977179
transform 1 0 2116 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_17
timestamp 1649977179
transform 1 0 2668 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_23
timestamp 1649977179
transform 1 0 3220 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_29
timestamp 1649977179
transform 1 0 3772 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_41
timestamp 1649977179
transform 1 0 4876 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_52
timestamp 1649977179
transform 1 0 5888 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_59
timestamp 1649977179
transform 1 0 6532 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_67
timestamp 1649977179
transform 1 0 7268 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_72
timestamp 1649977179
transform 1 0 7728 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_87
timestamp 1649977179
transform 1 0 9108 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_91
timestamp 1649977179
transform 1 0 9476 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_108
timestamp 1649977179
transform 1 0 11040 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_113
timestamp 1649977179
transform 1 0 11500 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_119
timestamp 1649977179
transform 1 0 12052 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_125
timestamp 1649977179
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_137
timestamp 1649977179
transform 1 0 13708 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_146
timestamp 1649977179
transform 1 0 14536 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_155
timestamp 1649977179
transform 1 0 15364 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_164
timestamp 1649977179
transform 1 0 16192 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_169
timestamp 1649977179
transform 1 0 16652 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_173
timestamp 1649977179
transform 1 0 17020 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_182
timestamp 1649977179
transform 1 0 17848 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_194
timestamp 1649977179
transform 1 0 18952 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_206
timestamp 1649977179
transform 1 0 20056 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_218
timestamp 1649977179
transform 1 0 21160 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_37_225
timestamp 1649977179
transform 1 0 21804 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_231
timestamp 1649977179
transform 1 0 22356 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_240
timestamp 1649977179
transform 1 0 23184 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_252
timestamp 1649977179
transform 1 0 24288 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_256
timestamp 1649977179
transform 1 0 24656 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_264
timestamp 1649977179
transform 1 0 25392 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_275
timestamp 1649977179
transform 1 0 26404 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1649977179
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_286
timestamp 1649977179
transform 1 0 27416 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_292
timestamp 1649977179
transform 1 0 27968 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_304
timestamp 1649977179
transform 1 0 29072 0 -1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_37_320
timestamp 1649977179
transform 1 0 30544 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_332
timestamp 1649977179
transform 1 0 31648 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_337
timestamp 1649977179
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_349
timestamp 1649977179
transform 1 0 33212 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_355
timestamp 1649977179
transform 1 0 33764 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_367
timestamp 1649977179
transform 1 0 34868 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_37_384
timestamp 1649977179
transform 1 0 36432 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_393
timestamp 1649977179
transform 1 0 37260 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_413
timestamp 1649977179
transform 1 0 39100 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_421
timestamp 1649977179
transform 1 0 39836 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_426
timestamp 1649977179
transform 1 0 40296 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_438
timestamp 1649977179
transform 1 0 41400 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_444
timestamp 1649977179
transform 1 0 41952 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_454
timestamp 1649977179
transform 1 0 42872 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_466
timestamp 1649977179
transform 1 0 43976 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_478
timestamp 1649977179
transform 1 0 45080 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_490
timestamp 1649977179
transform 1 0 46184 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_502
timestamp 1649977179
transform 1 0 47288 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_505
timestamp 1649977179
transform 1 0 47564 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_517
timestamp 1649977179
transform 1 0 48668 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_529
timestamp 1649977179
transform 1 0 49772 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_541
timestamp 1649977179
transform 1 0 50876 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_553
timestamp 1649977179
transform 1 0 51980 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_559
timestamp 1649977179
transform 1 0 52532 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_561
timestamp 1649977179
transform 1 0 52716 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_573
timestamp 1649977179
transform 1 0 53820 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_585
timestamp 1649977179
transform 1 0 54924 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_597
timestamp 1649977179
transform 1 0 56028 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_609
timestamp 1649977179
transform 1 0 57132 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_615
timestamp 1649977179
transform 1 0 57684 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_617
timestamp 1649977179
transform 1 0 57868 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_629
timestamp 1649977179
transform 1 0 58972 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_641
timestamp 1649977179
transform 1 0 60076 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_653
timestamp 1649977179
transform 1 0 61180 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_665
timestamp 1649977179
transform 1 0 62284 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_671
timestamp 1649977179
transform 1 0 62836 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_673
timestamp 1649977179
transform 1 0 63020 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_685
timestamp 1649977179
transform 1 0 64124 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_697
timestamp 1649977179
transform 1 0 65228 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_709
timestamp 1649977179
transform 1 0 66332 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_721
timestamp 1649977179
transform 1 0 67436 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_727
timestamp 1649977179
transform 1 0 67988 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_729
timestamp 1649977179
transform 1 0 68172 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_3
timestamp 1649977179
transform 1 0 1380 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_38_16
timestamp 1649977179
transform 1 0 2576 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_22
timestamp 1649977179
transform 1 0 3128 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_38_29
timestamp 1649977179
transform 1 0 3772 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_37
timestamp 1649977179
transform 1 0 4508 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_45
timestamp 1649977179
transform 1 0 5244 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_51
timestamp 1649977179
transform 1 0 5796 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_55
timestamp 1649977179
transform 1 0 6164 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_72
timestamp 1649977179
transform 1 0 7728 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_80
timestamp 1649977179
transform 1 0 8464 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_95
timestamp 1649977179
transform 1 0 9844 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_38_107
timestamp 1649977179
transform 1 0 10948 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_112
timestamp 1649977179
transform 1 0 11408 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_124
timestamp 1649977179
transform 1 0 12512 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_136
timestamp 1649977179
transform 1 0 13616 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_141
timestamp 1649977179
transform 1 0 14076 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_156
timestamp 1649977179
transform 1 0 15456 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_38_169
timestamp 1649977179
transform 1 0 16652 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_175
timestamp 1649977179
transform 1 0 17204 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_192
timestamp 1649977179
transform 1 0 18768 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_197
timestamp 1649977179
transform 1 0 19228 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_38_221
timestamp 1649977179
transform 1 0 21436 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_235
timestamp 1649977179
transform 1 0 22724 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_244
timestamp 1649977179
transform 1 0 23552 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_38_253
timestamp 1649977179
transform 1 0 24380 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_261
timestamp 1649977179
transform 1 0 25116 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_273
timestamp 1649977179
transform 1 0 26220 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_277
timestamp 1649977179
transform 1 0 26588 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_289
timestamp 1649977179
transform 1 0 27692 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_304
timestamp 1649977179
transform 1 0 29072 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_314
timestamp 1649977179
transform 1 0 29992 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_323
timestamp 1649977179
transform 1 0 30820 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_329
timestamp 1649977179
transform 1 0 31372 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_346
timestamp 1649977179
transform 1 0 32936 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_360
timestamp 1649977179
transform 1 0 34224 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_365
timestamp 1649977179
transform 1 0 34684 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_383
timestamp 1649977179
transform 1 0 36340 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_392
timestamp 1649977179
transform 1 0 37168 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_398
timestamp 1649977179
transform 1 0 37720 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_410
timestamp 1649977179
transform 1 0 38824 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_418
timestamp 1649977179
transform 1 0 39560 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_441
timestamp 1649977179
transform 1 0 41676 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_449
timestamp 1649977179
transform 1 0 42412 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_463
timestamp 1649977179
transform 1 0 43700 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_475
timestamp 1649977179
transform 1 0 44804 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_477
timestamp 1649977179
transform 1 0 44988 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_489
timestamp 1649977179
transform 1 0 46092 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_501
timestamp 1649977179
transform 1 0 47196 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_513
timestamp 1649977179
transform 1 0 48300 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_525
timestamp 1649977179
transform 1 0 49404 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_531
timestamp 1649977179
transform 1 0 49956 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_533
timestamp 1649977179
transform 1 0 50140 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_545
timestamp 1649977179
transform 1 0 51244 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_557
timestamp 1649977179
transform 1 0 52348 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_569
timestamp 1649977179
transform 1 0 53452 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_581
timestamp 1649977179
transform 1 0 54556 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_587
timestamp 1649977179
transform 1 0 55108 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_589
timestamp 1649977179
transform 1 0 55292 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_601
timestamp 1649977179
transform 1 0 56396 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_613
timestamp 1649977179
transform 1 0 57500 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_625
timestamp 1649977179
transform 1 0 58604 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_637
timestamp 1649977179
transform 1 0 59708 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_643
timestamp 1649977179
transform 1 0 60260 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_645
timestamp 1649977179
transform 1 0 60444 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_657
timestamp 1649977179
transform 1 0 61548 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_669
timestamp 1649977179
transform 1 0 62652 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_681
timestamp 1649977179
transform 1 0 63756 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_693
timestamp 1649977179
transform 1 0 64860 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_699
timestamp 1649977179
transform 1 0 65412 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_701
timestamp 1649977179
transform 1 0 65596 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_713
timestamp 1649977179
transform 1 0 66700 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_725
timestamp 1649977179
transform 1 0 67804 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_3
timestamp 1649977179
transform 1 0 1380 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_7
timestamp 1649977179
transform 1 0 1748 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_16
timestamp 1649977179
transform 1 0 2576 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_36
timestamp 1649977179
transform 1 0 4416 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_40
timestamp 1649977179
transform 1 0 4784 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_49
timestamp 1649977179
transform 1 0 5612 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1649977179
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1649977179
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_69
timestamp 1649977179
transform 1 0 7452 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_79
timestamp 1649977179
transform 1 0 8372 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_91
timestamp 1649977179
transform 1 0 9476 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_97
timestamp 1649977179
transform 1 0 10028 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_39_106
timestamp 1649977179
transform 1 0 10856 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_39_113
timestamp 1649977179
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_125
timestamp 1649977179
transform 1 0 12604 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_128
timestamp 1649977179
transform 1 0 12880 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_139
timestamp 1649977179
transform 1 0 13892 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_145
timestamp 1649977179
transform 1 0 14444 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_159
timestamp 1649977179
transform 1 0 15732 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1649977179
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_177
timestamp 1649977179
transform 1 0 17388 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_183
timestamp 1649977179
transform 1 0 17940 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_191
timestamp 1649977179
transform 1 0 18676 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_195
timestamp 1649977179
transform 1 0 19044 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_207
timestamp 1649977179
transform 1 0 20148 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_219
timestamp 1649977179
transform 1 0 21252 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1649977179
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_39_225
timestamp 1649977179
transform 1 0 21804 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_232
timestamp 1649977179
transform 1 0 22448 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_240
timestamp 1649977179
transform 1 0 23184 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_247
timestamp 1649977179
transform 1 0 23828 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_259
timestamp 1649977179
transform 1 0 24932 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_265
timestamp 1649977179
transform 1 0 25484 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_39_277
timestamp 1649977179
transform 1 0 26588 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_39_281
timestamp 1649977179
transform 1 0 26956 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_289
timestamp 1649977179
transform 1 0 27692 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_293
timestamp 1649977179
transform 1 0 28060 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_301
timestamp 1649977179
transform 1 0 28796 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_306
timestamp 1649977179
transform 1 0 29256 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_318
timestamp 1649977179
transform 1 0 30360 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_330
timestamp 1649977179
transform 1 0 31464 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_39_337
timestamp 1649977179
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_349
timestamp 1649977179
transform 1 0 33212 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_352
timestamp 1649977179
transform 1 0 33488 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_361
timestamp 1649977179
transform 1 0 34316 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_373
timestamp 1649977179
transform 1 0 35420 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_381
timestamp 1649977179
transform 1 0 36156 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_387
timestamp 1649977179
transform 1 0 36708 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1649977179
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_401
timestamp 1649977179
transform 1 0 37996 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_413
timestamp 1649977179
transform 1 0 39100 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_425
timestamp 1649977179
transform 1 0 40204 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_437
timestamp 1649977179
transform 1 0 41308 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_444
timestamp 1649977179
transform 1 0 41952 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_452
timestamp 1649977179
transform 1 0 42688 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_464
timestamp 1649977179
transform 1 0 43792 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_476
timestamp 1649977179
transform 1 0 44896 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_488
timestamp 1649977179
transform 1 0 46000 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_500
timestamp 1649977179
transform 1 0 47104 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_505
timestamp 1649977179
transform 1 0 47564 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_517
timestamp 1649977179
transform 1 0 48668 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_529
timestamp 1649977179
transform 1 0 49772 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_541
timestamp 1649977179
transform 1 0 50876 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_553
timestamp 1649977179
transform 1 0 51980 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_559
timestamp 1649977179
transform 1 0 52532 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_561
timestamp 1649977179
transform 1 0 52716 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_573
timestamp 1649977179
transform 1 0 53820 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_585
timestamp 1649977179
transform 1 0 54924 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_597
timestamp 1649977179
transform 1 0 56028 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_609
timestamp 1649977179
transform 1 0 57132 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_615
timestamp 1649977179
transform 1 0 57684 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_617
timestamp 1649977179
transform 1 0 57868 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_629
timestamp 1649977179
transform 1 0 58972 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_641
timestamp 1649977179
transform 1 0 60076 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_653
timestamp 1649977179
transform 1 0 61180 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_665
timestamp 1649977179
transform 1 0 62284 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_671
timestamp 1649977179
transform 1 0 62836 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_673
timestamp 1649977179
transform 1 0 63020 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_685
timestamp 1649977179
transform 1 0 64124 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_697
timestamp 1649977179
transform 1 0 65228 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_709
timestamp 1649977179
transform 1 0 66332 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_724
timestamp 1649977179
transform 1 0 67712 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_729
timestamp 1649977179
transform 1 0 68172 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_3
timestamp 1649977179
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_15
timestamp 1649977179
transform 1 0 2484 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_23
timestamp 1649977179
transform 1 0 3220 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1649977179
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_29
timestamp 1649977179
transform 1 0 3772 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_37
timestamp 1649977179
transform 1 0 4508 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_41
timestamp 1649977179
transform 1 0 4876 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_61
timestamp 1649977179
transform 1 0 6716 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_70
timestamp 1649977179
transform 1 0 7544 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1649977179
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1649977179
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_88
timestamp 1649977179
transform 1 0 9200 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_110
timestamp 1649977179
transform 1 0 11224 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_114
timestamp 1649977179
transform 1 0 11592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_131
timestamp 1649977179
transform 1 0 13156 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1649977179
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_157
timestamp 1649977179
transform 1 0 15548 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_163
timestamp 1649977179
transform 1 0 16100 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_172
timestamp 1649977179
transform 1 0 16928 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_184
timestamp 1649977179
transform 1 0 18032 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_190
timestamp 1649977179
transform 1 0 18584 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_40_197
timestamp 1649977179
transform 1 0 19228 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_206
timestamp 1649977179
transform 1 0 20056 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_212
timestamp 1649977179
transform 1 0 20608 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_218
timestamp 1649977179
transform 1 0 21160 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_224
timestamp 1649977179
transform 1 0 21712 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_244
timestamp 1649977179
transform 1 0 23552 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_255
timestamp 1649977179
transform 1 0 24564 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_275
timestamp 1649977179
transform 1 0 26404 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_295
timestamp 1649977179
transform 1 0 28244 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 1649977179
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_40_309
timestamp 1649977179
transform 1 0 29532 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_40_328
timestamp 1649977179
transform 1 0 31280 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_340
timestamp 1649977179
transform 1 0 32384 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_345
timestamp 1649977179
transform 1 0 32844 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_351
timestamp 1649977179
transform 1 0 33396 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 1649977179
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_365
timestamp 1649977179
transform 1 0 34684 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_373
timestamp 1649977179
transform 1 0 35420 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_385
timestamp 1649977179
transform 1 0 36524 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_40_409
timestamp 1649977179
transform 1 0 38732 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_417
timestamp 1649977179
transform 1 0 39468 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_40_424
timestamp 1649977179
transform 1 0 40112 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_432
timestamp 1649977179
transform 1 0 40848 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_438
timestamp 1649977179
transform 1 0 41400 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_454
timestamp 1649977179
transform 1 0 42872 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_462
timestamp 1649977179
transform 1 0 43608 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_474
timestamp 1649977179
transform 1 0 44712 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_477
timestamp 1649977179
transform 1 0 44988 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_489
timestamp 1649977179
transform 1 0 46092 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_501
timestamp 1649977179
transform 1 0 47196 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_513
timestamp 1649977179
transform 1 0 48300 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_525
timestamp 1649977179
transform 1 0 49404 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_531
timestamp 1649977179
transform 1 0 49956 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_533
timestamp 1649977179
transform 1 0 50140 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_545
timestamp 1649977179
transform 1 0 51244 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_557
timestamp 1649977179
transform 1 0 52348 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_569
timestamp 1649977179
transform 1 0 53452 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_581
timestamp 1649977179
transform 1 0 54556 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_587
timestamp 1649977179
transform 1 0 55108 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_589
timestamp 1649977179
transform 1 0 55292 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_601
timestamp 1649977179
transform 1 0 56396 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_613
timestamp 1649977179
transform 1 0 57500 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_625
timestamp 1649977179
transform 1 0 58604 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_637
timestamp 1649977179
transform 1 0 59708 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_643
timestamp 1649977179
transform 1 0 60260 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_645
timestamp 1649977179
transform 1 0 60444 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_657
timestamp 1649977179
transform 1 0 61548 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_669
timestamp 1649977179
transform 1 0 62652 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_681
timestamp 1649977179
transform 1 0 63756 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_693
timestamp 1649977179
transform 1 0 64860 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_699
timestamp 1649977179
transform 1 0 65412 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_701
timestamp 1649977179
transform 1 0 65596 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_713
timestamp 1649977179
transform 1 0 66700 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_725
timestamp 1649977179
transform 1 0 67804 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_41_3
timestamp 1649977179
transform 1 0 1380 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_11
timestamp 1649977179
transform 1 0 2116 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_19
timestamp 1649977179
transform 1 0 2852 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_31
timestamp 1649977179
transform 1 0 3956 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_37
timestamp 1649977179
transform 1 0 4508 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_49
timestamp 1649977179
transform 1 0 5612 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_52
timestamp 1649977179
transform 1 0 5888 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_57
timestamp 1649977179
transform 1 0 6348 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_60
timestamp 1649977179
transform 1 0 6624 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_69
timestamp 1649977179
transform 1 0 7452 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_41_82
timestamp 1649977179
transform 1 0 8648 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_88
timestamp 1649977179
transform 1 0 9200 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_100
timestamp 1649977179
transform 1 0 10304 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_118
timestamp 1649977179
transform 1 0 11960 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_140
timestamp 1649977179
transform 1 0 13984 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_149
timestamp 1649977179
transform 1 0 14812 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 1649977179
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1649977179
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_41_169
timestamp 1649977179
transform 1 0 16652 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_41_177
timestamp 1649977179
transform 1 0 17388 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_185
timestamp 1649977179
transform 1 0 18124 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_203
timestamp 1649977179
transform 1 0 19780 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_215
timestamp 1649977179
transform 1 0 20884 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1649977179
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_233
timestamp 1649977179
transform 1 0 22540 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_241
timestamp 1649977179
transform 1 0 23276 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_247
timestamp 1649977179
transform 1 0 23828 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_251
timestamp 1649977179
transform 1 0 24196 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_260
timestamp 1649977179
transform 1 0 25024 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_272
timestamp 1649977179
transform 1 0 26128 0 -1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_41_281
timestamp 1649977179
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_293
timestamp 1649977179
transform 1 0 28060 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_41_312
timestamp 1649977179
transform 1 0 29808 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_324
timestamp 1649977179
transform 1 0 30912 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_337
timestamp 1649977179
transform 1 0 32108 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_343
timestamp 1649977179
transform 1 0 32660 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_354
timestamp 1649977179
transform 1 0 33672 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_358
timestamp 1649977179
transform 1 0 34040 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_365
timestamp 1649977179
transform 1 0 34684 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_381
timestamp 1649977179
transform 1 0 36156 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_389
timestamp 1649977179
transform 1 0 36892 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_41_393
timestamp 1649977179
transform 1 0 37260 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_41_399
timestamp 1649977179
transform 1 0 37812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_411
timestamp 1649977179
transform 1 0 38916 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_432
timestamp 1649977179
transform 1 0 40848 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_444
timestamp 1649977179
transform 1 0 41952 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_449
timestamp 1649977179
transform 1 0 42412 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_453
timestamp 1649977179
transform 1 0 42780 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_466
timestamp 1649977179
transform 1 0 43976 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_478
timestamp 1649977179
transform 1 0 45080 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_490
timestamp 1649977179
transform 1 0 46184 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_502
timestamp 1649977179
transform 1 0 47288 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_505
timestamp 1649977179
transform 1 0 47564 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_517
timestamp 1649977179
transform 1 0 48668 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_529
timestamp 1649977179
transform 1 0 49772 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_541
timestamp 1649977179
transform 1 0 50876 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_553
timestamp 1649977179
transform 1 0 51980 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_559
timestamp 1649977179
transform 1 0 52532 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_561
timestamp 1649977179
transform 1 0 52716 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_573
timestamp 1649977179
transform 1 0 53820 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_585
timestamp 1649977179
transform 1 0 54924 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_597
timestamp 1649977179
transform 1 0 56028 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_609
timestamp 1649977179
transform 1 0 57132 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_615
timestamp 1649977179
transform 1 0 57684 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_617
timestamp 1649977179
transform 1 0 57868 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_629
timestamp 1649977179
transform 1 0 58972 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_641
timestamp 1649977179
transform 1 0 60076 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_653
timestamp 1649977179
transform 1 0 61180 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_665
timestamp 1649977179
transform 1 0 62284 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_671
timestamp 1649977179
transform 1 0 62836 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_673
timestamp 1649977179
transform 1 0 63020 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_685
timestamp 1649977179
transform 1 0 64124 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_697
timestamp 1649977179
transform 1 0 65228 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_709
timestamp 1649977179
transform 1 0 66332 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_724
timestamp 1649977179
transform 1 0 67712 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_729
timestamp 1649977179
transform 1 0 68172 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1649977179
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_15
timestamp 1649977179
transform 1 0 2484 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_42_20
timestamp 1649977179
transform 1 0 2944 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_29
timestamp 1649977179
transform 1 0 3772 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_47
timestamp 1649977179
transform 1 0 5428 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_55
timestamp 1649977179
transform 1 0 6164 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_67
timestamp 1649977179
transform 1 0 7268 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_71
timestamp 1649977179
transform 1 0 7636 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_80
timestamp 1649977179
transform 1 0 8464 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_95
timestamp 1649977179
transform 1 0 9844 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_103
timestamp 1649977179
transform 1 0 10580 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_114
timestamp 1649977179
transform 1 0 11592 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_42_132
timestamp 1649977179
transform 1 0 13248 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_141
timestamp 1649977179
transform 1 0 14076 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_153
timestamp 1649977179
transform 1 0 15180 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_165
timestamp 1649977179
transform 1 0 16284 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_173
timestamp 1649977179
transform 1 0 17020 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_182
timestamp 1649977179
transform 1 0 17848 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_188
timestamp 1649977179
transform 1 0 18400 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_42_197
timestamp 1649977179
transform 1 0 19228 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_205
timestamp 1649977179
transform 1 0 19964 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_217
timestamp 1649977179
transform 1 0 21068 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_221
timestamp 1649977179
transform 1 0 21436 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_225
timestamp 1649977179
transform 1 0 21804 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_42_235
timestamp 1649977179
transform 1 0 22724 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_248
timestamp 1649977179
transform 1 0 23920 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_253
timestamp 1649977179
transform 1 0 24380 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_262
timestamp 1649977179
transform 1 0 25208 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_274
timestamp 1649977179
transform 1 0 26312 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_292
timestamp 1649977179
transform 1 0 27968 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_304
timestamp 1649977179
transform 1 0 29072 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_309
timestamp 1649977179
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_321
timestamp 1649977179
transform 1 0 30636 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_338
timestamp 1649977179
transform 1 0 32200 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_346
timestamp 1649977179
transform 1 0 32936 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_353
timestamp 1649977179
transform 1 0 33580 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_360
timestamp 1649977179
transform 1 0 34224 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_365
timestamp 1649977179
transform 1 0 34684 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_371
timestamp 1649977179
transform 1 0 35236 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_375
timestamp 1649977179
transform 1 0 35604 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_383
timestamp 1649977179
transform 1 0 36340 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_404
timestamp 1649977179
transform 1 0 38272 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_416
timestamp 1649977179
transform 1 0 39376 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_421
timestamp 1649977179
transform 1 0 39836 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_433
timestamp 1649977179
transform 1 0 40940 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_445
timestamp 1649977179
transform 1 0 42044 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_457
timestamp 1649977179
transform 1 0 43148 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_469
timestamp 1649977179
transform 1 0 44252 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_475
timestamp 1649977179
transform 1 0 44804 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_477
timestamp 1649977179
transform 1 0 44988 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_489
timestamp 1649977179
transform 1 0 46092 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_501
timestamp 1649977179
transform 1 0 47196 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_513
timestamp 1649977179
transform 1 0 48300 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_525
timestamp 1649977179
transform 1 0 49404 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_531
timestamp 1649977179
transform 1 0 49956 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_533
timestamp 1649977179
transform 1 0 50140 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_545
timestamp 1649977179
transform 1 0 51244 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_557
timestamp 1649977179
transform 1 0 52348 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_569
timestamp 1649977179
transform 1 0 53452 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_581
timestamp 1649977179
transform 1 0 54556 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_587
timestamp 1649977179
transform 1 0 55108 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_589
timestamp 1649977179
transform 1 0 55292 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_601
timestamp 1649977179
transform 1 0 56396 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_613
timestamp 1649977179
transform 1 0 57500 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_625
timestamp 1649977179
transform 1 0 58604 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_637
timestamp 1649977179
transform 1 0 59708 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_643
timestamp 1649977179
transform 1 0 60260 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_645
timestamp 1649977179
transform 1 0 60444 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_657
timestamp 1649977179
transform 1 0 61548 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_669
timestamp 1649977179
transform 1 0 62652 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_681
timestamp 1649977179
transform 1 0 63756 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_693
timestamp 1649977179
transform 1 0 64860 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_699
timestamp 1649977179
transform 1 0 65412 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_701
timestamp 1649977179
transform 1 0 65596 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_713
timestamp 1649977179
transform 1 0 66700 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_725
timestamp 1649977179
transform 1 0 67804 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_43_3
timestamp 1649977179
transform 1 0 1380 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_11
timestamp 1649977179
transform 1 0 2116 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_18
timestamp 1649977179
transform 1 0 2760 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_30
timestamp 1649977179
transform 1 0 3864 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_36
timestamp 1649977179
transform 1 0 4416 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_48
timestamp 1649977179
transform 1 0 5520 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_43_73
timestamp 1649977179
transform 1 0 7820 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_81
timestamp 1649977179
transform 1 0 8556 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_98
timestamp 1649977179
transform 1 0 10120 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_110
timestamp 1649977179
transform 1 0 11224 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_129
timestamp 1649977179
transform 1 0 12972 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_157
timestamp 1649977179
transform 1 0 15548 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_161
timestamp 1649977179
transform 1 0 15916 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_164
timestamp 1649977179
transform 1 0 16192 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_172
timestamp 1649977179
transform 1 0 16928 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_180
timestamp 1649977179
transform 1 0 17664 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_43_198
timestamp 1649977179
transform 1 0 19320 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_43_214
timestamp 1649977179
transform 1 0 20792 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_222
timestamp 1649977179
transform 1 0 21528 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_241
timestamp 1649977179
transform 1 0 23276 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_250
timestamp 1649977179
transform 1 0 24104 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_256
timestamp 1649977179
transform 1 0 24656 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_276
timestamp 1649977179
transform 1 0 26496 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_281
timestamp 1649977179
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_293
timestamp 1649977179
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_305
timestamp 1649977179
transform 1 0 29164 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_317
timestamp 1649977179
transform 1 0 30268 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_329
timestamp 1649977179
transform 1 0 31372 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1649977179
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_337
timestamp 1649977179
transform 1 0 32108 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_345
timestamp 1649977179
transform 1 0 32844 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_367
timestamp 1649977179
transform 1 0 34868 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_371
timestamp 1649977179
transform 1 0 35236 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_375
timestamp 1649977179
transform 1 0 35604 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_387
timestamp 1649977179
transform 1 0 36708 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1649977179
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_393
timestamp 1649977179
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_405
timestamp 1649977179
transform 1 0 38364 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_417
timestamp 1649977179
transform 1 0 39468 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_429
timestamp 1649977179
transform 1 0 40572 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_441
timestamp 1649977179
transform 1 0 41676 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_447
timestamp 1649977179
transform 1 0 42228 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_449
timestamp 1649977179
transform 1 0 42412 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_461
timestamp 1649977179
transform 1 0 43516 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_473
timestamp 1649977179
transform 1 0 44620 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_485
timestamp 1649977179
transform 1 0 45724 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_497
timestamp 1649977179
transform 1 0 46828 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_503
timestamp 1649977179
transform 1 0 47380 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_505
timestamp 1649977179
transform 1 0 47564 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_517
timestamp 1649977179
transform 1 0 48668 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_529
timestamp 1649977179
transform 1 0 49772 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_541
timestamp 1649977179
transform 1 0 50876 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_553
timestamp 1649977179
transform 1 0 51980 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_559
timestamp 1649977179
transform 1 0 52532 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_561
timestamp 1649977179
transform 1 0 52716 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_573
timestamp 1649977179
transform 1 0 53820 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_585
timestamp 1649977179
transform 1 0 54924 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_597
timestamp 1649977179
transform 1 0 56028 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_609
timestamp 1649977179
transform 1 0 57132 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_615
timestamp 1649977179
transform 1 0 57684 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_617
timestamp 1649977179
transform 1 0 57868 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_629
timestamp 1649977179
transform 1 0 58972 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_641
timestamp 1649977179
transform 1 0 60076 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_653
timestamp 1649977179
transform 1 0 61180 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_665
timestamp 1649977179
transform 1 0 62284 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_671
timestamp 1649977179
transform 1 0 62836 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_673
timestamp 1649977179
transform 1 0 63020 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_685
timestamp 1649977179
transform 1 0 64124 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_697
timestamp 1649977179
transform 1 0 65228 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_709
timestamp 1649977179
transform 1 0 66332 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_721
timestamp 1649977179
transform 1 0 67436 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_727
timestamp 1649977179
transform 1 0 67988 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_729
timestamp 1649977179
transform 1 0 68172 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1649977179
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_15
timestamp 1649977179
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1649977179
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1649977179
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_41
timestamp 1649977179
transform 1 0 4876 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_44_49
timestamp 1649977179
transform 1 0 5612 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_61
timestamp 1649977179
transform 1 0 6716 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_67
timestamp 1649977179
transform 1 0 7268 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_73
timestamp 1649977179
transform 1 0 7820 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_81
timestamp 1649977179
transform 1 0 8556 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_85
timestamp 1649977179
transform 1 0 8924 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_93
timestamp 1649977179
transform 1 0 9660 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_99
timestamp 1649977179
transform 1 0 10212 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_113
timestamp 1649977179
transform 1 0 11500 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_119
timestamp 1649977179
transform 1 0 12052 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_127
timestamp 1649977179
transform 1 0 12788 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_134
timestamp 1649977179
transform 1 0 13432 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_44_151
timestamp 1649977179
transform 1 0 14996 0 1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_44_175
timestamp 1649977179
transform 1 0 17204 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_187
timestamp 1649977179
transform 1 0 18308 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1649977179
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_197
timestamp 1649977179
transform 1 0 19228 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_203
timestamp 1649977179
transform 1 0 19780 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_215
timestamp 1649977179
transform 1 0 20884 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_220
timestamp 1649977179
transform 1 0 21344 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_232
timestamp 1649977179
transform 1 0 22448 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_244
timestamp 1649977179
transform 1 0 23552 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_44_253
timestamp 1649977179
transform 1 0 24380 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_44_264
timestamp 1649977179
transform 1 0 25392 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_270
timestamp 1649977179
transform 1 0 25944 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_282
timestamp 1649977179
transform 1 0 27048 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_294
timestamp 1649977179
transform 1 0 28152 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_306
timestamp 1649977179
transform 1 0 29256 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_309
timestamp 1649977179
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_321
timestamp 1649977179
transform 1 0 30636 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_333
timestamp 1649977179
transform 1 0 31740 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_337
timestamp 1649977179
transform 1 0 32108 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_350
timestamp 1649977179
transform 1 0 33304 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_356
timestamp 1649977179
transform 1 0 33856 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_360
timestamp 1649977179
transform 1 0 34224 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_44_365
timestamp 1649977179
transform 1 0 34684 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_373
timestamp 1649977179
transform 1 0 35420 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_389
timestamp 1649977179
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_401
timestamp 1649977179
transform 1 0 37996 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_413
timestamp 1649977179
transform 1 0 39100 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_419
timestamp 1649977179
transform 1 0 39652 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_421
timestamp 1649977179
transform 1 0 39836 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_433
timestamp 1649977179
transform 1 0 40940 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_445
timestamp 1649977179
transform 1 0 42044 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_457
timestamp 1649977179
transform 1 0 43148 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_469
timestamp 1649977179
transform 1 0 44252 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_475
timestamp 1649977179
transform 1 0 44804 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_477
timestamp 1649977179
transform 1 0 44988 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_489
timestamp 1649977179
transform 1 0 46092 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_501
timestamp 1649977179
transform 1 0 47196 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_513
timestamp 1649977179
transform 1 0 48300 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_525
timestamp 1649977179
transform 1 0 49404 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_531
timestamp 1649977179
transform 1 0 49956 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_533
timestamp 1649977179
transform 1 0 50140 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_545
timestamp 1649977179
transform 1 0 51244 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_557
timestamp 1649977179
transform 1 0 52348 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_569
timestamp 1649977179
transform 1 0 53452 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_581
timestamp 1649977179
transform 1 0 54556 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_587
timestamp 1649977179
transform 1 0 55108 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_589
timestamp 1649977179
transform 1 0 55292 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_601
timestamp 1649977179
transform 1 0 56396 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_613
timestamp 1649977179
transform 1 0 57500 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_625
timestamp 1649977179
transform 1 0 58604 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_637
timestamp 1649977179
transform 1 0 59708 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_643
timestamp 1649977179
transform 1 0 60260 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_645
timestamp 1649977179
transform 1 0 60444 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_657
timestamp 1649977179
transform 1 0 61548 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_669
timestamp 1649977179
transform 1 0 62652 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_681
timestamp 1649977179
transform 1 0 63756 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_693
timestamp 1649977179
transform 1 0 64860 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_699
timestamp 1649977179
transform 1 0 65412 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_701
timestamp 1649977179
transform 1 0 65596 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_713
timestamp 1649977179
transform 1 0 66700 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_725
timestamp 1649977179
transform 1 0 67804 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_729
timestamp 1649977179
transform 1 0 68172 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_3
timestamp 1649977179
transform 1 0 1380 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_11
timestamp 1649977179
transform 1 0 2116 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_17
timestamp 1649977179
transform 1 0 2668 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_37
timestamp 1649977179
transform 1 0 4508 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_43
timestamp 1649977179
transform 1 0 5060 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_47
timestamp 1649977179
transform 1 0 5428 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1649977179
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_77
timestamp 1649977179
transform 1 0 8188 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_81
timestamp 1649977179
transform 1 0 8556 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_84
timestamp 1649977179
transform 1 0 8832 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_93
timestamp 1649977179
transform 1 0 9660 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_99
timestamp 1649977179
transform 1 0 10212 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_102
timestamp 1649977179
transform 1 0 10488 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_108
timestamp 1649977179
transform 1 0 11040 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_117
timestamp 1649977179
transform 1 0 11868 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_123
timestamp 1649977179
transform 1 0 12420 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_127
timestamp 1649977179
transform 1 0 12788 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_130
timestamp 1649977179
transform 1 0 13064 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_142
timestamp 1649977179
transform 1 0 14168 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_148
timestamp 1649977179
transform 1 0 14720 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_160
timestamp 1649977179
transform 1 0 15824 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_45_169
timestamp 1649977179
transform 1 0 16652 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_177
timestamp 1649977179
transform 1 0 17388 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_45_196
timestamp 1649977179
transform 1 0 19136 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_202
timestamp 1649977179
transform 1 0 19688 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_211
timestamp 1649977179
transform 1 0 20516 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_220
timestamp 1649977179
transform 1 0 21344 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_225
timestamp 1649977179
transform 1 0 21804 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_245
timestamp 1649977179
transform 1 0 23644 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_269
timestamp 1649977179
transform 1 0 25852 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_277
timestamp 1649977179
transform 1 0 26588 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_284
timestamp 1649977179
transform 1 0 27232 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_290
timestamp 1649977179
transform 1 0 27784 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_302
timestamp 1649977179
transform 1 0 28888 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_314
timestamp 1649977179
transform 1 0 29992 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_326
timestamp 1649977179
transform 1 0 31096 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_334
timestamp 1649977179
transform 1 0 31832 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_337
timestamp 1649977179
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_349
timestamp 1649977179
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_361
timestamp 1649977179
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_373
timestamp 1649977179
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_385
timestamp 1649977179
transform 1 0 36524 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1649977179
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_393
timestamp 1649977179
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_405
timestamp 1649977179
transform 1 0 38364 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_417
timestamp 1649977179
transform 1 0 39468 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_429
timestamp 1649977179
transform 1 0 40572 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_441
timestamp 1649977179
transform 1 0 41676 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_447
timestamp 1649977179
transform 1 0 42228 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_449
timestamp 1649977179
transform 1 0 42412 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_461
timestamp 1649977179
transform 1 0 43516 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_473
timestamp 1649977179
transform 1 0 44620 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_485
timestamp 1649977179
transform 1 0 45724 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_497
timestamp 1649977179
transform 1 0 46828 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_503
timestamp 1649977179
transform 1 0 47380 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_505
timestamp 1649977179
transform 1 0 47564 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_517
timestamp 1649977179
transform 1 0 48668 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_529
timestamp 1649977179
transform 1 0 49772 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_541
timestamp 1649977179
transform 1 0 50876 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_553
timestamp 1649977179
transform 1 0 51980 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_559
timestamp 1649977179
transform 1 0 52532 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_561
timestamp 1649977179
transform 1 0 52716 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_573
timestamp 1649977179
transform 1 0 53820 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_585
timestamp 1649977179
transform 1 0 54924 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_597
timestamp 1649977179
transform 1 0 56028 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_609
timestamp 1649977179
transform 1 0 57132 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_615
timestamp 1649977179
transform 1 0 57684 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_617
timestamp 1649977179
transform 1 0 57868 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_629
timestamp 1649977179
transform 1 0 58972 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_641
timestamp 1649977179
transform 1 0 60076 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_653
timestamp 1649977179
transform 1 0 61180 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_665
timestamp 1649977179
transform 1 0 62284 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_671
timestamp 1649977179
transform 1 0 62836 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_673
timestamp 1649977179
transform 1 0 63020 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_685
timestamp 1649977179
transform 1 0 64124 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_697
timestamp 1649977179
transform 1 0 65228 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_709
timestamp 1649977179
transform 1 0 66332 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_721
timestamp 1649977179
transform 1 0 67436 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_727
timestamp 1649977179
transform 1 0 67988 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_729
timestamp 1649977179
transform 1 0 68172 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_3
timestamp 1649977179
transform 1 0 1380 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_7
timestamp 1649977179
transform 1 0 1748 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_15
timestamp 1649977179
transform 1 0 2484 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_21
timestamp 1649977179
transform 1 0 3036 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1649977179
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_29
timestamp 1649977179
transform 1 0 3772 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_53
timestamp 1649977179
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_65
timestamp 1649977179
transform 1 0 7084 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_68
timestamp 1649977179
transform 1 0 7360 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_80
timestamp 1649977179
transform 1 0 8464 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_87
timestamp 1649977179
transform 1 0 9108 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_91
timestamp 1649977179
transform 1 0 9476 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_100
timestamp 1649977179
transform 1 0 10304 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_109
timestamp 1649977179
transform 1 0 11132 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_115
timestamp 1649977179
transform 1 0 11684 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_132
timestamp 1649977179
transform 1 0 13248 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_141
timestamp 1649977179
transform 1 0 14076 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_152
timestamp 1649977179
transform 1 0 15088 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_172
timestamp 1649977179
transform 1 0 16928 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_46_186
timestamp 1649977179
transform 1 0 18216 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_194
timestamp 1649977179
transform 1 0 18952 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_46_197
timestamp 1649977179
transform 1 0 19228 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_200
timestamp 1649977179
transform 1 0 19504 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_212
timestamp 1649977179
transform 1 0 20608 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_216
timestamp 1649977179
transform 1 0 20976 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_233
timestamp 1649977179
transform 1 0 22540 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_245
timestamp 1649977179
transform 1 0 23644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1649977179
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_253
timestamp 1649977179
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_265
timestamp 1649977179
transform 1 0 25484 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_269
timestamp 1649977179
transform 1 0 25852 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_290
timestamp 1649977179
transform 1 0 27784 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_302
timestamp 1649977179
transform 1 0 28888 0 1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_46_309
timestamp 1649977179
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_321
timestamp 1649977179
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_333
timestamp 1649977179
transform 1 0 31740 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_345
timestamp 1649977179
transform 1 0 32844 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_357
timestamp 1649977179
transform 1 0 33948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1649977179
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_365
timestamp 1649977179
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_377
timestamp 1649977179
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_389
timestamp 1649977179
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_401
timestamp 1649977179
transform 1 0 37996 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_413
timestamp 1649977179
transform 1 0 39100 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_419
timestamp 1649977179
transform 1 0 39652 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_421
timestamp 1649977179
transform 1 0 39836 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_433
timestamp 1649977179
transform 1 0 40940 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_445
timestamp 1649977179
transform 1 0 42044 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_457
timestamp 1649977179
transform 1 0 43148 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_469
timestamp 1649977179
transform 1 0 44252 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_475
timestamp 1649977179
transform 1 0 44804 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_477
timestamp 1649977179
transform 1 0 44988 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_489
timestamp 1649977179
transform 1 0 46092 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_501
timestamp 1649977179
transform 1 0 47196 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_513
timestamp 1649977179
transform 1 0 48300 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_525
timestamp 1649977179
transform 1 0 49404 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_531
timestamp 1649977179
transform 1 0 49956 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_533
timestamp 1649977179
transform 1 0 50140 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_545
timestamp 1649977179
transform 1 0 51244 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_557
timestamp 1649977179
transform 1 0 52348 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_569
timestamp 1649977179
transform 1 0 53452 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_581
timestamp 1649977179
transform 1 0 54556 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_587
timestamp 1649977179
transform 1 0 55108 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_589
timestamp 1649977179
transform 1 0 55292 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_601
timestamp 1649977179
transform 1 0 56396 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_613
timestamp 1649977179
transform 1 0 57500 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_625
timestamp 1649977179
transform 1 0 58604 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_637
timestamp 1649977179
transform 1 0 59708 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_643
timestamp 1649977179
transform 1 0 60260 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_645
timestamp 1649977179
transform 1 0 60444 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_657
timestamp 1649977179
transform 1 0 61548 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_669
timestamp 1649977179
transform 1 0 62652 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_681
timestamp 1649977179
transform 1 0 63756 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_693
timestamp 1649977179
transform 1 0 64860 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_699
timestamp 1649977179
transform 1 0 65412 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_701
timestamp 1649977179
transform 1 0 65596 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_713
timestamp 1649977179
transform 1 0 66700 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_725
timestamp 1649977179
transform 1 0 67804 0 1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_47_3
timestamp 1649977179
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_15
timestamp 1649977179
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_27
timestamp 1649977179
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_39
timestamp 1649977179
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1649977179
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1649977179
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_57
timestamp 1649977179
transform 1 0 6348 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_65
timestamp 1649977179
transform 1 0 7084 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_47_76
timestamp 1649977179
transform 1 0 8096 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_84
timestamp 1649977179
transform 1 0 8832 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_93
timestamp 1649977179
transform 1 0 9660 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_101
timestamp 1649977179
transform 1 0 10396 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_104
timestamp 1649977179
transform 1 0 10672 0 -1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_47_116
timestamp 1649977179
transform 1 0 11776 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_128
timestamp 1649977179
transform 1 0 12880 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_47_141
timestamp 1649977179
transform 1 0 14076 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_149
timestamp 1649977179
transform 1 0 14812 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_155
timestamp 1649977179
transform 1 0 15364 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1649977179
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_47_169
timestamp 1649977179
transform 1 0 16652 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_175
timestamp 1649977179
transform 1 0 17204 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_178
timestamp 1649977179
transform 1 0 17480 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_182
timestamp 1649977179
transform 1 0 17848 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_188
timestamp 1649977179
transform 1 0 18400 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_196
timestamp 1649977179
transform 1 0 19136 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_203
timestamp 1649977179
transform 1 0 19780 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_212
timestamp 1649977179
transform 1 0 20608 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_225
timestamp 1649977179
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_237
timestamp 1649977179
transform 1 0 22908 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_47_249
timestamp 1649977179
transform 1 0 24012 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_256
timestamp 1649977179
transform 1 0 24656 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_264
timestamp 1649977179
transform 1 0 25392 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_47_269
timestamp 1649977179
transform 1 0 25852 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_277
timestamp 1649977179
transform 1 0 26588 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_47_281
timestamp 1649977179
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_293
timestamp 1649977179
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_305
timestamp 1649977179
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_317
timestamp 1649977179
transform 1 0 30268 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_329
timestamp 1649977179
transform 1 0 31372 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 1649977179
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_337
timestamp 1649977179
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_349
timestamp 1649977179
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_361
timestamp 1649977179
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_373
timestamp 1649977179
transform 1 0 35420 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_385
timestamp 1649977179
transform 1 0 36524 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_391
timestamp 1649977179
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_393
timestamp 1649977179
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_405
timestamp 1649977179
transform 1 0 38364 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_417
timestamp 1649977179
transform 1 0 39468 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_429
timestamp 1649977179
transform 1 0 40572 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_441
timestamp 1649977179
transform 1 0 41676 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_447
timestamp 1649977179
transform 1 0 42228 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_449
timestamp 1649977179
transform 1 0 42412 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_461
timestamp 1649977179
transform 1 0 43516 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_473
timestamp 1649977179
transform 1 0 44620 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_485
timestamp 1649977179
transform 1 0 45724 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_497
timestamp 1649977179
transform 1 0 46828 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_503
timestamp 1649977179
transform 1 0 47380 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_505
timestamp 1649977179
transform 1 0 47564 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_517
timestamp 1649977179
transform 1 0 48668 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_529
timestamp 1649977179
transform 1 0 49772 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_541
timestamp 1649977179
transform 1 0 50876 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_553
timestamp 1649977179
transform 1 0 51980 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_559
timestamp 1649977179
transform 1 0 52532 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_561
timestamp 1649977179
transform 1 0 52716 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_573
timestamp 1649977179
transform 1 0 53820 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_585
timestamp 1649977179
transform 1 0 54924 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_597
timestamp 1649977179
transform 1 0 56028 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_609
timestamp 1649977179
transform 1 0 57132 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_615
timestamp 1649977179
transform 1 0 57684 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_617
timestamp 1649977179
transform 1 0 57868 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_629
timestamp 1649977179
transform 1 0 58972 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_641
timestamp 1649977179
transform 1 0 60076 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_653
timestamp 1649977179
transform 1 0 61180 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_665
timestamp 1649977179
transform 1 0 62284 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_671
timestamp 1649977179
transform 1 0 62836 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_673
timestamp 1649977179
transform 1 0 63020 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_685
timestamp 1649977179
transform 1 0 64124 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_697
timestamp 1649977179
transform 1 0 65228 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_709
timestamp 1649977179
transform 1 0 66332 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_724
timestamp 1649977179
transform 1 0 67712 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_729
timestamp 1649977179
transform 1 0 68172 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1649977179
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1649977179
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1649977179
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_41
timestamp 1649977179
transform 1 0 4876 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_50
timestamp 1649977179
transform 1 0 5704 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_57
timestamp 1649977179
transform 1 0 6348 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_64
timestamp 1649977179
transform 1 0 6992 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_48_80
timestamp 1649977179
transform 1 0 8464 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_85
timestamp 1649977179
transform 1 0 8924 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_97
timestamp 1649977179
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_109
timestamp 1649977179
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_121
timestamp 1649977179
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1649977179
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1649977179
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_141
timestamp 1649977179
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_153
timestamp 1649977179
transform 1 0 15180 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_48_160
timestamp 1649977179
transform 1 0 15824 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_166
timestamp 1649977179
transform 1 0 16376 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_174
timestamp 1649977179
transform 1 0 17112 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_180
timestamp 1649977179
transform 1 0 17664 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_187
timestamp 1649977179
transform 1 0 18308 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1649977179
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_197
timestamp 1649977179
transform 1 0 19228 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_201
timestamp 1649977179
transform 1 0 19596 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_208
timestamp 1649977179
transform 1 0 20240 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_220
timestamp 1649977179
transform 1 0 21344 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_236
timestamp 1649977179
transform 1 0 22816 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_248
timestamp 1649977179
transform 1 0 23920 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_253
timestamp 1649977179
transform 1 0 24380 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_264
timestamp 1649977179
transform 1 0 25392 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_280
timestamp 1649977179
transform 1 0 26864 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_292
timestamp 1649977179
transform 1 0 27968 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_304
timestamp 1649977179
transform 1 0 29072 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_309
timestamp 1649977179
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_321
timestamp 1649977179
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_333
timestamp 1649977179
transform 1 0 31740 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_345
timestamp 1649977179
transform 1 0 32844 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_357
timestamp 1649977179
transform 1 0 33948 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 1649977179
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_365
timestamp 1649977179
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_377
timestamp 1649977179
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_389
timestamp 1649977179
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_401
timestamp 1649977179
transform 1 0 37996 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_413
timestamp 1649977179
transform 1 0 39100 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_419
timestamp 1649977179
transform 1 0 39652 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_421
timestamp 1649977179
transform 1 0 39836 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_433
timestamp 1649977179
transform 1 0 40940 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_445
timestamp 1649977179
transform 1 0 42044 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_457
timestamp 1649977179
transform 1 0 43148 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_469
timestamp 1649977179
transform 1 0 44252 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_475
timestamp 1649977179
transform 1 0 44804 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_477
timestamp 1649977179
transform 1 0 44988 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_489
timestamp 1649977179
transform 1 0 46092 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_501
timestamp 1649977179
transform 1 0 47196 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_513
timestamp 1649977179
transform 1 0 48300 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_525
timestamp 1649977179
transform 1 0 49404 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_531
timestamp 1649977179
transform 1 0 49956 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_533
timestamp 1649977179
transform 1 0 50140 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_545
timestamp 1649977179
transform 1 0 51244 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_557
timestamp 1649977179
transform 1 0 52348 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_569
timestamp 1649977179
transform 1 0 53452 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_581
timestamp 1649977179
transform 1 0 54556 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_587
timestamp 1649977179
transform 1 0 55108 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_589
timestamp 1649977179
transform 1 0 55292 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_601
timestamp 1649977179
transform 1 0 56396 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_613
timestamp 1649977179
transform 1 0 57500 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_625
timestamp 1649977179
transform 1 0 58604 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_637
timestamp 1649977179
transform 1 0 59708 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_643
timestamp 1649977179
transform 1 0 60260 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_645
timestamp 1649977179
transform 1 0 60444 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_657
timestamp 1649977179
transform 1 0 61548 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_669
timestamp 1649977179
transform 1 0 62652 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_681
timestamp 1649977179
transform 1 0 63756 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_693
timestamp 1649977179
transform 1 0 64860 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_699
timestamp 1649977179
transform 1 0 65412 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_701
timestamp 1649977179
transform 1 0 65596 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_713
timestamp 1649977179
transform 1 0 66700 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_725
timestamp 1649977179
transform 1 0 67804 0 1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1649977179
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 1649977179
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_27
timestamp 1649977179
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_39
timestamp 1649977179
transform 1 0 4692 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_52
timestamp 1649977179
transform 1 0 5888 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_57
timestamp 1649977179
transform 1 0 6348 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_49_64
timestamp 1649977179
transform 1 0 6992 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_70
timestamp 1649977179
transform 1 0 7544 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_74
timestamp 1649977179
transform 1 0 7912 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_80
timestamp 1649977179
transform 1 0 8464 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_86
timestamp 1649977179
transform 1 0 9016 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_89
timestamp 1649977179
transform 1 0 9292 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_101
timestamp 1649977179
transform 1 0 10396 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_109
timestamp 1649977179
transform 1 0 11132 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_49_113
timestamp 1649977179
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_125
timestamp 1649977179
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_137
timestamp 1649977179
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_149
timestamp 1649977179
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_161
timestamp 1649977179
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1649977179
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_169
timestamp 1649977179
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_181
timestamp 1649977179
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_193
timestamp 1649977179
transform 1 0 18860 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_201
timestamp 1649977179
transform 1 0 19596 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_213
timestamp 1649977179
transform 1 0 20700 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_221
timestamp 1649977179
transform 1 0 21436 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_49_225
timestamp 1649977179
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_237
timestamp 1649977179
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_249
timestamp 1649977179
transform 1 0 24012 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_49_255
timestamp 1649977179
transform 1 0 24564 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_267
timestamp 1649977179
transform 1 0 25668 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1649977179
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_281
timestamp 1649977179
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_293
timestamp 1649977179
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_305
timestamp 1649977179
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_317
timestamp 1649977179
transform 1 0 30268 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_329
timestamp 1649977179
transform 1 0 31372 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1649977179
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_337
timestamp 1649977179
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_349
timestamp 1649977179
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_361
timestamp 1649977179
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_373
timestamp 1649977179
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_385
timestamp 1649977179
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 1649977179
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_393
timestamp 1649977179
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_405
timestamp 1649977179
transform 1 0 38364 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_417
timestamp 1649977179
transform 1 0 39468 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_429
timestamp 1649977179
transform 1 0 40572 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_441
timestamp 1649977179
transform 1 0 41676 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_447
timestamp 1649977179
transform 1 0 42228 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_449
timestamp 1649977179
transform 1 0 42412 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_461
timestamp 1649977179
transform 1 0 43516 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_473
timestamp 1649977179
transform 1 0 44620 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_485
timestamp 1649977179
transform 1 0 45724 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_497
timestamp 1649977179
transform 1 0 46828 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_503
timestamp 1649977179
transform 1 0 47380 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_505
timestamp 1649977179
transform 1 0 47564 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_517
timestamp 1649977179
transform 1 0 48668 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_529
timestamp 1649977179
transform 1 0 49772 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_541
timestamp 1649977179
transform 1 0 50876 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_553
timestamp 1649977179
transform 1 0 51980 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_559
timestamp 1649977179
transform 1 0 52532 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_561
timestamp 1649977179
transform 1 0 52716 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_573
timestamp 1649977179
transform 1 0 53820 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_585
timestamp 1649977179
transform 1 0 54924 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_597
timestamp 1649977179
transform 1 0 56028 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_609
timestamp 1649977179
transform 1 0 57132 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_615
timestamp 1649977179
transform 1 0 57684 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_617
timestamp 1649977179
transform 1 0 57868 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_629
timestamp 1649977179
transform 1 0 58972 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_641
timestamp 1649977179
transform 1 0 60076 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_653
timestamp 1649977179
transform 1 0 61180 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_665
timestamp 1649977179
transform 1 0 62284 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_671
timestamp 1649977179
transform 1 0 62836 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_673
timestamp 1649977179
transform 1 0 63020 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_685
timestamp 1649977179
transform 1 0 64124 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_697
timestamp 1649977179
transform 1 0 65228 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_709
timestamp 1649977179
transform 1 0 66332 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_721
timestamp 1649977179
transform 1 0 67436 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_727
timestamp 1649977179
transform 1 0 67988 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_729
timestamp 1649977179
transform 1 0 68172 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_3
timestamp 1649977179
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_15
timestamp 1649977179
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1649977179
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1649977179
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_41
timestamp 1649977179
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_53
timestamp 1649977179
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_65
timestamp 1649977179
transform 1 0 7084 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_70
timestamp 1649977179
transform 1 0 7544 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_82
timestamp 1649977179
transform 1 0 8648 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_85
timestamp 1649977179
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_97
timestamp 1649977179
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_109
timestamp 1649977179
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_121
timestamp 1649977179
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1649977179
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1649977179
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_141
timestamp 1649977179
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_153
timestamp 1649977179
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_165
timestamp 1649977179
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_177
timestamp 1649977179
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_189
timestamp 1649977179
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1649977179
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_197
timestamp 1649977179
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_209
timestamp 1649977179
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_221
timestamp 1649977179
transform 1 0 21436 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_233
timestamp 1649977179
transform 1 0 22540 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_245
timestamp 1649977179
transform 1 0 23644 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1649977179
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_253
timestamp 1649977179
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_265
timestamp 1649977179
transform 1 0 25484 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_271
timestamp 1649977179
transform 1 0 26036 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_284
timestamp 1649977179
transform 1 0 27232 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_296
timestamp 1649977179
transform 1 0 28336 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_309
timestamp 1649977179
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_321
timestamp 1649977179
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_333
timestamp 1649977179
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_345
timestamp 1649977179
transform 1 0 32844 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_357
timestamp 1649977179
transform 1 0 33948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1649977179
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_365
timestamp 1649977179
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_377
timestamp 1649977179
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_389
timestamp 1649977179
transform 1 0 36892 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_401
timestamp 1649977179
transform 1 0 37996 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_413
timestamp 1649977179
transform 1 0 39100 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_419
timestamp 1649977179
transform 1 0 39652 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_421
timestamp 1649977179
transform 1 0 39836 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_433
timestamp 1649977179
transform 1 0 40940 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_445
timestamp 1649977179
transform 1 0 42044 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_457
timestamp 1649977179
transform 1 0 43148 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_469
timestamp 1649977179
transform 1 0 44252 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_475
timestamp 1649977179
transform 1 0 44804 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_477
timestamp 1649977179
transform 1 0 44988 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_489
timestamp 1649977179
transform 1 0 46092 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_501
timestamp 1649977179
transform 1 0 47196 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_513
timestamp 1649977179
transform 1 0 48300 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_525
timestamp 1649977179
transform 1 0 49404 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_531
timestamp 1649977179
transform 1 0 49956 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_533
timestamp 1649977179
transform 1 0 50140 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_545
timestamp 1649977179
transform 1 0 51244 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_557
timestamp 1649977179
transform 1 0 52348 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_569
timestamp 1649977179
transform 1 0 53452 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_581
timestamp 1649977179
transform 1 0 54556 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_587
timestamp 1649977179
transform 1 0 55108 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_589
timestamp 1649977179
transform 1 0 55292 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_601
timestamp 1649977179
transform 1 0 56396 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_613
timestamp 1649977179
transform 1 0 57500 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_625
timestamp 1649977179
transform 1 0 58604 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_637
timestamp 1649977179
transform 1 0 59708 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_643
timestamp 1649977179
transform 1 0 60260 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_645
timestamp 1649977179
transform 1 0 60444 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_657
timestamp 1649977179
transform 1 0 61548 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_669
timestamp 1649977179
transform 1 0 62652 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_681
timestamp 1649977179
transform 1 0 63756 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_693
timestamp 1649977179
transform 1 0 64860 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_699
timestamp 1649977179
transform 1 0 65412 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_701
timestamp 1649977179
transform 1 0 65596 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_713
timestamp 1649977179
transform 1 0 66700 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_725
timestamp 1649977179
transform 1 0 67804 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_729
timestamp 1649977179
transform 1 0 68172 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1649977179
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1649977179
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_27
timestamp 1649977179
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_39
timestamp 1649977179
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1649977179
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1649977179
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_57
timestamp 1649977179
transform 1 0 6348 0 -1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_51_76
timestamp 1649977179
transform 1 0 8096 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_88
timestamp 1649977179
transform 1 0 9200 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_100
timestamp 1649977179
transform 1 0 10304 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_113
timestamp 1649977179
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_125
timestamp 1649977179
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_137
timestamp 1649977179
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_149
timestamp 1649977179
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_161
timestamp 1649977179
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1649977179
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_169
timestamp 1649977179
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_181
timestamp 1649977179
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_193
timestamp 1649977179
transform 1 0 18860 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_205
timestamp 1649977179
transform 1 0 19964 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_217
timestamp 1649977179
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1649977179
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_225
timestamp 1649977179
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_237
timestamp 1649977179
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_249
timestamp 1649977179
transform 1 0 24012 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_261
timestamp 1649977179
transform 1 0 25116 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_273
timestamp 1649977179
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1649977179
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_281
timestamp 1649977179
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_293
timestamp 1649977179
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_305
timestamp 1649977179
transform 1 0 29164 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_317
timestamp 1649977179
transform 1 0 30268 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_329
timestamp 1649977179
transform 1 0 31372 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_335
timestamp 1649977179
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_337
timestamp 1649977179
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_349
timestamp 1649977179
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_361
timestamp 1649977179
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_373
timestamp 1649977179
transform 1 0 35420 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_385
timestamp 1649977179
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1649977179
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_393
timestamp 1649977179
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_405
timestamp 1649977179
transform 1 0 38364 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_417
timestamp 1649977179
transform 1 0 39468 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_429
timestamp 1649977179
transform 1 0 40572 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_441
timestamp 1649977179
transform 1 0 41676 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_447
timestamp 1649977179
transform 1 0 42228 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_449
timestamp 1649977179
transform 1 0 42412 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_461
timestamp 1649977179
transform 1 0 43516 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_473
timestamp 1649977179
transform 1 0 44620 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_485
timestamp 1649977179
transform 1 0 45724 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_497
timestamp 1649977179
transform 1 0 46828 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_503
timestamp 1649977179
transform 1 0 47380 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_505
timestamp 1649977179
transform 1 0 47564 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_517
timestamp 1649977179
transform 1 0 48668 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_529
timestamp 1649977179
transform 1 0 49772 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_541
timestamp 1649977179
transform 1 0 50876 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_553
timestamp 1649977179
transform 1 0 51980 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_559
timestamp 1649977179
transform 1 0 52532 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_561
timestamp 1649977179
transform 1 0 52716 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_573
timestamp 1649977179
transform 1 0 53820 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_585
timestamp 1649977179
transform 1 0 54924 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_597
timestamp 1649977179
transform 1 0 56028 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_609
timestamp 1649977179
transform 1 0 57132 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_615
timestamp 1649977179
transform 1 0 57684 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_617
timestamp 1649977179
transform 1 0 57868 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_629
timestamp 1649977179
transform 1 0 58972 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_641
timestamp 1649977179
transform 1 0 60076 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_653
timestamp 1649977179
transform 1 0 61180 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_665
timestamp 1649977179
transform 1 0 62284 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_671
timestamp 1649977179
transform 1 0 62836 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_673
timestamp 1649977179
transform 1 0 63020 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_685
timestamp 1649977179
transform 1 0 64124 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_697
timestamp 1649977179
transform 1 0 65228 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_709
timestamp 1649977179
transform 1 0 66332 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_721
timestamp 1649977179
transform 1 0 67436 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_727
timestamp 1649977179
transform 1 0 67988 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_729
timestamp 1649977179
transform 1 0 68172 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_3
timestamp 1649977179
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_15
timestamp 1649977179
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1649977179
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1649977179
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1649977179
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_53
timestamp 1649977179
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_65
timestamp 1649977179
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1649977179
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1649977179
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_85
timestamp 1649977179
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_97
timestamp 1649977179
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_109
timestamp 1649977179
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_121
timestamp 1649977179
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1649977179
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1649977179
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_141
timestamp 1649977179
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_153
timestamp 1649977179
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_165
timestamp 1649977179
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_177
timestamp 1649977179
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_189
timestamp 1649977179
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1649977179
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_197
timestamp 1649977179
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_209
timestamp 1649977179
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_221
timestamp 1649977179
transform 1 0 21436 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_233
timestamp 1649977179
transform 1 0 22540 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_245
timestamp 1649977179
transform 1 0 23644 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1649977179
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_253
timestamp 1649977179
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_265
timestamp 1649977179
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_277
timestamp 1649977179
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_289
timestamp 1649977179
transform 1 0 27692 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_301
timestamp 1649977179
transform 1 0 28796 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1649977179
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_309
timestamp 1649977179
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_321
timestamp 1649977179
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_333
timestamp 1649977179
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_345
timestamp 1649977179
transform 1 0 32844 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_357
timestamp 1649977179
transform 1 0 33948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_363
timestamp 1649977179
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_365
timestamp 1649977179
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_377
timestamp 1649977179
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_389
timestamp 1649977179
transform 1 0 36892 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_401
timestamp 1649977179
transform 1 0 37996 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_413
timestamp 1649977179
transform 1 0 39100 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_419
timestamp 1649977179
transform 1 0 39652 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_421
timestamp 1649977179
transform 1 0 39836 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_433
timestamp 1649977179
transform 1 0 40940 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_445
timestamp 1649977179
transform 1 0 42044 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_457
timestamp 1649977179
transform 1 0 43148 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_469
timestamp 1649977179
transform 1 0 44252 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_475
timestamp 1649977179
transform 1 0 44804 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_477
timestamp 1649977179
transform 1 0 44988 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_489
timestamp 1649977179
transform 1 0 46092 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_501
timestamp 1649977179
transform 1 0 47196 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_513
timestamp 1649977179
transform 1 0 48300 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_525
timestamp 1649977179
transform 1 0 49404 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_531
timestamp 1649977179
transform 1 0 49956 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_533
timestamp 1649977179
transform 1 0 50140 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_545
timestamp 1649977179
transform 1 0 51244 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_557
timestamp 1649977179
transform 1 0 52348 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_569
timestamp 1649977179
transform 1 0 53452 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_581
timestamp 1649977179
transform 1 0 54556 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_587
timestamp 1649977179
transform 1 0 55108 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_589
timestamp 1649977179
transform 1 0 55292 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_601
timestamp 1649977179
transform 1 0 56396 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_613
timestamp 1649977179
transform 1 0 57500 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_625
timestamp 1649977179
transform 1 0 58604 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_637
timestamp 1649977179
transform 1 0 59708 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_643
timestamp 1649977179
transform 1 0 60260 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_645
timestamp 1649977179
transform 1 0 60444 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_657
timestamp 1649977179
transform 1 0 61548 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_669
timestamp 1649977179
transform 1 0 62652 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_681
timestamp 1649977179
transform 1 0 63756 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_693
timestamp 1649977179
transform 1 0 64860 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_699
timestamp 1649977179
transform 1 0 65412 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_701
timestamp 1649977179
transform 1 0 65596 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_713
timestamp 1649977179
transform 1 0 66700 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_725
timestamp 1649977179
transform 1 0 67804 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_729
timestamp 1649977179
transform 1 0 68172 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1649977179
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 1649977179
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_27
timestamp 1649977179
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_39
timestamp 1649977179
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1649977179
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1649977179
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1649977179
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_69
timestamp 1649977179
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_81
timestamp 1649977179
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_93
timestamp 1649977179
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1649977179
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1649977179
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_113
timestamp 1649977179
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_125
timestamp 1649977179
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_137
timestamp 1649977179
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_149
timestamp 1649977179
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 1649977179
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1649977179
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_169
timestamp 1649977179
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_181
timestamp 1649977179
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_193
timestamp 1649977179
transform 1 0 18860 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_205
timestamp 1649977179
transform 1 0 19964 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_217
timestamp 1649977179
transform 1 0 21068 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1649977179
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_225
timestamp 1649977179
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_237
timestamp 1649977179
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_249
timestamp 1649977179
transform 1 0 24012 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_261
timestamp 1649977179
transform 1 0 25116 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_273
timestamp 1649977179
transform 1 0 26220 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1649977179
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_281
timestamp 1649977179
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_293
timestamp 1649977179
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_305
timestamp 1649977179
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_317
timestamp 1649977179
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_329
timestamp 1649977179
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1649977179
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_337
timestamp 1649977179
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_349
timestamp 1649977179
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_361
timestamp 1649977179
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_373
timestamp 1649977179
transform 1 0 35420 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_385
timestamp 1649977179
transform 1 0 36524 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 1649977179
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_393
timestamp 1649977179
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_405
timestamp 1649977179
transform 1 0 38364 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_417
timestamp 1649977179
transform 1 0 39468 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_429
timestamp 1649977179
transform 1 0 40572 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_441
timestamp 1649977179
transform 1 0 41676 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_447
timestamp 1649977179
transform 1 0 42228 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_449
timestamp 1649977179
transform 1 0 42412 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_461
timestamp 1649977179
transform 1 0 43516 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_473
timestamp 1649977179
transform 1 0 44620 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_485
timestamp 1649977179
transform 1 0 45724 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_497
timestamp 1649977179
transform 1 0 46828 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_503
timestamp 1649977179
transform 1 0 47380 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_505
timestamp 1649977179
transform 1 0 47564 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_517
timestamp 1649977179
transform 1 0 48668 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_529
timestamp 1649977179
transform 1 0 49772 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_541
timestamp 1649977179
transform 1 0 50876 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_553
timestamp 1649977179
transform 1 0 51980 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_559
timestamp 1649977179
transform 1 0 52532 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_561
timestamp 1649977179
transform 1 0 52716 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_573
timestamp 1649977179
transform 1 0 53820 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_585
timestamp 1649977179
transform 1 0 54924 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_597
timestamp 1649977179
transform 1 0 56028 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_609
timestamp 1649977179
transform 1 0 57132 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_615
timestamp 1649977179
transform 1 0 57684 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_617
timestamp 1649977179
transform 1 0 57868 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_629
timestamp 1649977179
transform 1 0 58972 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_641
timestamp 1649977179
transform 1 0 60076 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_653
timestamp 1649977179
transform 1 0 61180 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_665
timestamp 1649977179
transform 1 0 62284 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_671
timestamp 1649977179
transform 1 0 62836 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_673
timestamp 1649977179
transform 1 0 63020 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_685
timestamp 1649977179
transform 1 0 64124 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_697
timestamp 1649977179
transform 1 0 65228 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_709
timestamp 1649977179
transform 1 0 66332 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_721
timestamp 1649977179
transform 1 0 67436 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_727
timestamp 1649977179
transform 1 0 67988 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_729
timestamp 1649977179
transform 1 0 68172 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1649977179
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1649977179
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1649977179
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1649977179
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1649977179
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_53
timestamp 1649977179
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_65
timestamp 1649977179
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1649977179
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1649977179
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_85
timestamp 1649977179
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_97
timestamp 1649977179
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_109
timestamp 1649977179
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_121
timestamp 1649977179
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1649977179
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1649977179
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_141
timestamp 1649977179
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_153
timestamp 1649977179
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_165
timestamp 1649977179
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_177
timestamp 1649977179
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_189
timestamp 1649977179
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1649977179
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_197
timestamp 1649977179
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_209
timestamp 1649977179
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_221
timestamp 1649977179
transform 1 0 21436 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_233
timestamp 1649977179
transform 1 0 22540 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_245
timestamp 1649977179
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1649977179
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_253
timestamp 1649977179
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_265
timestamp 1649977179
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_277
timestamp 1649977179
transform 1 0 26588 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_289
timestamp 1649977179
transform 1 0 27692 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_301
timestamp 1649977179
transform 1 0 28796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1649977179
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_309
timestamp 1649977179
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_321
timestamp 1649977179
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_333
timestamp 1649977179
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_345
timestamp 1649977179
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_357
timestamp 1649977179
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1649977179
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_365
timestamp 1649977179
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_377
timestamp 1649977179
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_389
timestamp 1649977179
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_401
timestamp 1649977179
transform 1 0 37996 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_413
timestamp 1649977179
transform 1 0 39100 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_419
timestamp 1649977179
transform 1 0 39652 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_421
timestamp 1649977179
transform 1 0 39836 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_433
timestamp 1649977179
transform 1 0 40940 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_445
timestamp 1649977179
transform 1 0 42044 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_457
timestamp 1649977179
transform 1 0 43148 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_469
timestamp 1649977179
transform 1 0 44252 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_475
timestamp 1649977179
transform 1 0 44804 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_477
timestamp 1649977179
transform 1 0 44988 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_489
timestamp 1649977179
transform 1 0 46092 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_501
timestamp 1649977179
transform 1 0 47196 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_513
timestamp 1649977179
transform 1 0 48300 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_525
timestamp 1649977179
transform 1 0 49404 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_531
timestamp 1649977179
transform 1 0 49956 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_533
timestamp 1649977179
transform 1 0 50140 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_545
timestamp 1649977179
transform 1 0 51244 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_557
timestamp 1649977179
transform 1 0 52348 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_569
timestamp 1649977179
transform 1 0 53452 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_581
timestamp 1649977179
transform 1 0 54556 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_587
timestamp 1649977179
transform 1 0 55108 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_589
timestamp 1649977179
transform 1 0 55292 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_601
timestamp 1649977179
transform 1 0 56396 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_613
timestamp 1649977179
transform 1 0 57500 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_625
timestamp 1649977179
transform 1 0 58604 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_637
timestamp 1649977179
transform 1 0 59708 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_643
timestamp 1649977179
transform 1 0 60260 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_645
timestamp 1649977179
transform 1 0 60444 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_657
timestamp 1649977179
transform 1 0 61548 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_669
timestamp 1649977179
transform 1 0 62652 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_681
timestamp 1649977179
transform 1 0 63756 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_693
timestamp 1649977179
transform 1 0 64860 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_699
timestamp 1649977179
transform 1 0 65412 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_701
timestamp 1649977179
transform 1 0 65596 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_713
timestamp 1649977179
transform 1 0 66700 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_725
timestamp 1649977179
transform 1 0 67804 0 1 31552
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_55_3
timestamp 1649977179
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_15
timestamp 1649977179
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_27
timestamp 1649977179
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_39
timestamp 1649977179
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 1649977179
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1649977179
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 1649977179
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_69
timestamp 1649977179
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_81
timestamp 1649977179
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_93
timestamp 1649977179
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1649977179
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1649977179
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_113
timestamp 1649977179
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_125
timestamp 1649977179
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_137
timestamp 1649977179
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_149
timestamp 1649977179
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1649977179
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1649977179
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_169
timestamp 1649977179
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_181
timestamp 1649977179
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_193
timestamp 1649977179
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_205
timestamp 1649977179
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_217
timestamp 1649977179
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1649977179
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_225
timestamp 1649977179
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_237
timestamp 1649977179
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_249
timestamp 1649977179
transform 1 0 24012 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_261
timestamp 1649977179
transform 1 0 25116 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_273
timestamp 1649977179
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1649977179
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_281
timestamp 1649977179
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_293
timestamp 1649977179
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_305
timestamp 1649977179
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_317
timestamp 1649977179
transform 1 0 30268 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_329
timestamp 1649977179
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 1649977179
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_337
timestamp 1649977179
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_349
timestamp 1649977179
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_361
timestamp 1649977179
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_373
timestamp 1649977179
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_385
timestamp 1649977179
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1649977179
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_393
timestamp 1649977179
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_405
timestamp 1649977179
transform 1 0 38364 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_417
timestamp 1649977179
transform 1 0 39468 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_429
timestamp 1649977179
transform 1 0 40572 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_441
timestamp 1649977179
transform 1 0 41676 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_447
timestamp 1649977179
transform 1 0 42228 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_449
timestamp 1649977179
transform 1 0 42412 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_461
timestamp 1649977179
transform 1 0 43516 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_473
timestamp 1649977179
transform 1 0 44620 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_485
timestamp 1649977179
transform 1 0 45724 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_497
timestamp 1649977179
transform 1 0 46828 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_503
timestamp 1649977179
transform 1 0 47380 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_505
timestamp 1649977179
transform 1 0 47564 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_517
timestamp 1649977179
transform 1 0 48668 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_529
timestamp 1649977179
transform 1 0 49772 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_541
timestamp 1649977179
transform 1 0 50876 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_553
timestamp 1649977179
transform 1 0 51980 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_559
timestamp 1649977179
transform 1 0 52532 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_561
timestamp 1649977179
transform 1 0 52716 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_573
timestamp 1649977179
transform 1 0 53820 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_585
timestamp 1649977179
transform 1 0 54924 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_597
timestamp 1649977179
transform 1 0 56028 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_609
timestamp 1649977179
transform 1 0 57132 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_615
timestamp 1649977179
transform 1 0 57684 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_617
timestamp 1649977179
transform 1 0 57868 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_629
timestamp 1649977179
transform 1 0 58972 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_641
timestamp 1649977179
transform 1 0 60076 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_653
timestamp 1649977179
transform 1 0 61180 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_665
timestamp 1649977179
transform 1 0 62284 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_671
timestamp 1649977179
transform 1 0 62836 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_673
timestamp 1649977179
transform 1 0 63020 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_685
timestamp 1649977179
transform 1 0 64124 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_697
timestamp 1649977179
transform 1 0 65228 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_709
timestamp 1649977179
transform 1 0 66332 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_724
timestamp 1649977179
transform 1 0 67712 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_729
timestamp 1649977179
transform 1 0 68172 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1649977179
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1649977179
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1649977179
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1649977179
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1649977179
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_53
timestamp 1649977179
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_65
timestamp 1649977179
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1649977179
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1649977179
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_85
timestamp 1649977179
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_97
timestamp 1649977179
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_109
timestamp 1649977179
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_121
timestamp 1649977179
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1649977179
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1649977179
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_141
timestamp 1649977179
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_153
timestamp 1649977179
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_165
timestamp 1649977179
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_177
timestamp 1649977179
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_189
timestamp 1649977179
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1649977179
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_197
timestamp 1649977179
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_209
timestamp 1649977179
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_221
timestamp 1649977179
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_233
timestamp 1649977179
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_245
timestamp 1649977179
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1649977179
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_253
timestamp 1649977179
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_265
timestamp 1649977179
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_277
timestamp 1649977179
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_289
timestamp 1649977179
transform 1 0 27692 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_301
timestamp 1649977179
transform 1 0 28796 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_307
timestamp 1649977179
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_309
timestamp 1649977179
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_321
timestamp 1649977179
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_333
timestamp 1649977179
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_345
timestamp 1649977179
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_357
timestamp 1649977179
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1649977179
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_365
timestamp 1649977179
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_377
timestamp 1649977179
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_389
timestamp 1649977179
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_401
timestamp 1649977179
transform 1 0 37996 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_413
timestamp 1649977179
transform 1 0 39100 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_419
timestamp 1649977179
transform 1 0 39652 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_421
timestamp 1649977179
transform 1 0 39836 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_433
timestamp 1649977179
transform 1 0 40940 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_445
timestamp 1649977179
transform 1 0 42044 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_457
timestamp 1649977179
transform 1 0 43148 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_469
timestamp 1649977179
transform 1 0 44252 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_475
timestamp 1649977179
transform 1 0 44804 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_477
timestamp 1649977179
transform 1 0 44988 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_489
timestamp 1649977179
transform 1 0 46092 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_501
timestamp 1649977179
transform 1 0 47196 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_513
timestamp 1649977179
transform 1 0 48300 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_525
timestamp 1649977179
transform 1 0 49404 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_531
timestamp 1649977179
transform 1 0 49956 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_533
timestamp 1649977179
transform 1 0 50140 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_545
timestamp 1649977179
transform 1 0 51244 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_557
timestamp 1649977179
transform 1 0 52348 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_569
timestamp 1649977179
transform 1 0 53452 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_581
timestamp 1649977179
transform 1 0 54556 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_587
timestamp 1649977179
transform 1 0 55108 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_589
timestamp 1649977179
transform 1 0 55292 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_601
timestamp 1649977179
transform 1 0 56396 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_613
timestamp 1649977179
transform 1 0 57500 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_625
timestamp 1649977179
transform 1 0 58604 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_637
timestamp 1649977179
transform 1 0 59708 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_643
timestamp 1649977179
transform 1 0 60260 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_645
timestamp 1649977179
transform 1 0 60444 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_657
timestamp 1649977179
transform 1 0 61548 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_669
timestamp 1649977179
transform 1 0 62652 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_681
timestamp 1649977179
transform 1 0 63756 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_693
timestamp 1649977179
transform 1 0 64860 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_699
timestamp 1649977179
transform 1 0 65412 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_701
timestamp 1649977179
transform 1 0 65596 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_713
timestamp 1649977179
transform 1 0 66700 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_725
timestamp 1649977179
transform 1 0 67804 0 1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1649977179
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_15
timestamp 1649977179
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_27
timestamp 1649977179
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_39
timestamp 1649977179
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1649977179
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1649977179
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1649977179
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_69
timestamp 1649977179
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_81
timestamp 1649977179
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_93
timestamp 1649977179
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1649977179
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1649977179
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_113
timestamp 1649977179
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_125
timestamp 1649977179
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_137
timestamp 1649977179
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_149
timestamp 1649977179
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1649977179
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1649977179
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_169
timestamp 1649977179
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_181
timestamp 1649977179
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_193
timestamp 1649977179
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_205
timestamp 1649977179
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_217
timestamp 1649977179
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1649977179
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_225
timestamp 1649977179
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_237
timestamp 1649977179
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_249
timestamp 1649977179
transform 1 0 24012 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_261
timestamp 1649977179
transform 1 0 25116 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_273
timestamp 1649977179
transform 1 0 26220 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1649977179
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_281
timestamp 1649977179
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_293
timestamp 1649977179
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_305
timestamp 1649977179
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_317
timestamp 1649977179
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_329
timestamp 1649977179
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1649977179
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_337
timestamp 1649977179
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_349
timestamp 1649977179
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_361
timestamp 1649977179
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_373
timestamp 1649977179
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_385
timestamp 1649977179
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1649977179
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_393
timestamp 1649977179
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_405
timestamp 1649977179
transform 1 0 38364 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_417
timestamp 1649977179
transform 1 0 39468 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_429
timestamp 1649977179
transform 1 0 40572 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_441
timestamp 1649977179
transform 1 0 41676 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_447
timestamp 1649977179
transform 1 0 42228 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_449
timestamp 1649977179
transform 1 0 42412 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_461
timestamp 1649977179
transform 1 0 43516 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_473
timestamp 1649977179
transform 1 0 44620 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_485
timestamp 1649977179
transform 1 0 45724 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_497
timestamp 1649977179
transform 1 0 46828 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_503
timestamp 1649977179
transform 1 0 47380 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_505
timestamp 1649977179
transform 1 0 47564 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_517
timestamp 1649977179
transform 1 0 48668 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_529
timestamp 1649977179
transform 1 0 49772 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_541
timestamp 1649977179
transform 1 0 50876 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_553
timestamp 1649977179
transform 1 0 51980 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_559
timestamp 1649977179
transform 1 0 52532 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_561
timestamp 1649977179
transform 1 0 52716 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_573
timestamp 1649977179
transform 1 0 53820 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_585
timestamp 1649977179
transform 1 0 54924 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_597
timestamp 1649977179
transform 1 0 56028 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_609
timestamp 1649977179
transform 1 0 57132 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_615
timestamp 1649977179
transform 1 0 57684 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_617
timestamp 1649977179
transform 1 0 57868 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_629
timestamp 1649977179
transform 1 0 58972 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_641
timestamp 1649977179
transform 1 0 60076 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_653
timestamp 1649977179
transform 1 0 61180 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_665
timestamp 1649977179
transform 1 0 62284 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_671
timestamp 1649977179
transform 1 0 62836 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_673
timestamp 1649977179
transform 1 0 63020 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_685
timestamp 1649977179
transform 1 0 64124 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_697
timestamp 1649977179
transform 1 0 65228 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_709
timestamp 1649977179
transform 1 0 66332 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_721
timestamp 1649977179
transform 1 0 67436 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_727
timestamp 1649977179
transform 1 0 67988 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_729
timestamp 1649977179
transform 1 0 68172 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1649977179
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1649977179
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1649977179
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1649977179
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1649977179
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_53
timestamp 1649977179
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_65
timestamp 1649977179
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1649977179
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1649977179
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_85
timestamp 1649977179
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_97
timestamp 1649977179
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_109
timestamp 1649977179
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_121
timestamp 1649977179
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1649977179
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1649977179
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_141
timestamp 1649977179
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_153
timestamp 1649977179
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_165
timestamp 1649977179
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_177
timestamp 1649977179
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1649977179
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1649977179
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_197
timestamp 1649977179
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_209
timestamp 1649977179
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_221
timestamp 1649977179
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_233
timestamp 1649977179
transform 1 0 22540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_245
timestamp 1649977179
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1649977179
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_253
timestamp 1649977179
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_265
timestamp 1649977179
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_277
timestamp 1649977179
transform 1 0 26588 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_289
timestamp 1649977179
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_301
timestamp 1649977179
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1649977179
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_309
timestamp 1649977179
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_321
timestamp 1649977179
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_333
timestamp 1649977179
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_345
timestamp 1649977179
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_357
timestamp 1649977179
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1649977179
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_365
timestamp 1649977179
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_377
timestamp 1649977179
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_389
timestamp 1649977179
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_401
timestamp 1649977179
transform 1 0 37996 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_413
timestamp 1649977179
transform 1 0 39100 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_419
timestamp 1649977179
transform 1 0 39652 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_421
timestamp 1649977179
transform 1 0 39836 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_433
timestamp 1649977179
transform 1 0 40940 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_445
timestamp 1649977179
transform 1 0 42044 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_457
timestamp 1649977179
transform 1 0 43148 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_469
timestamp 1649977179
transform 1 0 44252 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_475
timestamp 1649977179
transform 1 0 44804 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_477
timestamp 1649977179
transform 1 0 44988 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_489
timestamp 1649977179
transform 1 0 46092 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_501
timestamp 1649977179
transform 1 0 47196 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_513
timestamp 1649977179
transform 1 0 48300 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_525
timestamp 1649977179
transform 1 0 49404 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_531
timestamp 1649977179
transform 1 0 49956 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_533
timestamp 1649977179
transform 1 0 50140 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_545
timestamp 1649977179
transform 1 0 51244 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_557
timestamp 1649977179
transform 1 0 52348 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_569
timestamp 1649977179
transform 1 0 53452 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_581
timestamp 1649977179
transform 1 0 54556 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_587
timestamp 1649977179
transform 1 0 55108 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_589
timestamp 1649977179
transform 1 0 55292 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_601
timestamp 1649977179
transform 1 0 56396 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_613
timestamp 1649977179
transform 1 0 57500 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_625
timestamp 1649977179
transform 1 0 58604 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_637
timestamp 1649977179
transform 1 0 59708 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_643
timestamp 1649977179
transform 1 0 60260 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_645
timestamp 1649977179
transform 1 0 60444 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_657
timestamp 1649977179
transform 1 0 61548 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_669
timestamp 1649977179
transform 1 0 62652 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_681
timestamp 1649977179
transform 1 0 63756 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_693
timestamp 1649977179
transform 1 0 64860 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_699
timestamp 1649977179
transform 1 0 65412 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_701
timestamp 1649977179
transform 1 0 65596 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_713
timestamp 1649977179
transform 1 0 66700 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_725
timestamp 1649977179
transform 1 0 67804 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_729
timestamp 1649977179
transform 1 0 68172 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_3
timestamp 1649977179
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_15
timestamp 1649977179
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_27
timestamp 1649977179
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_39
timestamp 1649977179
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1649977179
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1649977179
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1649977179
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_69
timestamp 1649977179
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_81
timestamp 1649977179
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_93
timestamp 1649977179
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1649977179
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1649977179
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_113
timestamp 1649977179
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_125
timestamp 1649977179
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_137
timestamp 1649977179
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_149
timestamp 1649977179
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1649977179
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1649977179
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_169
timestamp 1649977179
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_181
timestamp 1649977179
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_193
timestamp 1649977179
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_205
timestamp 1649977179
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 1649977179
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1649977179
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_225
timestamp 1649977179
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_237
timestamp 1649977179
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_249
timestamp 1649977179
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_261
timestamp 1649977179
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_273
timestamp 1649977179
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1649977179
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_281
timestamp 1649977179
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_293
timestamp 1649977179
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_305
timestamp 1649977179
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_317
timestamp 1649977179
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_329
timestamp 1649977179
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1649977179
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_337
timestamp 1649977179
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_349
timestamp 1649977179
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_361
timestamp 1649977179
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_373
timestamp 1649977179
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_385
timestamp 1649977179
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 1649977179
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_393
timestamp 1649977179
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_405
timestamp 1649977179
transform 1 0 38364 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_417
timestamp 1649977179
transform 1 0 39468 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_429
timestamp 1649977179
transform 1 0 40572 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_441
timestamp 1649977179
transform 1 0 41676 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_447
timestamp 1649977179
transform 1 0 42228 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_449
timestamp 1649977179
transform 1 0 42412 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_461
timestamp 1649977179
transform 1 0 43516 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_473
timestamp 1649977179
transform 1 0 44620 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_485
timestamp 1649977179
transform 1 0 45724 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_497
timestamp 1649977179
transform 1 0 46828 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_503
timestamp 1649977179
transform 1 0 47380 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_505
timestamp 1649977179
transform 1 0 47564 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_517
timestamp 1649977179
transform 1 0 48668 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_529
timestamp 1649977179
transform 1 0 49772 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_541
timestamp 1649977179
transform 1 0 50876 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_553
timestamp 1649977179
transform 1 0 51980 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_559
timestamp 1649977179
transform 1 0 52532 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_561
timestamp 1649977179
transform 1 0 52716 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_573
timestamp 1649977179
transform 1 0 53820 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_585
timestamp 1649977179
transform 1 0 54924 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_597
timestamp 1649977179
transform 1 0 56028 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_609
timestamp 1649977179
transform 1 0 57132 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_615
timestamp 1649977179
transform 1 0 57684 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_617
timestamp 1649977179
transform 1 0 57868 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_629
timestamp 1649977179
transform 1 0 58972 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_641
timestamp 1649977179
transform 1 0 60076 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_653
timestamp 1649977179
transform 1 0 61180 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_665
timestamp 1649977179
transform 1 0 62284 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_671
timestamp 1649977179
transform 1 0 62836 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_673
timestamp 1649977179
transform 1 0 63020 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_685
timestamp 1649977179
transform 1 0 64124 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_697
timestamp 1649977179
transform 1 0 65228 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_709
timestamp 1649977179
transform 1 0 66332 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_721
timestamp 1649977179
transform 1 0 67436 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_727
timestamp 1649977179
transform 1 0 67988 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_729
timestamp 1649977179
transform 1 0 68172 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 1649977179
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_15
timestamp 1649977179
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1649977179
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1649977179
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1649977179
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_53
timestamp 1649977179
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_65
timestamp 1649977179
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1649977179
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1649977179
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_85
timestamp 1649977179
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_97
timestamp 1649977179
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_109
timestamp 1649977179
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_121
timestamp 1649977179
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1649977179
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1649977179
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_141
timestamp 1649977179
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_153
timestamp 1649977179
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_165
timestamp 1649977179
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_177
timestamp 1649977179
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_189
timestamp 1649977179
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1649977179
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_197
timestamp 1649977179
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_209
timestamp 1649977179
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_221
timestamp 1649977179
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_233
timestamp 1649977179
transform 1 0 22540 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_245
timestamp 1649977179
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1649977179
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_253
timestamp 1649977179
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_265
timestamp 1649977179
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_277
timestamp 1649977179
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_289
timestamp 1649977179
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_301
timestamp 1649977179
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1649977179
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_309
timestamp 1649977179
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_321
timestamp 1649977179
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_333
timestamp 1649977179
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_345
timestamp 1649977179
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_357
timestamp 1649977179
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 1649977179
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_365
timestamp 1649977179
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_377
timestamp 1649977179
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_389
timestamp 1649977179
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_401
timestamp 1649977179
transform 1 0 37996 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_413
timestamp 1649977179
transform 1 0 39100 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_419
timestamp 1649977179
transform 1 0 39652 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_421
timestamp 1649977179
transform 1 0 39836 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_433
timestamp 1649977179
transform 1 0 40940 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_445
timestamp 1649977179
transform 1 0 42044 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_457
timestamp 1649977179
transform 1 0 43148 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_469
timestamp 1649977179
transform 1 0 44252 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_475
timestamp 1649977179
transform 1 0 44804 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_477
timestamp 1649977179
transform 1 0 44988 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_489
timestamp 1649977179
transform 1 0 46092 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_501
timestamp 1649977179
transform 1 0 47196 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_513
timestamp 1649977179
transform 1 0 48300 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_525
timestamp 1649977179
transform 1 0 49404 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_531
timestamp 1649977179
transform 1 0 49956 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_533
timestamp 1649977179
transform 1 0 50140 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_545
timestamp 1649977179
transform 1 0 51244 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_557
timestamp 1649977179
transform 1 0 52348 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_569
timestamp 1649977179
transform 1 0 53452 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_581
timestamp 1649977179
transform 1 0 54556 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_587
timestamp 1649977179
transform 1 0 55108 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_589
timestamp 1649977179
transform 1 0 55292 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_601
timestamp 1649977179
transform 1 0 56396 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_613
timestamp 1649977179
transform 1 0 57500 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_625
timestamp 1649977179
transform 1 0 58604 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_637
timestamp 1649977179
transform 1 0 59708 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_643
timestamp 1649977179
transform 1 0 60260 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_645
timestamp 1649977179
transform 1 0 60444 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_657
timestamp 1649977179
transform 1 0 61548 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_669
timestamp 1649977179
transform 1 0 62652 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_681
timestamp 1649977179
transform 1 0 63756 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_693
timestamp 1649977179
transform 1 0 64860 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_699
timestamp 1649977179
transform 1 0 65412 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_701
timestamp 1649977179
transform 1 0 65596 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_713
timestamp 1649977179
transform 1 0 66700 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_725
timestamp 1649977179
transform 1 0 67804 0 1 34816
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_61_3
timestamp 1649977179
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_15
timestamp 1649977179
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_27
timestamp 1649977179
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_39
timestamp 1649977179
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 1649977179
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1649977179
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1649977179
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_69
timestamp 1649977179
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_81
timestamp 1649977179
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_93
timestamp 1649977179
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1649977179
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1649977179
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_113
timestamp 1649977179
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_125
timestamp 1649977179
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_137
timestamp 1649977179
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_149
timestamp 1649977179
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1649977179
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1649977179
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_169
timestamp 1649977179
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_181
timestamp 1649977179
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_193
timestamp 1649977179
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_205
timestamp 1649977179
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_217
timestamp 1649977179
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1649977179
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_225
timestamp 1649977179
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_237
timestamp 1649977179
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_249
timestamp 1649977179
transform 1 0 24012 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_261
timestamp 1649977179
transform 1 0 25116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_273
timestamp 1649977179
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1649977179
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_281
timestamp 1649977179
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_293
timestamp 1649977179
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_305
timestamp 1649977179
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_317
timestamp 1649977179
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_329
timestamp 1649977179
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1649977179
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_337
timestamp 1649977179
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_349
timestamp 1649977179
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_361
timestamp 1649977179
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_373
timestamp 1649977179
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_385
timestamp 1649977179
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_391
timestamp 1649977179
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_393
timestamp 1649977179
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_405
timestamp 1649977179
transform 1 0 38364 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_417
timestamp 1649977179
transform 1 0 39468 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_429
timestamp 1649977179
transform 1 0 40572 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_441
timestamp 1649977179
transform 1 0 41676 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_447
timestamp 1649977179
transform 1 0 42228 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_449
timestamp 1649977179
transform 1 0 42412 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_461
timestamp 1649977179
transform 1 0 43516 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_473
timestamp 1649977179
transform 1 0 44620 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_485
timestamp 1649977179
transform 1 0 45724 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_497
timestamp 1649977179
transform 1 0 46828 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_503
timestamp 1649977179
transform 1 0 47380 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_505
timestamp 1649977179
transform 1 0 47564 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_517
timestamp 1649977179
transform 1 0 48668 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_529
timestamp 1649977179
transform 1 0 49772 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_541
timestamp 1649977179
transform 1 0 50876 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_553
timestamp 1649977179
transform 1 0 51980 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_559
timestamp 1649977179
transform 1 0 52532 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_561
timestamp 1649977179
transform 1 0 52716 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_573
timestamp 1649977179
transform 1 0 53820 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_585
timestamp 1649977179
transform 1 0 54924 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_597
timestamp 1649977179
transform 1 0 56028 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_609
timestamp 1649977179
transform 1 0 57132 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_615
timestamp 1649977179
transform 1 0 57684 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_617
timestamp 1649977179
transform 1 0 57868 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_629
timestamp 1649977179
transform 1 0 58972 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_641
timestamp 1649977179
transform 1 0 60076 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_653
timestamp 1649977179
transform 1 0 61180 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_665
timestamp 1649977179
transform 1 0 62284 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_671
timestamp 1649977179
transform 1 0 62836 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_673
timestamp 1649977179
transform 1 0 63020 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_685
timestamp 1649977179
transform 1 0 64124 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_697
timestamp 1649977179
transform 1 0 65228 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_709
timestamp 1649977179
transform 1 0 66332 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_724
timestamp 1649977179
transform 1 0 67712 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_729
timestamp 1649977179
transform 1 0 68172 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_3
timestamp 1649977179
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_15
timestamp 1649977179
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1649977179
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1649977179
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_41
timestamp 1649977179
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_53
timestamp 1649977179
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_65
timestamp 1649977179
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1649977179
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1649977179
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_85
timestamp 1649977179
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_97
timestamp 1649977179
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_109
timestamp 1649977179
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_121
timestamp 1649977179
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1649977179
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1649977179
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_141
timestamp 1649977179
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_153
timestamp 1649977179
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_165
timestamp 1649977179
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_177
timestamp 1649977179
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1649977179
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1649977179
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_197
timestamp 1649977179
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_209
timestamp 1649977179
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_221
timestamp 1649977179
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_233
timestamp 1649977179
transform 1 0 22540 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_245
timestamp 1649977179
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1649977179
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_253
timestamp 1649977179
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_265
timestamp 1649977179
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_277
timestamp 1649977179
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_289
timestamp 1649977179
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_301
timestamp 1649977179
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 1649977179
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_309
timestamp 1649977179
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_321
timestamp 1649977179
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_333
timestamp 1649977179
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_345
timestamp 1649977179
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 1649977179
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1649977179
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_365
timestamp 1649977179
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_377
timestamp 1649977179
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_389
timestamp 1649977179
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_401
timestamp 1649977179
transform 1 0 37996 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_413
timestamp 1649977179
transform 1 0 39100 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_419
timestamp 1649977179
transform 1 0 39652 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_421
timestamp 1649977179
transform 1 0 39836 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_433
timestamp 1649977179
transform 1 0 40940 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_445
timestamp 1649977179
transform 1 0 42044 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_457
timestamp 1649977179
transform 1 0 43148 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_469
timestamp 1649977179
transform 1 0 44252 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_475
timestamp 1649977179
transform 1 0 44804 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_477
timestamp 1649977179
transform 1 0 44988 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_489
timestamp 1649977179
transform 1 0 46092 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_501
timestamp 1649977179
transform 1 0 47196 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_513
timestamp 1649977179
transform 1 0 48300 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_525
timestamp 1649977179
transform 1 0 49404 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_531
timestamp 1649977179
transform 1 0 49956 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_533
timestamp 1649977179
transform 1 0 50140 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_545
timestamp 1649977179
transform 1 0 51244 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_557
timestamp 1649977179
transform 1 0 52348 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_569
timestamp 1649977179
transform 1 0 53452 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_581
timestamp 1649977179
transform 1 0 54556 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_587
timestamp 1649977179
transform 1 0 55108 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_589
timestamp 1649977179
transform 1 0 55292 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_601
timestamp 1649977179
transform 1 0 56396 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_613
timestamp 1649977179
transform 1 0 57500 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_625
timestamp 1649977179
transform 1 0 58604 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_637
timestamp 1649977179
transform 1 0 59708 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_643
timestamp 1649977179
transform 1 0 60260 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_645
timestamp 1649977179
transform 1 0 60444 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_657
timestamp 1649977179
transform 1 0 61548 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_669
timestamp 1649977179
transform 1 0 62652 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_681
timestamp 1649977179
transform 1 0 63756 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_693
timestamp 1649977179
transform 1 0 64860 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_699
timestamp 1649977179
transform 1 0 65412 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_701
timestamp 1649977179
transform 1 0 65596 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_713
timestamp 1649977179
transform 1 0 66700 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_725
timestamp 1649977179
transform 1 0 67804 0 1 35904
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_63_3
timestamp 1649977179
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_15
timestamp 1649977179
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_27
timestamp 1649977179
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_39
timestamp 1649977179
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_51
timestamp 1649977179
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1649977179
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_57
timestamp 1649977179
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_69
timestamp 1649977179
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_81
timestamp 1649977179
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_93
timestamp 1649977179
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1649977179
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1649977179
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_113
timestamp 1649977179
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_125
timestamp 1649977179
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_137
timestamp 1649977179
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_149
timestamp 1649977179
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1649977179
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1649977179
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_169
timestamp 1649977179
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_181
timestamp 1649977179
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_193
timestamp 1649977179
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_205
timestamp 1649977179
transform 1 0 19964 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_217
timestamp 1649977179
transform 1 0 21068 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1649977179
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_225
timestamp 1649977179
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_237
timestamp 1649977179
transform 1 0 22908 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_249
timestamp 1649977179
transform 1 0 24012 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_261
timestamp 1649977179
transform 1 0 25116 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_273
timestamp 1649977179
transform 1 0 26220 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_279
timestamp 1649977179
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_281
timestamp 1649977179
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_293
timestamp 1649977179
transform 1 0 28060 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_305
timestamp 1649977179
transform 1 0 29164 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_317
timestamp 1649977179
transform 1 0 30268 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_329
timestamp 1649977179
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_335
timestamp 1649977179
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_337
timestamp 1649977179
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_349
timestamp 1649977179
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_361
timestamp 1649977179
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_373
timestamp 1649977179
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_385
timestamp 1649977179
transform 1 0 36524 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_391
timestamp 1649977179
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_393
timestamp 1649977179
transform 1 0 37260 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_405
timestamp 1649977179
transform 1 0 38364 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_417
timestamp 1649977179
transform 1 0 39468 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_429
timestamp 1649977179
transform 1 0 40572 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_441
timestamp 1649977179
transform 1 0 41676 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_447
timestamp 1649977179
transform 1 0 42228 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_449
timestamp 1649977179
transform 1 0 42412 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_461
timestamp 1649977179
transform 1 0 43516 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_473
timestamp 1649977179
transform 1 0 44620 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_485
timestamp 1649977179
transform 1 0 45724 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_497
timestamp 1649977179
transform 1 0 46828 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_503
timestamp 1649977179
transform 1 0 47380 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_505
timestamp 1649977179
transform 1 0 47564 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_517
timestamp 1649977179
transform 1 0 48668 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_529
timestamp 1649977179
transform 1 0 49772 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_541
timestamp 1649977179
transform 1 0 50876 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_553
timestamp 1649977179
transform 1 0 51980 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_559
timestamp 1649977179
transform 1 0 52532 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_561
timestamp 1649977179
transform 1 0 52716 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_573
timestamp 1649977179
transform 1 0 53820 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_585
timestamp 1649977179
transform 1 0 54924 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_597
timestamp 1649977179
transform 1 0 56028 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_609
timestamp 1649977179
transform 1 0 57132 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_615
timestamp 1649977179
transform 1 0 57684 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_617
timestamp 1649977179
transform 1 0 57868 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_629
timestamp 1649977179
transform 1 0 58972 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_641
timestamp 1649977179
transform 1 0 60076 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_653
timestamp 1649977179
transform 1 0 61180 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_665
timestamp 1649977179
transform 1 0 62284 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_671
timestamp 1649977179
transform 1 0 62836 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_673
timestamp 1649977179
transform 1 0 63020 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_685
timestamp 1649977179
transform 1 0 64124 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_697
timestamp 1649977179
transform 1 0 65228 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_709
timestamp 1649977179
transform 1 0 66332 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_724
timestamp 1649977179
transform 1 0 67712 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_729
timestamp 1649977179
transform 1 0 68172 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_3
timestamp 1649977179
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_15
timestamp 1649977179
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1649977179
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_29
timestamp 1649977179
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_41
timestamp 1649977179
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_53
timestamp 1649977179
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_65
timestamp 1649977179
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1649977179
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1649977179
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_85
timestamp 1649977179
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_97
timestamp 1649977179
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_109
timestamp 1649977179
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_121
timestamp 1649977179
transform 1 0 12236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_133
timestamp 1649977179
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1649977179
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_141
timestamp 1649977179
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_153
timestamp 1649977179
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_165
timestamp 1649977179
transform 1 0 16284 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_177
timestamp 1649977179
transform 1 0 17388 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_189
timestamp 1649977179
transform 1 0 18492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 1649977179
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_197
timestamp 1649977179
transform 1 0 19228 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_209
timestamp 1649977179
transform 1 0 20332 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_221
timestamp 1649977179
transform 1 0 21436 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_233
timestamp 1649977179
transform 1 0 22540 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_245
timestamp 1649977179
transform 1 0 23644 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_251
timestamp 1649977179
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_253
timestamp 1649977179
transform 1 0 24380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_265
timestamp 1649977179
transform 1 0 25484 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_277
timestamp 1649977179
transform 1 0 26588 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_289
timestamp 1649977179
transform 1 0 27692 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_301
timestamp 1649977179
transform 1 0 28796 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_307
timestamp 1649977179
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_309
timestamp 1649977179
transform 1 0 29532 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_321
timestamp 1649977179
transform 1 0 30636 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_333
timestamp 1649977179
transform 1 0 31740 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_345
timestamp 1649977179
transform 1 0 32844 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_357
timestamp 1649977179
transform 1 0 33948 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_363
timestamp 1649977179
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_365
timestamp 1649977179
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_377
timestamp 1649977179
transform 1 0 35788 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_389
timestamp 1649977179
transform 1 0 36892 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_401
timestamp 1649977179
transform 1 0 37996 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_413
timestamp 1649977179
transform 1 0 39100 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_419
timestamp 1649977179
transform 1 0 39652 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_421
timestamp 1649977179
transform 1 0 39836 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_433
timestamp 1649977179
transform 1 0 40940 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_445
timestamp 1649977179
transform 1 0 42044 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_457
timestamp 1649977179
transform 1 0 43148 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_469
timestamp 1649977179
transform 1 0 44252 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_475
timestamp 1649977179
transform 1 0 44804 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_477
timestamp 1649977179
transform 1 0 44988 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_489
timestamp 1649977179
transform 1 0 46092 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_501
timestamp 1649977179
transform 1 0 47196 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_513
timestamp 1649977179
transform 1 0 48300 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_525
timestamp 1649977179
transform 1 0 49404 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_531
timestamp 1649977179
transform 1 0 49956 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_533
timestamp 1649977179
transform 1 0 50140 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_545
timestamp 1649977179
transform 1 0 51244 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_557
timestamp 1649977179
transform 1 0 52348 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_569
timestamp 1649977179
transform 1 0 53452 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_581
timestamp 1649977179
transform 1 0 54556 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_587
timestamp 1649977179
transform 1 0 55108 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_589
timestamp 1649977179
transform 1 0 55292 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_601
timestamp 1649977179
transform 1 0 56396 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_613
timestamp 1649977179
transform 1 0 57500 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_625
timestamp 1649977179
transform 1 0 58604 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_637
timestamp 1649977179
transform 1 0 59708 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_643
timestamp 1649977179
transform 1 0 60260 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_645
timestamp 1649977179
transform 1 0 60444 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_657
timestamp 1649977179
transform 1 0 61548 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_669
timestamp 1649977179
transform 1 0 62652 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_681
timestamp 1649977179
transform 1 0 63756 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_693
timestamp 1649977179
transform 1 0 64860 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_699
timestamp 1649977179
transform 1 0 65412 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_701
timestamp 1649977179
transform 1 0 65596 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_713
timestamp 1649977179
transform 1 0 66700 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_725
timestamp 1649977179
transform 1 0 67804 0 1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_65_3
timestamp 1649977179
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_15
timestamp 1649977179
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_27
timestamp 1649977179
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_39
timestamp 1649977179
transform 1 0 4692 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_51
timestamp 1649977179
transform 1 0 5796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1649977179
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_57
timestamp 1649977179
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_69
timestamp 1649977179
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_81
timestamp 1649977179
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_93
timestamp 1649977179
transform 1 0 9660 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_105
timestamp 1649977179
transform 1 0 10764 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_111
timestamp 1649977179
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_113
timestamp 1649977179
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_125
timestamp 1649977179
transform 1 0 12604 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_137
timestamp 1649977179
transform 1 0 13708 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_149
timestamp 1649977179
transform 1 0 14812 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_161
timestamp 1649977179
transform 1 0 15916 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_167
timestamp 1649977179
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_169
timestamp 1649977179
transform 1 0 16652 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_181
timestamp 1649977179
transform 1 0 17756 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_193
timestamp 1649977179
transform 1 0 18860 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_205
timestamp 1649977179
transform 1 0 19964 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_217
timestamp 1649977179
transform 1 0 21068 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_223
timestamp 1649977179
transform 1 0 21620 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_225
timestamp 1649977179
transform 1 0 21804 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_237
timestamp 1649977179
transform 1 0 22908 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_249
timestamp 1649977179
transform 1 0 24012 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_261
timestamp 1649977179
transform 1 0 25116 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_273
timestamp 1649977179
transform 1 0 26220 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_279
timestamp 1649977179
transform 1 0 26772 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_281
timestamp 1649977179
transform 1 0 26956 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_293
timestamp 1649977179
transform 1 0 28060 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_305
timestamp 1649977179
transform 1 0 29164 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_317
timestamp 1649977179
transform 1 0 30268 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_329
timestamp 1649977179
transform 1 0 31372 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_335
timestamp 1649977179
transform 1 0 31924 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_337
timestamp 1649977179
transform 1 0 32108 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_349
timestamp 1649977179
transform 1 0 33212 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_361
timestamp 1649977179
transform 1 0 34316 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_373
timestamp 1649977179
transform 1 0 35420 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_385
timestamp 1649977179
transform 1 0 36524 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_391
timestamp 1649977179
transform 1 0 37076 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_393
timestamp 1649977179
transform 1 0 37260 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_405
timestamp 1649977179
transform 1 0 38364 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_417
timestamp 1649977179
transform 1 0 39468 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_429
timestamp 1649977179
transform 1 0 40572 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_441
timestamp 1649977179
transform 1 0 41676 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_447
timestamp 1649977179
transform 1 0 42228 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_449
timestamp 1649977179
transform 1 0 42412 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_461
timestamp 1649977179
transform 1 0 43516 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_473
timestamp 1649977179
transform 1 0 44620 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_485
timestamp 1649977179
transform 1 0 45724 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_497
timestamp 1649977179
transform 1 0 46828 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_503
timestamp 1649977179
transform 1 0 47380 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_505
timestamp 1649977179
transform 1 0 47564 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_517
timestamp 1649977179
transform 1 0 48668 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_529
timestamp 1649977179
transform 1 0 49772 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_541
timestamp 1649977179
transform 1 0 50876 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_553
timestamp 1649977179
transform 1 0 51980 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_559
timestamp 1649977179
transform 1 0 52532 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_561
timestamp 1649977179
transform 1 0 52716 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_573
timestamp 1649977179
transform 1 0 53820 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_585
timestamp 1649977179
transform 1 0 54924 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_597
timestamp 1649977179
transform 1 0 56028 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_609
timestamp 1649977179
transform 1 0 57132 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_615
timestamp 1649977179
transform 1 0 57684 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_617
timestamp 1649977179
transform 1 0 57868 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_629
timestamp 1649977179
transform 1 0 58972 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_641
timestamp 1649977179
transform 1 0 60076 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_653
timestamp 1649977179
transform 1 0 61180 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_665
timestamp 1649977179
transform 1 0 62284 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_671
timestamp 1649977179
transform 1 0 62836 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_673
timestamp 1649977179
transform 1 0 63020 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_685
timestamp 1649977179
transform 1 0 64124 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_697
timestamp 1649977179
transform 1 0 65228 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_709
timestamp 1649977179
transform 1 0 66332 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_721
timestamp 1649977179
transform 1 0 67436 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_727
timestamp 1649977179
transform 1 0 67988 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_729
timestamp 1649977179
transform 1 0 68172 0 -1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_66_3
timestamp 1649977179
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_15
timestamp 1649977179
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1649977179
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_29
timestamp 1649977179
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_41
timestamp 1649977179
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_53
timestamp 1649977179
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_65
timestamp 1649977179
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_77
timestamp 1649977179
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1649977179
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_85
timestamp 1649977179
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_97
timestamp 1649977179
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_109
timestamp 1649977179
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_121
timestamp 1649977179
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_133
timestamp 1649977179
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 1649977179
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_141
timestamp 1649977179
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_153
timestamp 1649977179
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_165
timestamp 1649977179
transform 1 0 16284 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_177
timestamp 1649977179
transform 1 0 17388 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_189
timestamp 1649977179
transform 1 0 18492 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_195
timestamp 1649977179
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_197
timestamp 1649977179
transform 1 0 19228 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_209
timestamp 1649977179
transform 1 0 20332 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_221
timestamp 1649977179
transform 1 0 21436 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_233
timestamp 1649977179
transform 1 0 22540 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_245
timestamp 1649977179
transform 1 0 23644 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_251
timestamp 1649977179
transform 1 0 24196 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_253
timestamp 1649977179
transform 1 0 24380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_265
timestamp 1649977179
transform 1 0 25484 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_277
timestamp 1649977179
transform 1 0 26588 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_289
timestamp 1649977179
transform 1 0 27692 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_301
timestamp 1649977179
transform 1 0 28796 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_307
timestamp 1649977179
transform 1 0 29348 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_309
timestamp 1649977179
transform 1 0 29532 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_321
timestamp 1649977179
transform 1 0 30636 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_333
timestamp 1649977179
transform 1 0 31740 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_345
timestamp 1649977179
transform 1 0 32844 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_357
timestamp 1649977179
transform 1 0 33948 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_363
timestamp 1649977179
transform 1 0 34500 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_365
timestamp 1649977179
transform 1 0 34684 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_377
timestamp 1649977179
transform 1 0 35788 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_389
timestamp 1649977179
transform 1 0 36892 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_401
timestamp 1649977179
transform 1 0 37996 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_413
timestamp 1649977179
transform 1 0 39100 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_419
timestamp 1649977179
transform 1 0 39652 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_421
timestamp 1649977179
transform 1 0 39836 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_433
timestamp 1649977179
transform 1 0 40940 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_445
timestamp 1649977179
transform 1 0 42044 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_457
timestamp 1649977179
transform 1 0 43148 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_469
timestamp 1649977179
transform 1 0 44252 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_475
timestamp 1649977179
transform 1 0 44804 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_477
timestamp 1649977179
transform 1 0 44988 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_489
timestamp 1649977179
transform 1 0 46092 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_501
timestamp 1649977179
transform 1 0 47196 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_513
timestamp 1649977179
transform 1 0 48300 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_525
timestamp 1649977179
transform 1 0 49404 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_531
timestamp 1649977179
transform 1 0 49956 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_533
timestamp 1649977179
transform 1 0 50140 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_545
timestamp 1649977179
transform 1 0 51244 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_557
timestamp 1649977179
transform 1 0 52348 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_569
timestamp 1649977179
transform 1 0 53452 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_581
timestamp 1649977179
transform 1 0 54556 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_587
timestamp 1649977179
transform 1 0 55108 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_589
timestamp 1649977179
transform 1 0 55292 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_601
timestamp 1649977179
transform 1 0 56396 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_613
timestamp 1649977179
transform 1 0 57500 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_625
timestamp 1649977179
transform 1 0 58604 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_637
timestamp 1649977179
transform 1 0 59708 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_643
timestamp 1649977179
transform 1 0 60260 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_645
timestamp 1649977179
transform 1 0 60444 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_657
timestamp 1649977179
transform 1 0 61548 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_669
timestamp 1649977179
transform 1 0 62652 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_681
timestamp 1649977179
transform 1 0 63756 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_693
timestamp 1649977179
transform 1 0 64860 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_699
timestamp 1649977179
transform 1 0 65412 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_701
timestamp 1649977179
transform 1 0 65596 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_713
timestamp 1649977179
transform 1 0 66700 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_725
timestamp 1649977179
transform 1 0 67804 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_729
timestamp 1649977179
transform 1 0 68172 0 1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_67_3
timestamp 1649977179
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_15
timestamp 1649977179
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_27
timestamp 1649977179
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_39
timestamp 1649977179
transform 1 0 4692 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_51
timestamp 1649977179
transform 1 0 5796 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_55
timestamp 1649977179
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_57
timestamp 1649977179
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_69
timestamp 1649977179
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_81
timestamp 1649977179
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_93
timestamp 1649977179
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_105
timestamp 1649977179
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 1649977179
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_113
timestamp 1649977179
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_125
timestamp 1649977179
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_137
timestamp 1649977179
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_149
timestamp 1649977179
transform 1 0 14812 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_161
timestamp 1649977179
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_167
timestamp 1649977179
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_169
timestamp 1649977179
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_181
timestamp 1649977179
transform 1 0 17756 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_193
timestamp 1649977179
transform 1 0 18860 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_205
timestamp 1649977179
transform 1 0 19964 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_217
timestamp 1649977179
transform 1 0 21068 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_223
timestamp 1649977179
transform 1 0 21620 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_225
timestamp 1649977179
transform 1 0 21804 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_237
timestamp 1649977179
transform 1 0 22908 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_249
timestamp 1649977179
transform 1 0 24012 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_261
timestamp 1649977179
transform 1 0 25116 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_273
timestamp 1649977179
transform 1 0 26220 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_279
timestamp 1649977179
transform 1 0 26772 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_281
timestamp 1649977179
transform 1 0 26956 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_293
timestamp 1649977179
transform 1 0 28060 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_305
timestamp 1649977179
transform 1 0 29164 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_317
timestamp 1649977179
transform 1 0 30268 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_329
timestamp 1649977179
transform 1 0 31372 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_335
timestamp 1649977179
transform 1 0 31924 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_337
timestamp 1649977179
transform 1 0 32108 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_349
timestamp 1649977179
transform 1 0 33212 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_361
timestamp 1649977179
transform 1 0 34316 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_373
timestamp 1649977179
transform 1 0 35420 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_385
timestamp 1649977179
transform 1 0 36524 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_391
timestamp 1649977179
transform 1 0 37076 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_393
timestamp 1649977179
transform 1 0 37260 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_405
timestamp 1649977179
transform 1 0 38364 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_417
timestamp 1649977179
transform 1 0 39468 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_429
timestamp 1649977179
transform 1 0 40572 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_441
timestamp 1649977179
transform 1 0 41676 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_447
timestamp 1649977179
transform 1 0 42228 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_449
timestamp 1649977179
transform 1 0 42412 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_461
timestamp 1649977179
transform 1 0 43516 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_473
timestamp 1649977179
transform 1 0 44620 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_485
timestamp 1649977179
transform 1 0 45724 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_497
timestamp 1649977179
transform 1 0 46828 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_503
timestamp 1649977179
transform 1 0 47380 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_505
timestamp 1649977179
transform 1 0 47564 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_517
timestamp 1649977179
transform 1 0 48668 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_529
timestamp 1649977179
transform 1 0 49772 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_541
timestamp 1649977179
transform 1 0 50876 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_553
timestamp 1649977179
transform 1 0 51980 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_559
timestamp 1649977179
transform 1 0 52532 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_561
timestamp 1649977179
transform 1 0 52716 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_573
timestamp 1649977179
transform 1 0 53820 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_585
timestamp 1649977179
transform 1 0 54924 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_597
timestamp 1649977179
transform 1 0 56028 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_609
timestamp 1649977179
transform 1 0 57132 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_615
timestamp 1649977179
transform 1 0 57684 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_617
timestamp 1649977179
transform 1 0 57868 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_629
timestamp 1649977179
transform 1 0 58972 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_641
timestamp 1649977179
transform 1 0 60076 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_653
timestamp 1649977179
transform 1 0 61180 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_665
timestamp 1649977179
transform 1 0 62284 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_671
timestamp 1649977179
transform 1 0 62836 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_673
timestamp 1649977179
transform 1 0 63020 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_685
timestamp 1649977179
transform 1 0 64124 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_697
timestamp 1649977179
transform 1 0 65228 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_709
timestamp 1649977179
transform 1 0 66332 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_721
timestamp 1649977179
transform 1 0 67436 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_727
timestamp 1649977179
transform 1 0 67988 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_729
timestamp 1649977179
transform 1 0 68172 0 -1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_68_3
timestamp 1649977179
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_15
timestamp 1649977179
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1649977179
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_29
timestamp 1649977179
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_41
timestamp 1649977179
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_53
timestamp 1649977179
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_65
timestamp 1649977179
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_77
timestamp 1649977179
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 1649977179
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_85
timestamp 1649977179
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_97
timestamp 1649977179
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_109
timestamp 1649977179
transform 1 0 11132 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_121
timestamp 1649977179
transform 1 0 12236 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_133
timestamp 1649977179
transform 1 0 13340 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_139
timestamp 1649977179
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_141
timestamp 1649977179
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_153
timestamp 1649977179
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_165
timestamp 1649977179
transform 1 0 16284 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_177
timestamp 1649977179
transform 1 0 17388 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_189
timestamp 1649977179
transform 1 0 18492 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_195
timestamp 1649977179
transform 1 0 19044 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_197
timestamp 1649977179
transform 1 0 19228 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_209
timestamp 1649977179
transform 1 0 20332 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_221
timestamp 1649977179
transform 1 0 21436 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_233
timestamp 1649977179
transform 1 0 22540 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_245
timestamp 1649977179
transform 1 0 23644 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_251
timestamp 1649977179
transform 1 0 24196 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_253
timestamp 1649977179
transform 1 0 24380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_265
timestamp 1649977179
transform 1 0 25484 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_277
timestamp 1649977179
transform 1 0 26588 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_289
timestamp 1649977179
transform 1 0 27692 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_301
timestamp 1649977179
transform 1 0 28796 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_307
timestamp 1649977179
transform 1 0 29348 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_309
timestamp 1649977179
transform 1 0 29532 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_321
timestamp 1649977179
transform 1 0 30636 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_333
timestamp 1649977179
transform 1 0 31740 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_345
timestamp 1649977179
transform 1 0 32844 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_357
timestamp 1649977179
transform 1 0 33948 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_363
timestamp 1649977179
transform 1 0 34500 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_365
timestamp 1649977179
transform 1 0 34684 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_377
timestamp 1649977179
transform 1 0 35788 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_389
timestamp 1649977179
transform 1 0 36892 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_401
timestamp 1649977179
transform 1 0 37996 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_413
timestamp 1649977179
transform 1 0 39100 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_419
timestamp 1649977179
transform 1 0 39652 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_421
timestamp 1649977179
transform 1 0 39836 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_433
timestamp 1649977179
transform 1 0 40940 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_445
timestamp 1649977179
transform 1 0 42044 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_457
timestamp 1649977179
transform 1 0 43148 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_469
timestamp 1649977179
transform 1 0 44252 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_475
timestamp 1649977179
transform 1 0 44804 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_477
timestamp 1649977179
transform 1 0 44988 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_489
timestamp 1649977179
transform 1 0 46092 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_501
timestamp 1649977179
transform 1 0 47196 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_513
timestamp 1649977179
transform 1 0 48300 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_525
timestamp 1649977179
transform 1 0 49404 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_531
timestamp 1649977179
transform 1 0 49956 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_533
timestamp 1649977179
transform 1 0 50140 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_545
timestamp 1649977179
transform 1 0 51244 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_557
timestamp 1649977179
transform 1 0 52348 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_569
timestamp 1649977179
transform 1 0 53452 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_581
timestamp 1649977179
transform 1 0 54556 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_587
timestamp 1649977179
transform 1 0 55108 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_589
timestamp 1649977179
transform 1 0 55292 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_601
timestamp 1649977179
transform 1 0 56396 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_613
timestamp 1649977179
transform 1 0 57500 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_625
timestamp 1649977179
transform 1 0 58604 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_637
timestamp 1649977179
transform 1 0 59708 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_643
timestamp 1649977179
transform 1 0 60260 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_645
timestamp 1649977179
transform 1 0 60444 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_657
timestamp 1649977179
transform 1 0 61548 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_669
timestamp 1649977179
transform 1 0 62652 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_681
timestamp 1649977179
transform 1 0 63756 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_693
timestamp 1649977179
transform 1 0 64860 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_699
timestamp 1649977179
transform 1 0 65412 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_701
timestamp 1649977179
transform 1 0 65596 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_713
timestamp 1649977179
transform 1 0 66700 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_725
timestamp 1649977179
transform 1 0 67804 0 1 39168
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_69_3
timestamp 1649977179
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_15
timestamp 1649977179
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_27
timestamp 1649977179
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_39
timestamp 1649977179
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_51
timestamp 1649977179
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1649977179
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_57
timestamp 1649977179
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_69
timestamp 1649977179
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_81
timestamp 1649977179
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_93
timestamp 1649977179
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_105
timestamp 1649977179
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_111
timestamp 1649977179
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_113
timestamp 1649977179
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_125
timestamp 1649977179
transform 1 0 12604 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_137
timestamp 1649977179
transform 1 0 13708 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_149
timestamp 1649977179
transform 1 0 14812 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_161
timestamp 1649977179
transform 1 0 15916 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_167
timestamp 1649977179
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_169
timestamp 1649977179
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_181
timestamp 1649977179
transform 1 0 17756 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_193
timestamp 1649977179
transform 1 0 18860 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_205
timestamp 1649977179
transform 1 0 19964 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_217
timestamp 1649977179
transform 1 0 21068 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_223
timestamp 1649977179
transform 1 0 21620 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_225
timestamp 1649977179
transform 1 0 21804 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_237
timestamp 1649977179
transform 1 0 22908 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_249
timestamp 1649977179
transform 1 0 24012 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_261
timestamp 1649977179
transform 1 0 25116 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_273
timestamp 1649977179
transform 1 0 26220 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_279
timestamp 1649977179
transform 1 0 26772 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_281
timestamp 1649977179
transform 1 0 26956 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_293
timestamp 1649977179
transform 1 0 28060 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_305
timestamp 1649977179
transform 1 0 29164 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_317
timestamp 1649977179
transform 1 0 30268 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_329
timestamp 1649977179
transform 1 0 31372 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_335
timestamp 1649977179
transform 1 0 31924 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_337
timestamp 1649977179
transform 1 0 32108 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_349
timestamp 1649977179
transform 1 0 33212 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_361
timestamp 1649977179
transform 1 0 34316 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_373
timestamp 1649977179
transform 1 0 35420 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_385
timestamp 1649977179
transform 1 0 36524 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_391
timestamp 1649977179
transform 1 0 37076 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_393
timestamp 1649977179
transform 1 0 37260 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_405
timestamp 1649977179
transform 1 0 38364 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_417
timestamp 1649977179
transform 1 0 39468 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_429
timestamp 1649977179
transform 1 0 40572 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_441
timestamp 1649977179
transform 1 0 41676 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_447
timestamp 1649977179
transform 1 0 42228 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_449
timestamp 1649977179
transform 1 0 42412 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_461
timestamp 1649977179
transform 1 0 43516 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_473
timestamp 1649977179
transform 1 0 44620 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_485
timestamp 1649977179
transform 1 0 45724 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_497
timestamp 1649977179
transform 1 0 46828 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_503
timestamp 1649977179
transform 1 0 47380 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_505
timestamp 1649977179
transform 1 0 47564 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_517
timestamp 1649977179
transform 1 0 48668 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_529
timestamp 1649977179
transform 1 0 49772 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_541
timestamp 1649977179
transform 1 0 50876 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_553
timestamp 1649977179
transform 1 0 51980 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_559
timestamp 1649977179
transform 1 0 52532 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_561
timestamp 1649977179
transform 1 0 52716 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_573
timestamp 1649977179
transform 1 0 53820 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_585
timestamp 1649977179
transform 1 0 54924 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_597
timestamp 1649977179
transform 1 0 56028 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_609
timestamp 1649977179
transform 1 0 57132 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_615
timestamp 1649977179
transform 1 0 57684 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_617
timestamp 1649977179
transform 1 0 57868 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_629
timestamp 1649977179
transform 1 0 58972 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_641
timestamp 1649977179
transform 1 0 60076 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_653
timestamp 1649977179
transform 1 0 61180 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_665
timestamp 1649977179
transform 1 0 62284 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_671
timestamp 1649977179
transform 1 0 62836 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_673
timestamp 1649977179
transform 1 0 63020 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_685
timestamp 1649977179
transform 1 0 64124 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_697
timestamp 1649977179
transform 1 0 65228 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_709
timestamp 1649977179
transform 1 0 66332 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_724
timestamp 1649977179
transform 1 0 67712 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_729
timestamp 1649977179
transform 1 0 68172 0 -1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_70_3
timestamp 1649977179
transform 1 0 1380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_15
timestamp 1649977179
transform 1 0 2484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1649977179
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_29
timestamp 1649977179
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_41
timestamp 1649977179
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_53
timestamp 1649977179
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_65
timestamp 1649977179
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_77
timestamp 1649977179
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1649977179
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_85
timestamp 1649977179
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_97
timestamp 1649977179
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_109
timestamp 1649977179
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_121
timestamp 1649977179
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_133
timestamp 1649977179
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_139
timestamp 1649977179
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_141
timestamp 1649977179
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_153
timestamp 1649977179
transform 1 0 15180 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_165
timestamp 1649977179
transform 1 0 16284 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_177
timestamp 1649977179
transform 1 0 17388 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_189
timestamp 1649977179
transform 1 0 18492 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_195
timestamp 1649977179
transform 1 0 19044 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_197
timestamp 1649977179
transform 1 0 19228 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_209
timestamp 1649977179
transform 1 0 20332 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_221
timestamp 1649977179
transform 1 0 21436 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_233
timestamp 1649977179
transform 1 0 22540 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_245
timestamp 1649977179
transform 1 0 23644 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_251
timestamp 1649977179
transform 1 0 24196 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_253
timestamp 1649977179
transform 1 0 24380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_265
timestamp 1649977179
transform 1 0 25484 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_277
timestamp 1649977179
transform 1 0 26588 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_289
timestamp 1649977179
transform 1 0 27692 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_301
timestamp 1649977179
transform 1 0 28796 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_307
timestamp 1649977179
transform 1 0 29348 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_309
timestamp 1649977179
transform 1 0 29532 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_321
timestamp 1649977179
transform 1 0 30636 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_333
timestamp 1649977179
transform 1 0 31740 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_345
timestamp 1649977179
transform 1 0 32844 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_357
timestamp 1649977179
transform 1 0 33948 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_363
timestamp 1649977179
transform 1 0 34500 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_365
timestamp 1649977179
transform 1 0 34684 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_377
timestamp 1649977179
transform 1 0 35788 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_389
timestamp 1649977179
transform 1 0 36892 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_401
timestamp 1649977179
transform 1 0 37996 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_413
timestamp 1649977179
transform 1 0 39100 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_419
timestamp 1649977179
transform 1 0 39652 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_421
timestamp 1649977179
transform 1 0 39836 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_433
timestamp 1649977179
transform 1 0 40940 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_445
timestamp 1649977179
transform 1 0 42044 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_457
timestamp 1649977179
transform 1 0 43148 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_469
timestamp 1649977179
transform 1 0 44252 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_475
timestamp 1649977179
transform 1 0 44804 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_477
timestamp 1649977179
transform 1 0 44988 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_489
timestamp 1649977179
transform 1 0 46092 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_501
timestamp 1649977179
transform 1 0 47196 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_513
timestamp 1649977179
transform 1 0 48300 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_525
timestamp 1649977179
transform 1 0 49404 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_531
timestamp 1649977179
transform 1 0 49956 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_533
timestamp 1649977179
transform 1 0 50140 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_545
timestamp 1649977179
transform 1 0 51244 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_557
timestamp 1649977179
transform 1 0 52348 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_569
timestamp 1649977179
transform 1 0 53452 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_581
timestamp 1649977179
transform 1 0 54556 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_587
timestamp 1649977179
transform 1 0 55108 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_589
timestamp 1649977179
transform 1 0 55292 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_601
timestamp 1649977179
transform 1 0 56396 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_613
timestamp 1649977179
transform 1 0 57500 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_625
timestamp 1649977179
transform 1 0 58604 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_637
timestamp 1649977179
transform 1 0 59708 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_643
timestamp 1649977179
transform 1 0 60260 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_645
timestamp 1649977179
transform 1 0 60444 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_657
timestamp 1649977179
transform 1 0 61548 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_669
timestamp 1649977179
transform 1 0 62652 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_681
timestamp 1649977179
transform 1 0 63756 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_693
timestamp 1649977179
transform 1 0 64860 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_699
timestamp 1649977179
transform 1 0 65412 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_701
timestamp 1649977179
transform 1 0 65596 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_713
timestamp 1649977179
transform 1 0 66700 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_725
timestamp 1649977179
transform 1 0 67804 0 1 40256
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_71_3
timestamp 1649977179
transform 1 0 1380 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_15
timestamp 1649977179
transform 1 0 2484 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_27
timestamp 1649977179
transform 1 0 3588 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_39
timestamp 1649977179
transform 1 0 4692 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_51
timestamp 1649977179
transform 1 0 5796 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_55
timestamp 1649977179
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_57
timestamp 1649977179
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_69
timestamp 1649977179
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_81
timestamp 1649977179
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_93
timestamp 1649977179
transform 1 0 9660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_105
timestamp 1649977179
transform 1 0 10764 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_111
timestamp 1649977179
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_113
timestamp 1649977179
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_125
timestamp 1649977179
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_137
timestamp 1649977179
transform 1 0 13708 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_149
timestamp 1649977179
transform 1 0 14812 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_161
timestamp 1649977179
transform 1 0 15916 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_167
timestamp 1649977179
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_169
timestamp 1649977179
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_181
timestamp 1649977179
transform 1 0 17756 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_193
timestamp 1649977179
transform 1 0 18860 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_205
timestamp 1649977179
transform 1 0 19964 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_217
timestamp 1649977179
transform 1 0 21068 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_223
timestamp 1649977179
transform 1 0 21620 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_225
timestamp 1649977179
transform 1 0 21804 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_237
timestamp 1649977179
transform 1 0 22908 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_249
timestamp 1649977179
transform 1 0 24012 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_261
timestamp 1649977179
transform 1 0 25116 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_273
timestamp 1649977179
transform 1 0 26220 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_279
timestamp 1649977179
transform 1 0 26772 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_281
timestamp 1649977179
transform 1 0 26956 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_293
timestamp 1649977179
transform 1 0 28060 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_305
timestamp 1649977179
transform 1 0 29164 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_317
timestamp 1649977179
transform 1 0 30268 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_329
timestamp 1649977179
transform 1 0 31372 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_335
timestamp 1649977179
transform 1 0 31924 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_337
timestamp 1649977179
transform 1 0 32108 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_349
timestamp 1649977179
transform 1 0 33212 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_361
timestamp 1649977179
transform 1 0 34316 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_373
timestamp 1649977179
transform 1 0 35420 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_385
timestamp 1649977179
transform 1 0 36524 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_391
timestamp 1649977179
transform 1 0 37076 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_393
timestamp 1649977179
transform 1 0 37260 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_405
timestamp 1649977179
transform 1 0 38364 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_417
timestamp 1649977179
transform 1 0 39468 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_429
timestamp 1649977179
transform 1 0 40572 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_441
timestamp 1649977179
transform 1 0 41676 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_447
timestamp 1649977179
transform 1 0 42228 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_449
timestamp 1649977179
transform 1 0 42412 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_461
timestamp 1649977179
transform 1 0 43516 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_473
timestamp 1649977179
transform 1 0 44620 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_485
timestamp 1649977179
transform 1 0 45724 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_497
timestamp 1649977179
transform 1 0 46828 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_503
timestamp 1649977179
transform 1 0 47380 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_505
timestamp 1649977179
transform 1 0 47564 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_517
timestamp 1649977179
transform 1 0 48668 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_529
timestamp 1649977179
transform 1 0 49772 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_541
timestamp 1649977179
transform 1 0 50876 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_553
timestamp 1649977179
transform 1 0 51980 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_559
timestamp 1649977179
transform 1 0 52532 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_561
timestamp 1649977179
transform 1 0 52716 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_573
timestamp 1649977179
transform 1 0 53820 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_585
timestamp 1649977179
transform 1 0 54924 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_597
timestamp 1649977179
transform 1 0 56028 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_609
timestamp 1649977179
transform 1 0 57132 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_615
timestamp 1649977179
transform 1 0 57684 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_617
timestamp 1649977179
transform 1 0 57868 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_629
timestamp 1649977179
transform 1 0 58972 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_641
timestamp 1649977179
transform 1 0 60076 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_653
timestamp 1649977179
transform 1 0 61180 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_665
timestamp 1649977179
transform 1 0 62284 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_671
timestamp 1649977179
transform 1 0 62836 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_673
timestamp 1649977179
transform 1 0 63020 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_685
timestamp 1649977179
transform 1 0 64124 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_697
timestamp 1649977179
transform 1 0 65228 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_709
timestamp 1649977179
transform 1 0 66332 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_721
timestamp 1649977179
transform 1 0 67436 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_727
timestamp 1649977179
transform 1 0 67988 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_729
timestamp 1649977179
transform 1 0 68172 0 -1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_72_3
timestamp 1649977179
transform 1 0 1380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_15
timestamp 1649977179
transform 1 0 2484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_27
timestamp 1649977179
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_29
timestamp 1649977179
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_41
timestamp 1649977179
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_53
timestamp 1649977179
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_65
timestamp 1649977179
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_77
timestamp 1649977179
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1649977179
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_85
timestamp 1649977179
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_97
timestamp 1649977179
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_109
timestamp 1649977179
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_121
timestamp 1649977179
transform 1 0 12236 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_133
timestamp 1649977179
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 1649977179
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_141
timestamp 1649977179
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_153
timestamp 1649977179
transform 1 0 15180 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_165
timestamp 1649977179
transform 1 0 16284 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_177
timestamp 1649977179
transform 1 0 17388 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_189
timestamp 1649977179
transform 1 0 18492 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_195
timestamp 1649977179
transform 1 0 19044 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_197
timestamp 1649977179
transform 1 0 19228 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_209
timestamp 1649977179
transform 1 0 20332 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_221
timestamp 1649977179
transform 1 0 21436 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_233
timestamp 1649977179
transform 1 0 22540 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_245
timestamp 1649977179
transform 1 0 23644 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_251
timestamp 1649977179
transform 1 0 24196 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_253
timestamp 1649977179
transform 1 0 24380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_265
timestamp 1649977179
transform 1 0 25484 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_277
timestamp 1649977179
transform 1 0 26588 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_289
timestamp 1649977179
transform 1 0 27692 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_301
timestamp 1649977179
transform 1 0 28796 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_307
timestamp 1649977179
transform 1 0 29348 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_309
timestamp 1649977179
transform 1 0 29532 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_321
timestamp 1649977179
transform 1 0 30636 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_333
timestamp 1649977179
transform 1 0 31740 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_345
timestamp 1649977179
transform 1 0 32844 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_357
timestamp 1649977179
transform 1 0 33948 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_363
timestamp 1649977179
transform 1 0 34500 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_365
timestamp 1649977179
transform 1 0 34684 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_377
timestamp 1649977179
transform 1 0 35788 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_389
timestamp 1649977179
transform 1 0 36892 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_401
timestamp 1649977179
transform 1 0 37996 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_413
timestamp 1649977179
transform 1 0 39100 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_419
timestamp 1649977179
transform 1 0 39652 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_421
timestamp 1649977179
transform 1 0 39836 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_433
timestamp 1649977179
transform 1 0 40940 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_445
timestamp 1649977179
transform 1 0 42044 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_457
timestamp 1649977179
transform 1 0 43148 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_469
timestamp 1649977179
transform 1 0 44252 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_475
timestamp 1649977179
transform 1 0 44804 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_477
timestamp 1649977179
transform 1 0 44988 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_489
timestamp 1649977179
transform 1 0 46092 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_501
timestamp 1649977179
transform 1 0 47196 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_513
timestamp 1649977179
transform 1 0 48300 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_525
timestamp 1649977179
transform 1 0 49404 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_531
timestamp 1649977179
transform 1 0 49956 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_533
timestamp 1649977179
transform 1 0 50140 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_545
timestamp 1649977179
transform 1 0 51244 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_557
timestamp 1649977179
transform 1 0 52348 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_569
timestamp 1649977179
transform 1 0 53452 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_581
timestamp 1649977179
transform 1 0 54556 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_587
timestamp 1649977179
transform 1 0 55108 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_589
timestamp 1649977179
transform 1 0 55292 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_601
timestamp 1649977179
transform 1 0 56396 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_613
timestamp 1649977179
transform 1 0 57500 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_625
timestamp 1649977179
transform 1 0 58604 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_637
timestamp 1649977179
transform 1 0 59708 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_643
timestamp 1649977179
transform 1 0 60260 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_645
timestamp 1649977179
transform 1 0 60444 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_657
timestamp 1649977179
transform 1 0 61548 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_669
timestamp 1649977179
transform 1 0 62652 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_681
timestamp 1649977179
transform 1 0 63756 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_693
timestamp 1649977179
transform 1 0 64860 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_699
timestamp 1649977179
transform 1 0 65412 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_701
timestamp 1649977179
transform 1 0 65596 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_713
timestamp 1649977179
transform 1 0 66700 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_725
timestamp 1649977179
transform 1 0 67804 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_729
timestamp 1649977179
transform 1 0 68172 0 1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_73_3
timestamp 1649977179
transform 1 0 1380 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_15
timestamp 1649977179
transform 1 0 2484 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_27
timestamp 1649977179
transform 1 0 3588 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_39
timestamp 1649977179
transform 1 0 4692 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_51
timestamp 1649977179
transform 1 0 5796 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 1649977179
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_57
timestamp 1649977179
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_69
timestamp 1649977179
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_81
timestamp 1649977179
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_93
timestamp 1649977179
transform 1 0 9660 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_105
timestamp 1649977179
transform 1 0 10764 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_111
timestamp 1649977179
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_113
timestamp 1649977179
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_125
timestamp 1649977179
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_137
timestamp 1649977179
transform 1 0 13708 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_149
timestamp 1649977179
transform 1 0 14812 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_161
timestamp 1649977179
transform 1 0 15916 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_167
timestamp 1649977179
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_169
timestamp 1649977179
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_181
timestamp 1649977179
transform 1 0 17756 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_193
timestamp 1649977179
transform 1 0 18860 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_205
timestamp 1649977179
transform 1 0 19964 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_217
timestamp 1649977179
transform 1 0 21068 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_223
timestamp 1649977179
transform 1 0 21620 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_225
timestamp 1649977179
transform 1 0 21804 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_237
timestamp 1649977179
transform 1 0 22908 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_249
timestamp 1649977179
transform 1 0 24012 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_261
timestamp 1649977179
transform 1 0 25116 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_273
timestamp 1649977179
transform 1 0 26220 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_279
timestamp 1649977179
transform 1 0 26772 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_281
timestamp 1649977179
transform 1 0 26956 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_293
timestamp 1649977179
transform 1 0 28060 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_305
timestamp 1649977179
transform 1 0 29164 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_317
timestamp 1649977179
transform 1 0 30268 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_329
timestamp 1649977179
transform 1 0 31372 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_335
timestamp 1649977179
transform 1 0 31924 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_337
timestamp 1649977179
transform 1 0 32108 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_349
timestamp 1649977179
transform 1 0 33212 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_361
timestamp 1649977179
transform 1 0 34316 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_373
timestamp 1649977179
transform 1 0 35420 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_385
timestamp 1649977179
transform 1 0 36524 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_391
timestamp 1649977179
transform 1 0 37076 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_393
timestamp 1649977179
transform 1 0 37260 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_405
timestamp 1649977179
transform 1 0 38364 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_417
timestamp 1649977179
transform 1 0 39468 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_429
timestamp 1649977179
transform 1 0 40572 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_441
timestamp 1649977179
transform 1 0 41676 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_447
timestamp 1649977179
transform 1 0 42228 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_449
timestamp 1649977179
transform 1 0 42412 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_461
timestamp 1649977179
transform 1 0 43516 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_473
timestamp 1649977179
transform 1 0 44620 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_485
timestamp 1649977179
transform 1 0 45724 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_497
timestamp 1649977179
transform 1 0 46828 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_503
timestamp 1649977179
transform 1 0 47380 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_505
timestamp 1649977179
transform 1 0 47564 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_517
timestamp 1649977179
transform 1 0 48668 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_529
timestamp 1649977179
transform 1 0 49772 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_541
timestamp 1649977179
transform 1 0 50876 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_553
timestamp 1649977179
transform 1 0 51980 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_559
timestamp 1649977179
transform 1 0 52532 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_561
timestamp 1649977179
transform 1 0 52716 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_573
timestamp 1649977179
transform 1 0 53820 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_585
timestamp 1649977179
transform 1 0 54924 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_597
timestamp 1649977179
transform 1 0 56028 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_609
timestamp 1649977179
transform 1 0 57132 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_615
timestamp 1649977179
transform 1 0 57684 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_617
timestamp 1649977179
transform 1 0 57868 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_629
timestamp 1649977179
transform 1 0 58972 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_641
timestamp 1649977179
transform 1 0 60076 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_653
timestamp 1649977179
transform 1 0 61180 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_665
timestamp 1649977179
transform 1 0 62284 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_671
timestamp 1649977179
transform 1 0 62836 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_673
timestamp 1649977179
transform 1 0 63020 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_685
timestamp 1649977179
transform 1 0 64124 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_697
timestamp 1649977179
transform 1 0 65228 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_709
timestamp 1649977179
transform 1 0 66332 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_721
timestamp 1649977179
transform 1 0 67436 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_727
timestamp 1649977179
transform 1 0 67988 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_729
timestamp 1649977179
transform 1 0 68172 0 -1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_74_3
timestamp 1649977179
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_15
timestamp 1649977179
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1649977179
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_29
timestamp 1649977179
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_41
timestamp 1649977179
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_53
timestamp 1649977179
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_65
timestamp 1649977179
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_77
timestamp 1649977179
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 1649977179
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_85
timestamp 1649977179
transform 1 0 8924 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_97
timestamp 1649977179
transform 1 0 10028 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_109
timestamp 1649977179
transform 1 0 11132 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_121
timestamp 1649977179
transform 1 0 12236 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_133
timestamp 1649977179
transform 1 0 13340 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_139
timestamp 1649977179
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_141
timestamp 1649977179
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_153
timestamp 1649977179
transform 1 0 15180 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_165
timestamp 1649977179
transform 1 0 16284 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_177
timestamp 1649977179
transform 1 0 17388 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_189
timestamp 1649977179
transform 1 0 18492 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_195
timestamp 1649977179
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_197
timestamp 1649977179
transform 1 0 19228 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_209
timestamp 1649977179
transform 1 0 20332 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_221
timestamp 1649977179
transform 1 0 21436 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_233
timestamp 1649977179
transform 1 0 22540 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_245
timestamp 1649977179
transform 1 0 23644 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_251
timestamp 1649977179
transform 1 0 24196 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_253
timestamp 1649977179
transform 1 0 24380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_265
timestamp 1649977179
transform 1 0 25484 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_277
timestamp 1649977179
transform 1 0 26588 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_289
timestamp 1649977179
transform 1 0 27692 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_301
timestamp 1649977179
transform 1 0 28796 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_307
timestamp 1649977179
transform 1 0 29348 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_309
timestamp 1649977179
transform 1 0 29532 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_321
timestamp 1649977179
transform 1 0 30636 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_333
timestamp 1649977179
transform 1 0 31740 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_345
timestamp 1649977179
transform 1 0 32844 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_357
timestamp 1649977179
transform 1 0 33948 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_363
timestamp 1649977179
transform 1 0 34500 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_365
timestamp 1649977179
transform 1 0 34684 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_377
timestamp 1649977179
transform 1 0 35788 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_389
timestamp 1649977179
transform 1 0 36892 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_401
timestamp 1649977179
transform 1 0 37996 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_413
timestamp 1649977179
transform 1 0 39100 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_419
timestamp 1649977179
transform 1 0 39652 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_421
timestamp 1649977179
transform 1 0 39836 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_433
timestamp 1649977179
transform 1 0 40940 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_445
timestamp 1649977179
transform 1 0 42044 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_457
timestamp 1649977179
transform 1 0 43148 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_469
timestamp 1649977179
transform 1 0 44252 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_475
timestamp 1649977179
transform 1 0 44804 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_477
timestamp 1649977179
transform 1 0 44988 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_489
timestamp 1649977179
transform 1 0 46092 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_501
timestamp 1649977179
transform 1 0 47196 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_513
timestamp 1649977179
transform 1 0 48300 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_525
timestamp 1649977179
transform 1 0 49404 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_531
timestamp 1649977179
transform 1 0 49956 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_533
timestamp 1649977179
transform 1 0 50140 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_545
timestamp 1649977179
transform 1 0 51244 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_557
timestamp 1649977179
transform 1 0 52348 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_569
timestamp 1649977179
transform 1 0 53452 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_581
timestamp 1649977179
transform 1 0 54556 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_587
timestamp 1649977179
transform 1 0 55108 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_589
timestamp 1649977179
transform 1 0 55292 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_601
timestamp 1649977179
transform 1 0 56396 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_613
timestamp 1649977179
transform 1 0 57500 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_625
timestamp 1649977179
transform 1 0 58604 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_637
timestamp 1649977179
transform 1 0 59708 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_643
timestamp 1649977179
transform 1 0 60260 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_645
timestamp 1649977179
transform 1 0 60444 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_657
timestamp 1649977179
transform 1 0 61548 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_669
timestamp 1649977179
transform 1 0 62652 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_681
timestamp 1649977179
transform 1 0 63756 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_693
timestamp 1649977179
transform 1 0 64860 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_699
timestamp 1649977179
transform 1 0 65412 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_701
timestamp 1649977179
transform 1 0 65596 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_713
timestamp 1649977179
transform 1 0 66700 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_725
timestamp 1649977179
transform 1 0 67804 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_729
timestamp 1649977179
transform 1 0 68172 0 1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_75_3
timestamp 1649977179
transform 1 0 1380 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_15
timestamp 1649977179
transform 1 0 2484 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_27
timestamp 1649977179
transform 1 0 3588 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_39
timestamp 1649977179
transform 1 0 4692 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_51
timestamp 1649977179
transform 1 0 5796 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_55
timestamp 1649977179
transform 1 0 6164 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_57
timestamp 1649977179
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_69
timestamp 1649977179
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_81
timestamp 1649977179
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_93
timestamp 1649977179
transform 1 0 9660 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_105
timestamp 1649977179
transform 1 0 10764 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_111
timestamp 1649977179
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_113
timestamp 1649977179
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_125
timestamp 1649977179
transform 1 0 12604 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_137
timestamp 1649977179
transform 1 0 13708 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_149
timestamp 1649977179
transform 1 0 14812 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_161
timestamp 1649977179
transform 1 0 15916 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_167
timestamp 1649977179
transform 1 0 16468 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_169
timestamp 1649977179
transform 1 0 16652 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_181
timestamp 1649977179
transform 1 0 17756 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_193
timestamp 1649977179
transform 1 0 18860 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_205
timestamp 1649977179
transform 1 0 19964 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_217
timestamp 1649977179
transform 1 0 21068 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_223
timestamp 1649977179
transform 1 0 21620 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_225
timestamp 1649977179
transform 1 0 21804 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_237
timestamp 1649977179
transform 1 0 22908 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_249
timestamp 1649977179
transform 1 0 24012 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_261
timestamp 1649977179
transform 1 0 25116 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_273
timestamp 1649977179
transform 1 0 26220 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_279
timestamp 1649977179
transform 1 0 26772 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_281
timestamp 1649977179
transform 1 0 26956 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_293
timestamp 1649977179
transform 1 0 28060 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_305
timestamp 1649977179
transform 1 0 29164 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_317
timestamp 1649977179
transform 1 0 30268 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_329
timestamp 1649977179
transform 1 0 31372 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_335
timestamp 1649977179
transform 1 0 31924 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_337
timestamp 1649977179
transform 1 0 32108 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_349
timestamp 1649977179
transform 1 0 33212 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_361
timestamp 1649977179
transform 1 0 34316 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_373
timestamp 1649977179
transform 1 0 35420 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_385
timestamp 1649977179
transform 1 0 36524 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_391
timestamp 1649977179
transform 1 0 37076 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_393
timestamp 1649977179
transform 1 0 37260 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_405
timestamp 1649977179
transform 1 0 38364 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_417
timestamp 1649977179
transform 1 0 39468 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_429
timestamp 1649977179
transform 1 0 40572 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_441
timestamp 1649977179
transform 1 0 41676 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_447
timestamp 1649977179
transform 1 0 42228 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_449
timestamp 1649977179
transform 1 0 42412 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_461
timestamp 1649977179
transform 1 0 43516 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_473
timestamp 1649977179
transform 1 0 44620 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_485
timestamp 1649977179
transform 1 0 45724 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_497
timestamp 1649977179
transform 1 0 46828 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_503
timestamp 1649977179
transform 1 0 47380 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_505
timestamp 1649977179
transform 1 0 47564 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_517
timestamp 1649977179
transform 1 0 48668 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_529
timestamp 1649977179
transform 1 0 49772 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_541
timestamp 1649977179
transform 1 0 50876 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_553
timestamp 1649977179
transform 1 0 51980 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_559
timestamp 1649977179
transform 1 0 52532 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_561
timestamp 1649977179
transform 1 0 52716 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_573
timestamp 1649977179
transform 1 0 53820 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_585
timestamp 1649977179
transform 1 0 54924 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_597
timestamp 1649977179
transform 1 0 56028 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_609
timestamp 1649977179
transform 1 0 57132 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_615
timestamp 1649977179
transform 1 0 57684 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_617
timestamp 1649977179
transform 1 0 57868 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_629
timestamp 1649977179
transform 1 0 58972 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_641
timestamp 1649977179
transform 1 0 60076 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_653
timestamp 1649977179
transform 1 0 61180 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_665
timestamp 1649977179
transform 1 0 62284 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_671
timestamp 1649977179
transform 1 0 62836 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_673
timestamp 1649977179
transform 1 0 63020 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_685
timestamp 1649977179
transform 1 0 64124 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_697
timestamp 1649977179
transform 1 0 65228 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_709
timestamp 1649977179
transform 1 0 66332 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_721
timestamp 1649977179
transform 1 0 67436 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_727
timestamp 1649977179
transform 1 0 67988 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_729
timestamp 1649977179
transform 1 0 68172 0 -1 43520
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_76_3
timestamp 1649977179
transform 1 0 1380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_15
timestamp 1649977179
transform 1 0 2484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 1649977179
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_29
timestamp 1649977179
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_41
timestamp 1649977179
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_53
timestamp 1649977179
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_65
timestamp 1649977179
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_77
timestamp 1649977179
transform 1 0 8188 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_83
timestamp 1649977179
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_85
timestamp 1649977179
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_97
timestamp 1649977179
transform 1 0 10028 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_109
timestamp 1649977179
transform 1 0 11132 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_121
timestamp 1649977179
transform 1 0 12236 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_133
timestamp 1649977179
transform 1 0 13340 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_139
timestamp 1649977179
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_141
timestamp 1649977179
transform 1 0 14076 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_153
timestamp 1649977179
transform 1 0 15180 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_165
timestamp 1649977179
transform 1 0 16284 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_177
timestamp 1649977179
transform 1 0 17388 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_189
timestamp 1649977179
transform 1 0 18492 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_195
timestamp 1649977179
transform 1 0 19044 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_197
timestamp 1649977179
transform 1 0 19228 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_209
timestamp 1649977179
transform 1 0 20332 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_221
timestamp 1649977179
transform 1 0 21436 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_233
timestamp 1649977179
transform 1 0 22540 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_245
timestamp 1649977179
transform 1 0 23644 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_251
timestamp 1649977179
transform 1 0 24196 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_253
timestamp 1649977179
transform 1 0 24380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_265
timestamp 1649977179
transform 1 0 25484 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_277
timestamp 1649977179
transform 1 0 26588 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_289
timestamp 1649977179
transform 1 0 27692 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_301
timestamp 1649977179
transform 1 0 28796 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_307
timestamp 1649977179
transform 1 0 29348 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_309
timestamp 1649977179
transform 1 0 29532 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_321
timestamp 1649977179
transform 1 0 30636 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_333
timestamp 1649977179
transform 1 0 31740 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_345
timestamp 1649977179
transform 1 0 32844 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_357
timestamp 1649977179
transform 1 0 33948 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_363
timestamp 1649977179
transform 1 0 34500 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_365
timestamp 1649977179
transform 1 0 34684 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_377
timestamp 1649977179
transform 1 0 35788 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_389
timestamp 1649977179
transform 1 0 36892 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_401
timestamp 1649977179
transform 1 0 37996 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_413
timestamp 1649977179
transform 1 0 39100 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_419
timestamp 1649977179
transform 1 0 39652 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_421
timestamp 1649977179
transform 1 0 39836 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_433
timestamp 1649977179
transform 1 0 40940 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_445
timestamp 1649977179
transform 1 0 42044 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_457
timestamp 1649977179
transform 1 0 43148 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_469
timestamp 1649977179
transform 1 0 44252 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_475
timestamp 1649977179
transform 1 0 44804 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_477
timestamp 1649977179
transform 1 0 44988 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_489
timestamp 1649977179
transform 1 0 46092 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_501
timestamp 1649977179
transform 1 0 47196 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_513
timestamp 1649977179
transform 1 0 48300 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_525
timestamp 1649977179
transform 1 0 49404 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_531
timestamp 1649977179
transform 1 0 49956 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_533
timestamp 1649977179
transform 1 0 50140 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_545
timestamp 1649977179
transform 1 0 51244 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_557
timestamp 1649977179
transform 1 0 52348 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_569
timestamp 1649977179
transform 1 0 53452 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_581
timestamp 1649977179
transform 1 0 54556 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_587
timestamp 1649977179
transform 1 0 55108 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_589
timestamp 1649977179
transform 1 0 55292 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_601
timestamp 1649977179
transform 1 0 56396 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_613
timestamp 1649977179
transform 1 0 57500 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_625
timestamp 1649977179
transform 1 0 58604 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_637
timestamp 1649977179
transform 1 0 59708 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_643
timestamp 1649977179
transform 1 0 60260 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_645
timestamp 1649977179
transform 1 0 60444 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_657
timestamp 1649977179
transform 1 0 61548 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_669
timestamp 1649977179
transform 1 0 62652 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_681
timestamp 1649977179
transform 1 0 63756 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_693
timestamp 1649977179
transform 1 0 64860 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_699
timestamp 1649977179
transform 1 0 65412 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_701
timestamp 1649977179
transform 1 0 65596 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_713
timestamp 1649977179
transform 1 0 66700 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_725
timestamp 1649977179
transform 1 0 67804 0 1 43520
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_77_3
timestamp 1649977179
transform 1 0 1380 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_15
timestamp 1649977179
transform 1 0 2484 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_27
timestamp 1649977179
transform 1 0 3588 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_39
timestamp 1649977179
transform 1 0 4692 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_51
timestamp 1649977179
transform 1 0 5796 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_55
timestamp 1649977179
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_57
timestamp 1649977179
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_69
timestamp 1649977179
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_81
timestamp 1649977179
transform 1 0 8556 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_93
timestamp 1649977179
transform 1 0 9660 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_105
timestamp 1649977179
transform 1 0 10764 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_111
timestamp 1649977179
transform 1 0 11316 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_113
timestamp 1649977179
transform 1 0 11500 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_125
timestamp 1649977179
transform 1 0 12604 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_137
timestamp 1649977179
transform 1 0 13708 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_149
timestamp 1649977179
transform 1 0 14812 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_161
timestamp 1649977179
transform 1 0 15916 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_167
timestamp 1649977179
transform 1 0 16468 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_169
timestamp 1649977179
transform 1 0 16652 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_181
timestamp 1649977179
transform 1 0 17756 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_193
timestamp 1649977179
transform 1 0 18860 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_205
timestamp 1649977179
transform 1 0 19964 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_217
timestamp 1649977179
transform 1 0 21068 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_223
timestamp 1649977179
transform 1 0 21620 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_225
timestamp 1649977179
transform 1 0 21804 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_237
timestamp 1649977179
transform 1 0 22908 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_249
timestamp 1649977179
transform 1 0 24012 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_261
timestamp 1649977179
transform 1 0 25116 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_273
timestamp 1649977179
transform 1 0 26220 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_279
timestamp 1649977179
transform 1 0 26772 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_281
timestamp 1649977179
transform 1 0 26956 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_293
timestamp 1649977179
transform 1 0 28060 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_305
timestamp 1649977179
transform 1 0 29164 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_317
timestamp 1649977179
transform 1 0 30268 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_329
timestamp 1649977179
transform 1 0 31372 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_335
timestamp 1649977179
transform 1 0 31924 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_337
timestamp 1649977179
transform 1 0 32108 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_349
timestamp 1649977179
transform 1 0 33212 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_361
timestamp 1649977179
transform 1 0 34316 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_373
timestamp 1649977179
transform 1 0 35420 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_385
timestamp 1649977179
transform 1 0 36524 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_391
timestamp 1649977179
transform 1 0 37076 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_393
timestamp 1649977179
transform 1 0 37260 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_405
timestamp 1649977179
transform 1 0 38364 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_417
timestamp 1649977179
transform 1 0 39468 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_429
timestamp 1649977179
transform 1 0 40572 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_441
timestamp 1649977179
transform 1 0 41676 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_447
timestamp 1649977179
transform 1 0 42228 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_449
timestamp 1649977179
transform 1 0 42412 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_461
timestamp 1649977179
transform 1 0 43516 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_473
timestamp 1649977179
transform 1 0 44620 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_485
timestamp 1649977179
transform 1 0 45724 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_497
timestamp 1649977179
transform 1 0 46828 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_503
timestamp 1649977179
transform 1 0 47380 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_505
timestamp 1649977179
transform 1 0 47564 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_517
timestamp 1649977179
transform 1 0 48668 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_529
timestamp 1649977179
transform 1 0 49772 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_541
timestamp 1649977179
transform 1 0 50876 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_553
timestamp 1649977179
transform 1 0 51980 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_559
timestamp 1649977179
transform 1 0 52532 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_561
timestamp 1649977179
transform 1 0 52716 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_573
timestamp 1649977179
transform 1 0 53820 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_585
timestamp 1649977179
transform 1 0 54924 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_597
timestamp 1649977179
transform 1 0 56028 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_609
timestamp 1649977179
transform 1 0 57132 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_615
timestamp 1649977179
transform 1 0 57684 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_617
timestamp 1649977179
transform 1 0 57868 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_629
timestamp 1649977179
transform 1 0 58972 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_641
timestamp 1649977179
transform 1 0 60076 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_653
timestamp 1649977179
transform 1 0 61180 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_665
timestamp 1649977179
transform 1 0 62284 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_671
timestamp 1649977179
transform 1 0 62836 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_673
timestamp 1649977179
transform 1 0 63020 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_685
timestamp 1649977179
transform 1 0 64124 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_697
timestamp 1649977179
transform 1 0 65228 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_709
timestamp 1649977179
transform 1 0 66332 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_724
timestamp 1649977179
transform 1 0 67712 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_729
timestamp 1649977179
transform 1 0 68172 0 -1 44608
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_78_3
timestamp 1649977179
transform 1 0 1380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_15
timestamp 1649977179
transform 1 0 2484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 1649977179
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_29
timestamp 1649977179
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_41
timestamp 1649977179
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_53
timestamp 1649977179
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_65
timestamp 1649977179
transform 1 0 7084 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_77
timestamp 1649977179
transform 1 0 8188 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_83
timestamp 1649977179
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_85
timestamp 1649977179
transform 1 0 8924 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_97
timestamp 1649977179
transform 1 0 10028 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_109
timestamp 1649977179
transform 1 0 11132 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_121
timestamp 1649977179
transform 1 0 12236 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_133
timestamp 1649977179
transform 1 0 13340 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_139
timestamp 1649977179
transform 1 0 13892 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_141
timestamp 1649977179
transform 1 0 14076 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_153
timestamp 1649977179
transform 1 0 15180 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_165
timestamp 1649977179
transform 1 0 16284 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_177
timestamp 1649977179
transform 1 0 17388 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_189
timestamp 1649977179
transform 1 0 18492 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_195
timestamp 1649977179
transform 1 0 19044 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_197
timestamp 1649977179
transform 1 0 19228 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_209
timestamp 1649977179
transform 1 0 20332 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_221
timestamp 1649977179
transform 1 0 21436 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_233
timestamp 1649977179
transform 1 0 22540 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_245
timestamp 1649977179
transform 1 0 23644 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_251
timestamp 1649977179
transform 1 0 24196 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_253
timestamp 1649977179
transform 1 0 24380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_265
timestamp 1649977179
transform 1 0 25484 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_277
timestamp 1649977179
transform 1 0 26588 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_289
timestamp 1649977179
transform 1 0 27692 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_301
timestamp 1649977179
transform 1 0 28796 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_307
timestamp 1649977179
transform 1 0 29348 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_309
timestamp 1649977179
transform 1 0 29532 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_321
timestamp 1649977179
transform 1 0 30636 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_333
timestamp 1649977179
transform 1 0 31740 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_345
timestamp 1649977179
transform 1 0 32844 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_357
timestamp 1649977179
transform 1 0 33948 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_363
timestamp 1649977179
transform 1 0 34500 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_365
timestamp 1649977179
transform 1 0 34684 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_377
timestamp 1649977179
transform 1 0 35788 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_389
timestamp 1649977179
transform 1 0 36892 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_401
timestamp 1649977179
transform 1 0 37996 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_413
timestamp 1649977179
transform 1 0 39100 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_419
timestamp 1649977179
transform 1 0 39652 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_421
timestamp 1649977179
transform 1 0 39836 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_433
timestamp 1649977179
transform 1 0 40940 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_445
timestamp 1649977179
transform 1 0 42044 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_457
timestamp 1649977179
transform 1 0 43148 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_469
timestamp 1649977179
transform 1 0 44252 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_475
timestamp 1649977179
transform 1 0 44804 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_477
timestamp 1649977179
transform 1 0 44988 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_489
timestamp 1649977179
transform 1 0 46092 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_501
timestamp 1649977179
transform 1 0 47196 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_513
timestamp 1649977179
transform 1 0 48300 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_525
timestamp 1649977179
transform 1 0 49404 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_531
timestamp 1649977179
transform 1 0 49956 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_533
timestamp 1649977179
transform 1 0 50140 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_545
timestamp 1649977179
transform 1 0 51244 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_557
timestamp 1649977179
transform 1 0 52348 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_569
timestamp 1649977179
transform 1 0 53452 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_581
timestamp 1649977179
transform 1 0 54556 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_587
timestamp 1649977179
transform 1 0 55108 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_589
timestamp 1649977179
transform 1 0 55292 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_601
timestamp 1649977179
transform 1 0 56396 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_613
timestamp 1649977179
transform 1 0 57500 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_625
timestamp 1649977179
transform 1 0 58604 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_637
timestamp 1649977179
transform 1 0 59708 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_643
timestamp 1649977179
transform 1 0 60260 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_645
timestamp 1649977179
transform 1 0 60444 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_657
timestamp 1649977179
transform 1 0 61548 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_669
timestamp 1649977179
transform 1 0 62652 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_681
timestamp 1649977179
transform 1 0 63756 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_693
timestamp 1649977179
transform 1 0 64860 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_699
timestamp 1649977179
transform 1 0 65412 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_701
timestamp 1649977179
transform 1 0 65596 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_713
timestamp 1649977179
transform 1 0 66700 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_725
timestamp 1649977179
transform 1 0 67804 0 1 44608
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_79_3
timestamp 1649977179
transform 1 0 1380 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_15
timestamp 1649977179
transform 1 0 2484 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_27
timestamp 1649977179
transform 1 0 3588 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_39
timestamp 1649977179
transform 1 0 4692 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_51
timestamp 1649977179
transform 1 0 5796 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_55
timestamp 1649977179
transform 1 0 6164 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_57
timestamp 1649977179
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_69
timestamp 1649977179
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_81
timestamp 1649977179
transform 1 0 8556 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_93
timestamp 1649977179
transform 1 0 9660 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_105
timestamp 1649977179
transform 1 0 10764 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_111
timestamp 1649977179
transform 1 0 11316 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_113
timestamp 1649977179
transform 1 0 11500 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_125
timestamp 1649977179
transform 1 0 12604 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_137
timestamp 1649977179
transform 1 0 13708 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_149
timestamp 1649977179
transform 1 0 14812 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_161
timestamp 1649977179
transform 1 0 15916 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_167
timestamp 1649977179
transform 1 0 16468 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_169
timestamp 1649977179
transform 1 0 16652 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_181
timestamp 1649977179
transform 1 0 17756 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_193
timestamp 1649977179
transform 1 0 18860 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_205
timestamp 1649977179
transform 1 0 19964 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_217
timestamp 1649977179
transform 1 0 21068 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_223
timestamp 1649977179
transform 1 0 21620 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_225
timestamp 1649977179
transform 1 0 21804 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_237
timestamp 1649977179
transform 1 0 22908 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_249
timestamp 1649977179
transform 1 0 24012 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_261
timestamp 1649977179
transform 1 0 25116 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_273
timestamp 1649977179
transform 1 0 26220 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_279
timestamp 1649977179
transform 1 0 26772 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_281
timestamp 1649977179
transform 1 0 26956 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_293
timestamp 1649977179
transform 1 0 28060 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_305
timestamp 1649977179
transform 1 0 29164 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_317
timestamp 1649977179
transform 1 0 30268 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_329
timestamp 1649977179
transform 1 0 31372 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_335
timestamp 1649977179
transform 1 0 31924 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_337
timestamp 1649977179
transform 1 0 32108 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_349
timestamp 1649977179
transform 1 0 33212 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_361
timestamp 1649977179
transform 1 0 34316 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_373
timestamp 1649977179
transform 1 0 35420 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_385
timestamp 1649977179
transform 1 0 36524 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_391
timestamp 1649977179
transform 1 0 37076 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_393
timestamp 1649977179
transform 1 0 37260 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_405
timestamp 1649977179
transform 1 0 38364 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_417
timestamp 1649977179
transform 1 0 39468 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_429
timestamp 1649977179
transform 1 0 40572 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_441
timestamp 1649977179
transform 1 0 41676 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_447
timestamp 1649977179
transform 1 0 42228 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_449
timestamp 1649977179
transform 1 0 42412 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_461
timestamp 1649977179
transform 1 0 43516 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_473
timestamp 1649977179
transform 1 0 44620 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_485
timestamp 1649977179
transform 1 0 45724 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_497
timestamp 1649977179
transform 1 0 46828 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_503
timestamp 1649977179
transform 1 0 47380 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_505
timestamp 1649977179
transform 1 0 47564 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_517
timestamp 1649977179
transform 1 0 48668 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_529
timestamp 1649977179
transform 1 0 49772 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_541
timestamp 1649977179
transform 1 0 50876 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_553
timestamp 1649977179
transform 1 0 51980 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_559
timestamp 1649977179
transform 1 0 52532 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_561
timestamp 1649977179
transform 1 0 52716 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_573
timestamp 1649977179
transform 1 0 53820 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_585
timestamp 1649977179
transform 1 0 54924 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_597
timestamp 1649977179
transform 1 0 56028 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_609
timestamp 1649977179
transform 1 0 57132 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_615
timestamp 1649977179
transform 1 0 57684 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_617
timestamp 1649977179
transform 1 0 57868 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_629
timestamp 1649977179
transform 1 0 58972 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_641
timestamp 1649977179
transform 1 0 60076 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_653
timestamp 1649977179
transform 1 0 61180 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_665
timestamp 1649977179
transform 1 0 62284 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_671
timestamp 1649977179
transform 1 0 62836 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_673
timestamp 1649977179
transform 1 0 63020 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_685
timestamp 1649977179
transform 1 0 64124 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_697
timestamp 1649977179
transform 1 0 65228 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_709
timestamp 1649977179
transform 1 0 66332 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_721
timestamp 1649977179
transform 1 0 67436 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_727
timestamp 1649977179
transform 1 0 67988 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_729
timestamp 1649977179
transform 1 0 68172 0 -1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_80_3
timestamp 1649977179
transform 1 0 1380 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_15
timestamp 1649977179
transform 1 0 2484 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 1649977179
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_29
timestamp 1649977179
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_41
timestamp 1649977179
transform 1 0 4876 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_53
timestamp 1649977179
transform 1 0 5980 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_65
timestamp 1649977179
transform 1 0 7084 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_77
timestamp 1649977179
transform 1 0 8188 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_83
timestamp 1649977179
transform 1 0 8740 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_85
timestamp 1649977179
transform 1 0 8924 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_97
timestamp 1649977179
transform 1 0 10028 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_109
timestamp 1649977179
transform 1 0 11132 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_121
timestamp 1649977179
transform 1 0 12236 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_133
timestamp 1649977179
transform 1 0 13340 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_139
timestamp 1649977179
transform 1 0 13892 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_141
timestamp 1649977179
transform 1 0 14076 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_153
timestamp 1649977179
transform 1 0 15180 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_165
timestamp 1649977179
transform 1 0 16284 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_177
timestamp 1649977179
transform 1 0 17388 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_189
timestamp 1649977179
transform 1 0 18492 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_195
timestamp 1649977179
transform 1 0 19044 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_197
timestamp 1649977179
transform 1 0 19228 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_209
timestamp 1649977179
transform 1 0 20332 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_221
timestamp 1649977179
transform 1 0 21436 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_233
timestamp 1649977179
transform 1 0 22540 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_245
timestamp 1649977179
transform 1 0 23644 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_251
timestamp 1649977179
transform 1 0 24196 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_253
timestamp 1649977179
transform 1 0 24380 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_265
timestamp 1649977179
transform 1 0 25484 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_277
timestamp 1649977179
transform 1 0 26588 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_289
timestamp 1649977179
transform 1 0 27692 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_301
timestamp 1649977179
transform 1 0 28796 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_307
timestamp 1649977179
transform 1 0 29348 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_309
timestamp 1649977179
transform 1 0 29532 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_321
timestamp 1649977179
transform 1 0 30636 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_333
timestamp 1649977179
transform 1 0 31740 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_345
timestamp 1649977179
transform 1 0 32844 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_357
timestamp 1649977179
transform 1 0 33948 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_363
timestamp 1649977179
transform 1 0 34500 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_365
timestamp 1649977179
transform 1 0 34684 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_377
timestamp 1649977179
transform 1 0 35788 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_389
timestamp 1649977179
transform 1 0 36892 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_401
timestamp 1649977179
transform 1 0 37996 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_413
timestamp 1649977179
transform 1 0 39100 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_419
timestamp 1649977179
transform 1 0 39652 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_421
timestamp 1649977179
transform 1 0 39836 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_433
timestamp 1649977179
transform 1 0 40940 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_445
timestamp 1649977179
transform 1 0 42044 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_457
timestamp 1649977179
transform 1 0 43148 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_469
timestamp 1649977179
transform 1 0 44252 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_475
timestamp 1649977179
transform 1 0 44804 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_477
timestamp 1649977179
transform 1 0 44988 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_489
timestamp 1649977179
transform 1 0 46092 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_501
timestamp 1649977179
transform 1 0 47196 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_513
timestamp 1649977179
transform 1 0 48300 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_525
timestamp 1649977179
transform 1 0 49404 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_531
timestamp 1649977179
transform 1 0 49956 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_533
timestamp 1649977179
transform 1 0 50140 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_545
timestamp 1649977179
transform 1 0 51244 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_557
timestamp 1649977179
transform 1 0 52348 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_569
timestamp 1649977179
transform 1 0 53452 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_581
timestamp 1649977179
transform 1 0 54556 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_587
timestamp 1649977179
transform 1 0 55108 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_589
timestamp 1649977179
transform 1 0 55292 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_601
timestamp 1649977179
transform 1 0 56396 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_613
timestamp 1649977179
transform 1 0 57500 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_625
timestamp 1649977179
transform 1 0 58604 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_637
timestamp 1649977179
transform 1 0 59708 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_643
timestamp 1649977179
transform 1 0 60260 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_645
timestamp 1649977179
transform 1 0 60444 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_657
timestamp 1649977179
transform 1 0 61548 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_669
timestamp 1649977179
transform 1 0 62652 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_681
timestamp 1649977179
transform 1 0 63756 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_693
timestamp 1649977179
transform 1 0 64860 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_699
timestamp 1649977179
transform 1 0 65412 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_701
timestamp 1649977179
transform 1 0 65596 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_713
timestamp 1649977179
transform 1 0 66700 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_725
timestamp 1649977179
transform 1 0 67804 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_729
timestamp 1649977179
transform 1 0 68172 0 1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_81_3
timestamp 1649977179
transform 1 0 1380 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_15
timestamp 1649977179
transform 1 0 2484 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_27
timestamp 1649977179
transform 1 0 3588 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_39
timestamp 1649977179
transform 1 0 4692 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_51
timestamp 1649977179
transform 1 0 5796 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_55
timestamp 1649977179
transform 1 0 6164 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_57
timestamp 1649977179
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_69
timestamp 1649977179
transform 1 0 7452 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_81
timestamp 1649977179
transform 1 0 8556 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_93
timestamp 1649977179
transform 1 0 9660 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_105
timestamp 1649977179
transform 1 0 10764 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_111
timestamp 1649977179
transform 1 0 11316 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_113
timestamp 1649977179
transform 1 0 11500 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_125
timestamp 1649977179
transform 1 0 12604 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_137
timestamp 1649977179
transform 1 0 13708 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_149
timestamp 1649977179
transform 1 0 14812 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_161
timestamp 1649977179
transform 1 0 15916 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_167
timestamp 1649977179
transform 1 0 16468 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_169
timestamp 1649977179
transform 1 0 16652 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_181
timestamp 1649977179
transform 1 0 17756 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_193
timestamp 1649977179
transform 1 0 18860 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_205
timestamp 1649977179
transform 1 0 19964 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_217
timestamp 1649977179
transform 1 0 21068 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_223
timestamp 1649977179
transform 1 0 21620 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_225
timestamp 1649977179
transform 1 0 21804 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_237
timestamp 1649977179
transform 1 0 22908 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_249
timestamp 1649977179
transform 1 0 24012 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_261
timestamp 1649977179
transform 1 0 25116 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_273
timestamp 1649977179
transform 1 0 26220 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_279
timestamp 1649977179
transform 1 0 26772 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_281
timestamp 1649977179
transform 1 0 26956 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_293
timestamp 1649977179
transform 1 0 28060 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_305
timestamp 1649977179
transform 1 0 29164 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_317
timestamp 1649977179
transform 1 0 30268 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_329
timestamp 1649977179
transform 1 0 31372 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_335
timestamp 1649977179
transform 1 0 31924 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_337
timestamp 1649977179
transform 1 0 32108 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_349
timestamp 1649977179
transform 1 0 33212 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_361
timestamp 1649977179
transform 1 0 34316 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_373
timestamp 1649977179
transform 1 0 35420 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_385
timestamp 1649977179
transform 1 0 36524 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_391
timestamp 1649977179
transform 1 0 37076 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_393
timestamp 1649977179
transform 1 0 37260 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_405
timestamp 1649977179
transform 1 0 38364 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_417
timestamp 1649977179
transform 1 0 39468 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_429
timestamp 1649977179
transform 1 0 40572 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_441
timestamp 1649977179
transform 1 0 41676 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_447
timestamp 1649977179
transform 1 0 42228 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_449
timestamp 1649977179
transform 1 0 42412 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_461
timestamp 1649977179
transform 1 0 43516 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_473
timestamp 1649977179
transform 1 0 44620 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_485
timestamp 1649977179
transform 1 0 45724 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_497
timestamp 1649977179
transform 1 0 46828 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_503
timestamp 1649977179
transform 1 0 47380 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_505
timestamp 1649977179
transform 1 0 47564 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_517
timestamp 1649977179
transform 1 0 48668 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_529
timestamp 1649977179
transform 1 0 49772 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_541
timestamp 1649977179
transform 1 0 50876 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_553
timestamp 1649977179
transform 1 0 51980 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_559
timestamp 1649977179
transform 1 0 52532 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_561
timestamp 1649977179
transform 1 0 52716 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_573
timestamp 1649977179
transform 1 0 53820 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_585
timestamp 1649977179
transform 1 0 54924 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_597
timestamp 1649977179
transform 1 0 56028 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_609
timestamp 1649977179
transform 1 0 57132 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_615
timestamp 1649977179
transform 1 0 57684 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_617
timestamp 1649977179
transform 1 0 57868 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_629
timestamp 1649977179
transform 1 0 58972 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_641
timestamp 1649977179
transform 1 0 60076 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_653
timestamp 1649977179
transform 1 0 61180 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_665
timestamp 1649977179
transform 1 0 62284 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_671
timestamp 1649977179
transform 1 0 62836 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_673
timestamp 1649977179
transform 1 0 63020 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_685
timestamp 1649977179
transform 1 0 64124 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_697
timestamp 1649977179
transform 1 0 65228 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_709
timestamp 1649977179
transform 1 0 66332 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_721
timestamp 1649977179
transform 1 0 67436 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_727
timestamp 1649977179
transform 1 0 67988 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_729
timestamp 1649977179
transform 1 0 68172 0 -1 46784
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_82_3
timestamp 1649977179
transform 1 0 1380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_15
timestamp 1649977179
transform 1 0 2484 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 1649977179
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_29
timestamp 1649977179
transform 1 0 3772 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_41
timestamp 1649977179
transform 1 0 4876 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_53
timestamp 1649977179
transform 1 0 5980 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_65
timestamp 1649977179
transform 1 0 7084 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_77
timestamp 1649977179
transform 1 0 8188 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_83
timestamp 1649977179
transform 1 0 8740 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_85
timestamp 1649977179
transform 1 0 8924 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_97
timestamp 1649977179
transform 1 0 10028 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_109
timestamp 1649977179
transform 1 0 11132 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_121
timestamp 1649977179
transform 1 0 12236 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_133
timestamp 1649977179
transform 1 0 13340 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_139
timestamp 1649977179
transform 1 0 13892 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_141
timestamp 1649977179
transform 1 0 14076 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_153
timestamp 1649977179
transform 1 0 15180 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_165
timestamp 1649977179
transform 1 0 16284 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_177
timestamp 1649977179
transform 1 0 17388 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_189
timestamp 1649977179
transform 1 0 18492 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_195
timestamp 1649977179
transform 1 0 19044 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_197
timestamp 1649977179
transform 1 0 19228 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_209
timestamp 1649977179
transform 1 0 20332 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_221
timestamp 1649977179
transform 1 0 21436 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_233
timestamp 1649977179
transform 1 0 22540 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_245
timestamp 1649977179
transform 1 0 23644 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_251
timestamp 1649977179
transform 1 0 24196 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_253
timestamp 1649977179
transform 1 0 24380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_265
timestamp 1649977179
transform 1 0 25484 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_277
timestamp 1649977179
transform 1 0 26588 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_289
timestamp 1649977179
transform 1 0 27692 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_301
timestamp 1649977179
transform 1 0 28796 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_307
timestamp 1649977179
transform 1 0 29348 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_309
timestamp 1649977179
transform 1 0 29532 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_321
timestamp 1649977179
transform 1 0 30636 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_333
timestamp 1649977179
transform 1 0 31740 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_345
timestamp 1649977179
transform 1 0 32844 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_357
timestamp 1649977179
transform 1 0 33948 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_363
timestamp 1649977179
transform 1 0 34500 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_365
timestamp 1649977179
transform 1 0 34684 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_377
timestamp 1649977179
transform 1 0 35788 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_389
timestamp 1649977179
transform 1 0 36892 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_401
timestamp 1649977179
transform 1 0 37996 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_413
timestamp 1649977179
transform 1 0 39100 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_419
timestamp 1649977179
transform 1 0 39652 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_421
timestamp 1649977179
transform 1 0 39836 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_433
timestamp 1649977179
transform 1 0 40940 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_445
timestamp 1649977179
transform 1 0 42044 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_457
timestamp 1649977179
transform 1 0 43148 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_469
timestamp 1649977179
transform 1 0 44252 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_475
timestamp 1649977179
transform 1 0 44804 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_477
timestamp 1649977179
transform 1 0 44988 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_489
timestamp 1649977179
transform 1 0 46092 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_501
timestamp 1649977179
transform 1 0 47196 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_513
timestamp 1649977179
transform 1 0 48300 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_525
timestamp 1649977179
transform 1 0 49404 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_531
timestamp 1649977179
transform 1 0 49956 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_533
timestamp 1649977179
transform 1 0 50140 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_545
timestamp 1649977179
transform 1 0 51244 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_557
timestamp 1649977179
transform 1 0 52348 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_569
timestamp 1649977179
transform 1 0 53452 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_581
timestamp 1649977179
transform 1 0 54556 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_587
timestamp 1649977179
transform 1 0 55108 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_589
timestamp 1649977179
transform 1 0 55292 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_601
timestamp 1649977179
transform 1 0 56396 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_613
timestamp 1649977179
transform 1 0 57500 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_625
timestamp 1649977179
transform 1 0 58604 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_637
timestamp 1649977179
transform 1 0 59708 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_643
timestamp 1649977179
transform 1 0 60260 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_645
timestamp 1649977179
transform 1 0 60444 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_657
timestamp 1649977179
transform 1 0 61548 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_669
timestamp 1649977179
transform 1 0 62652 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_681
timestamp 1649977179
transform 1 0 63756 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_693
timestamp 1649977179
transform 1 0 64860 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_699
timestamp 1649977179
transform 1 0 65412 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_701
timestamp 1649977179
transform 1 0 65596 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_713
timestamp 1649977179
transform 1 0 66700 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_725
timestamp 1649977179
transform 1 0 67804 0 1 46784
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_83_3
timestamp 1649977179
transform 1 0 1380 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_15
timestamp 1649977179
transform 1 0 2484 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_27
timestamp 1649977179
transform 1 0 3588 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_39
timestamp 1649977179
transform 1 0 4692 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_51
timestamp 1649977179
transform 1 0 5796 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_55
timestamp 1649977179
transform 1 0 6164 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_57
timestamp 1649977179
transform 1 0 6348 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_69
timestamp 1649977179
transform 1 0 7452 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_81
timestamp 1649977179
transform 1 0 8556 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_93
timestamp 1649977179
transform 1 0 9660 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_105
timestamp 1649977179
transform 1 0 10764 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_111
timestamp 1649977179
transform 1 0 11316 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_113
timestamp 1649977179
transform 1 0 11500 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_125
timestamp 1649977179
transform 1 0 12604 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_137
timestamp 1649977179
transform 1 0 13708 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_149
timestamp 1649977179
transform 1 0 14812 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_161
timestamp 1649977179
transform 1 0 15916 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_167
timestamp 1649977179
transform 1 0 16468 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_169
timestamp 1649977179
transform 1 0 16652 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_181
timestamp 1649977179
transform 1 0 17756 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_193
timestamp 1649977179
transform 1 0 18860 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_205
timestamp 1649977179
transform 1 0 19964 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_217
timestamp 1649977179
transform 1 0 21068 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_223
timestamp 1649977179
transform 1 0 21620 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_225
timestamp 1649977179
transform 1 0 21804 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_237
timestamp 1649977179
transform 1 0 22908 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_249
timestamp 1649977179
transform 1 0 24012 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_261
timestamp 1649977179
transform 1 0 25116 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_273
timestamp 1649977179
transform 1 0 26220 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_279
timestamp 1649977179
transform 1 0 26772 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_281
timestamp 1649977179
transform 1 0 26956 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_293
timestamp 1649977179
transform 1 0 28060 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_305
timestamp 1649977179
transform 1 0 29164 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_317
timestamp 1649977179
transform 1 0 30268 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_329
timestamp 1649977179
transform 1 0 31372 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_335
timestamp 1649977179
transform 1 0 31924 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_337
timestamp 1649977179
transform 1 0 32108 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_349
timestamp 1649977179
transform 1 0 33212 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_361
timestamp 1649977179
transform 1 0 34316 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_373
timestamp 1649977179
transform 1 0 35420 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_385
timestamp 1649977179
transform 1 0 36524 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_391
timestamp 1649977179
transform 1 0 37076 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_393
timestamp 1649977179
transform 1 0 37260 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_405
timestamp 1649977179
transform 1 0 38364 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_417
timestamp 1649977179
transform 1 0 39468 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_429
timestamp 1649977179
transform 1 0 40572 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_441
timestamp 1649977179
transform 1 0 41676 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_447
timestamp 1649977179
transform 1 0 42228 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_449
timestamp 1649977179
transform 1 0 42412 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_461
timestamp 1649977179
transform 1 0 43516 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_473
timestamp 1649977179
transform 1 0 44620 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_485
timestamp 1649977179
transform 1 0 45724 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_497
timestamp 1649977179
transform 1 0 46828 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_503
timestamp 1649977179
transform 1 0 47380 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_505
timestamp 1649977179
transform 1 0 47564 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_517
timestamp 1649977179
transform 1 0 48668 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_529
timestamp 1649977179
transform 1 0 49772 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_541
timestamp 1649977179
transform 1 0 50876 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_553
timestamp 1649977179
transform 1 0 51980 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_559
timestamp 1649977179
transform 1 0 52532 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_561
timestamp 1649977179
transform 1 0 52716 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_573
timestamp 1649977179
transform 1 0 53820 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_585
timestamp 1649977179
transform 1 0 54924 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_597
timestamp 1649977179
transform 1 0 56028 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_609
timestamp 1649977179
transform 1 0 57132 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_615
timestamp 1649977179
transform 1 0 57684 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_617
timestamp 1649977179
transform 1 0 57868 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_629
timestamp 1649977179
transform 1 0 58972 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_641
timestamp 1649977179
transform 1 0 60076 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_653
timestamp 1649977179
transform 1 0 61180 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_665
timestamp 1649977179
transform 1 0 62284 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_671
timestamp 1649977179
transform 1 0 62836 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_673
timestamp 1649977179
transform 1 0 63020 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_685
timestamp 1649977179
transform 1 0 64124 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_697
timestamp 1649977179
transform 1 0 65228 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_709
timestamp 1649977179
transform 1 0 66332 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_724
timestamp 1649977179
transform 1 0 67712 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_729
timestamp 1649977179
transform 1 0 68172 0 -1 47872
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_84_3
timestamp 1649977179
transform 1 0 1380 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_15
timestamp 1649977179
transform 1 0 2484 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_84_27
timestamp 1649977179
transform 1 0 3588 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_29
timestamp 1649977179
transform 1 0 3772 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_41
timestamp 1649977179
transform 1 0 4876 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_53
timestamp 1649977179
transform 1 0 5980 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_65
timestamp 1649977179
transform 1 0 7084 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_77
timestamp 1649977179
transform 1 0 8188 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_83
timestamp 1649977179
transform 1 0 8740 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_85
timestamp 1649977179
transform 1 0 8924 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_97
timestamp 1649977179
transform 1 0 10028 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_109
timestamp 1649977179
transform 1 0 11132 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_121
timestamp 1649977179
transform 1 0 12236 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_133
timestamp 1649977179
transform 1 0 13340 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_139
timestamp 1649977179
transform 1 0 13892 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_141
timestamp 1649977179
transform 1 0 14076 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_153
timestamp 1649977179
transform 1 0 15180 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_165
timestamp 1649977179
transform 1 0 16284 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_177
timestamp 1649977179
transform 1 0 17388 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_189
timestamp 1649977179
transform 1 0 18492 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_195
timestamp 1649977179
transform 1 0 19044 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_197
timestamp 1649977179
transform 1 0 19228 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_209
timestamp 1649977179
transform 1 0 20332 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_221
timestamp 1649977179
transform 1 0 21436 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_233
timestamp 1649977179
transform 1 0 22540 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_245
timestamp 1649977179
transform 1 0 23644 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_251
timestamp 1649977179
transform 1 0 24196 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_253
timestamp 1649977179
transform 1 0 24380 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_265
timestamp 1649977179
transform 1 0 25484 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_277
timestamp 1649977179
transform 1 0 26588 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_289
timestamp 1649977179
transform 1 0 27692 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_301
timestamp 1649977179
transform 1 0 28796 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_307
timestamp 1649977179
transform 1 0 29348 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_309
timestamp 1649977179
transform 1 0 29532 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_321
timestamp 1649977179
transform 1 0 30636 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_333
timestamp 1649977179
transform 1 0 31740 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_345
timestamp 1649977179
transform 1 0 32844 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_357
timestamp 1649977179
transform 1 0 33948 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_363
timestamp 1649977179
transform 1 0 34500 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_365
timestamp 1649977179
transform 1 0 34684 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_377
timestamp 1649977179
transform 1 0 35788 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_389
timestamp 1649977179
transform 1 0 36892 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_401
timestamp 1649977179
transform 1 0 37996 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_413
timestamp 1649977179
transform 1 0 39100 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_419
timestamp 1649977179
transform 1 0 39652 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_421
timestamp 1649977179
transform 1 0 39836 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_433
timestamp 1649977179
transform 1 0 40940 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_445
timestamp 1649977179
transform 1 0 42044 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_457
timestamp 1649977179
transform 1 0 43148 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_469
timestamp 1649977179
transform 1 0 44252 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_475
timestamp 1649977179
transform 1 0 44804 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_477
timestamp 1649977179
transform 1 0 44988 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_489
timestamp 1649977179
transform 1 0 46092 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_501
timestamp 1649977179
transform 1 0 47196 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_513
timestamp 1649977179
transform 1 0 48300 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_525
timestamp 1649977179
transform 1 0 49404 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_531
timestamp 1649977179
transform 1 0 49956 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_533
timestamp 1649977179
transform 1 0 50140 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_545
timestamp 1649977179
transform 1 0 51244 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_557
timestamp 1649977179
transform 1 0 52348 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_569
timestamp 1649977179
transform 1 0 53452 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_581
timestamp 1649977179
transform 1 0 54556 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_587
timestamp 1649977179
transform 1 0 55108 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_589
timestamp 1649977179
transform 1 0 55292 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_601
timestamp 1649977179
transform 1 0 56396 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_613
timestamp 1649977179
transform 1 0 57500 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_625
timestamp 1649977179
transform 1 0 58604 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_637
timestamp 1649977179
transform 1 0 59708 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_643
timestamp 1649977179
transform 1 0 60260 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_645
timestamp 1649977179
transform 1 0 60444 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_657
timestamp 1649977179
transform 1 0 61548 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_669
timestamp 1649977179
transform 1 0 62652 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_681
timestamp 1649977179
transform 1 0 63756 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_693
timestamp 1649977179
transform 1 0 64860 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_699
timestamp 1649977179
transform 1 0 65412 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_701
timestamp 1649977179
transform 1 0 65596 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_713
timestamp 1649977179
transform 1 0 66700 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_84_725
timestamp 1649977179
transform 1 0 67804 0 1 47872
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_85_3
timestamp 1649977179
transform 1 0 1380 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_15
timestamp 1649977179
transform 1 0 2484 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_27
timestamp 1649977179
transform 1 0 3588 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_39
timestamp 1649977179
transform 1 0 4692 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_51
timestamp 1649977179
transform 1 0 5796 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_55
timestamp 1649977179
transform 1 0 6164 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_57
timestamp 1649977179
transform 1 0 6348 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_69
timestamp 1649977179
transform 1 0 7452 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_81
timestamp 1649977179
transform 1 0 8556 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_93
timestamp 1649977179
transform 1 0 9660 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_105
timestamp 1649977179
transform 1 0 10764 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_111
timestamp 1649977179
transform 1 0 11316 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_113
timestamp 1649977179
transform 1 0 11500 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_125
timestamp 1649977179
transform 1 0 12604 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_137
timestamp 1649977179
transform 1 0 13708 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_149
timestamp 1649977179
transform 1 0 14812 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_161
timestamp 1649977179
transform 1 0 15916 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_167
timestamp 1649977179
transform 1 0 16468 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_169
timestamp 1649977179
transform 1 0 16652 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_181
timestamp 1649977179
transform 1 0 17756 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_193
timestamp 1649977179
transform 1 0 18860 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_205
timestamp 1649977179
transform 1 0 19964 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_217
timestamp 1649977179
transform 1 0 21068 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_223
timestamp 1649977179
transform 1 0 21620 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_225
timestamp 1649977179
transform 1 0 21804 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_237
timestamp 1649977179
transform 1 0 22908 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_249
timestamp 1649977179
transform 1 0 24012 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_261
timestamp 1649977179
transform 1 0 25116 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_273
timestamp 1649977179
transform 1 0 26220 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_279
timestamp 1649977179
transform 1 0 26772 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_281
timestamp 1649977179
transform 1 0 26956 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_293
timestamp 1649977179
transform 1 0 28060 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_305
timestamp 1649977179
transform 1 0 29164 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_317
timestamp 1649977179
transform 1 0 30268 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_329
timestamp 1649977179
transform 1 0 31372 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_335
timestamp 1649977179
transform 1 0 31924 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_337
timestamp 1649977179
transform 1 0 32108 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_349
timestamp 1649977179
transform 1 0 33212 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_361
timestamp 1649977179
transform 1 0 34316 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_373
timestamp 1649977179
transform 1 0 35420 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_385
timestamp 1649977179
transform 1 0 36524 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_391
timestamp 1649977179
transform 1 0 37076 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_393
timestamp 1649977179
transform 1 0 37260 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_405
timestamp 1649977179
transform 1 0 38364 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_417
timestamp 1649977179
transform 1 0 39468 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_429
timestamp 1649977179
transform 1 0 40572 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_441
timestamp 1649977179
transform 1 0 41676 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_447
timestamp 1649977179
transform 1 0 42228 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_449
timestamp 1649977179
transform 1 0 42412 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_461
timestamp 1649977179
transform 1 0 43516 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_473
timestamp 1649977179
transform 1 0 44620 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_485
timestamp 1649977179
transform 1 0 45724 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_497
timestamp 1649977179
transform 1 0 46828 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_503
timestamp 1649977179
transform 1 0 47380 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_505
timestamp 1649977179
transform 1 0 47564 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_517
timestamp 1649977179
transform 1 0 48668 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_529
timestamp 1649977179
transform 1 0 49772 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_541
timestamp 1649977179
transform 1 0 50876 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_553
timestamp 1649977179
transform 1 0 51980 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_559
timestamp 1649977179
transform 1 0 52532 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_561
timestamp 1649977179
transform 1 0 52716 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_573
timestamp 1649977179
transform 1 0 53820 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_585
timestamp 1649977179
transform 1 0 54924 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_597
timestamp 1649977179
transform 1 0 56028 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_609
timestamp 1649977179
transform 1 0 57132 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_615
timestamp 1649977179
transform 1 0 57684 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_617
timestamp 1649977179
transform 1 0 57868 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_629
timestamp 1649977179
transform 1 0 58972 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_641
timestamp 1649977179
transform 1 0 60076 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_653
timestamp 1649977179
transform 1 0 61180 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_665
timestamp 1649977179
transform 1 0 62284 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_671
timestamp 1649977179
transform 1 0 62836 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_673
timestamp 1649977179
transform 1 0 63020 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_685
timestamp 1649977179
transform 1 0 64124 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_697
timestamp 1649977179
transform 1 0 65228 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_709
timestamp 1649977179
transform 1 0 66332 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_724
timestamp 1649977179
transform 1 0 67712 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_729
timestamp 1649977179
transform 1 0 68172 0 -1 48960
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_86_3
timestamp 1649977179
transform 1 0 1380 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_15
timestamp 1649977179
transform 1 0 2484 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_86_27
timestamp 1649977179
transform 1 0 3588 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_29
timestamp 1649977179
transform 1 0 3772 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_41
timestamp 1649977179
transform 1 0 4876 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_53
timestamp 1649977179
transform 1 0 5980 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_65
timestamp 1649977179
transform 1 0 7084 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_77
timestamp 1649977179
transform 1 0 8188 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_83
timestamp 1649977179
transform 1 0 8740 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_85
timestamp 1649977179
transform 1 0 8924 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_97
timestamp 1649977179
transform 1 0 10028 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_109
timestamp 1649977179
transform 1 0 11132 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_121
timestamp 1649977179
transform 1 0 12236 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_133
timestamp 1649977179
transform 1 0 13340 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_139
timestamp 1649977179
transform 1 0 13892 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_141
timestamp 1649977179
transform 1 0 14076 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_153
timestamp 1649977179
transform 1 0 15180 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_165
timestamp 1649977179
transform 1 0 16284 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_177
timestamp 1649977179
transform 1 0 17388 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_189
timestamp 1649977179
transform 1 0 18492 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_195
timestamp 1649977179
transform 1 0 19044 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_197
timestamp 1649977179
transform 1 0 19228 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_209
timestamp 1649977179
transform 1 0 20332 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_221
timestamp 1649977179
transform 1 0 21436 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_233
timestamp 1649977179
transform 1 0 22540 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_245
timestamp 1649977179
transform 1 0 23644 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_251
timestamp 1649977179
transform 1 0 24196 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_253
timestamp 1649977179
transform 1 0 24380 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_265
timestamp 1649977179
transform 1 0 25484 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_277
timestamp 1649977179
transform 1 0 26588 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_289
timestamp 1649977179
transform 1 0 27692 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_301
timestamp 1649977179
transform 1 0 28796 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_307
timestamp 1649977179
transform 1 0 29348 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_309
timestamp 1649977179
transform 1 0 29532 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_321
timestamp 1649977179
transform 1 0 30636 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_333
timestamp 1649977179
transform 1 0 31740 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_345
timestamp 1649977179
transform 1 0 32844 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_357
timestamp 1649977179
transform 1 0 33948 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_363
timestamp 1649977179
transform 1 0 34500 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_365
timestamp 1649977179
transform 1 0 34684 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_377
timestamp 1649977179
transform 1 0 35788 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_389
timestamp 1649977179
transform 1 0 36892 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_401
timestamp 1649977179
transform 1 0 37996 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_413
timestamp 1649977179
transform 1 0 39100 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_419
timestamp 1649977179
transform 1 0 39652 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_421
timestamp 1649977179
transform 1 0 39836 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_433
timestamp 1649977179
transform 1 0 40940 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_445
timestamp 1649977179
transform 1 0 42044 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_457
timestamp 1649977179
transform 1 0 43148 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_469
timestamp 1649977179
transform 1 0 44252 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_475
timestamp 1649977179
transform 1 0 44804 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_477
timestamp 1649977179
transform 1 0 44988 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_489
timestamp 1649977179
transform 1 0 46092 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_501
timestamp 1649977179
transform 1 0 47196 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_513
timestamp 1649977179
transform 1 0 48300 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_525
timestamp 1649977179
transform 1 0 49404 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_531
timestamp 1649977179
transform 1 0 49956 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_533
timestamp 1649977179
transform 1 0 50140 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_545
timestamp 1649977179
transform 1 0 51244 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_557
timestamp 1649977179
transform 1 0 52348 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_569
timestamp 1649977179
transform 1 0 53452 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_581
timestamp 1649977179
transform 1 0 54556 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_587
timestamp 1649977179
transform 1 0 55108 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_589
timestamp 1649977179
transform 1 0 55292 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_601
timestamp 1649977179
transform 1 0 56396 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_613
timestamp 1649977179
transform 1 0 57500 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_625
timestamp 1649977179
transform 1 0 58604 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_637
timestamp 1649977179
transform 1 0 59708 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_643
timestamp 1649977179
transform 1 0 60260 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_645
timestamp 1649977179
transform 1 0 60444 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_657
timestamp 1649977179
transform 1 0 61548 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_669
timestamp 1649977179
transform 1 0 62652 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_681
timestamp 1649977179
transform 1 0 63756 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_693
timestamp 1649977179
transform 1 0 64860 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_699
timestamp 1649977179
transform 1 0 65412 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_701
timestamp 1649977179
transform 1 0 65596 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_713
timestamp 1649977179
transform 1 0 66700 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_725
timestamp 1649977179
transform 1 0 67804 0 1 48960
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_87_3
timestamp 1649977179
transform 1 0 1380 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_15
timestamp 1649977179
transform 1 0 2484 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_27
timestamp 1649977179
transform 1 0 3588 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_39
timestamp 1649977179
transform 1 0 4692 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_51
timestamp 1649977179
transform 1 0 5796 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_55
timestamp 1649977179
transform 1 0 6164 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_57
timestamp 1649977179
transform 1 0 6348 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_69
timestamp 1649977179
transform 1 0 7452 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_81
timestamp 1649977179
transform 1 0 8556 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_93
timestamp 1649977179
transform 1 0 9660 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_105
timestamp 1649977179
transform 1 0 10764 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_111
timestamp 1649977179
transform 1 0 11316 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_113
timestamp 1649977179
transform 1 0 11500 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_125
timestamp 1649977179
transform 1 0 12604 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_137
timestamp 1649977179
transform 1 0 13708 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_149
timestamp 1649977179
transform 1 0 14812 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_161
timestamp 1649977179
transform 1 0 15916 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_167
timestamp 1649977179
transform 1 0 16468 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_169
timestamp 1649977179
transform 1 0 16652 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_181
timestamp 1649977179
transform 1 0 17756 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_193
timestamp 1649977179
transform 1 0 18860 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_205
timestamp 1649977179
transform 1 0 19964 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_217
timestamp 1649977179
transform 1 0 21068 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_223
timestamp 1649977179
transform 1 0 21620 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_225
timestamp 1649977179
transform 1 0 21804 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_237
timestamp 1649977179
transform 1 0 22908 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_249
timestamp 1649977179
transform 1 0 24012 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_261
timestamp 1649977179
transform 1 0 25116 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_273
timestamp 1649977179
transform 1 0 26220 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_279
timestamp 1649977179
transform 1 0 26772 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_281
timestamp 1649977179
transform 1 0 26956 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_293
timestamp 1649977179
transform 1 0 28060 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_305
timestamp 1649977179
transform 1 0 29164 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_317
timestamp 1649977179
transform 1 0 30268 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_329
timestamp 1649977179
transform 1 0 31372 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_335
timestamp 1649977179
transform 1 0 31924 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_337
timestamp 1649977179
transform 1 0 32108 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_349
timestamp 1649977179
transform 1 0 33212 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_361
timestamp 1649977179
transform 1 0 34316 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_373
timestamp 1649977179
transform 1 0 35420 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_385
timestamp 1649977179
transform 1 0 36524 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_391
timestamp 1649977179
transform 1 0 37076 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_393
timestamp 1649977179
transform 1 0 37260 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_405
timestamp 1649977179
transform 1 0 38364 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_417
timestamp 1649977179
transform 1 0 39468 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_429
timestamp 1649977179
transform 1 0 40572 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_441
timestamp 1649977179
transform 1 0 41676 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_447
timestamp 1649977179
transform 1 0 42228 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_449
timestamp 1649977179
transform 1 0 42412 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_461
timestamp 1649977179
transform 1 0 43516 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_473
timestamp 1649977179
transform 1 0 44620 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_485
timestamp 1649977179
transform 1 0 45724 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_497
timestamp 1649977179
transform 1 0 46828 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_503
timestamp 1649977179
transform 1 0 47380 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_505
timestamp 1649977179
transform 1 0 47564 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_517
timestamp 1649977179
transform 1 0 48668 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_529
timestamp 1649977179
transform 1 0 49772 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_541
timestamp 1649977179
transform 1 0 50876 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_553
timestamp 1649977179
transform 1 0 51980 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_559
timestamp 1649977179
transform 1 0 52532 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_561
timestamp 1649977179
transform 1 0 52716 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_573
timestamp 1649977179
transform 1 0 53820 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_585
timestamp 1649977179
transform 1 0 54924 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_597
timestamp 1649977179
transform 1 0 56028 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_609
timestamp 1649977179
transform 1 0 57132 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_615
timestamp 1649977179
transform 1 0 57684 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_617
timestamp 1649977179
transform 1 0 57868 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_629
timestamp 1649977179
transform 1 0 58972 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_641
timestamp 1649977179
transform 1 0 60076 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_653
timestamp 1649977179
transform 1 0 61180 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_665
timestamp 1649977179
transform 1 0 62284 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_671
timestamp 1649977179
transform 1 0 62836 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_673
timestamp 1649977179
transform 1 0 63020 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_685
timestamp 1649977179
transform 1 0 64124 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_697
timestamp 1649977179
transform 1 0 65228 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_709
timestamp 1649977179
transform 1 0 66332 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_721
timestamp 1649977179
transform 1 0 67436 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_727
timestamp 1649977179
transform 1 0 67988 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_87_729
timestamp 1649977179
transform 1 0 68172 0 -1 50048
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_88_3
timestamp 1649977179
transform 1 0 1380 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_15
timestamp 1649977179
transform 1 0 2484 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_88_27
timestamp 1649977179
transform 1 0 3588 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_29
timestamp 1649977179
transform 1 0 3772 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_41
timestamp 1649977179
transform 1 0 4876 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_53
timestamp 1649977179
transform 1 0 5980 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_65
timestamp 1649977179
transform 1 0 7084 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_77
timestamp 1649977179
transform 1 0 8188 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_83
timestamp 1649977179
transform 1 0 8740 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_85
timestamp 1649977179
transform 1 0 8924 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_97
timestamp 1649977179
transform 1 0 10028 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_109
timestamp 1649977179
transform 1 0 11132 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_121
timestamp 1649977179
transform 1 0 12236 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_133
timestamp 1649977179
transform 1 0 13340 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_139
timestamp 1649977179
transform 1 0 13892 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_141
timestamp 1649977179
transform 1 0 14076 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_153
timestamp 1649977179
transform 1 0 15180 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_165
timestamp 1649977179
transform 1 0 16284 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_177
timestamp 1649977179
transform 1 0 17388 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_189
timestamp 1649977179
transform 1 0 18492 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_195
timestamp 1649977179
transform 1 0 19044 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_197
timestamp 1649977179
transform 1 0 19228 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_209
timestamp 1649977179
transform 1 0 20332 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_221
timestamp 1649977179
transform 1 0 21436 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_233
timestamp 1649977179
transform 1 0 22540 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_245
timestamp 1649977179
transform 1 0 23644 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_251
timestamp 1649977179
transform 1 0 24196 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_253
timestamp 1649977179
transform 1 0 24380 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_265
timestamp 1649977179
transform 1 0 25484 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_277
timestamp 1649977179
transform 1 0 26588 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_289
timestamp 1649977179
transform 1 0 27692 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_301
timestamp 1649977179
transform 1 0 28796 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_307
timestamp 1649977179
transform 1 0 29348 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_309
timestamp 1649977179
transform 1 0 29532 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_321
timestamp 1649977179
transform 1 0 30636 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_333
timestamp 1649977179
transform 1 0 31740 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_345
timestamp 1649977179
transform 1 0 32844 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_357
timestamp 1649977179
transform 1 0 33948 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_363
timestamp 1649977179
transform 1 0 34500 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_365
timestamp 1649977179
transform 1 0 34684 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_377
timestamp 1649977179
transform 1 0 35788 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_389
timestamp 1649977179
transform 1 0 36892 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_401
timestamp 1649977179
transform 1 0 37996 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_413
timestamp 1649977179
transform 1 0 39100 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_419
timestamp 1649977179
transform 1 0 39652 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_421
timestamp 1649977179
transform 1 0 39836 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_433
timestamp 1649977179
transform 1 0 40940 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_445
timestamp 1649977179
transform 1 0 42044 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_457
timestamp 1649977179
transform 1 0 43148 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_469
timestamp 1649977179
transform 1 0 44252 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_475
timestamp 1649977179
transform 1 0 44804 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_477
timestamp 1649977179
transform 1 0 44988 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_489
timestamp 1649977179
transform 1 0 46092 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_501
timestamp 1649977179
transform 1 0 47196 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_513
timestamp 1649977179
transform 1 0 48300 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_525
timestamp 1649977179
transform 1 0 49404 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_531
timestamp 1649977179
transform 1 0 49956 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_533
timestamp 1649977179
transform 1 0 50140 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_545
timestamp 1649977179
transform 1 0 51244 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_557
timestamp 1649977179
transform 1 0 52348 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_569
timestamp 1649977179
transform 1 0 53452 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_581
timestamp 1649977179
transform 1 0 54556 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_587
timestamp 1649977179
transform 1 0 55108 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_589
timestamp 1649977179
transform 1 0 55292 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_601
timestamp 1649977179
transform 1 0 56396 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_613
timestamp 1649977179
transform 1 0 57500 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_625
timestamp 1649977179
transform 1 0 58604 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_637
timestamp 1649977179
transform 1 0 59708 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_643
timestamp 1649977179
transform 1 0 60260 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_645
timestamp 1649977179
transform 1 0 60444 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_657
timestamp 1649977179
transform 1 0 61548 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_669
timestamp 1649977179
transform 1 0 62652 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_681
timestamp 1649977179
transform 1 0 63756 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_693
timestamp 1649977179
transform 1 0 64860 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_699
timestamp 1649977179
transform 1 0 65412 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_701
timestamp 1649977179
transform 1 0 65596 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_713
timestamp 1649977179
transform 1 0 66700 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_88_725
timestamp 1649977179
transform 1 0 67804 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_88_729
timestamp 1649977179
transform 1 0 68172 0 1 50048
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_89_3
timestamp 1649977179
transform 1 0 1380 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_15
timestamp 1649977179
transform 1 0 2484 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_27
timestamp 1649977179
transform 1 0 3588 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_39
timestamp 1649977179
transform 1 0 4692 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_51
timestamp 1649977179
transform 1 0 5796 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_55
timestamp 1649977179
transform 1 0 6164 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_57
timestamp 1649977179
transform 1 0 6348 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_69
timestamp 1649977179
transform 1 0 7452 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_81
timestamp 1649977179
transform 1 0 8556 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_93
timestamp 1649977179
transform 1 0 9660 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_105
timestamp 1649977179
transform 1 0 10764 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_111
timestamp 1649977179
transform 1 0 11316 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_113
timestamp 1649977179
transform 1 0 11500 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_125
timestamp 1649977179
transform 1 0 12604 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_137
timestamp 1649977179
transform 1 0 13708 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_149
timestamp 1649977179
transform 1 0 14812 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_161
timestamp 1649977179
transform 1 0 15916 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_167
timestamp 1649977179
transform 1 0 16468 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_169
timestamp 1649977179
transform 1 0 16652 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_181
timestamp 1649977179
transform 1 0 17756 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_193
timestamp 1649977179
transform 1 0 18860 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_205
timestamp 1649977179
transform 1 0 19964 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_217
timestamp 1649977179
transform 1 0 21068 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_223
timestamp 1649977179
transform 1 0 21620 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_225
timestamp 1649977179
transform 1 0 21804 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_237
timestamp 1649977179
transform 1 0 22908 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_249
timestamp 1649977179
transform 1 0 24012 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_261
timestamp 1649977179
transform 1 0 25116 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_273
timestamp 1649977179
transform 1 0 26220 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_279
timestamp 1649977179
transform 1 0 26772 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_281
timestamp 1649977179
transform 1 0 26956 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_293
timestamp 1649977179
transform 1 0 28060 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_305
timestamp 1649977179
transform 1 0 29164 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_317
timestamp 1649977179
transform 1 0 30268 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_329
timestamp 1649977179
transform 1 0 31372 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_335
timestamp 1649977179
transform 1 0 31924 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_337
timestamp 1649977179
transform 1 0 32108 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_349
timestamp 1649977179
transform 1 0 33212 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_361
timestamp 1649977179
transform 1 0 34316 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_373
timestamp 1649977179
transform 1 0 35420 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_385
timestamp 1649977179
transform 1 0 36524 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_391
timestamp 1649977179
transform 1 0 37076 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_393
timestamp 1649977179
transform 1 0 37260 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_405
timestamp 1649977179
transform 1 0 38364 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_417
timestamp 1649977179
transform 1 0 39468 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_429
timestamp 1649977179
transform 1 0 40572 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_441
timestamp 1649977179
transform 1 0 41676 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_447
timestamp 1649977179
transform 1 0 42228 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_449
timestamp 1649977179
transform 1 0 42412 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_461
timestamp 1649977179
transform 1 0 43516 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_473
timestamp 1649977179
transform 1 0 44620 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_485
timestamp 1649977179
transform 1 0 45724 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_497
timestamp 1649977179
transform 1 0 46828 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_503
timestamp 1649977179
transform 1 0 47380 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_505
timestamp 1649977179
transform 1 0 47564 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_517
timestamp 1649977179
transform 1 0 48668 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_529
timestamp 1649977179
transform 1 0 49772 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_541
timestamp 1649977179
transform 1 0 50876 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_553
timestamp 1649977179
transform 1 0 51980 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_559
timestamp 1649977179
transform 1 0 52532 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_561
timestamp 1649977179
transform 1 0 52716 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_573
timestamp 1649977179
transform 1 0 53820 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_585
timestamp 1649977179
transform 1 0 54924 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_597
timestamp 1649977179
transform 1 0 56028 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_609
timestamp 1649977179
transform 1 0 57132 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_615
timestamp 1649977179
transform 1 0 57684 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_617
timestamp 1649977179
transform 1 0 57868 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_629
timestamp 1649977179
transform 1 0 58972 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_641
timestamp 1649977179
transform 1 0 60076 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_653
timestamp 1649977179
transform 1 0 61180 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_665
timestamp 1649977179
transform 1 0 62284 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_671
timestamp 1649977179
transform 1 0 62836 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_673
timestamp 1649977179
transform 1 0 63020 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_685
timestamp 1649977179
transform 1 0 64124 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_697
timestamp 1649977179
transform 1 0 65228 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_709
timestamp 1649977179
transform 1 0 66332 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_721
timestamp 1649977179
transform 1 0 67436 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_727
timestamp 1649977179
transform 1 0 67988 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_89_729
timestamp 1649977179
transform 1 0 68172 0 -1 51136
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_90_3
timestamp 1649977179
transform 1 0 1380 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_15
timestamp 1649977179
transform 1 0 2484 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_90_27
timestamp 1649977179
transform 1 0 3588 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_29
timestamp 1649977179
transform 1 0 3772 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_41
timestamp 1649977179
transform 1 0 4876 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_53
timestamp 1649977179
transform 1 0 5980 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_65
timestamp 1649977179
transform 1 0 7084 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_77
timestamp 1649977179
transform 1 0 8188 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_83
timestamp 1649977179
transform 1 0 8740 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_85
timestamp 1649977179
transform 1 0 8924 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_97
timestamp 1649977179
transform 1 0 10028 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_109
timestamp 1649977179
transform 1 0 11132 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_121
timestamp 1649977179
transform 1 0 12236 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_133
timestamp 1649977179
transform 1 0 13340 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_139
timestamp 1649977179
transform 1 0 13892 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_141
timestamp 1649977179
transform 1 0 14076 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_153
timestamp 1649977179
transform 1 0 15180 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_165
timestamp 1649977179
transform 1 0 16284 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_177
timestamp 1649977179
transform 1 0 17388 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_189
timestamp 1649977179
transform 1 0 18492 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_195
timestamp 1649977179
transform 1 0 19044 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_197
timestamp 1649977179
transform 1 0 19228 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_209
timestamp 1649977179
transform 1 0 20332 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_221
timestamp 1649977179
transform 1 0 21436 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_233
timestamp 1649977179
transform 1 0 22540 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_245
timestamp 1649977179
transform 1 0 23644 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_251
timestamp 1649977179
transform 1 0 24196 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_253
timestamp 1649977179
transform 1 0 24380 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_265
timestamp 1649977179
transform 1 0 25484 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_277
timestamp 1649977179
transform 1 0 26588 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_289
timestamp 1649977179
transform 1 0 27692 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_301
timestamp 1649977179
transform 1 0 28796 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_307
timestamp 1649977179
transform 1 0 29348 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_309
timestamp 1649977179
transform 1 0 29532 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_321
timestamp 1649977179
transform 1 0 30636 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_333
timestamp 1649977179
transform 1 0 31740 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_345
timestamp 1649977179
transform 1 0 32844 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_357
timestamp 1649977179
transform 1 0 33948 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_363
timestamp 1649977179
transform 1 0 34500 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_365
timestamp 1649977179
transform 1 0 34684 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_377
timestamp 1649977179
transform 1 0 35788 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_389
timestamp 1649977179
transform 1 0 36892 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_401
timestamp 1649977179
transform 1 0 37996 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_413
timestamp 1649977179
transform 1 0 39100 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_419
timestamp 1649977179
transform 1 0 39652 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_421
timestamp 1649977179
transform 1 0 39836 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_433
timestamp 1649977179
transform 1 0 40940 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_445
timestamp 1649977179
transform 1 0 42044 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_457
timestamp 1649977179
transform 1 0 43148 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_469
timestamp 1649977179
transform 1 0 44252 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_475
timestamp 1649977179
transform 1 0 44804 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_477
timestamp 1649977179
transform 1 0 44988 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_489
timestamp 1649977179
transform 1 0 46092 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_501
timestamp 1649977179
transform 1 0 47196 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_513
timestamp 1649977179
transform 1 0 48300 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_525
timestamp 1649977179
transform 1 0 49404 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_531
timestamp 1649977179
transform 1 0 49956 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_533
timestamp 1649977179
transform 1 0 50140 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_545
timestamp 1649977179
transform 1 0 51244 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_557
timestamp 1649977179
transform 1 0 52348 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_569
timestamp 1649977179
transform 1 0 53452 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_581
timestamp 1649977179
transform 1 0 54556 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_587
timestamp 1649977179
transform 1 0 55108 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_589
timestamp 1649977179
transform 1 0 55292 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_601
timestamp 1649977179
transform 1 0 56396 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_613
timestamp 1649977179
transform 1 0 57500 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_625
timestamp 1649977179
transform 1 0 58604 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_637
timestamp 1649977179
transform 1 0 59708 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_643
timestamp 1649977179
transform 1 0 60260 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_645
timestamp 1649977179
transform 1 0 60444 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_657
timestamp 1649977179
transform 1 0 61548 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_669
timestamp 1649977179
transform 1 0 62652 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_681
timestamp 1649977179
transform 1 0 63756 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_693
timestamp 1649977179
transform 1 0 64860 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_699
timestamp 1649977179
transform 1 0 65412 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_701
timestamp 1649977179
transform 1 0 65596 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_713
timestamp 1649977179
transform 1 0 66700 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_90_725
timestamp 1649977179
transform 1 0 67804 0 1 51136
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_91_3
timestamp 1649977179
transform 1 0 1380 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_15
timestamp 1649977179
transform 1 0 2484 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_27
timestamp 1649977179
transform 1 0 3588 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_39
timestamp 1649977179
transform 1 0 4692 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_91_51
timestamp 1649977179
transform 1 0 5796 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_91_55
timestamp 1649977179
transform 1 0 6164 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_57
timestamp 1649977179
transform 1 0 6348 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_69
timestamp 1649977179
transform 1 0 7452 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_81
timestamp 1649977179
transform 1 0 8556 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_93
timestamp 1649977179
transform 1 0 9660 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_105
timestamp 1649977179
transform 1 0 10764 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_111
timestamp 1649977179
transform 1 0 11316 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_113
timestamp 1649977179
transform 1 0 11500 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_125
timestamp 1649977179
transform 1 0 12604 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_137
timestamp 1649977179
transform 1 0 13708 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_149
timestamp 1649977179
transform 1 0 14812 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_161
timestamp 1649977179
transform 1 0 15916 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_167
timestamp 1649977179
transform 1 0 16468 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_169
timestamp 1649977179
transform 1 0 16652 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_181
timestamp 1649977179
transform 1 0 17756 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_193
timestamp 1649977179
transform 1 0 18860 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_205
timestamp 1649977179
transform 1 0 19964 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_217
timestamp 1649977179
transform 1 0 21068 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_223
timestamp 1649977179
transform 1 0 21620 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_225
timestamp 1649977179
transform 1 0 21804 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_237
timestamp 1649977179
transform 1 0 22908 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_249
timestamp 1649977179
transform 1 0 24012 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_261
timestamp 1649977179
transform 1 0 25116 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_273
timestamp 1649977179
transform 1 0 26220 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_279
timestamp 1649977179
transform 1 0 26772 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_281
timestamp 1649977179
transform 1 0 26956 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_293
timestamp 1649977179
transform 1 0 28060 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_305
timestamp 1649977179
transform 1 0 29164 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_317
timestamp 1649977179
transform 1 0 30268 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_329
timestamp 1649977179
transform 1 0 31372 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_335
timestamp 1649977179
transform 1 0 31924 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_337
timestamp 1649977179
transform 1 0 32108 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_349
timestamp 1649977179
transform 1 0 33212 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_361
timestamp 1649977179
transform 1 0 34316 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_373
timestamp 1649977179
transform 1 0 35420 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_385
timestamp 1649977179
transform 1 0 36524 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_391
timestamp 1649977179
transform 1 0 37076 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_393
timestamp 1649977179
transform 1 0 37260 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_405
timestamp 1649977179
transform 1 0 38364 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_417
timestamp 1649977179
transform 1 0 39468 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_429
timestamp 1649977179
transform 1 0 40572 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_441
timestamp 1649977179
transform 1 0 41676 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_447
timestamp 1649977179
transform 1 0 42228 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_449
timestamp 1649977179
transform 1 0 42412 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_461
timestamp 1649977179
transform 1 0 43516 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_473
timestamp 1649977179
transform 1 0 44620 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_485
timestamp 1649977179
transform 1 0 45724 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_497
timestamp 1649977179
transform 1 0 46828 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_503
timestamp 1649977179
transform 1 0 47380 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_505
timestamp 1649977179
transform 1 0 47564 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_517
timestamp 1649977179
transform 1 0 48668 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_529
timestamp 1649977179
transform 1 0 49772 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_541
timestamp 1649977179
transform 1 0 50876 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_553
timestamp 1649977179
transform 1 0 51980 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_559
timestamp 1649977179
transform 1 0 52532 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_561
timestamp 1649977179
transform 1 0 52716 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_573
timestamp 1649977179
transform 1 0 53820 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_585
timestamp 1649977179
transform 1 0 54924 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_597
timestamp 1649977179
transform 1 0 56028 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_609
timestamp 1649977179
transform 1 0 57132 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_615
timestamp 1649977179
transform 1 0 57684 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_617
timestamp 1649977179
transform 1 0 57868 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_629
timestamp 1649977179
transform 1 0 58972 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_641
timestamp 1649977179
transform 1 0 60076 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_653
timestamp 1649977179
transform 1 0 61180 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_665
timestamp 1649977179
transform 1 0 62284 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_671
timestamp 1649977179
transform 1 0 62836 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_673
timestamp 1649977179
transform 1 0 63020 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_685
timestamp 1649977179
transform 1 0 64124 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_697
timestamp 1649977179
transform 1 0 65228 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_709
timestamp 1649977179
transform 1 0 66332 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_91_724
timestamp 1649977179
transform 1 0 67712 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_91_729
timestamp 1649977179
transform 1 0 68172 0 -1 52224
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_92_3
timestamp 1649977179
transform 1 0 1380 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_15
timestamp 1649977179
transform 1 0 2484 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_92_27
timestamp 1649977179
transform 1 0 3588 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_29
timestamp 1649977179
transform 1 0 3772 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_41
timestamp 1649977179
transform 1 0 4876 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_53
timestamp 1649977179
transform 1 0 5980 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_65
timestamp 1649977179
transform 1 0 7084 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_77
timestamp 1649977179
transform 1 0 8188 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_83
timestamp 1649977179
transform 1 0 8740 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_85
timestamp 1649977179
transform 1 0 8924 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_97
timestamp 1649977179
transform 1 0 10028 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_109
timestamp 1649977179
transform 1 0 11132 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_121
timestamp 1649977179
transform 1 0 12236 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_133
timestamp 1649977179
transform 1 0 13340 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_139
timestamp 1649977179
transform 1 0 13892 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_141
timestamp 1649977179
transform 1 0 14076 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_153
timestamp 1649977179
transform 1 0 15180 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_165
timestamp 1649977179
transform 1 0 16284 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_177
timestamp 1649977179
transform 1 0 17388 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_189
timestamp 1649977179
transform 1 0 18492 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_195
timestamp 1649977179
transform 1 0 19044 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_197
timestamp 1649977179
transform 1 0 19228 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_209
timestamp 1649977179
transform 1 0 20332 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_221
timestamp 1649977179
transform 1 0 21436 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_233
timestamp 1649977179
transform 1 0 22540 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_245
timestamp 1649977179
transform 1 0 23644 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_251
timestamp 1649977179
transform 1 0 24196 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_253
timestamp 1649977179
transform 1 0 24380 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_265
timestamp 1649977179
transform 1 0 25484 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_277
timestamp 1649977179
transform 1 0 26588 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_289
timestamp 1649977179
transform 1 0 27692 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_301
timestamp 1649977179
transform 1 0 28796 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_307
timestamp 1649977179
transform 1 0 29348 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_309
timestamp 1649977179
transform 1 0 29532 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_321
timestamp 1649977179
transform 1 0 30636 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_333
timestamp 1649977179
transform 1 0 31740 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_345
timestamp 1649977179
transform 1 0 32844 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_357
timestamp 1649977179
transform 1 0 33948 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_363
timestamp 1649977179
transform 1 0 34500 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_365
timestamp 1649977179
transform 1 0 34684 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_377
timestamp 1649977179
transform 1 0 35788 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_389
timestamp 1649977179
transform 1 0 36892 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_401
timestamp 1649977179
transform 1 0 37996 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_413
timestamp 1649977179
transform 1 0 39100 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_419
timestamp 1649977179
transform 1 0 39652 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_421
timestamp 1649977179
transform 1 0 39836 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_433
timestamp 1649977179
transform 1 0 40940 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_445
timestamp 1649977179
transform 1 0 42044 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_457
timestamp 1649977179
transform 1 0 43148 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_469
timestamp 1649977179
transform 1 0 44252 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_475
timestamp 1649977179
transform 1 0 44804 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_477
timestamp 1649977179
transform 1 0 44988 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_489
timestamp 1649977179
transform 1 0 46092 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_501
timestamp 1649977179
transform 1 0 47196 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_513
timestamp 1649977179
transform 1 0 48300 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_525
timestamp 1649977179
transform 1 0 49404 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_531
timestamp 1649977179
transform 1 0 49956 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_533
timestamp 1649977179
transform 1 0 50140 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_545
timestamp 1649977179
transform 1 0 51244 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_557
timestamp 1649977179
transform 1 0 52348 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_569
timestamp 1649977179
transform 1 0 53452 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_581
timestamp 1649977179
transform 1 0 54556 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_587
timestamp 1649977179
transform 1 0 55108 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_589
timestamp 1649977179
transform 1 0 55292 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_601
timestamp 1649977179
transform 1 0 56396 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_613
timestamp 1649977179
transform 1 0 57500 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_625
timestamp 1649977179
transform 1 0 58604 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_637
timestamp 1649977179
transform 1 0 59708 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_643
timestamp 1649977179
transform 1 0 60260 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_645
timestamp 1649977179
transform 1 0 60444 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_657
timestamp 1649977179
transform 1 0 61548 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_669
timestamp 1649977179
transform 1 0 62652 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_681
timestamp 1649977179
transform 1 0 63756 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_693
timestamp 1649977179
transform 1 0 64860 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_699
timestamp 1649977179
transform 1 0 65412 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_701
timestamp 1649977179
transform 1 0 65596 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_713
timestamp 1649977179
transform 1 0 66700 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_92_725
timestamp 1649977179
transform 1 0 67804 0 1 52224
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_93_3
timestamp 1649977179
transform 1 0 1380 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_15
timestamp 1649977179
transform 1 0 2484 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_27
timestamp 1649977179
transform 1 0 3588 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_39
timestamp 1649977179
transform 1 0 4692 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_51
timestamp 1649977179
transform 1 0 5796 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_55
timestamp 1649977179
transform 1 0 6164 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_57
timestamp 1649977179
transform 1 0 6348 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_69
timestamp 1649977179
transform 1 0 7452 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_81
timestamp 1649977179
transform 1 0 8556 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_93
timestamp 1649977179
transform 1 0 9660 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_105
timestamp 1649977179
transform 1 0 10764 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_111
timestamp 1649977179
transform 1 0 11316 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_113
timestamp 1649977179
transform 1 0 11500 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_125
timestamp 1649977179
transform 1 0 12604 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_137
timestamp 1649977179
transform 1 0 13708 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_149
timestamp 1649977179
transform 1 0 14812 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_161
timestamp 1649977179
transform 1 0 15916 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_167
timestamp 1649977179
transform 1 0 16468 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_169
timestamp 1649977179
transform 1 0 16652 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_181
timestamp 1649977179
transform 1 0 17756 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_193
timestamp 1649977179
transform 1 0 18860 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_205
timestamp 1649977179
transform 1 0 19964 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_217
timestamp 1649977179
transform 1 0 21068 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_223
timestamp 1649977179
transform 1 0 21620 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_225
timestamp 1649977179
transform 1 0 21804 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_237
timestamp 1649977179
transform 1 0 22908 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_249
timestamp 1649977179
transform 1 0 24012 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_261
timestamp 1649977179
transform 1 0 25116 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_273
timestamp 1649977179
transform 1 0 26220 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_279
timestamp 1649977179
transform 1 0 26772 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_281
timestamp 1649977179
transform 1 0 26956 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_293
timestamp 1649977179
transform 1 0 28060 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_305
timestamp 1649977179
transform 1 0 29164 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_317
timestamp 1649977179
transform 1 0 30268 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_329
timestamp 1649977179
transform 1 0 31372 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_335
timestamp 1649977179
transform 1 0 31924 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_337
timestamp 1649977179
transform 1 0 32108 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_349
timestamp 1649977179
transform 1 0 33212 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_361
timestamp 1649977179
transform 1 0 34316 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_373
timestamp 1649977179
transform 1 0 35420 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_385
timestamp 1649977179
transform 1 0 36524 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_391
timestamp 1649977179
transform 1 0 37076 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_393
timestamp 1649977179
transform 1 0 37260 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_405
timestamp 1649977179
transform 1 0 38364 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_417
timestamp 1649977179
transform 1 0 39468 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_429
timestamp 1649977179
transform 1 0 40572 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_441
timestamp 1649977179
transform 1 0 41676 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_447
timestamp 1649977179
transform 1 0 42228 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_449
timestamp 1649977179
transform 1 0 42412 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_461
timestamp 1649977179
transform 1 0 43516 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_473
timestamp 1649977179
transform 1 0 44620 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_485
timestamp 1649977179
transform 1 0 45724 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_497
timestamp 1649977179
transform 1 0 46828 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_503
timestamp 1649977179
transform 1 0 47380 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_505
timestamp 1649977179
transform 1 0 47564 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_517
timestamp 1649977179
transform 1 0 48668 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_529
timestamp 1649977179
transform 1 0 49772 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_541
timestamp 1649977179
transform 1 0 50876 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_553
timestamp 1649977179
transform 1 0 51980 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_559
timestamp 1649977179
transform 1 0 52532 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_561
timestamp 1649977179
transform 1 0 52716 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_573
timestamp 1649977179
transform 1 0 53820 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_585
timestamp 1649977179
transform 1 0 54924 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_597
timestamp 1649977179
transform 1 0 56028 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_609
timestamp 1649977179
transform 1 0 57132 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_615
timestamp 1649977179
transform 1 0 57684 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_617
timestamp 1649977179
transform 1 0 57868 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_629
timestamp 1649977179
transform 1 0 58972 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_641
timestamp 1649977179
transform 1 0 60076 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_653
timestamp 1649977179
transform 1 0 61180 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_665
timestamp 1649977179
transform 1 0 62284 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_671
timestamp 1649977179
transform 1 0 62836 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_673
timestamp 1649977179
transform 1 0 63020 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_685
timestamp 1649977179
transform 1 0 64124 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_697
timestamp 1649977179
transform 1 0 65228 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_709
timestamp 1649977179
transform 1 0 66332 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_721
timestamp 1649977179
transform 1 0 67436 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_727
timestamp 1649977179
transform 1 0 67988 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_93_729
timestamp 1649977179
transform 1 0 68172 0 -1 53312
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_94_3
timestamp 1649977179
transform 1 0 1380 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_15
timestamp 1649977179
transform 1 0 2484 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_94_27
timestamp 1649977179
transform 1 0 3588 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_29
timestamp 1649977179
transform 1 0 3772 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_41
timestamp 1649977179
transform 1 0 4876 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_53
timestamp 1649977179
transform 1 0 5980 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_65
timestamp 1649977179
transform 1 0 7084 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_77
timestamp 1649977179
transform 1 0 8188 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_83
timestamp 1649977179
transform 1 0 8740 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_85
timestamp 1649977179
transform 1 0 8924 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_97
timestamp 1649977179
transform 1 0 10028 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_109
timestamp 1649977179
transform 1 0 11132 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_121
timestamp 1649977179
transform 1 0 12236 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_133
timestamp 1649977179
transform 1 0 13340 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_139
timestamp 1649977179
transform 1 0 13892 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_141
timestamp 1649977179
transform 1 0 14076 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_153
timestamp 1649977179
transform 1 0 15180 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_165
timestamp 1649977179
transform 1 0 16284 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_177
timestamp 1649977179
transform 1 0 17388 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_189
timestamp 1649977179
transform 1 0 18492 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_195
timestamp 1649977179
transform 1 0 19044 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_197
timestamp 1649977179
transform 1 0 19228 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_209
timestamp 1649977179
transform 1 0 20332 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_221
timestamp 1649977179
transform 1 0 21436 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_233
timestamp 1649977179
transform 1 0 22540 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_245
timestamp 1649977179
transform 1 0 23644 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_251
timestamp 1649977179
transform 1 0 24196 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_253
timestamp 1649977179
transform 1 0 24380 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_265
timestamp 1649977179
transform 1 0 25484 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_277
timestamp 1649977179
transform 1 0 26588 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_289
timestamp 1649977179
transform 1 0 27692 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_301
timestamp 1649977179
transform 1 0 28796 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_307
timestamp 1649977179
transform 1 0 29348 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_309
timestamp 1649977179
transform 1 0 29532 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_321
timestamp 1649977179
transform 1 0 30636 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_333
timestamp 1649977179
transform 1 0 31740 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_345
timestamp 1649977179
transform 1 0 32844 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_357
timestamp 1649977179
transform 1 0 33948 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_363
timestamp 1649977179
transform 1 0 34500 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_365
timestamp 1649977179
transform 1 0 34684 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_377
timestamp 1649977179
transform 1 0 35788 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_389
timestamp 1649977179
transform 1 0 36892 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_401
timestamp 1649977179
transform 1 0 37996 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_413
timestamp 1649977179
transform 1 0 39100 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_419
timestamp 1649977179
transform 1 0 39652 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_421
timestamp 1649977179
transform 1 0 39836 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_433
timestamp 1649977179
transform 1 0 40940 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_445
timestamp 1649977179
transform 1 0 42044 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_457
timestamp 1649977179
transform 1 0 43148 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_469
timestamp 1649977179
transform 1 0 44252 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_475
timestamp 1649977179
transform 1 0 44804 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_477
timestamp 1649977179
transform 1 0 44988 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_489
timestamp 1649977179
transform 1 0 46092 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_501
timestamp 1649977179
transform 1 0 47196 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_513
timestamp 1649977179
transform 1 0 48300 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_525
timestamp 1649977179
transform 1 0 49404 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_531
timestamp 1649977179
transform 1 0 49956 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_533
timestamp 1649977179
transform 1 0 50140 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_545
timestamp 1649977179
transform 1 0 51244 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_557
timestamp 1649977179
transform 1 0 52348 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_569
timestamp 1649977179
transform 1 0 53452 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_581
timestamp 1649977179
transform 1 0 54556 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_587
timestamp 1649977179
transform 1 0 55108 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_589
timestamp 1649977179
transform 1 0 55292 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_601
timestamp 1649977179
transform 1 0 56396 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_613
timestamp 1649977179
transform 1 0 57500 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_625
timestamp 1649977179
transform 1 0 58604 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_637
timestamp 1649977179
transform 1 0 59708 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_643
timestamp 1649977179
transform 1 0 60260 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_645
timestamp 1649977179
transform 1 0 60444 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_657
timestamp 1649977179
transform 1 0 61548 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_669
timestamp 1649977179
transform 1 0 62652 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_681
timestamp 1649977179
transform 1 0 63756 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_693
timestamp 1649977179
transform 1 0 64860 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_699
timestamp 1649977179
transform 1 0 65412 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_701
timestamp 1649977179
transform 1 0 65596 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_713
timestamp 1649977179
transform 1 0 66700 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_94_725
timestamp 1649977179
transform 1 0 67804 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_94_729
timestamp 1649977179
transform 1 0 68172 0 1 53312
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_95_3
timestamp 1649977179
transform 1 0 1380 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_15
timestamp 1649977179
transform 1 0 2484 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_27
timestamp 1649977179
transform 1 0 3588 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_39
timestamp 1649977179
transform 1 0 4692 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_95_51
timestamp 1649977179
transform 1 0 5796 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_55
timestamp 1649977179
transform 1 0 6164 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_57
timestamp 1649977179
transform 1 0 6348 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_69
timestamp 1649977179
transform 1 0 7452 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_81
timestamp 1649977179
transform 1 0 8556 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_93
timestamp 1649977179
transform 1 0 9660 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_105
timestamp 1649977179
transform 1 0 10764 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_111
timestamp 1649977179
transform 1 0 11316 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_113
timestamp 1649977179
transform 1 0 11500 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_125
timestamp 1649977179
transform 1 0 12604 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_137
timestamp 1649977179
transform 1 0 13708 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_149
timestamp 1649977179
transform 1 0 14812 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_161
timestamp 1649977179
transform 1 0 15916 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_167
timestamp 1649977179
transform 1 0 16468 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_169
timestamp 1649977179
transform 1 0 16652 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_181
timestamp 1649977179
transform 1 0 17756 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_193
timestamp 1649977179
transform 1 0 18860 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_205
timestamp 1649977179
transform 1 0 19964 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_217
timestamp 1649977179
transform 1 0 21068 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_223
timestamp 1649977179
transform 1 0 21620 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_225
timestamp 1649977179
transform 1 0 21804 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_237
timestamp 1649977179
transform 1 0 22908 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_249
timestamp 1649977179
transform 1 0 24012 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_261
timestamp 1649977179
transform 1 0 25116 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_273
timestamp 1649977179
transform 1 0 26220 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_279
timestamp 1649977179
transform 1 0 26772 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_281
timestamp 1649977179
transform 1 0 26956 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_293
timestamp 1649977179
transform 1 0 28060 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_305
timestamp 1649977179
transform 1 0 29164 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_317
timestamp 1649977179
transform 1 0 30268 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_329
timestamp 1649977179
transform 1 0 31372 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_335
timestamp 1649977179
transform 1 0 31924 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_337
timestamp 1649977179
transform 1 0 32108 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_349
timestamp 1649977179
transform 1 0 33212 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_361
timestamp 1649977179
transform 1 0 34316 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_373
timestamp 1649977179
transform 1 0 35420 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_385
timestamp 1649977179
transform 1 0 36524 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_391
timestamp 1649977179
transform 1 0 37076 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_393
timestamp 1649977179
transform 1 0 37260 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_405
timestamp 1649977179
transform 1 0 38364 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_417
timestamp 1649977179
transform 1 0 39468 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_429
timestamp 1649977179
transform 1 0 40572 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_441
timestamp 1649977179
transform 1 0 41676 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_447
timestamp 1649977179
transform 1 0 42228 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_449
timestamp 1649977179
transform 1 0 42412 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_461
timestamp 1649977179
transform 1 0 43516 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_473
timestamp 1649977179
transform 1 0 44620 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_485
timestamp 1649977179
transform 1 0 45724 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_497
timestamp 1649977179
transform 1 0 46828 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_503
timestamp 1649977179
transform 1 0 47380 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_505
timestamp 1649977179
transform 1 0 47564 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_517
timestamp 1649977179
transform 1 0 48668 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_529
timestamp 1649977179
transform 1 0 49772 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_541
timestamp 1649977179
transform 1 0 50876 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_553
timestamp 1649977179
transform 1 0 51980 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_559
timestamp 1649977179
transform 1 0 52532 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_561
timestamp 1649977179
transform 1 0 52716 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_573
timestamp 1649977179
transform 1 0 53820 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_585
timestamp 1649977179
transform 1 0 54924 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_597
timestamp 1649977179
transform 1 0 56028 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_609
timestamp 1649977179
transform 1 0 57132 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_615
timestamp 1649977179
transform 1 0 57684 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_617
timestamp 1649977179
transform 1 0 57868 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_629
timestamp 1649977179
transform 1 0 58972 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_641
timestamp 1649977179
transform 1 0 60076 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_653
timestamp 1649977179
transform 1 0 61180 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_665
timestamp 1649977179
transform 1 0 62284 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_671
timestamp 1649977179
transform 1 0 62836 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_673
timestamp 1649977179
transform 1 0 63020 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_685
timestamp 1649977179
transform 1 0 64124 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_697
timestamp 1649977179
transform 1 0 65228 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_709
timestamp 1649977179
transform 1 0 66332 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_721
timestamp 1649977179
transform 1 0 67436 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_727
timestamp 1649977179
transform 1 0 67988 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_95_729
timestamp 1649977179
transform 1 0 68172 0 -1 54400
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_96_3
timestamp 1649977179
transform 1 0 1380 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_15
timestamp 1649977179
transform 1 0 2484 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_96_27
timestamp 1649977179
transform 1 0 3588 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_29
timestamp 1649977179
transform 1 0 3772 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_41
timestamp 1649977179
transform 1 0 4876 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_53
timestamp 1649977179
transform 1 0 5980 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_65
timestamp 1649977179
transform 1 0 7084 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_77
timestamp 1649977179
transform 1 0 8188 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_83
timestamp 1649977179
transform 1 0 8740 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_85
timestamp 1649977179
transform 1 0 8924 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_97
timestamp 1649977179
transform 1 0 10028 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_109
timestamp 1649977179
transform 1 0 11132 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_121
timestamp 1649977179
transform 1 0 12236 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_133
timestamp 1649977179
transform 1 0 13340 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_139
timestamp 1649977179
transform 1 0 13892 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_141
timestamp 1649977179
transform 1 0 14076 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_153
timestamp 1649977179
transform 1 0 15180 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_165
timestamp 1649977179
transform 1 0 16284 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_177
timestamp 1649977179
transform 1 0 17388 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_189
timestamp 1649977179
transform 1 0 18492 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_195
timestamp 1649977179
transform 1 0 19044 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_197
timestamp 1649977179
transform 1 0 19228 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_209
timestamp 1649977179
transform 1 0 20332 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_221
timestamp 1649977179
transform 1 0 21436 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_233
timestamp 1649977179
transform 1 0 22540 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_245
timestamp 1649977179
transform 1 0 23644 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_251
timestamp 1649977179
transform 1 0 24196 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_253
timestamp 1649977179
transform 1 0 24380 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_265
timestamp 1649977179
transform 1 0 25484 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_277
timestamp 1649977179
transform 1 0 26588 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_289
timestamp 1649977179
transform 1 0 27692 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_301
timestamp 1649977179
transform 1 0 28796 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_307
timestamp 1649977179
transform 1 0 29348 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_309
timestamp 1649977179
transform 1 0 29532 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_321
timestamp 1649977179
transform 1 0 30636 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_333
timestamp 1649977179
transform 1 0 31740 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_345
timestamp 1649977179
transform 1 0 32844 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_357
timestamp 1649977179
transform 1 0 33948 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_363
timestamp 1649977179
transform 1 0 34500 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_365
timestamp 1649977179
transform 1 0 34684 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_377
timestamp 1649977179
transform 1 0 35788 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_389
timestamp 1649977179
transform 1 0 36892 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_401
timestamp 1649977179
transform 1 0 37996 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_413
timestamp 1649977179
transform 1 0 39100 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_419
timestamp 1649977179
transform 1 0 39652 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_421
timestamp 1649977179
transform 1 0 39836 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_433
timestamp 1649977179
transform 1 0 40940 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_445
timestamp 1649977179
transform 1 0 42044 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_457
timestamp 1649977179
transform 1 0 43148 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_469
timestamp 1649977179
transform 1 0 44252 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_475
timestamp 1649977179
transform 1 0 44804 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_477
timestamp 1649977179
transform 1 0 44988 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_489
timestamp 1649977179
transform 1 0 46092 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_501
timestamp 1649977179
transform 1 0 47196 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_513
timestamp 1649977179
transform 1 0 48300 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_525
timestamp 1649977179
transform 1 0 49404 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_531
timestamp 1649977179
transform 1 0 49956 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_533
timestamp 1649977179
transform 1 0 50140 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_545
timestamp 1649977179
transform 1 0 51244 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_557
timestamp 1649977179
transform 1 0 52348 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_569
timestamp 1649977179
transform 1 0 53452 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_581
timestamp 1649977179
transform 1 0 54556 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_587
timestamp 1649977179
transform 1 0 55108 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_589
timestamp 1649977179
transform 1 0 55292 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_601
timestamp 1649977179
transform 1 0 56396 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_613
timestamp 1649977179
transform 1 0 57500 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_625
timestamp 1649977179
transform 1 0 58604 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_637
timestamp 1649977179
transform 1 0 59708 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_643
timestamp 1649977179
transform 1 0 60260 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_645
timestamp 1649977179
transform 1 0 60444 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_657
timestamp 1649977179
transform 1 0 61548 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_669
timestamp 1649977179
transform 1 0 62652 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_681
timestamp 1649977179
transform 1 0 63756 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_693
timestamp 1649977179
transform 1 0 64860 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_699
timestamp 1649977179
transform 1 0 65412 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_701
timestamp 1649977179
transform 1 0 65596 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_713
timestamp 1649977179
transform 1 0 66700 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_96_725
timestamp 1649977179
transform 1 0 67804 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_96_729
timestamp 1649977179
transform 1 0 68172 0 1 54400
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_97_3
timestamp 1649977179
transform 1 0 1380 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_15
timestamp 1649977179
transform 1 0 2484 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_27
timestamp 1649977179
transform 1 0 3588 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_39
timestamp 1649977179
transform 1 0 4692 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_97_51
timestamp 1649977179
transform 1 0 5796 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_97_55
timestamp 1649977179
transform 1 0 6164 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_57
timestamp 1649977179
transform 1 0 6348 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_69
timestamp 1649977179
transform 1 0 7452 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_81
timestamp 1649977179
transform 1 0 8556 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_93
timestamp 1649977179
transform 1 0 9660 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_105
timestamp 1649977179
transform 1 0 10764 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_111
timestamp 1649977179
transform 1 0 11316 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_113
timestamp 1649977179
transform 1 0 11500 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_125
timestamp 1649977179
transform 1 0 12604 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_137
timestamp 1649977179
transform 1 0 13708 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_149
timestamp 1649977179
transform 1 0 14812 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_161
timestamp 1649977179
transform 1 0 15916 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_167
timestamp 1649977179
transform 1 0 16468 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_169
timestamp 1649977179
transform 1 0 16652 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_181
timestamp 1649977179
transform 1 0 17756 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_193
timestamp 1649977179
transform 1 0 18860 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_205
timestamp 1649977179
transform 1 0 19964 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_217
timestamp 1649977179
transform 1 0 21068 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_223
timestamp 1649977179
transform 1 0 21620 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_225
timestamp 1649977179
transform 1 0 21804 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_237
timestamp 1649977179
transform 1 0 22908 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_249
timestamp 1649977179
transform 1 0 24012 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_261
timestamp 1649977179
transform 1 0 25116 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_273
timestamp 1649977179
transform 1 0 26220 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_279
timestamp 1649977179
transform 1 0 26772 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_281
timestamp 1649977179
transform 1 0 26956 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_293
timestamp 1649977179
transform 1 0 28060 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_305
timestamp 1649977179
transform 1 0 29164 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_317
timestamp 1649977179
transform 1 0 30268 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_329
timestamp 1649977179
transform 1 0 31372 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_335
timestamp 1649977179
transform 1 0 31924 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_337
timestamp 1649977179
transform 1 0 32108 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_349
timestamp 1649977179
transform 1 0 33212 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_361
timestamp 1649977179
transform 1 0 34316 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_373
timestamp 1649977179
transform 1 0 35420 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_385
timestamp 1649977179
transform 1 0 36524 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_391
timestamp 1649977179
transform 1 0 37076 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_393
timestamp 1649977179
transform 1 0 37260 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_405
timestamp 1649977179
transform 1 0 38364 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_417
timestamp 1649977179
transform 1 0 39468 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_429
timestamp 1649977179
transform 1 0 40572 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_441
timestamp 1649977179
transform 1 0 41676 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_447
timestamp 1649977179
transform 1 0 42228 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_449
timestamp 1649977179
transform 1 0 42412 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_461
timestamp 1649977179
transform 1 0 43516 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_473
timestamp 1649977179
transform 1 0 44620 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_485
timestamp 1649977179
transform 1 0 45724 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_497
timestamp 1649977179
transform 1 0 46828 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_503
timestamp 1649977179
transform 1 0 47380 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_505
timestamp 1649977179
transform 1 0 47564 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_517
timestamp 1649977179
transform 1 0 48668 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_529
timestamp 1649977179
transform 1 0 49772 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_541
timestamp 1649977179
transform 1 0 50876 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_553
timestamp 1649977179
transform 1 0 51980 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_559
timestamp 1649977179
transform 1 0 52532 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_561
timestamp 1649977179
transform 1 0 52716 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_573
timestamp 1649977179
transform 1 0 53820 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_585
timestamp 1649977179
transform 1 0 54924 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_597
timestamp 1649977179
transform 1 0 56028 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_609
timestamp 1649977179
transform 1 0 57132 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_615
timestamp 1649977179
transform 1 0 57684 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_617
timestamp 1649977179
transform 1 0 57868 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_629
timestamp 1649977179
transform 1 0 58972 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_641
timestamp 1649977179
transform 1 0 60076 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_653
timestamp 1649977179
transform 1 0 61180 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_665
timestamp 1649977179
transform 1 0 62284 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_671
timestamp 1649977179
transform 1 0 62836 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_673
timestamp 1649977179
transform 1 0 63020 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_685
timestamp 1649977179
transform 1 0 64124 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_697
timestamp 1649977179
transform 1 0 65228 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_709
timestamp 1649977179
transform 1 0 66332 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_721
timestamp 1649977179
transform 1 0 67436 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_727
timestamp 1649977179
transform 1 0 67988 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_97_729
timestamp 1649977179
transform 1 0 68172 0 -1 55488
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_98_3
timestamp 1649977179
transform 1 0 1380 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_15
timestamp 1649977179
transform 1 0 2484 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_98_27
timestamp 1649977179
transform 1 0 3588 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_29
timestamp 1649977179
transform 1 0 3772 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_41
timestamp 1649977179
transform 1 0 4876 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_53
timestamp 1649977179
transform 1 0 5980 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_65
timestamp 1649977179
transform 1 0 7084 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_77
timestamp 1649977179
transform 1 0 8188 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_83
timestamp 1649977179
transform 1 0 8740 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_85
timestamp 1649977179
transform 1 0 8924 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_97
timestamp 1649977179
transform 1 0 10028 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_109
timestamp 1649977179
transform 1 0 11132 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_121
timestamp 1649977179
transform 1 0 12236 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_133
timestamp 1649977179
transform 1 0 13340 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_139
timestamp 1649977179
transform 1 0 13892 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_141
timestamp 1649977179
transform 1 0 14076 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_153
timestamp 1649977179
transform 1 0 15180 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_165
timestamp 1649977179
transform 1 0 16284 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_177
timestamp 1649977179
transform 1 0 17388 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_189
timestamp 1649977179
transform 1 0 18492 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_195
timestamp 1649977179
transform 1 0 19044 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_197
timestamp 1649977179
transform 1 0 19228 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_209
timestamp 1649977179
transform 1 0 20332 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_221
timestamp 1649977179
transform 1 0 21436 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_233
timestamp 1649977179
transform 1 0 22540 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_245
timestamp 1649977179
transform 1 0 23644 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_251
timestamp 1649977179
transform 1 0 24196 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_253
timestamp 1649977179
transform 1 0 24380 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_265
timestamp 1649977179
transform 1 0 25484 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_277
timestamp 1649977179
transform 1 0 26588 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_289
timestamp 1649977179
transform 1 0 27692 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_301
timestamp 1649977179
transform 1 0 28796 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_307
timestamp 1649977179
transform 1 0 29348 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_309
timestamp 1649977179
transform 1 0 29532 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_321
timestamp 1649977179
transform 1 0 30636 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_333
timestamp 1649977179
transform 1 0 31740 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_345
timestamp 1649977179
transform 1 0 32844 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_357
timestamp 1649977179
transform 1 0 33948 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_363
timestamp 1649977179
transform 1 0 34500 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_365
timestamp 1649977179
transform 1 0 34684 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_377
timestamp 1649977179
transform 1 0 35788 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_389
timestamp 1649977179
transform 1 0 36892 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_401
timestamp 1649977179
transform 1 0 37996 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_413
timestamp 1649977179
transform 1 0 39100 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_419
timestamp 1649977179
transform 1 0 39652 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_421
timestamp 1649977179
transform 1 0 39836 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_433
timestamp 1649977179
transform 1 0 40940 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_445
timestamp 1649977179
transform 1 0 42044 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_457
timestamp 1649977179
transform 1 0 43148 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_469
timestamp 1649977179
transform 1 0 44252 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_475
timestamp 1649977179
transform 1 0 44804 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_477
timestamp 1649977179
transform 1 0 44988 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_489
timestamp 1649977179
transform 1 0 46092 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_501
timestamp 1649977179
transform 1 0 47196 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_513
timestamp 1649977179
transform 1 0 48300 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_525
timestamp 1649977179
transform 1 0 49404 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_531
timestamp 1649977179
transform 1 0 49956 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_533
timestamp 1649977179
transform 1 0 50140 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_545
timestamp 1649977179
transform 1 0 51244 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_557
timestamp 1649977179
transform 1 0 52348 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_569
timestamp 1649977179
transform 1 0 53452 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_581
timestamp 1649977179
transform 1 0 54556 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_587
timestamp 1649977179
transform 1 0 55108 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_589
timestamp 1649977179
transform 1 0 55292 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_601
timestamp 1649977179
transform 1 0 56396 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_613
timestamp 1649977179
transform 1 0 57500 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_625
timestamp 1649977179
transform 1 0 58604 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_637
timestamp 1649977179
transform 1 0 59708 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_643
timestamp 1649977179
transform 1 0 60260 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_645
timestamp 1649977179
transform 1 0 60444 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_657
timestamp 1649977179
transform 1 0 61548 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_669
timestamp 1649977179
transform 1 0 62652 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_681
timestamp 1649977179
transform 1 0 63756 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_693
timestamp 1649977179
transform 1 0 64860 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_699
timestamp 1649977179
transform 1 0 65412 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_701
timestamp 1649977179
transform 1 0 65596 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_713
timestamp 1649977179
transform 1 0 66700 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_98_725
timestamp 1649977179
transform 1 0 67804 0 1 55488
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_99_3
timestamp 1649977179
transform 1 0 1380 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_15
timestamp 1649977179
transform 1 0 2484 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_27
timestamp 1649977179
transform 1 0 3588 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_39
timestamp 1649977179
transform 1 0 4692 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_99_51
timestamp 1649977179
transform 1 0 5796 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_99_55
timestamp 1649977179
transform 1 0 6164 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_57
timestamp 1649977179
transform 1 0 6348 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_69
timestamp 1649977179
transform 1 0 7452 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_81
timestamp 1649977179
transform 1 0 8556 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_93
timestamp 1649977179
transform 1 0 9660 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_105
timestamp 1649977179
transform 1 0 10764 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_111
timestamp 1649977179
transform 1 0 11316 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_113
timestamp 1649977179
transform 1 0 11500 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_125
timestamp 1649977179
transform 1 0 12604 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_137
timestamp 1649977179
transform 1 0 13708 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_149
timestamp 1649977179
transform 1 0 14812 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_161
timestamp 1649977179
transform 1 0 15916 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_167
timestamp 1649977179
transform 1 0 16468 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_169
timestamp 1649977179
transform 1 0 16652 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_181
timestamp 1649977179
transform 1 0 17756 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_193
timestamp 1649977179
transform 1 0 18860 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_205
timestamp 1649977179
transform 1 0 19964 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_217
timestamp 1649977179
transform 1 0 21068 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_223
timestamp 1649977179
transform 1 0 21620 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_225
timestamp 1649977179
transform 1 0 21804 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_237
timestamp 1649977179
transform 1 0 22908 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_249
timestamp 1649977179
transform 1 0 24012 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_261
timestamp 1649977179
transform 1 0 25116 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_273
timestamp 1649977179
transform 1 0 26220 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_279
timestamp 1649977179
transform 1 0 26772 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_281
timestamp 1649977179
transform 1 0 26956 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_293
timestamp 1649977179
transform 1 0 28060 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_305
timestamp 1649977179
transform 1 0 29164 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_317
timestamp 1649977179
transform 1 0 30268 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_329
timestamp 1649977179
transform 1 0 31372 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_335
timestamp 1649977179
transform 1 0 31924 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_337
timestamp 1649977179
transform 1 0 32108 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_349
timestamp 1649977179
transform 1 0 33212 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_361
timestamp 1649977179
transform 1 0 34316 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_373
timestamp 1649977179
transform 1 0 35420 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_385
timestamp 1649977179
transform 1 0 36524 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_391
timestamp 1649977179
transform 1 0 37076 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_393
timestamp 1649977179
transform 1 0 37260 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_405
timestamp 1649977179
transform 1 0 38364 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_417
timestamp 1649977179
transform 1 0 39468 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_429
timestamp 1649977179
transform 1 0 40572 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_441
timestamp 1649977179
transform 1 0 41676 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_447
timestamp 1649977179
transform 1 0 42228 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_449
timestamp 1649977179
transform 1 0 42412 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_461
timestamp 1649977179
transform 1 0 43516 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_473
timestamp 1649977179
transform 1 0 44620 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_485
timestamp 1649977179
transform 1 0 45724 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_497
timestamp 1649977179
transform 1 0 46828 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_503
timestamp 1649977179
transform 1 0 47380 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_505
timestamp 1649977179
transform 1 0 47564 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_517
timestamp 1649977179
transform 1 0 48668 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_529
timestamp 1649977179
transform 1 0 49772 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_541
timestamp 1649977179
transform 1 0 50876 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_553
timestamp 1649977179
transform 1 0 51980 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_559
timestamp 1649977179
transform 1 0 52532 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_561
timestamp 1649977179
transform 1 0 52716 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_573
timestamp 1649977179
transform 1 0 53820 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_585
timestamp 1649977179
transform 1 0 54924 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_597
timestamp 1649977179
transform 1 0 56028 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_609
timestamp 1649977179
transform 1 0 57132 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_615
timestamp 1649977179
transform 1 0 57684 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_617
timestamp 1649977179
transform 1 0 57868 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_629
timestamp 1649977179
transform 1 0 58972 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_641
timestamp 1649977179
transform 1 0 60076 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_653
timestamp 1649977179
transform 1 0 61180 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_665
timestamp 1649977179
transform 1 0 62284 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_671
timestamp 1649977179
transform 1 0 62836 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_673
timestamp 1649977179
transform 1 0 63020 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_685
timestamp 1649977179
transform 1 0 64124 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_697
timestamp 1649977179
transform 1 0 65228 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_709
timestamp 1649977179
transform 1 0 66332 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_99_724
timestamp 1649977179
transform 1 0 67712 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_729
timestamp 1649977179
transform 1 0 68172 0 -1 56576
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_100_3
timestamp 1649977179
transform 1 0 1380 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_15
timestamp 1649977179
transform 1 0 2484 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_100_27
timestamp 1649977179
transform 1 0 3588 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_29
timestamp 1649977179
transform 1 0 3772 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_41
timestamp 1649977179
transform 1 0 4876 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_53
timestamp 1649977179
transform 1 0 5980 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_65
timestamp 1649977179
transform 1 0 7084 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_77
timestamp 1649977179
transform 1 0 8188 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_83
timestamp 1649977179
transform 1 0 8740 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_85
timestamp 1649977179
transform 1 0 8924 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_97
timestamp 1649977179
transform 1 0 10028 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_109
timestamp 1649977179
transform 1 0 11132 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_121
timestamp 1649977179
transform 1 0 12236 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_133
timestamp 1649977179
transform 1 0 13340 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_139
timestamp 1649977179
transform 1 0 13892 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_141
timestamp 1649977179
transform 1 0 14076 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_153
timestamp 1649977179
transform 1 0 15180 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_165
timestamp 1649977179
transform 1 0 16284 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_177
timestamp 1649977179
transform 1 0 17388 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_189
timestamp 1649977179
transform 1 0 18492 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_195
timestamp 1649977179
transform 1 0 19044 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_197
timestamp 1649977179
transform 1 0 19228 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_209
timestamp 1649977179
transform 1 0 20332 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_100_221
timestamp 1649977179
transform 1 0 21436 0 1 56576
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_100_226
timestamp 1649977179
transform 1 0 21896 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_238
timestamp 1649977179
transform 1 0 23000 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_100_250
timestamp 1649977179
transform 1 0 24104 0 1 56576
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_100_253
timestamp 1649977179
transform 1 0 24380 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_265
timestamp 1649977179
transform 1 0 25484 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_277
timestamp 1649977179
transform 1 0 26588 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_289
timestamp 1649977179
transform 1 0 27692 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_301
timestamp 1649977179
transform 1 0 28796 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_307
timestamp 1649977179
transform 1 0 29348 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_309
timestamp 1649977179
transform 1 0 29532 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_321
timestamp 1649977179
transform 1 0 30636 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_333
timestamp 1649977179
transform 1 0 31740 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_345
timestamp 1649977179
transform 1 0 32844 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_357
timestamp 1649977179
transform 1 0 33948 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_363
timestamp 1649977179
transform 1 0 34500 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_365
timestamp 1649977179
transform 1 0 34684 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_377
timestamp 1649977179
transform 1 0 35788 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_389
timestamp 1649977179
transform 1 0 36892 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_401
timestamp 1649977179
transform 1 0 37996 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_413
timestamp 1649977179
transform 1 0 39100 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_419
timestamp 1649977179
transform 1 0 39652 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_421
timestamp 1649977179
transform 1 0 39836 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_433
timestamp 1649977179
transform 1 0 40940 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_445
timestamp 1649977179
transform 1 0 42044 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_457
timestamp 1649977179
transform 1 0 43148 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_469
timestamp 1649977179
transform 1 0 44252 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_475
timestamp 1649977179
transform 1 0 44804 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_477
timestamp 1649977179
transform 1 0 44988 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_489
timestamp 1649977179
transform 1 0 46092 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_501
timestamp 1649977179
transform 1 0 47196 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_513
timestamp 1649977179
transform 1 0 48300 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_525
timestamp 1649977179
transform 1 0 49404 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_531
timestamp 1649977179
transform 1 0 49956 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_533
timestamp 1649977179
transform 1 0 50140 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_545
timestamp 1649977179
transform 1 0 51244 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_557
timestamp 1649977179
transform 1 0 52348 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_569
timestamp 1649977179
transform 1 0 53452 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_581
timestamp 1649977179
transform 1 0 54556 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_587
timestamp 1649977179
transform 1 0 55108 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_589
timestamp 1649977179
transform 1 0 55292 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_601
timestamp 1649977179
transform 1 0 56396 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_613
timestamp 1649977179
transform 1 0 57500 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_625
timestamp 1649977179
transform 1 0 58604 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_637
timestamp 1649977179
transform 1 0 59708 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_643
timestamp 1649977179
transform 1 0 60260 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_645
timestamp 1649977179
transform 1 0 60444 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_657
timestamp 1649977179
transform 1 0 61548 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_669
timestamp 1649977179
transform 1 0 62652 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_681
timestamp 1649977179
transform 1 0 63756 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_693
timestamp 1649977179
transform 1 0 64860 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_699
timestamp 1649977179
transform 1 0 65412 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_701
timestamp 1649977179
transform 1 0 65596 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_713
timestamp 1649977179
transform 1 0 66700 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_725
timestamp 1649977179
transform 1 0 67804 0 1 56576
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_101_3
timestamp 1649977179
transform 1 0 1380 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_15
timestamp 1649977179
transform 1 0 2484 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_101_27
timestamp 1649977179
transform 1 0 3588 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_101_29
timestamp 1649977179
transform 1 0 3772 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_35
timestamp 1649977179
transform 1 0 4324 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_39
timestamp 1649977179
transform 1 0 4692 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_101_51
timestamp 1649977179
transform 1 0 5796 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_55
timestamp 1649977179
transform 1 0 6164 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_57
timestamp 1649977179
transform 1 0 6348 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_69
timestamp 1649977179
transform 1 0 7452 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_81
timestamp 1649977179
transform 1 0 8556 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_85
timestamp 1649977179
transform 1 0 8924 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_97
timestamp 1649977179
transform 1 0 10028 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_109
timestamp 1649977179
transform 1 0 11132 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_113
timestamp 1649977179
transform 1 0 11500 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_125
timestamp 1649977179
transform 1 0 12604 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_101_134
timestamp 1649977179
transform 1 0 13432 0 -1 57664
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_101_141
timestamp 1649977179
transform 1 0 14076 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_153
timestamp 1649977179
transform 1 0 15180 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_165
timestamp 1649977179
transform 1 0 16284 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_169
timestamp 1649977179
transform 1 0 16652 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_181
timestamp 1649977179
transform 1 0 17756 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_193
timestamp 1649977179
transform 1 0 18860 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_197
timestamp 1649977179
transform 1 0 19228 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_209
timestamp 1649977179
transform 1 0 20332 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_221
timestamp 1649977179
transform 1 0 21436 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_101_225
timestamp 1649977179
transform 1 0 21804 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_230
timestamp 1649977179
transform 1 0 22264 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_101_242
timestamp 1649977179
transform 1 0 23368 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_101_250
timestamp 1649977179
transform 1 0 24104 0 -1 57664
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_101_253
timestamp 1649977179
transform 1 0 24380 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_265
timestamp 1649977179
transform 1 0 25484 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_277
timestamp 1649977179
transform 1 0 26588 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_281
timestamp 1649977179
transform 1 0 26956 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_293
timestamp 1649977179
transform 1 0 28060 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_305
timestamp 1649977179
transform 1 0 29164 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_101_309
timestamp 1649977179
transform 1 0 29532 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_101_317
timestamp 1649977179
transform 1 0 30268 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_101_325
timestamp 1649977179
transform 1 0 31004 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_101_333
timestamp 1649977179
transform 1 0 31740 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_337
timestamp 1649977179
transform 1 0 32108 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_349
timestamp 1649977179
transform 1 0 33212 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_361
timestamp 1649977179
transform 1 0 34316 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_365
timestamp 1649977179
transform 1 0 34684 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_377
timestamp 1649977179
transform 1 0 35788 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_389
timestamp 1649977179
transform 1 0 36892 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_393
timestamp 1649977179
transform 1 0 37260 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_101_405
timestamp 1649977179
transform 1 0 38364 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_101_413
timestamp 1649977179
transform 1 0 39100 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_416
timestamp 1649977179
transform 1 0 39376 0 -1 57664
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_101_425
timestamp 1649977179
transform 1 0 40204 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_101_437
timestamp 1649977179
transform 1 0 41308 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_101_445
timestamp 1649977179
transform 1 0 42044 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_449
timestamp 1649977179
transform 1 0 42412 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_461
timestamp 1649977179
transform 1 0 43516 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_473
timestamp 1649977179
transform 1 0 44620 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_477
timestamp 1649977179
transform 1 0 44988 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_489
timestamp 1649977179
transform 1 0 46092 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_501
timestamp 1649977179
transform 1 0 47196 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_101_507
timestamp 1649977179
transform 1 0 47748 0 -1 57664
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_101_515
timestamp 1649977179
transform 1 0 48484 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_101_527
timestamp 1649977179
transform 1 0 49588 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_531
timestamp 1649977179
transform 1 0 49956 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_533
timestamp 1649977179
transform 1 0 50140 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_545
timestamp 1649977179
transform 1 0 51244 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_557
timestamp 1649977179
transform 1 0 52348 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_561
timestamp 1649977179
transform 1 0 52716 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_573
timestamp 1649977179
transform 1 0 53820 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_585
timestamp 1649977179
transform 1 0 54924 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_101_589
timestamp 1649977179
transform 1 0 55292 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_101_597
timestamp 1649977179
transform 1 0 56028 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_101_602
timestamp 1649977179
transform 1 0 56488 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_101_610
timestamp 1649977179
transform 1 0 57224 0 -1 57664
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_101_617
timestamp 1649977179
transform 1 0 57868 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_629
timestamp 1649977179
transform 1 0 58972 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_641
timestamp 1649977179
transform 1 0 60076 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_645
timestamp 1649977179
transform 1 0 60444 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_657
timestamp 1649977179
transform 1 0 61548 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_669
timestamp 1649977179
transform 1 0 62652 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_673
timestamp 1649977179
transform 1 0 63020 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_101_685
timestamp 1649977179
transform 1 0 64124 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_101_693
timestamp 1649977179
transform 1 0 64860 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_696
timestamp 1649977179
transform 1 0 65136 0 -1 57664
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_101_705
timestamp 1649977179
transform 1 0 65964 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_101_717
timestamp 1649977179
transform 1 0 67068 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_724
timestamp 1649977179
transform 1 0 67712 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_729
timestamp 1649977179
transform 1 0 68172 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1649977179
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1649977179
transform -1 0 68816 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1649977179
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1649977179
transform -1 0 68816 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1649977179
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1649977179
transform -1 0 68816 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1649977179
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1649977179
transform -1 0 68816 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1649977179
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1649977179
transform -1 0 68816 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1649977179
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1649977179
transform -1 0 68816 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1649977179
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1649977179
transform -1 0 68816 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1649977179
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1649977179
transform -1 0 68816 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1649977179
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1649977179
transform -1 0 68816 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1649977179
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1649977179
transform -1 0 68816 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1649977179
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1649977179
transform -1 0 68816 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1649977179
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1649977179
transform -1 0 68816 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1649977179
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1649977179
transform -1 0 68816 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1649977179
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1649977179
transform -1 0 68816 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1649977179
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1649977179
transform -1 0 68816 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1649977179
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1649977179
transform -1 0 68816 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1649977179
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1649977179
transform -1 0 68816 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1649977179
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1649977179
transform -1 0 68816 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1649977179
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1649977179
transform -1 0 68816 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1649977179
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1649977179
transform -1 0 68816 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1649977179
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1649977179
transform -1 0 68816 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1649977179
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1649977179
transform -1 0 68816 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1649977179
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1649977179
transform -1 0 68816 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1649977179
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1649977179
transform -1 0 68816 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1649977179
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1649977179
transform -1 0 68816 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1649977179
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1649977179
transform -1 0 68816 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1649977179
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1649977179
transform -1 0 68816 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1649977179
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1649977179
transform -1 0 68816 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1649977179
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1649977179
transform -1 0 68816 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1649977179
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1649977179
transform -1 0 68816 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1649977179
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1649977179
transform -1 0 68816 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1649977179
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1649977179
transform -1 0 68816 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1649977179
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1649977179
transform -1 0 68816 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1649977179
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1649977179
transform -1 0 68816 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1649977179
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1649977179
transform -1 0 68816 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1649977179
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1649977179
transform -1 0 68816 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1649977179
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1649977179
transform -1 0 68816 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1649977179
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1649977179
transform -1 0 68816 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1649977179
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1649977179
transform -1 0 68816 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1649977179
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1649977179
transform -1 0 68816 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1649977179
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1649977179
transform -1 0 68816 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1649977179
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1649977179
transform -1 0 68816 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1649977179
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1649977179
transform -1 0 68816 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1649977179
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1649977179
transform -1 0 68816 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1649977179
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1649977179
transform -1 0 68816 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1649977179
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1649977179
transform -1 0 68816 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1649977179
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1649977179
transform -1 0 68816 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1649977179
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1649977179
transform -1 0 68816 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1649977179
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1649977179
transform -1 0 68816 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1649977179
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1649977179
transform -1 0 68816 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1649977179
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1649977179
transform -1 0 68816 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1649977179
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1649977179
transform -1 0 68816 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1649977179
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1649977179
transform -1 0 68816 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1649977179
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1649977179
transform -1 0 68816 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1649977179
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1649977179
transform -1 0 68816 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1649977179
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1649977179
transform -1 0 68816 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1649977179
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1649977179
transform -1 0 68816 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1649977179
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1649977179
transform -1 0 68816 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1649977179
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1649977179
transform -1 0 68816 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1649977179
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1649977179
transform -1 0 68816 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1649977179
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1649977179
transform -1 0 68816 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1649977179
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1649977179
transform -1 0 68816 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1649977179
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1649977179
transform -1 0 68816 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1649977179
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1649977179
transform -1 0 68816 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1649977179
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1649977179
transform -1 0 68816 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1649977179
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1649977179
transform -1 0 68816 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1649977179
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1649977179
transform -1 0 68816 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1649977179
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1649977179
transform -1 0 68816 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1649977179
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1649977179
transform -1 0 68816 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1649977179
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1649977179
transform -1 0 68816 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1649977179
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1649977179
transform -1 0 68816 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1649977179
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1649977179
transform -1 0 68816 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1649977179
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1649977179
transform -1 0 68816 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1649977179
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1649977179
transform -1 0 68816 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1649977179
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1649977179
transform -1 0 68816 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1649977179
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1649977179
transform -1 0 68816 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1649977179
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1649977179
transform -1 0 68816 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1649977179
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1649977179
transform -1 0 68816 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1649977179
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1649977179
transform -1 0 68816 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1649977179
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1649977179
transform -1 0 68816 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1649977179
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1649977179
transform -1 0 68816 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1649977179
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1649977179
transform -1 0 68816 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1649977179
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1649977179
transform -1 0 68816 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_166
timestamp 1649977179
transform 1 0 1104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 1649977179
transform -1 0 68816 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_168
timestamp 1649977179
transform 1 0 1104 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_169
timestamp 1649977179
transform -1 0 68816 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_170
timestamp 1649977179
transform 1 0 1104 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_171
timestamp 1649977179
transform -1 0 68816 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_172
timestamp 1649977179
transform 1 0 1104 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_173
timestamp 1649977179
transform -1 0 68816 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_174
timestamp 1649977179
transform 1 0 1104 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_175
timestamp 1649977179
transform -1 0 68816 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_176
timestamp 1649977179
transform 1 0 1104 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_177
timestamp 1649977179
transform -1 0 68816 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_178
timestamp 1649977179
transform 1 0 1104 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_179
timestamp 1649977179
transform -1 0 68816 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_180
timestamp 1649977179
transform 1 0 1104 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_181
timestamp 1649977179
transform -1 0 68816 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_182
timestamp 1649977179
transform 1 0 1104 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_183
timestamp 1649977179
transform -1 0 68816 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_184
timestamp 1649977179
transform 1 0 1104 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_185
timestamp 1649977179
transform -1 0 68816 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_186
timestamp 1649977179
transform 1 0 1104 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_187
timestamp 1649977179
transform -1 0 68816 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_188
timestamp 1649977179
transform 1 0 1104 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_189
timestamp 1649977179
transform -1 0 68816 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_190
timestamp 1649977179
transform 1 0 1104 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_191
timestamp 1649977179
transform -1 0 68816 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_192
timestamp 1649977179
transform 1 0 1104 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_193
timestamp 1649977179
transform -1 0 68816 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_194
timestamp 1649977179
transform 1 0 1104 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_195
timestamp 1649977179
transform -1 0 68816 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_196
timestamp 1649977179
transform 1 0 1104 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_197
timestamp 1649977179
transform -1 0 68816 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_198
timestamp 1649977179
transform 1 0 1104 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_199
timestamp 1649977179
transform -1 0 68816 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_200
timestamp 1649977179
transform 1 0 1104 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_201
timestamp 1649977179
transform -1 0 68816 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_202
timestamp 1649977179
transform 1 0 1104 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_203
timestamp 1649977179
transform -1 0 68816 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1649977179
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1649977179
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1649977179
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1649977179
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1649977179
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1649977179
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1649977179
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1649977179
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1649977179
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1649977179
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1649977179
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1649977179
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1649977179
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1649977179
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1649977179
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1649977179
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1649977179
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1649977179
transform 1 0 50048 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1649977179
transform 1 0 52624 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1649977179
transform 1 0 55200 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1649977179
transform 1 0 57776 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1649977179
transform 1 0 60352 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1649977179
transform 1 0 62928 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1649977179
transform 1 0 65504 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1649977179
transform 1 0 68080 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1649977179
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1649977179
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1649977179
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1649977179
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1649977179
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1649977179
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1649977179
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1649977179
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1649977179
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1649977179
transform 1 0 52624 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1649977179
transform 1 0 57776 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1649977179
transform 1 0 62928 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1649977179
transform 1 0 68080 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1649977179
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1649977179
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1649977179
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1649977179
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1649977179
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1649977179
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1649977179
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1649977179
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1649977179
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1649977179
transform 1 0 50048 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1649977179
transform 1 0 55200 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1649977179
transform 1 0 60352 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1649977179
transform 1 0 65504 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1649977179
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1649977179
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1649977179
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1649977179
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1649977179
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1649977179
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1649977179
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1649977179
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1649977179
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1649977179
transform 1 0 52624 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1649977179
transform 1 0 57776 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1649977179
transform 1 0 62928 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1649977179
transform 1 0 68080 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1649977179
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1649977179
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1649977179
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1649977179
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1649977179
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1649977179
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1649977179
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1649977179
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1649977179
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1649977179
transform 1 0 50048 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1649977179
transform 1 0 55200 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1649977179
transform 1 0 60352 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1649977179
transform 1 0 65504 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1649977179
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1649977179
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1649977179
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1649977179
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1649977179
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1649977179
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1649977179
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1649977179
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1649977179
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1649977179
transform 1 0 52624 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1649977179
transform 1 0 57776 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1649977179
transform 1 0 62928 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1649977179
transform 1 0 68080 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1649977179
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1649977179
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1649977179
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1649977179
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1649977179
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1649977179
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1649977179
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1649977179
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1649977179
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1649977179
transform 1 0 50048 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1649977179
transform 1 0 55200 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1649977179
transform 1 0 60352 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1649977179
transform 1 0 65504 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1649977179
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1649977179
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1649977179
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1649977179
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1649977179
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1649977179
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1649977179
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1649977179
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1649977179
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1649977179
transform 1 0 52624 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1649977179
transform 1 0 57776 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1649977179
transform 1 0 62928 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1649977179
transform 1 0 68080 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1649977179
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1649977179
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1649977179
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1649977179
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1649977179
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1649977179
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1649977179
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1649977179
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1649977179
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1649977179
transform 1 0 50048 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1649977179
transform 1 0 55200 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1649977179
transform 1 0 60352 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1649977179
transform 1 0 65504 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1649977179
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1649977179
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1649977179
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1649977179
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1649977179
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1649977179
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1649977179
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1649977179
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1649977179
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1649977179
transform 1 0 52624 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1649977179
transform 1 0 57776 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1649977179
transform 1 0 62928 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1649977179
transform 1 0 68080 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1649977179
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1649977179
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1649977179
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1649977179
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1649977179
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1649977179
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1649977179
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1649977179
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1649977179
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1649977179
transform 1 0 50048 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1649977179
transform 1 0 55200 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1649977179
transform 1 0 60352 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1649977179
transform 1 0 65504 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1649977179
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1649977179
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1649977179
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1649977179
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1649977179
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1649977179
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1649977179
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1649977179
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1649977179
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1649977179
transform 1 0 52624 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1649977179
transform 1 0 57776 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1649977179
transform 1 0 62928 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1649977179
transform 1 0 68080 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1649977179
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1649977179
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1649977179
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1649977179
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1649977179
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1649977179
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1649977179
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1649977179
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1649977179
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1649977179
transform 1 0 50048 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1649977179
transform 1 0 55200 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1649977179
transform 1 0 60352 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1649977179
transform 1 0 65504 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1649977179
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1649977179
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1649977179
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1649977179
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1649977179
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1649977179
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1649977179
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1649977179
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1649977179
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1649977179
transform 1 0 52624 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1649977179
transform 1 0 57776 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1649977179
transform 1 0 62928 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1649977179
transform 1 0 68080 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1649977179
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1649977179
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1649977179
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1649977179
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1649977179
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1649977179
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1649977179
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1649977179
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1649977179
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1649977179
transform 1 0 50048 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1649977179
transform 1 0 55200 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1649977179
transform 1 0 60352 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1649977179
transform 1 0 65504 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1649977179
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1649977179
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1649977179
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1649977179
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1649977179
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1649977179
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1649977179
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1649977179
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1649977179
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1649977179
transform 1 0 52624 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1649977179
transform 1 0 57776 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1649977179
transform 1 0 62928 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1649977179
transform 1 0 68080 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1649977179
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1649977179
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1649977179
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1649977179
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1649977179
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1649977179
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1649977179
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1649977179
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1649977179
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1649977179
transform 1 0 50048 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1649977179
transform 1 0 55200 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1649977179
transform 1 0 60352 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1649977179
transform 1 0 65504 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1649977179
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1649977179
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1649977179
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1649977179
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1649977179
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1649977179
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1649977179
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1649977179
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1649977179
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1649977179
transform 1 0 52624 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1649977179
transform 1 0 57776 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1649977179
transform 1 0 62928 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1649977179
transform 1 0 68080 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1649977179
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1649977179
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1649977179
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1649977179
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1649977179
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1649977179
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1649977179
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1649977179
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1649977179
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1649977179
transform 1 0 50048 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1649977179
transform 1 0 55200 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1649977179
transform 1 0 60352 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1649977179
transform 1 0 65504 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1649977179
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1649977179
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1649977179
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1649977179
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1649977179
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1649977179
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1649977179
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1649977179
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1649977179
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1649977179
transform 1 0 52624 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1649977179
transform 1 0 57776 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1649977179
transform 1 0 62928 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1649977179
transform 1 0 68080 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1649977179
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1649977179
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1649977179
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1649977179
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1649977179
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1649977179
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1649977179
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1649977179
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1649977179
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1649977179
transform 1 0 50048 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1649977179
transform 1 0 55200 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1649977179
transform 1 0 60352 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1649977179
transform 1 0 65504 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1649977179
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1649977179
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1649977179
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1649977179
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1649977179
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1649977179
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1649977179
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1649977179
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1649977179
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1649977179
transform 1 0 52624 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1649977179
transform 1 0 57776 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1649977179
transform 1 0 62928 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1649977179
transform 1 0 68080 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1649977179
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1649977179
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1649977179
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1649977179
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1649977179
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1649977179
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1649977179
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1649977179
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1649977179
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1649977179
transform 1 0 50048 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1649977179
transform 1 0 55200 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1649977179
transform 1 0 60352 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1649977179
transform 1 0 65504 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1649977179
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1649977179
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1649977179
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1649977179
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1649977179
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1649977179
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1649977179
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1649977179
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1649977179
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1649977179
transform 1 0 52624 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1649977179
transform 1 0 57776 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1649977179
transform 1 0 62928 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1649977179
transform 1 0 68080 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1649977179
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1649977179
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1649977179
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1649977179
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1649977179
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1649977179
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1649977179
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1649977179
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1649977179
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1649977179
transform 1 0 50048 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1649977179
transform 1 0 55200 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1649977179
transform 1 0 60352 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1649977179
transform 1 0 65504 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1649977179
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1649977179
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1649977179
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1649977179
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1649977179
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1649977179
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1649977179
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1649977179
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1649977179
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1649977179
transform 1 0 52624 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1649977179
transform 1 0 57776 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1649977179
transform 1 0 62928 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1649977179
transform 1 0 68080 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1649977179
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1649977179
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1649977179
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1649977179
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1649977179
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1649977179
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1649977179
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1649977179
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1649977179
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1649977179
transform 1 0 50048 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1649977179
transform 1 0 55200 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1649977179
transform 1 0 60352 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1649977179
transform 1 0 65504 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1649977179
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1649977179
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1649977179
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1649977179
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1649977179
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1649977179
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1649977179
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1649977179
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1649977179
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1649977179
transform 1 0 52624 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1649977179
transform 1 0 57776 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1649977179
transform 1 0 62928 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1649977179
transform 1 0 68080 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1649977179
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1649977179
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1649977179
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1649977179
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1649977179
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1649977179
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1649977179
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1649977179
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1649977179
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1649977179
transform 1 0 50048 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1649977179
transform 1 0 55200 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1649977179
transform 1 0 60352 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1649977179
transform 1 0 65504 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1649977179
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1649977179
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1649977179
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1649977179
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1649977179
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1649977179
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1649977179
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1649977179
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1649977179
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1649977179
transform 1 0 52624 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1649977179
transform 1 0 57776 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1649977179
transform 1 0 62928 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1649977179
transform 1 0 68080 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1649977179
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1649977179
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1649977179
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1649977179
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1649977179
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1649977179
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1649977179
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1649977179
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1649977179
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1649977179
transform 1 0 50048 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1649977179
transform 1 0 55200 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1649977179
transform 1 0 60352 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1649977179
transform 1 0 65504 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1649977179
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1649977179
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1649977179
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1649977179
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1649977179
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1649977179
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1649977179
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1649977179
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1649977179
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1649977179
transform 1 0 52624 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1649977179
transform 1 0 57776 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1649977179
transform 1 0 62928 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1649977179
transform 1 0 68080 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1649977179
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1649977179
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1649977179
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1649977179
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1649977179
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1649977179
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1649977179
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1649977179
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1649977179
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1649977179
transform 1 0 50048 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1649977179
transform 1 0 55200 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1649977179
transform 1 0 60352 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1649977179
transform 1 0 65504 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1649977179
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1649977179
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1649977179
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1649977179
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1649977179
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1649977179
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1649977179
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1649977179
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1649977179
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1649977179
transform 1 0 52624 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1649977179
transform 1 0 57776 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1649977179
transform 1 0 62928 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1649977179
transform 1 0 68080 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1649977179
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1649977179
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1649977179
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1649977179
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1649977179
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1649977179
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1649977179
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1649977179
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1649977179
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1649977179
transform 1 0 50048 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1649977179
transform 1 0 55200 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1649977179
transform 1 0 60352 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1649977179
transform 1 0 65504 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1649977179
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1649977179
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1649977179
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1649977179
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1649977179
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1649977179
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1649977179
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1649977179
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1649977179
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1649977179
transform 1 0 52624 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1649977179
transform 1 0 57776 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1649977179
transform 1 0 62928 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1649977179
transform 1 0 68080 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1649977179
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1649977179
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1649977179
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1649977179
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1649977179
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1649977179
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1649977179
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1649977179
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1649977179
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1649977179
transform 1 0 50048 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1649977179
transform 1 0 55200 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1649977179
transform 1 0 60352 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1649977179
transform 1 0 65504 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1649977179
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1649977179
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1649977179
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1649977179
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1649977179
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1649977179
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1649977179
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1649977179
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1649977179
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1649977179
transform 1 0 52624 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1649977179
transform 1 0 57776 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1649977179
transform 1 0 62928 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1649977179
transform 1 0 68080 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1649977179
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1649977179
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1649977179
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1649977179
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1649977179
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1649977179
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1649977179
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1649977179
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1649977179
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1649977179
transform 1 0 50048 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1649977179
transform 1 0 55200 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1649977179
transform 1 0 60352 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1649977179
transform 1 0 65504 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1649977179
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1649977179
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1649977179
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1649977179
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1649977179
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1649977179
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1649977179
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1649977179
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1649977179
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1649977179
transform 1 0 52624 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1649977179
transform 1 0 57776 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1649977179
transform 1 0 62928 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1649977179
transform 1 0 68080 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1649977179
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1649977179
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1649977179
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1649977179
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1649977179
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1649977179
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1649977179
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1649977179
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1649977179
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1649977179
transform 1 0 50048 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1649977179
transform 1 0 55200 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1649977179
transform 1 0 60352 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1649977179
transform 1 0 65504 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1649977179
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1649977179
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1649977179
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1649977179
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1649977179
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1649977179
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1649977179
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1649977179
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1649977179
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1649977179
transform 1 0 52624 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1649977179
transform 1 0 57776 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1649977179
transform 1 0 62928 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1649977179
transform 1 0 68080 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1649977179
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1649977179
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1649977179
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1649977179
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1649977179
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1649977179
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1649977179
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1649977179
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1649977179
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1649977179
transform 1 0 50048 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1649977179
transform 1 0 55200 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1649977179
transform 1 0 60352 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1649977179
transform 1 0 65504 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1649977179
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1649977179
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1649977179
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1649977179
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1649977179
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1649977179
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1649977179
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1649977179
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1649977179
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1649977179
transform 1 0 52624 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1649977179
transform 1 0 57776 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1649977179
transform 1 0 62928 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1649977179
transform 1 0 68080 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1649977179
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1649977179
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1649977179
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1649977179
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1649977179
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1649977179
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1649977179
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1649977179
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1649977179
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1649977179
transform 1 0 50048 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1649977179
transform 1 0 55200 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1649977179
transform 1 0 60352 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1649977179
transform 1 0 65504 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1649977179
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1649977179
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1649977179
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1649977179
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1649977179
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1649977179
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1649977179
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1649977179
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1649977179
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1649977179
transform 1 0 52624 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1649977179
transform 1 0 57776 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1649977179
transform 1 0 62928 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1649977179
transform 1 0 68080 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1649977179
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1649977179
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1649977179
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1649977179
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1649977179
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1649977179
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1649977179
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1649977179
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1649977179
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1649977179
transform 1 0 50048 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1649977179
transform 1 0 55200 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1649977179
transform 1 0 60352 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1649977179
transform 1 0 65504 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1649977179
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1649977179
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1649977179
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1649977179
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1649977179
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1649977179
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1649977179
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1649977179
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1649977179
transform 1 0 47472 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1649977179
transform 1 0 52624 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1649977179
transform 1 0 57776 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1649977179
transform 1 0 62928 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1649977179
transform 1 0 68080 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1649977179
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1649977179
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1649977179
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1649977179
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1649977179
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1649977179
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1649977179
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1649977179
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1649977179
transform 1 0 44896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1649977179
transform 1 0 50048 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1649977179
transform 1 0 55200 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1649977179
transform 1 0 60352 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1649977179
transform 1 0 65504 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1649977179
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1649977179
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1649977179
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1649977179
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1649977179
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1649977179
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1649977179
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1649977179
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1649977179
transform 1 0 47472 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1649977179
transform 1 0 52624 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1649977179
transform 1 0 57776 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1649977179
transform 1 0 62928 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1649977179
transform 1 0 68080 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1649977179
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1649977179
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1649977179
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1649977179
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1649977179
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1649977179
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1649977179
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1649977179
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1649977179
transform 1 0 44896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1649977179
transform 1 0 50048 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1649977179
transform 1 0 55200 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1649977179
transform 1 0 60352 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1649977179
transform 1 0 65504 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1649977179
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1649977179
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1649977179
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1649977179
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1649977179
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1649977179
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1649977179
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1649977179
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1649977179
transform 1 0 47472 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1649977179
transform 1 0 52624 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1649977179
transform 1 0 57776 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1649977179
transform 1 0 62928 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1649977179
transform 1 0 68080 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1649977179
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1649977179
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1649977179
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1649977179
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1649977179
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1649977179
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1649977179
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1649977179
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1649977179
transform 1 0 44896 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1649977179
transform 1 0 50048 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1649977179
transform 1 0 55200 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1649977179
transform 1 0 60352 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1649977179
transform 1 0 65504 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1649977179
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1649977179
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1649977179
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1649977179
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1649977179
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1649977179
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1649977179
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1649977179
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1649977179
transform 1 0 47472 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1649977179
transform 1 0 52624 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1649977179
transform 1 0 57776 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1649977179
transform 1 0 62928 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1649977179
transform 1 0 68080 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_919
timestamp 1649977179
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_920
timestamp 1649977179
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_921
timestamp 1649977179
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_922
timestamp 1649977179
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_923
timestamp 1649977179
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_924
timestamp 1649977179
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_925
timestamp 1649977179
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_926
timestamp 1649977179
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_927
timestamp 1649977179
transform 1 0 44896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_928
timestamp 1649977179
transform 1 0 50048 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_929
timestamp 1649977179
transform 1 0 55200 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_930
timestamp 1649977179
transform 1 0 60352 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_931
timestamp 1649977179
transform 1 0 65504 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_932
timestamp 1649977179
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_933
timestamp 1649977179
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_934
timestamp 1649977179
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_935
timestamp 1649977179
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_936
timestamp 1649977179
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_937
timestamp 1649977179
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_938
timestamp 1649977179
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_939
timestamp 1649977179
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_940
timestamp 1649977179
transform 1 0 47472 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_941
timestamp 1649977179
transform 1 0 52624 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_942
timestamp 1649977179
transform 1 0 57776 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_943
timestamp 1649977179
transform 1 0 62928 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_944
timestamp 1649977179
transform 1 0 68080 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_945
timestamp 1649977179
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_946
timestamp 1649977179
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_947
timestamp 1649977179
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_948
timestamp 1649977179
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_949
timestamp 1649977179
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_950
timestamp 1649977179
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_951
timestamp 1649977179
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_952
timestamp 1649977179
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_953
timestamp 1649977179
transform 1 0 44896 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_954
timestamp 1649977179
transform 1 0 50048 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_955
timestamp 1649977179
transform 1 0 55200 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_956
timestamp 1649977179
transform 1 0 60352 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_957
timestamp 1649977179
transform 1 0 65504 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_958
timestamp 1649977179
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_959
timestamp 1649977179
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_960
timestamp 1649977179
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_961
timestamp 1649977179
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_962
timestamp 1649977179
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_963
timestamp 1649977179
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_964
timestamp 1649977179
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_965
timestamp 1649977179
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_966
timestamp 1649977179
transform 1 0 47472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_967
timestamp 1649977179
transform 1 0 52624 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_968
timestamp 1649977179
transform 1 0 57776 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_969
timestamp 1649977179
transform 1 0 62928 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_970
timestamp 1649977179
transform 1 0 68080 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_971
timestamp 1649977179
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_972
timestamp 1649977179
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_973
timestamp 1649977179
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_974
timestamp 1649977179
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_975
timestamp 1649977179
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_976
timestamp 1649977179
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_977
timestamp 1649977179
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_978
timestamp 1649977179
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_979
timestamp 1649977179
transform 1 0 44896 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_980
timestamp 1649977179
transform 1 0 50048 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_981
timestamp 1649977179
transform 1 0 55200 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_982
timestamp 1649977179
transform 1 0 60352 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_983
timestamp 1649977179
transform 1 0 65504 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_984
timestamp 1649977179
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_985
timestamp 1649977179
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_986
timestamp 1649977179
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_987
timestamp 1649977179
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_988
timestamp 1649977179
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_989
timestamp 1649977179
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_990
timestamp 1649977179
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_991
timestamp 1649977179
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_992
timestamp 1649977179
transform 1 0 47472 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_993
timestamp 1649977179
transform 1 0 52624 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_994
timestamp 1649977179
transform 1 0 57776 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_995
timestamp 1649977179
transform 1 0 62928 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_996
timestamp 1649977179
transform 1 0 68080 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_997
timestamp 1649977179
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_998
timestamp 1649977179
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_999
timestamp 1649977179
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1000
timestamp 1649977179
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1001
timestamp 1649977179
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1002
timestamp 1649977179
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1003
timestamp 1649977179
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1004
timestamp 1649977179
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1005
timestamp 1649977179
transform 1 0 44896 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1006
timestamp 1649977179
transform 1 0 50048 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1007
timestamp 1649977179
transform 1 0 55200 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1008
timestamp 1649977179
transform 1 0 60352 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1009
timestamp 1649977179
transform 1 0 65504 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1010
timestamp 1649977179
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1011
timestamp 1649977179
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1012
timestamp 1649977179
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1013
timestamp 1649977179
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1014
timestamp 1649977179
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1015
timestamp 1649977179
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1016
timestamp 1649977179
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1017
timestamp 1649977179
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1018
timestamp 1649977179
transform 1 0 47472 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1019
timestamp 1649977179
transform 1 0 52624 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1020
timestamp 1649977179
transform 1 0 57776 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1021
timestamp 1649977179
transform 1 0 62928 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1022
timestamp 1649977179
transform 1 0 68080 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1023
timestamp 1649977179
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1024
timestamp 1649977179
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1025
timestamp 1649977179
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1026
timestamp 1649977179
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1027
timestamp 1649977179
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1028
timestamp 1649977179
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1029
timestamp 1649977179
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1030
timestamp 1649977179
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1031
timestamp 1649977179
transform 1 0 44896 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1032
timestamp 1649977179
transform 1 0 50048 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1033
timestamp 1649977179
transform 1 0 55200 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1034
timestamp 1649977179
transform 1 0 60352 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1035
timestamp 1649977179
transform 1 0 65504 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1036
timestamp 1649977179
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1037
timestamp 1649977179
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1038
timestamp 1649977179
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1039
timestamp 1649977179
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1040
timestamp 1649977179
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1041
timestamp 1649977179
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1042
timestamp 1649977179
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1043
timestamp 1649977179
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1044
timestamp 1649977179
transform 1 0 47472 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1045
timestamp 1649977179
transform 1 0 52624 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1046
timestamp 1649977179
transform 1 0 57776 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1047
timestamp 1649977179
transform 1 0 62928 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1048
timestamp 1649977179
transform 1 0 68080 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1049
timestamp 1649977179
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1050
timestamp 1649977179
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1051
timestamp 1649977179
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1052
timestamp 1649977179
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1053
timestamp 1649977179
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1054
timestamp 1649977179
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1055
timestamp 1649977179
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1056
timestamp 1649977179
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1057
timestamp 1649977179
transform 1 0 44896 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1058
timestamp 1649977179
transform 1 0 50048 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1059
timestamp 1649977179
transform 1 0 55200 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1060
timestamp 1649977179
transform 1 0 60352 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1061
timestamp 1649977179
transform 1 0 65504 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1062
timestamp 1649977179
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1063
timestamp 1649977179
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1064
timestamp 1649977179
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1065
timestamp 1649977179
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1066
timestamp 1649977179
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1067
timestamp 1649977179
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1068
timestamp 1649977179
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1069
timestamp 1649977179
transform 1 0 42320 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1070
timestamp 1649977179
transform 1 0 47472 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1071
timestamp 1649977179
transform 1 0 52624 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1072
timestamp 1649977179
transform 1 0 57776 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1073
timestamp 1649977179
transform 1 0 62928 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1074
timestamp 1649977179
transform 1 0 68080 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1075
timestamp 1649977179
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1076
timestamp 1649977179
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1077
timestamp 1649977179
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1078
timestamp 1649977179
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1079
timestamp 1649977179
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1080
timestamp 1649977179
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1081
timestamp 1649977179
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1082
timestamp 1649977179
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1083
timestamp 1649977179
transform 1 0 44896 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1084
timestamp 1649977179
transform 1 0 50048 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1085
timestamp 1649977179
transform 1 0 55200 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1086
timestamp 1649977179
transform 1 0 60352 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1087
timestamp 1649977179
transform 1 0 65504 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1088
timestamp 1649977179
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1089
timestamp 1649977179
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1090
timestamp 1649977179
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1091
timestamp 1649977179
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1092
timestamp 1649977179
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1093
timestamp 1649977179
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1094
timestamp 1649977179
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1095
timestamp 1649977179
transform 1 0 42320 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1096
timestamp 1649977179
transform 1 0 47472 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1097
timestamp 1649977179
transform 1 0 52624 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1098
timestamp 1649977179
transform 1 0 57776 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1099
timestamp 1649977179
transform 1 0 62928 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1100
timestamp 1649977179
transform 1 0 68080 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1101
timestamp 1649977179
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1102
timestamp 1649977179
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1103
timestamp 1649977179
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1104
timestamp 1649977179
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1105
timestamp 1649977179
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1106
timestamp 1649977179
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1107
timestamp 1649977179
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1108
timestamp 1649977179
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1109
timestamp 1649977179
transform 1 0 44896 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1110
timestamp 1649977179
transform 1 0 50048 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1111
timestamp 1649977179
transform 1 0 55200 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1112
timestamp 1649977179
transform 1 0 60352 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1113
timestamp 1649977179
transform 1 0 65504 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1114
timestamp 1649977179
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1115
timestamp 1649977179
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1116
timestamp 1649977179
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1117
timestamp 1649977179
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1118
timestamp 1649977179
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1119
timestamp 1649977179
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1120
timestamp 1649977179
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1121
timestamp 1649977179
transform 1 0 42320 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1122
timestamp 1649977179
transform 1 0 47472 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1123
timestamp 1649977179
transform 1 0 52624 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1124
timestamp 1649977179
transform 1 0 57776 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1125
timestamp 1649977179
transform 1 0 62928 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1126
timestamp 1649977179
transform 1 0 68080 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1127
timestamp 1649977179
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1128
timestamp 1649977179
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1129
timestamp 1649977179
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1130
timestamp 1649977179
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1131
timestamp 1649977179
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1132
timestamp 1649977179
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1133
timestamp 1649977179
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1134
timestamp 1649977179
transform 1 0 39744 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1135
timestamp 1649977179
transform 1 0 44896 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1136
timestamp 1649977179
transform 1 0 50048 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1137
timestamp 1649977179
transform 1 0 55200 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1138
timestamp 1649977179
transform 1 0 60352 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1139
timestamp 1649977179
transform 1 0 65504 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1140
timestamp 1649977179
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1141
timestamp 1649977179
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1142
timestamp 1649977179
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1143
timestamp 1649977179
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1144
timestamp 1649977179
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1145
timestamp 1649977179
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1146
timestamp 1649977179
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1147
timestamp 1649977179
transform 1 0 42320 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1148
timestamp 1649977179
transform 1 0 47472 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1149
timestamp 1649977179
transform 1 0 52624 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1150
timestamp 1649977179
transform 1 0 57776 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1151
timestamp 1649977179
transform 1 0 62928 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1152
timestamp 1649977179
transform 1 0 68080 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1153
timestamp 1649977179
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1154
timestamp 1649977179
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1155
timestamp 1649977179
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1156
timestamp 1649977179
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1157
timestamp 1649977179
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1158
timestamp 1649977179
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1159
timestamp 1649977179
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1160
timestamp 1649977179
transform 1 0 39744 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1161
timestamp 1649977179
transform 1 0 44896 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1162
timestamp 1649977179
transform 1 0 50048 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1163
timestamp 1649977179
transform 1 0 55200 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1164
timestamp 1649977179
transform 1 0 60352 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1165
timestamp 1649977179
transform 1 0 65504 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1166
timestamp 1649977179
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1167
timestamp 1649977179
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1168
timestamp 1649977179
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1169
timestamp 1649977179
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1170
timestamp 1649977179
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1171
timestamp 1649977179
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1172
timestamp 1649977179
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1173
timestamp 1649977179
transform 1 0 42320 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1174
timestamp 1649977179
transform 1 0 47472 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1175
timestamp 1649977179
transform 1 0 52624 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1176
timestamp 1649977179
transform 1 0 57776 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1177
timestamp 1649977179
transform 1 0 62928 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1178
timestamp 1649977179
transform 1 0 68080 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1179
timestamp 1649977179
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1180
timestamp 1649977179
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1181
timestamp 1649977179
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1182
timestamp 1649977179
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1183
timestamp 1649977179
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1184
timestamp 1649977179
transform 1 0 29440 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1185
timestamp 1649977179
transform 1 0 34592 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1186
timestamp 1649977179
transform 1 0 39744 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1187
timestamp 1649977179
transform 1 0 44896 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1188
timestamp 1649977179
transform 1 0 50048 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1189
timestamp 1649977179
transform 1 0 55200 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1190
timestamp 1649977179
transform 1 0 60352 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1191
timestamp 1649977179
transform 1 0 65504 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1192
timestamp 1649977179
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1193
timestamp 1649977179
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1194
timestamp 1649977179
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1195
timestamp 1649977179
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1196
timestamp 1649977179
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1197
timestamp 1649977179
transform 1 0 32016 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1198
timestamp 1649977179
transform 1 0 37168 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1199
timestamp 1649977179
transform 1 0 42320 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1200
timestamp 1649977179
transform 1 0 47472 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1201
timestamp 1649977179
transform 1 0 52624 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1202
timestamp 1649977179
transform 1 0 57776 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1203
timestamp 1649977179
transform 1 0 62928 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1204
timestamp 1649977179
transform 1 0 68080 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1205
timestamp 1649977179
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1206
timestamp 1649977179
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1207
timestamp 1649977179
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1208
timestamp 1649977179
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1209
timestamp 1649977179
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1210
timestamp 1649977179
transform 1 0 29440 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1211
timestamp 1649977179
transform 1 0 34592 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1212
timestamp 1649977179
transform 1 0 39744 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1213
timestamp 1649977179
transform 1 0 44896 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1214
timestamp 1649977179
transform 1 0 50048 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1215
timestamp 1649977179
transform 1 0 55200 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1216
timestamp 1649977179
transform 1 0 60352 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1217
timestamp 1649977179
transform 1 0 65504 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1218
timestamp 1649977179
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1219
timestamp 1649977179
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1220
timestamp 1649977179
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1221
timestamp 1649977179
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1222
timestamp 1649977179
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1223
timestamp 1649977179
transform 1 0 32016 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1224
timestamp 1649977179
transform 1 0 37168 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1225
timestamp 1649977179
transform 1 0 42320 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1226
timestamp 1649977179
transform 1 0 47472 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1227
timestamp 1649977179
transform 1 0 52624 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1228
timestamp 1649977179
transform 1 0 57776 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1229
timestamp 1649977179
transform 1 0 62928 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1230
timestamp 1649977179
transform 1 0 68080 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1231
timestamp 1649977179
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1232
timestamp 1649977179
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1233
timestamp 1649977179
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1234
timestamp 1649977179
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1235
timestamp 1649977179
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1236
timestamp 1649977179
transform 1 0 29440 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1237
timestamp 1649977179
transform 1 0 34592 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1238
timestamp 1649977179
transform 1 0 39744 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1239
timestamp 1649977179
transform 1 0 44896 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1240
timestamp 1649977179
transform 1 0 50048 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1241
timestamp 1649977179
transform 1 0 55200 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1242
timestamp 1649977179
transform 1 0 60352 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1243
timestamp 1649977179
transform 1 0 65504 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1244
timestamp 1649977179
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1245
timestamp 1649977179
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1246
timestamp 1649977179
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1247
timestamp 1649977179
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1248
timestamp 1649977179
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1249
timestamp 1649977179
transform 1 0 32016 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1250
timestamp 1649977179
transform 1 0 37168 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1251
timestamp 1649977179
transform 1 0 42320 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1252
timestamp 1649977179
transform 1 0 47472 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1253
timestamp 1649977179
transform 1 0 52624 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1254
timestamp 1649977179
transform 1 0 57776 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1255
timestamp 1649977179
transform 1 0 62928 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1256
timestamp 1649977179
transform 1 0 68080 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1257
timestamp 1649977179
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1258
timestamp 1649977179
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1259
timestamp 1649977179
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1260
timestamp 1649977179
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1261
timestamp 1649977179
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1262
timestamp 1649977179
transform 1 0 29440 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1263
timestamp 1649977179
transform 1 0 34592 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1264
timestamp 1649977179
transform 1 0 39744 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1265
timestamp 1649977179
transform 1 0 44896 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1266
timestamp 1649977179
transform 1 0 50048 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1267
timestamp 1649977179
transform 1 0 55200 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1268
timestamp 1649977179
transform 1 0 60352 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1269
timestamp 1649977179
transform 1 0 65504 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1270
timestamp 1649977179
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1271
timestamp 1649977179
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1272
timestamp 1649977179
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1273
timestamp 1649977179
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1274
timestamp 1649977179
transform 1 0 26864 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1275
timestamp 1649977179
transform 1 0 32016 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1276
timestamp 1649977179
transform 1 0 37168 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1277
timestamp 1649977179
transform 1 0 42320 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1278
timestamp 1649977179
transform 1 0 47472 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1279
timestamp 1649977179
transform 1 0 52624 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1280
timestamp 1649977179
transform 1 0 57776 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1281
timestamp 1649977179
transform 1 0 62928 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1282
timestamp 1649977179
transform 1 0 68080 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1283
timestamp 1649977179
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1284
timestamp 1649977179
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1285
timestamp 1649977179
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1286
timestamp 1649977179
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1287
timestamp 1649977179
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1288
timestamp 1649977179
transform 1 0 29440 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1289
timestamp 1649977179
transform 1 0 34592 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1290
timestamp 1649977179
transform 1 0 39744 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1291
timestamp 1649977179
transform 1 0 44896 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1292
timestamp 1649977179
transform 1 0 50048 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1293
timestamp 1649977179
transform 1 0 55200 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1294
timestamp 1649977179
transform 1 0 60352 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1295
timestamp 1649977179
transform 1 0 65504 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1296
timestamp 1649977179
transform 1 0 6256 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1297
timestamp 1649977179
transform 1 0 11408 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1298
timestamp 1649977179
transform 1 0 16560 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1299
timestamp 1649977179
transform 1 0 21712 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1300
timestamp 1649977179
transform 1 0 26864 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1301
timestamp 1649977179
transform 1 0 32016 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1302
timestamp 1649977179
transform 1 0 37168 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1303
timestamp 1649977179
transform 1 0 42320 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1304
timestamp 1649977179
transform 1 0 47472 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1305
timestamp 1649977179
transform 1 0 52624 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1306
timestamp 1649977179
transform 1 0 57776 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1307
timestamp 1649977179
transform 1 0 62928 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1308
timestamp 1649977179
transform 1 0 68080 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1309
timestamp 1649977179
transform 1 0 3680 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1310
timestamp 1649977179
transform 1 0 8832 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1311
timestamp 1649977179
transform 1 0 13984 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1312
timestamp 1649977179
transform 1 0 19136 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1313
timestamp 1649977179
transform 1 0 24288 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1314
timestamp 1649977179
transform 1 0 29440 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1315
timestamp 1649977179
transform 1 0 34592 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1316
timestamp 1649977179
transform 1 0 39744 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1317
timestamp 1649977179
transform 1 0 44896 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1318
timestamp 1649977179
transform 1 0 50048 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1319
timestamp 1649977179
transform 1 0 55200 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1320
timestamp 1649977179
transform 1 0 60352 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1321
timestamp 1649977179
transform 1 0 65504 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1322
timestamp 1649977179
transform 1 0 6256 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1323
timestamp 1649977179
transform 1 0 11408 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1324
timestamp 1649977179
transform 1 0 16560 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1325
timestamp 1649977179
transform 1 0 21712 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1326
timestamp 1649977179
transform 1 0 26864 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1327
timestamp 1649977179
transform 1 0 32016 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1328
timestamp 1649977179
transform 1 0 37168 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1329
timestamp 1649977179
transform 1 0 42320 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1330
timestamp 1649977179
transform 1 0 47472 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1331
timestamp 1649977179
transform 1 0 52624 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1332
timestamp 1649977179
transform 1 0 57776 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1333
timestamp 1649977179
transform 1 0 62928 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1334
timestamp 1649977179
transform 1 0 68080 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1335
timestamp 1649977179
transform 1 0 3680 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1336
timestamp 1649977179
transform 1 0 8832 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1337
timestamp 1649977179
transform 1 0 13984 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1338
timestamp 1649977179
transform 1 0 19136 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1339
timestamp 1649977179
transform 1 0 24288 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1340
timestamp 1649977179
transform 1 0 29440 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1341
timestamp 1649977179
transform 1 0 34592 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1342
timestamp 1649977179
transform 1 0 39744 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1343
timestamp 1649977179
transform 1 0 44896 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1344
timestamp 1649977179
transform 1 0 50048 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1345
timestamp 1649977179
transform 1 0 55200 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1346
timestamp 1649977179
transform 1 0 60352 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1347
timestamp 1649977179
transform 1 0 65504 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1348
timestamp 1649977179
transform 1 0 6256 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1349
timestamp 1649977179
transform 1 0 11408 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1350
timestamp 1649977179
transform 1 0 16560 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1351
timestamp 1649977179
transform 1 0 21712 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1352
timestamp 1649977179
transform 1 0 26864 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1353
timestamp 1649977179
transform 1 0 32016 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1354
timestamp 1649977179
transform 1 0 37168 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1355
timestamp 1649977179
transform 1 0 42320 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1356
timestamp 1649977179
transform 1 0 47472 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1357
timestamp 1649977179
transform 1 0 52624 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1358
timestamp 1649977179
transform 1 0 57776 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1359
timestamp 1649977179
transform 1 0 62928 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1360
timestamp 1649977179
transform 1 0 68080 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1361
timestamp 1649977179
transform 1 0 3680 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1362
timestamp 1649977179
transform 1 0 8832 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1363
timestamp 1649977179
transform 1 0 13984 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1364
timestamp 1649977179
transform 1 0 19136 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1365
timestamp 1649977179
transform 1 0 24288 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1366
timestamp 1649977179
transform 1 0 29440 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1367
timestamp 1649977179
transform 1 0 34592 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1368
timestamp 1649977179
transform 1 0 39744 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1369
timestamp 1649977179
transform 1 0 44896 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1370
timestamp 1649977179
transform 1 0 50048 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1371
timestamp 1649977179
transform 1 0 55200 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1372
timestamp 1649977179
transform 1 0 60352 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1373
timestamp 1649977179
transform 1 0 65504 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1374
timestamp 1649977179
transform 1 0 6256 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1375
timestamp 1649977179
transform 1 0 11408 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1376
timestamp 1649977179
transform 1 0 16560 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1377
timestamp 1649977179
transform 1 0 21712 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1378
timestamp 1649977179
transform 1 0 26864 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1379
timestamp 1649977179
transform 1 0 32016 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1380
timestamp 1649977179
transform 1 0 37168 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1381
timestamp 1649977179
transform 1 0 42320 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1382
timestamp 1649977179
transform 1 0 47472 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1383
timestamp 1649977179
transform 1 0 52624 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1384
timestamp 1649977179
transform 1 0 57776 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1385
timestamp 1649977179
transform 1 0 62928 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1386
timestamp 1649977179
transform 1 0 68080 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1387
timestamp 1649977179
transform 1 0 3680 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1388
timestamp 1649977179
transform 1 0 8832 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1389
timestamp 1649977179
transform 1 0 13984 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1390
timestamp 1649977179
transform 1 0 19136 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1391
timestamp 1649977179
transform 1 0 24288 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1392
timestamp 1649977179
transform 1 0 29440 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1393
timestamp 1649977179
transform 1 0 34592 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1394
timestamp 1649977179
transform 1 0 39744 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1395
timestamp 1649977179
transform 1 0 44896 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1396
timestamp 1649977179
transform 1 0 50048 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1397
timestamp 1649977179
transform 1 0 55200 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1398
timestamp 1649977179
transform 1 0 60352 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1399
timestamp 1649977179
transform 1 0 65504 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1400
timestamp 1649977179
transform 1 0 6256 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1401
timestamp 1649977179
transform 1 0 11408 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1402
timestamp 1649977179
transform 1 0 16560 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1403
timestamp 1649977179
transform 1 0 21712 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1404
timestamp 1649977179
transform 1 0 26864 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1405
timestamp 1649977179
transform 1 0 32016 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1406
timestamp 1649977179
transform 1 0 37168 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1407
timestamp 1649977179
transform 1 0 42320 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1408
timestamp 1649977179
transform 1 0 47472 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1409
timestamp 1649977179
transform 1 0 52624 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1410
timestamp 1649977179
transform 1 0 57776 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1411
timestamp 1649977179
transform 1 0 62928 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1412
timestamp 1649977179
transform 1 0 68080 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1413
timestamp 1649977179
transform 1 0 3680 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1414
timestamp 1649977179
transform 1 0 8832 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1415
timestamp 1649977179
transform 1 0 13984 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1416
timestamp 1649977179
transform 1 0 19136 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1417
timestamp 1649977179
transform 1 0 24288 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1418
timestamp 1649977179
transform 1 0 29440 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1419
timestamp 1649977179
transform 1 0 34592 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1420
timestamp 1649977179
transform 1 0 39744 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1421
timestamp 1649977179
transform 1 0 44896 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1422
timestamp 1649977179
transform 1 0 50048 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1423
timestamp 1649977179
transform 1 0 55200 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1424
timestamp 1649977179
transform 1 0 60352 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1425
timestamp 1649977179
transform 1 0 65504 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1426
timestamp 1649977179
transform 1 0 6256 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1427
timestamp 1649977179
transform 1 0 11408 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1428
timestamp 1649977179
transform 1 0 16560 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1429
timestamp 1649977179
transform 1 0 21712 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1430
timestamp 1649977179
transform 1 0 26864 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1431
timestamp 1649977179
transform 1 0 32016 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1432
timestamp 1649977179
transform 1 0 37168 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1433
timestamp 1649977179
transform 1 0 42320 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1434
timestamp 1649977179
transform 1 0 47472 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1435
timestamp 1649977179
transform 1 0 52624 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1436
timestamp 1649977179
transform 1 0 57776 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1437
timestamp 1649977179
transform 1 0 62928 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1438
timestamp 1649977179
transform 1 0 68080 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1439
timestamp 1649977179
transform 1 0 3680 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1440
timestamp 1649977179
transform 1 0 8832 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1441
timestamp 1649977179
transform 1 0 13984 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1442
timestamp 1649977179
transform 1 0 19136 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1443
timestamp 1649977179
transform 1 0 24288 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1444
timestamp 1649977179
transform 1 0 29440 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1445
timestamp 1649977179
transform 1 0 34592 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1446
timestamp 1649977179
transform 1 0 39744 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1447
timestamp 1649977179
transform 1 0 44896 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1448
timestamp 1649977179
transform 1 0 50048 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1449
timestamp 1649977179
transform 1 0 55200 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1450
timestamp 1649977179
transform 1 0 60352 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1451
timestamp 1649977179
transform 1 0 65504 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1452
timestamp 1649977179
transform 1 0 6256 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1453
timestamp 1649977179
transform 1 0 11408 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1454
timestamp 1649977179
transform 1 0 16560 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1455
timestamp 1649977179
transform 1 0 21712 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1456
timestamp 1649977179
transform 1 0 26864 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1457
timestamp 1649977179
transform 1 0 32016 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1458
timestamp 1649977179
transform 1 0 37168 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1459
timestamp 1649977179
transform 1 0 42320 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1460
timestamp 1649977179
transform 1 0 47472 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1461
timestamp 1649977179
transform 1 0 52624 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1462
timestamp 1649977179
transform 1 0 57776 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1463
timestamp 1649977179
transform 1 0 62928 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1464
timestamp 1649977179
transform 1 0 68080 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1465
timestamp 1649977179
transform 1 0 3680 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1466
timestamp 1649977179
transform 1 0 8832 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1467
timestamp 1649977179
transform 1 0 13984 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1468
timestamp 1649977179
transform 1 0 19136 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1469
timestamp 1649977179
transform 1 0 24288 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1470
timestamp 1649977179
transform 1 0 29440 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1471
timestamp 1649977179
transform 1 0 34592 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1472
timestamp 1649977179
transform 1 0 39744 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1473
timestamp 1649977179
transform 1 0 44896 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1474
timestamp 1649977179
transform 1 0 50048 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1475
timestamp 1649977179
transform 1 0 55200 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1476
timestamp 1649977179
transform 1 0 60352 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1477
timestamp 1649977179
transform 1 0 65504 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1478
timestamp 1649977179
transform 1 0 6256 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1479
timestamp 1649977179
transform 1 0 11408 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1480
timestamp 1649977179
transform 1 0 16560 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1481
timestamp 1649977179
transform 1 0 21712 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1482
timestamp 1649977179
transform 1 0 26864 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1483
timestamp 1649977179
transform 1 0 32016 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1484
timestamp 1649977179
transform 1 0 37168 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1485
timestamp 1649977179
transform 1 0 42320 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1486
timestamp 1649977179
transform 1 0 47472 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1487
timestamp 1649977179
transform 1 0 52624 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1488
timestamp 1649977179
transform 1 0 57776 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1489
timestamp 1649977179
transform 1 0 62928 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1490
timestamp 1649977179
transform 1 0 68080 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1491
timestamp 1649977179
transform 1 0 3680 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1492
timestamp 1649977179
transform 1 0 8832 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1493
timestamp 1649977179
transform 1 0 13984 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1494
timestamp 1649977179
transform 1 0 19136 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1495
timestamp 1649977179
transform 1 0 24288 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1496
timestamp 1649977179
transform 1 0 29440 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1497
timestamp 1649977179
transform 1 0 34592 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1498
timestamp 1649977179
transform 1 0 39744 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1499
timestamp 1649977179
transform 1 0 44896 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1500
timestamp 1649977179
transform 1 0 50048 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1501
timestamp 1649977179
transform 1 0 55200 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1502
timestamp 1649977179
transform 1 0 60352 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1503
timestamp 1649977179
transform 1 0 65504 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1504
timestamp 1649977179
transform 1 0 6256 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1505
timestamp 1649977179
transform 1 0 11408 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1506
timestamp 1649977179
transform 1 0 16560 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1507
timestamp 1649977179
transform 1 0 21712 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1508
timestamp 1649977179
transform 1 0 26864 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1509
timestamp 1649977179
transform 1 0 32016 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1510
timestamp 1649977179
transform 1 0 37168 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1511
timestamp 1649977179
transform 1 0 42320 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1512
timestamp 1649977179
transform 1 0 47472 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1513
timestamp 1649977179
transform 1 0 52624 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1514
timestamp 1649977179
transform 1 0 57776 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1515
timestamp 1649977179
transform 1 0 62928 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1516
timestamp 1649977179
transform 1 0 68080 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1517
timestamp 1649977179
transform 1 0 3680 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1518
timestamp 1649977179
transform 1 0 8832 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1519
timestamp 1649977179
transform 1 0 13984 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1520
timestamp 1649977179
transform 1 0 19136 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1521
timestamp 1649977179
transform 1 0 24288 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1522
timestamp 1649977179
transform 1 0 29440 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1523
timestamp 1649977179
transform 1 0 34592 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1524
timestamp 1649977179
transform 1 0 39744 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1525
timestamp 1649977179
transform 1 0 44896 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1526
timestamp 1649977179
transform 1 0 50048 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1527
timestamp 1649977179
transform 1 0 55200 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1528
timestamp 1649977179
transform 1 0 60352 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1529
timestamp 1649977179
transform 1 0 65504 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1530
timestamp 1649977179
transform 1 0 3680 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1531
timestamp 1649977179
transform 1 0 6256 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1532
timestamp 1649977179
transform 1 0 8832 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1533
timestamp 1649977179
transform 1 0 11408 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1534
timestamp 1649977179
transform 1 0 13984 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1535
timestamp 1649977179
transform 1 0 16560 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1536
timestamp 1649977179
transform 1 0 19136 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1537
timestamp 1649977179
transform 1 0 21712 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1538
timestamp 1649977179
transform 1 0 24288 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1539
timestamp 1649977179
transform 1 0 26864 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1540
timestamp 1649977179
transform 1 0 29440 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1541
timestamp 1649977179
transform 1 0 32016 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1542
timestamp 1649977179
transform 1 0 34592 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1543
timestamp 1649977179
transform 1 0 37168 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1544
timestamp 1649977179
transform 1 0 39744 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1545
timestamp 1649977179
transform 1 0 42320 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1546
timestamp 1649977179
transform 1 0 44896 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1547
timestamp 1649977179
transform 1 0 47472 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1548
timestamp 1649977179
transform 1 0 50048 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1549
timestamp 1649977179
transform 1 0 52624 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1550
timestamp 1649977179
transform 1 0 55200 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1551
timestamp 1649977179
transform 1 0 57776 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1552
timestamp 1649977179
transform 1 0 60352 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1553
timestamp 1649977179
transform 1 0 62928 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1554
timestamp 1649977179
transform 1 0 65504 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1555
timestamp 1649977179
transform 1 0 68080 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__and2b_1  _0761_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 34868 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0762_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 35604 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0763_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 2484 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0764_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1932 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0765_
timestamp 1649977179
transform -1 0 7912 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0766_
timestamp 1649977179
transform 1 0 7268 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0767_
timestamp 1649977179
transform -1 0 24564 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0768_
timestamp 1649977179
transform -1 0 24656 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0769_
timestamp 1649977179
transform 1 0 36892 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0770_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 36432 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0771_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 37536 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0772_
timestamp 1649977179
transform 1 0 41124 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0773_
timestamp 1649977179
transform 1 0 42412 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0774_
timestamp 1649977179
transform 1 0 43240 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0775_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 2392 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0776_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 3128 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0777_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0778_
timestamp 1649977179
transform -1 0 12328 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0779_
timestamp 1649977179
transform -1 0 2576 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__o2bb2a_1  _0780_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0781_
timestamp 1649977179
transform 1 0 1748 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0782_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 2024 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0783_
timestamp 1649977179
transform 1 0 1380 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0784_
timestamp 1649977179
transform -1 0 5428 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0785_
timestamp 1649977179
transform -1 0 9568 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0786_
timestamp 1649977179
transform -1 0 7360 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o22ai_1  _0787_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 6992 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0788_
timestamp 1649977179
transform -1 0 11592 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _0789_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 6532 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0790_
timestamp 1649977179
transform 1 0 5980 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0791_
timestamp 1649977179
transform -1 0 3128 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _0792_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1472 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _0793_
timestamp 1649977179
transform 1 0 9200 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0794_
timestamp 1649977179
transform -1 0 13432 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _0795_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 18124 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _0796_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 8464 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _0797_
timestamp 1649977179
transform 1 0 7360 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _0798_
timestamp 1649977179
transform 1 0 6072 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0799_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 9292 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0800_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 11868 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0801_
timestamp 1649977179
transform 1 0 11500 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0802_
timestamp 1649977179
transform -1 0 10856 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0803_
timestamp 1649977179
transform -1 0 8464 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _0804_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 7728 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0805_
timestamp 1649977179
transform 1 0 7912 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a2111oi_1  _0806_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 8924 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0807_
timestamp 1649977179
transform -1 0 8188 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0808_
timestamp 1649977179
transform 1 0 1472 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0809_
timestamp 1649977179
transform 1 0 1840 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__o22ai_1  _0810_
timestamp 1649977179
transform 1 0 10672 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a2111oi_1  _0811_
timestamp 1649977179
transform -1 0 10304 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _0812_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 9292 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0813_
timestamp 1649977179
transform -1 0 5704 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0814_
timestamp 1649977179
transform 1 0 15364 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0815_
timestamp 1649977179
transform 1 0 20148 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0816_
timestamp 1649977179
transform 1 0 21896 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0817_
timestamp 1649977179
transform -1 0 23828 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0818_
timestamp 1649977179
transform 1 0 23460 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__o2bb2a_1  _0819_
timestamp 1649977179
transform -1 0 23920 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0820_
timestamp 1649977179
transform 1 0 19688 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0821_
timestamp 1649977179
transform -1 0 19596 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0822_
timestamp 1649977179
transform 1 0 16468 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0823_
timestamp 1649977179
transform -1 0 15824 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0824_
timestamp 1649977179
transform 1 0 18768 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0825_
timestamp 1649977179
transform 1 0 15732 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0826_
timestamp 1649977179
transform 1 0 15548 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0827_
timestamp 1649977179
transform 1 0 17664 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0828_
timestamp 1649977179
transform 1 0 17756 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _0829_
timestamp 1649977179
transform 1 0 17664 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0830_
timestamp 1649977179
transform 1 0 17112 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0831_
timestamp 1649977179
transform 1 0 17756 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _0832_
timestamp 1649977179
transform -1 0 21344 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0833_
timestamp 1649977179
transform 1 0 29900 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0834_
timestamp 1649977179
transform 1 0 30268 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0835_
timestamp 1649977179
transform -1 0 33212 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0836_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 33672 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _0837_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 32844 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0838_
timestamp 1649977179
transform 1 0 32384 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0839_
timestamp 1649977179
transform 1 0 33028 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0840_
timestamp 1649977179
transform 1 0 33948 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0841_
timestamp 1649977179
transform 1 0 27692 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0842_
timestamp 1649977179
transform -1 0 29072 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _0843_
timestamp 1649977179
transform -1 0 30176 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0844_
timestamp 1649977179
transform 1 0 27600 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0845_
timestamp 1649977179
transform 1 0 31004 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0846_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 29716 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a2111o_1  _0847_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 30176 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _0848_
timestamp 1649977179
transform 1 0 30544 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0849_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 34684 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0850_
timestamp 1649977179
transform 1 0 24472 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0851_
timestamp 1649977179
transform 1 0 28336 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0852_
timestamp 1649977179
transform 1 0 30176 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0853_
timestamp 1649977179
transform 1 0 31648 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0854_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 33764 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0855_
timestamp 1649977179
transform -1 0 34960 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0856_
timestamp 1649977179
transform 1 0 26956 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0857_
timestamp 1649977179
transform 1 0 28796 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0858_
timestamp 1649977179
transform 1 0 29716 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0859_
timestamp 1649977179
transform 1 0 30452 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0860_
timestamp 1649977179
transform 1 0 31004 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0861_
timestamp 1649977179
transform -1 0 34224 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0862_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 32568 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _0863_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 33120 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0864_
timestamp 1649977179
transform 1 0 31464 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0865_
timestamp 1649977179
transform 1 0 31832 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _0866_
timestamp 1649977179
transform 1 0 34684 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0867_
timestamp 1649977179
transform 1 0 35696 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0868_
timestamp 1649977179
transform 1 0 35696 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0869_
timestamp 1649977179
transform 1 0 40112 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0870_
timestamp 1649977179
transform 1 0 41216 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0871_
timestamp 1649977179
transform -1 0 42872 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0872_
timestamp 1649977179
transform -1 0 42320 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0873_
timestamp 1649977179
transform 1 0 37444 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0874_
timestamp 1649977179
transform 1 0 37536 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0875_
timestamp 1649977179
transform 1 0 38272 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0876_
timestamp 1649977179
transform 1 0 40572 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0877_
timestamp 1649977179
transform 1 0 41216 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0878_
timestamp 1649977179
transform 1 0 41216 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0879_
timestamp 1649977179
transform 1 0 41308 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _0880_
timestamp 1649977179
transform 1 0 41216 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0881_
timestamp 1649977179
transform 1 0 40848 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0882_
timestamp 1649977179
transform 1 0 42412 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _0883_
timestamp 1649977179
transform -1 0 43148 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0884_
timestamp 1649977179
transform 1 0 36248 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0885_
timestamp 1649977179
transform 1 0 36248 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0886_
timestamp 1649977179
transform 1 0 41676 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0887_
timestamp 1649977179
transform -1 0 41952 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0888_
timestamp 1649977179
transform 1 0 34960 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0889_
timestamp 1649977179
transform -1 0 35604 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0890_
timestamp 1649977179
transform 1 0 24932 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0891_
timestamp 1649977179
transform -1 0 25852 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0892_
timestamp 1649977179
transform 1 0 6532 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0893_
timestamp 1649977179
transform 1 0 6716 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0894_
timestamp 1649977179
transform -1 0 2668 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0895_
timestamp 1649977179
transform 1 0 2116 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nor4_2  _0896_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 20148 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__nor4_2  _0897_
timestamp 1649977179
transform -1 0 17204 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _0898_
timestamp 1649977179
transform -1 0 19688 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and4bb_1  _0899_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 20148 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _0900_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 11868 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0901_
timestamp 1649977179
transform 1 0 11408 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0902_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 12604 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0903_
timestamp 1649977179
transform 1 0 12696 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _0904_
timestamp 1649977179
transform -1 0 10212 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0905_
timestamp 1649977179
transform -1 0 6808 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _0906_
timestamp 1649977179
transform -1 0 10488 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0907_
timestamp 1649977179
transform 1 0 6440 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0908_
timestamp 1649977179
transform 1 0 1748 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0909_
timestamp 1649977179
transform 1 0 22540 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0910_
timestamp 1649977179
transform -1 0 22080 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0911_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 20976 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _0912_
timestamp 1649977179
transform -1 0 2484 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0913_
timestamp 1649977179
transform -1 0 3036 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0914_
timestamp 1649977179
transform 1 0 1840 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0915_
timestamp 1649977179
transform 1 0 1840 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0916_
timestamp 1649977179
transform 1 0 1656 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0917_
timestamp 1649977179
transform 1 0 1748 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0918_
timestamp 1649977179
transform 1 0 1840 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0919_
timestamp 1649977179
transform 1 0 5428 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0920_
timestamp 1649977179
transform -1 0 14996 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0921_
timestamp 1649977179
transform -1 0 11500 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _0922_
timestamp 1649977179
transform 1 0 5152 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0923_
timestamp 1649977179
transform -1 0 9844 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _0924_
timestamp 1649977179
transform -1 0 7084 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0925_
timestamp 1649977179
transform 1 0 11500 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0926_
timestamp 1649977179
transform -1 0 12604 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0927_
timestamp 1649977179
transform 1 0 10580 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0928_
timestamp 1649977179
transform -1 0 12236 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0929_
timestamp 1649977179
transform 1 0 7728 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0930_
timestamp 1649977179
transform -1 0 8464 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0931_
timestamp 1649977179
transform 1 0 11316 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0932_
timestamp 1649977179
transform -1 0 12880 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0933_
timestamp 1649977179
transform 1 0 10856 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0934_
timestamp 1649977179
transform 1 0 11500 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _0935_
timestamp 1649977179
transform -1 0 12420 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0936_
timestamp 1649977179
transform -1 0 10028 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0937_
timestamp 1649977179
transform -1 0 10304 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0938_
timestamp 1649977179
transform -1 0 12604 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__nor4b_2  _0939_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 20240 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_1  _0940_
timestamp 1649977179
transform -1 0 19688 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0941_
timestamp 1649977179
transform 1 0 16744 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0942_
timestamp 1649977179
transform -1 0 13708 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _0943_
timestamp 1649977179
transform -1 0 12052 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0944_
timestamp 1649977179
transform 1 0 5612 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _0945_
timestamp 1649977179
transform 1 0 5612 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0946_
timestamp 1649977179
transform -1 0 6164 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0947_
timestamp 1649977179
transform 1 0 1748 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0948_
timestamp 1649977179
transform -1 0 12420 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0949_
timestamp 1649977179
transform 1 0 5612 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0950_
timestamp 1649977179
transform -1 0 2576 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0951_
timestamp 1649977179
transform -1 0 3220 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0952_
timestamp 1649977179
transform 1 0 2484 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0953_
timestamp 1649977179
transform 1 0 2484 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0954_
timestamp 1649977179
transform -1 0 3220 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0955_
timestamp 1649977179
transform -1 0 17664 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0956_
timestamp 1649977179
transform 1 0 2944 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0957_
timestamp 1649977179
transform 1 0 11500 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _0958_
timestamp 1649977179
transform -1 0 3680 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0959_
timestamp 1649977179
transform -1 0 19596 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0960_
timestamp 1649977179
transform -1 0 4784 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0961_
timestamp 1649977179
transform 1 0 2484 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0962_
timestamp 1649977179
transform -1 0 21344 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0963_
timestamp 1649977179
transform -1 0 7728 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _0964_
timestamp 1649977179
transform 1 0 5428 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0965_
timestamp 1649977179
transform 1 0 6440 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0966_
timestamp 1649977179
transform -1 0 22172 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0967_
timestamp 1649977179
transform 1 0 11316 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0968_
timestamp 1649977179
transform -1 0 12328 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0969_
timestamp 1649977179
transform -1 0 16744 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0970_
timestamp 1649977179
transform 1 0 7452 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0971_
timestamp 1649977179
transform -1 0 8832 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0972_
timestamp 1649977179
transform -1 0 23828 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0973_
timestamp 1649977179
transform -1 0 9384 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0974_
timestamp 1649977179
transform -1 0 11040 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _0975_
timestamp 1649977179
transform -1 0 8096 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0976_
timestamp 1649977179
transform -1 0 22540 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0977_
timestamp 1649977179
transform 1 0 9936 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0978_
timestamp 1649977179
transform -1 0 10396 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0979_
timestamp 1649977179
transform -1 0 18768 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0980_
timestamp 1649977179
transform 1 0 10580 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0981_
timestamp 1649977179
transform -1 0 11776 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__nor4b_2  _0982_
timestamp 1649977179
transform 1 0 20240 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_1  _0983_
timestamp 1649977179
transform -1 0 21712 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0984_
timestamp 1649977179
transform -1 0 10396 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _0985_
timestamp 1649977179
transform 1 0 9384 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0986_
timestamp 1649977179
transform 1 0 8924 0 1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _0987_
timestamp 1649977179
transform -1 0 9200 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0988_
timestamp 1649977179
transform -1 0 9476 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0989_
timestamp 1649977179
transform -1 0 8648 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0990_
timestamp 1649977179
transform 1 0 6348 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0991_
timestamp 1649977179
transform 1 0 4784 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0992_
timestamp 1649977179
transform -1 0 5612 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0993_
timestamp 1649977179
transform -1 0 2576 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0994_
timestamp 1649977179
transform -1 0 17020 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0995_
timestamp 1649977179
transform -1 0 10212 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _0996_
timestamp 1649977179
transform 1 0 1840 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0997_
timestamp 1649977179
transform 1 0 2208 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0998_
timestamp 1649977179
transform -1 0 3128 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0999_
timestamp 1649977179
transform -1 0 6440 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1000_
timestamp 1649977179
transform 1 0 5152 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1001_
timestamp 1649977179
transform 1 0 8924 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1002_
timestamp 1649977179
transform 1 0 6348 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1003_
timestamp 1649977179
transform 1 0 6808 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1004_
timestamp 1649977179
transform 1 0 8372 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1005_
timestamp 1649977179
transform -1 0 9660 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1006_
timestamp 1649977179
transform 1 0 7268 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1007_
timestamp 1649977179
transform -1 0 9844 0 1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1008_
timestamp 1649977179
transform 1 0 7636 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1009_
timestamp 1649977179
transform -1 0 7636 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1010_
timestamp 1649977179
transform 1 0 6808 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1011_
timestamp 1649977179
transform 1 0 8188 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1012_
timestamp 1649977179
transform -1 0 9752 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1013_
timestamp 1649977179
transform 1 0 8004 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1014_
timestamp 1649977179
transform -1 0 10948 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1015_
timestamp 1649977179
transform 1 0 14076 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__and4bb_1  _1016_
timestamp 1649977179
transform 1 0 18952 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1017_
timestamp 1649977179
transform -1 0 20148 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1018_
timestamp 1649977179
transform 1 0 19320 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1019_
timestamp 1649977179
transform 1 0 18860 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1020_
timestamp 1649977179
transform -1 0 18124 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1021_
timestamp 1649977179
transform -1 0 13248 0 1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1022_
timestamp 1649977179
transform 1 0 16284 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1023_
timestamp 1649977179
transform -1 0 17112 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1024_
timestamp 1649977179
transform -1 0 13984 0 -1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1025_
timestamp 1649977179
transform -1 0 7452 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1026_
timestamp 1649977179
transform 1 0 6532 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1027_
timestamp 1649977179
transform 1 0 2392 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1028_
timestamp 1649977179
transform 1 0 10672 0 1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1029_
timestamp 1649977179
transform -1 0 3956 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1030_
timestamp 1649977179
transform -1 0 8648 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1031_
timestamp 1649977179
transform -1 0 8464 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1032_
timestamp 1649977179
transform -1 0 11960 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1033_
timestamp 1649977179
transform -1 0 11500 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1034_
timestamp 1649977179
transform 1 0 2300 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1035_
timestamp 1649977179
transform 1 0 3128 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1036_
timestamp 1649977179
transform -1 0 15180 0 1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1037_
timestamp 1649977179
transform -1 0 16928 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1038_
timestamp 1649977179
transform -1 0 13892 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1039_
timestamp 1649977179
transform -1 0 16284 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1040_
timestamp 1649977179
transform 1 0 16928 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1041_
timestamp 1649977179
transform -1 0 15732 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1042_
timestamp 1649977179
transform -1 0 17848 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1043_
timestamp 1649977179
transform 1 0 14352 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1044_
timestamp 1649977179
transform -1 0 15916 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1045_
timestamp 1649977179
transform 1 0 16192 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1046_
timestamp 1649977179
transform -1 0 17388 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1047_
timestamp 1649977179
transform 1 0 16468 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1048_
timestamp 1649977179
transform -1 0 18032 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1049_
timestamp 1649977179
transform 1 0 16652 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1050_
timestamp 1649977179
transform 1 0 15916 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__nor4b_4  _1051_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 17020 0 1 4352
box -38 -48 1786 592
use sky130_fd_sc_hd__and2_1  _1052_
timestamp 1649977179
transform 1 0 20148 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1053_
timestamp 1649977179
transform 1 0 21804 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1054_
timestamp 1649977179
transform -1 0 21160 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1055_
timestamp 1649977179
transform 1 0 19872 0 -1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1056_
timestamp 1649977179
transform 1 0 11960 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1057_
timestamp 1649977179
transform -1 0 21896 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1058_
timestamp 1649977179
transform 1 0 21068 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1059_
timestamp 1649977179
transform -1 0 15364 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1060_
timestamp 1649977179
transform -1 0 14996 0 1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1061_
timestamp 1649977179
transform -1 0 15088 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1062_
timestamp 1649977179
transform -1 0 14076 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1063_
timestamp 1649977179
transform 1 0 13432 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1064_
timestamp 1649977179
transform 1 0 19320 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1065_
timestamp 1649977179
transform -1 0 20608 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1066_
timestamp 1649977179
transform -1 0 18400 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1067_
timestamp 1649977179
transform 1 0 17480 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1068_
timestamp 1649977179
transform -1 0 21344 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1069_
timestamp 1649977179
transform -1 0 20516 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1070_
timestamp 1649977179
transform -1 0 21068 0 1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1071_
timestamp 1649977179
transform 1 0 21528 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1072_
timestamp 1649977179
transform 1 0 23460 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1073_
timestamp 1649977179
transform -1 0 20884 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1074_
timestamp 1649977179
transform -1 0 22724 0 1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1075_
timestamp 1649977179
transform -1 0 25208 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1076_
timestamp 1649977179
transform 1 0 23644 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1077_
timestamp 1649977179
transform -1 0 25024 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1078_
timestamp 1649977179
transform -1 0 20056 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1079_
timestamp 1649977179
transform -1 0 20884 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1080_
timestamp 1649977179
transform 1 0 23368 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1081_
timestamp 1649977179
transform -1 0 24932 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1082_
timestamp 1649977179
transform 1 0 21252 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1083_
timestamp 1649977179
transform -1 0 22540 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1084_
timestamp 1649977179
transform -1 0 23552 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1085_
timestamp 1649977179
transform -1 0 20056 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1086_
timestamp 1649977179
transform -1 0 20148 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1087_
timestamp 1649977179
transform -1 0 18584 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1088_
timestamp 1649977179
transform 1 0 15548 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1089_
timestamp 1649977179
transform 1 0 14720 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1090_
timestamp 1649977179
transform -1 0 15088 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1091_
timestamp 1649977179
transform -1 0 16376 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1092_
timestamp 1649977179
transform 1 0 15180 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1093_
timestamp 1649977179
transform 1 0 15456 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1094_
timestamp 1649977179
transform -1 0 15364 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1095_
timestamp 1649977179
transform -1 0 13248 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1096_
timestamp 1649977179
transform -1 0 14536 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1097_
timestamp 1649977179
transform -1 0 13616 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1098_
timestamp 1649977179
transform -1 0 12604 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1099_
timestamp 1649977179
transform 1 0 11776 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1100_
timestamp 1649977179
transform -1 0 12604 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1101_
timestamp 1649977179
transform 1 0 11500 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1102_
timestamp 1649977179
transform 1 0 14076 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1103_
timestamp 1649977179
transform 1 0 20148 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1104_
timestamp 1649977179
transform 1 0 14076 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1105_
timestamp 1649977179
transform 1 0 15916 0 1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1106_
timestamp 1649977179
transform -1 0 16284 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1107_
timestamp 1649977179
transform -1 0 15088 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1108_
timestamp 1649977179
transform 1 0 15456 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1109_
timestamp 1649977179
transform 1 0 19228 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1110_
timestamp 1649977179
transform -1 0 19504 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1111_
timestamp 1649977179
transform 1 0 17480 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1112_
timestamp 1649977179
transform -1 0 17664 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1113_
timestamp 1649977179
transform -1 0 16100 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1114_
timestamp 1649977179
transform -1 0 16192 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1115_
timestamp 1649977179
transform 1 0 18952 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1116_
timestamp 1649977179
transform 1 0 23184 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1117_
timestamp 1649977179
transform -1 0 19964 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1118_
timestamp 1649977179
transform 1 0 19228 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1119_
timestamp 1649977179
transform 1 0 19228 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1120_
timestamp 1649977179
transform 1 0 26220 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1121_
timestamp 1649977179
transform 1 0 21804 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1122_
timestamp 1649977179
transform -1 0 20976 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1123_
timestamp 1649977179
transform 1 0 20424 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1124_
timestamp 1649977179
transform 1 0 23000 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1125_
timestamp 1649977179
transform 1 0 24564 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1126_
timestamp 1649977179
transform 1 0 25300 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1127_
timestamp 1649977179
transform 1 0 22172 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1128_
timestamp 1649977179
transform -1 0 24656 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1129_
timestamp 1649977179
transform 1 0 24840 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1130_
timestamp 1649977179
transform 1 0 24840 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1131_
timestamp 1649977179
transform 1 0 26128 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1132_
timestamp 1649977179
transform 1 0 25576 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1133_
timestamp 1649977179
transform -1 0 26220 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1134_
timestamp 1649977179
transform 1 0 28152 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1135_
timestamp 1649977179
transform 1 0 25208 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1136_
timestamp 1649977179
transform -1 0 26220 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1137_
timestamp 1649977179
transform 1 0 23644 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1138_
timestamp 1649977179
transform 1 0 24380 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1139_
timestamp 1649977179
transform 1 0 24748 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1140_
timestamp 1649977179
transform 1 0 24380 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1141_
timestamp 1649977179
transform 1 0 23276 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1142_
timestamp 1649977179
transform 1 0 25392 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1143_
timestamp 1649977179
transform -1 0 26220 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1144_
timestamp 1649977179
transform 1 0 28520 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1145_
timestamp 1649977179
transform 1 0 27692 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1146_
timestamp 1649977179
transform -1 0 26864 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1147_
timestamp 1649977179
transform -1 0 29992 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1148_
timestamp 1649977179
transform 1 0 28336 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1149_
timestamp 1649977179
transform 1 0 25668 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1150_
timestamp 1649977179
transform 1 0 26956 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1151_
timestamp 1649977179
transform 1 0 26956 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1152_
timestamp 1649977179
transform 1 0 27876 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1153_
timestamp 1649977179
transform 1 0 28152 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1154_
timestamp 1649977179
transform -1 0 29348 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1155_
timestamp 1649977179
transform 1 0 26956 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1156_
timestamp 1649977179
transform 1 0 29532 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1157_
timestamp 1649977179
transform 1 0 30268 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1158_
timestamp 1649977179
transform -1 0 31096 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1159_
timestamp 1649977179
transform -1 0 30360 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1160_
timestamp 1649977179
transform 1 0 25208 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1161_
timestamp 1649977179
transform 1 0 30360 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1162_
timestamp 1649977179
transform -1 0 30544 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1163_
timestamp 1649977179
transform 1 0 24380 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1164_
timestamp 1649977179
transform 1 0 27232 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1165_
timestamp 1649977179
transform -1 0 28428 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1166_
timestamp 1649977179
transform 1 0 20700 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1167_
timestamp 1649977179
transform 1 0 21988 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1168_
timestamp 1649977179
transform 1 0 27968 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1169_
timestamp 1649977179
transform 1 0 31188 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1170_
timestamp 1649977179
transform 1 0 31464 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1171_
timestamp 1649977179
transform 1 0 28428 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1172_
timestamp 1649977179
transform -1 0 28060 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1173_
timestamp 1649977179
transform 1 0 28244 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1174_
timestamp 1649977179
transform -1 0 29072 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1175_
timestamp 1649977179
transform 1 0 28244 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1176_
timestamp 1649977179
transform 1 0 28152 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1177_
timestamp 1649977179
transform 1 0 31004 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1178_
timestamp 1649977179
transform -1 0 35144 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1179_
timestamp 1649977179
transform 1 0 29900 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1180_
timestamp 1649977179
transform 1 0 30820 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1181_
timestamp 1649977179
transform -1 0 32844 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1182_
timestamp 1649977179
transform 1 0 29256 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1183_
timestamp 1649977179
transform 1 0 29532 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1184_
timestamp 1649977179
transform 1 0 32936 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1185_
timestamp 1649977179
transform -1 0 33212 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1186_
timestamp 1649977179
transform -1 0 37720 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1187_
timestamp 1649977179
transform -1 0 37996 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1188_
timestamp 1649977179
transform 1 0 33764 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1189_
timestamp 1649977179
transform -1 0 35420 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1190_
timestamp 1649977179
transform -1 0 31556 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1191_
timestamp 1649977179
transform -1 0 35236 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1192_
timestamp 1649977179
transform 1 0 32660 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1193_
timestamp 1649977179
transform 1 0 37628 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1194_
timestamp 1649977179
transform -1 0 37996 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1195_
timestamp 1649977179
transform 1 0 36800 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1196_
timestamp 1649977179
transform -1 0 37996 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1197_
timestamp 1649977179
transform -1 0 35144 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1198_
timestamp 1649977179
transform 1 0 32844 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__nor4b_2  _1199_
timestamp 1649977179
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_1  _1200_
timestamp 1649977179
transform 1 0 22356 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1201_
timestamp 1649977179
transform 1 0 29256 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1202_
timestamp 1649977179
transform -1 0 34132 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1203_
timestamp 1649977179
transform -1 0 33672 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1204_
timestamp 1649977179
transform -1 0 36800 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1205_
timestamp 1649977179
transform 1 0 33304 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1206_
timestamp 1649977179
transform -1 0 35328 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1207_
timestamp 1649977179
transform 1 0 33488 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1208_
timestamp 1649977179
transform -1 0 36248 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1209_
timestamp 1649977179
transform 1 0 36892 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1210_
timestamp 1649977179
transform -1 0 35604 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1211_
timestamp 1649977179
transform -1 0 38456 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1212_
timestamp 1649977179
transform 1 0 37352 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1213_
timestamp 1649977179
transform -1 0 38364 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1214_
timestamp 1649977179
transform 1 0 33304 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1215_
timestamp 1649977179
transform -1 0 34868 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1216_
timestamp 1649977179
transform 1 0 34500 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1217_
timestamp 1649977179
transform -1 0 35696 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1218_
timestamp 1649977179
transform 1 0 37720 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1219_
timestamp 1649977179
transform -1 0 36708 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1220_
timestamp 1649977179
transform 1 0 36708 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1221_
timestamp 1649977179
transform -1 0 37352 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1222_
timestamp 1649977179
transform 1 0 38272 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1223_
timestamp 1649977179
transform 1 0 37260 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1224_
timestamp 1649977179
transform -1 0 38088 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1225_
timestamp 1649977179
transform 1 0 40572 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1226_
timestamp 1649977179
transform -1 0 38548 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1227_
timestamp 1649977179
transform 1 0 36340 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1228_
timestamp 1649977179
transform -1 0 37904 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1229_
timestamp 1649977179
transform 1 0 36340 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1230_
timestamp 1649977179
transform -1 0 38364 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1231_
timestamp 1649977179
transform -1 0 36340 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1232_
timestamp 1649977179
transform -1 0 37812 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _1233_
timestamp 1649977179
transform -1 0 22448 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1234_
timestamp 1649977179
transform 1 0 22356 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1235_
timestamp 1649977179
transform 1 0 20976 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1236_
timestamp 1649977179
transform 1 0 32568 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1237_
timestamp 1649977179
transform 1 0 34684 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1238_
timestamp 1649977179
transform 1 0 31740 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1239_
timestamp 1649977179
transform -1 0 33764 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1240_
timestamp 1649977179
transform 1 0 38088 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1241_
timestamp 1649977179
transform 1 0 30452 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1242_
timestamp 1649977179
transform 1 0 33396 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1243_
timestamp 1649977179
transform -1 0 37536 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1244_
timestamp 1649977179
transform 1 0 35972 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1245_
timestamp 1649977179
transform -1 0 38180 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1246_
timestamp 1649977179
transform -1 0 37720 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1247_
timestamp 1649977179
transform -1 0 37996 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1248_
timestamp 1649977179
transform 1 0 33764 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1249_
timestamp 1649977179
transform -1 0 35420 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1250_
timestamp 1649977179
transform -1 0 34592 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1251_
timestamp 1649977179
transform -1 0 34224 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1252_
timestamp 1649977179
transform 1 0 35144 0 -1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1253_
timestamp 1649977179
transform -1 0 34960 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1254_
timestamp 1649977179
transform -1 0 34316 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1255_
timestamp 1649977179
transform 1 0 33304 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1256_
timestamp 1649977179
transform 1 0 33488 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1257_
timestamp 1649977179
transform -1 0 33764 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1258_
timestamp 1649977179
transform -1 0 34868 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1259_
timestamp 1649977179
transform 1 0 37168 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1260_
timestamp 1649977179
transform -1 0 38272 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1261_
timestamp 1649977179
transform 1 0 36248 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1262_
timestamp 1649977179
transform -1 0 37996 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1263_
timestamp 1649977179
transform 1 0 36708 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1264_
timestamp 1649977179
transform -1 0 37904 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1265_
timestamp 1649977179
transform 1 0 32200 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1266_
timestamp 1649977179
transform 1 0 32476 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1267_
timestamp 1649977179
transform -1 0 33028 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1268_
timestamp 1649977179
transform 1 0 22172 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1269_
timestamp 1649977179
transform 1 0 23552 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1270_
timestamp 1649977179
transform -1 0 27692 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1271_
timestamp 1649977179
transform 1 0 30176 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1272_
timestamp 1649977179
transform -1 0 27968 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1273_
timestamp 1649977179
transform -1 0 27416 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1274_
timestamp 1649977179
transform 1 0 26312 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1275_
timestamp 1649977179
transform 1 0 25208 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1276_
timestamp 1649977179
transform 1 0 25392 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1277_
timestamp 1649977179
transform 1 0 27048 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1278_
timestamp 1649977179
transform -1 0 28060 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1279_
timestamp 1649977179
transform 1 0 27048 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1280_
timestamp 1649977179
transform -1 0 25852 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1281_
timestamp 1649977179
transform 1 0 25024 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1282_
timestamp 1649977179
transform 1 0 24932 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1283_
timestamp 1649977179
transform 1 0 25760 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1284_
timestamp 1649977179
transform 1 0 32016 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1285_
timestamp 1649977179
transform 1 0 25760 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1286_
timestamp 1649977179
transform -1 0 33396 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1287_
timestamp 1649977179
transform -1 0 28060 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1288_
timestamp 1649977179
transform 1 0 33672 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1289_
timestamp 1649977179
transform 1 0 34684 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1290_
timestamp 1649977179
transform 1 0 34684 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1291_
timestamp 1649977179
transform -1 0 34592 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1292_
timestamp 1649977179
transform 1 0 33304 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1293_
timestamp 1649977179
transform 1 0 32936 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1294_
timestamp 1649977179
transform 1 0 34684 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1295_
timestamp 1649977179
transform -1 0 35696 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1296_
timestamp 1649977179
transform 1 0 31096 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1297_
timestamp 1649977179
transform 1 0 30728 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1298_
timestamp 1649977179
transform -1 0 32476 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1299_
timestamp 1649977179
transform -1 0 29992 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1300_
timestamp 1649977179
transform -1 0 29808 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1301_
timestamp 1649977179
transform 1 0 20516 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1302_
timestamp 1649977179
transform 1 0 24288 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1303_
timestamp 1649977179
transform -1 0 24656 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1304_
timestamp 1649977179
transform 1 0 24472 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1305_
timestamp 1649977179
transform 1 0 24104 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1306_
timestamp 1649977179
transform 1 0 23368 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1307_
timestamp 1649977179
transform -1 0 25668 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1308_
timestamp 1649977179
transform 1 0 28796 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1309_
timestamp 1649977179
transform -1 0 30268 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1310_
timestamp 1649977179
transform 1 0 28520 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1311_
timestamp 1649977179
transform 1 0 28336 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1312_
timestamp 1649977179
transform 1 0 28060 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1313_
timestamp 1649977179
transform 1 0 28060 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1314_
timestamp 1649977179
transform -1 0 22632 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1315_
timestamp 1649977179
transform 1 0 21620 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1316_
timestamp 1649977179
transform 1 0 21804 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1317_
timestamp 1649977179
transform -1 0 23000 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1318_
timestamp 1649977179
transform -1 0 23552 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1319_
timestamp 1649977179
transform 1 0 21988 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1320_
timestamp 1649977179
transform 1 0 24380 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1321_
timestamp 1649977179
transform -1 0 24748 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1322_
timestamp 1649977179
transform -1 0 26220 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1323_
timestamp 1649977179
transform -1 0 26404 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1324_
timestamp 1649977179
transform 1 0 24564 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1325_
timestamp 1649977179
transform 1 0 24380 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1326_
timestamp 1649977179
transform 1 0 25392 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1327_
timestamp 1649977179
transform -1 0 26496 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1328_
timestamp 1649977179
transform 1 0 26220 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1329_
timestamp 1649977179
transform 1 0 20976 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1330_
timestamp 1649977179
transform -1 0 26496 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1331_
timestamp 1649977179
transform 1 0 25116 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1332_
timestamp 1649977179
transform -1 0 25760 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1333_
timestamp 1649977179
transform -1 0 24840 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1334_
timestamp 1649977179
transform 1 0 23828 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__and4bb_1  _1335_
timestamp 1649977179
transform 1 0 16652 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1336_
timestamp 1649977179
transform -1 0 18768 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1337_
timestamp 1649977179
transform -1 0 11776 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1338_
timestamp 1649977179
transform 1 0 10672 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1339_
timestamp 1649977179
transform 1 0 8924 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1340_
timestamp 1649977179
transform 1 0 6440 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1341_
timestamp 1649977179
transform 1 0 11500 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1342_
timestamp 1649977179
transform -1 0 8280 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1343_
timestamp 1649977179
transform 1 0 6440 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1344_
timestamp 1649977179
transform 1 0 7728 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1345_
timestamp 1649977179
transform -1 0 9292 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1346_
timestamp 1649977179
transform 1 0 6440 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1347_
timestamp 1649977179
transform -1 0 7636 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1348_
timestamp 1649977179
transform 1 0 7268 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1349_
timestamp 1649977179
transform 1 0 6532 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1350_
timestamp 1649977179
transform 1 0 7728 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1351_
timestamp 1649977179
transform -1 0 5980 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1352_
timestamp 1649977179
transform 1 0 5520 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1353_
timestamp 1649977179
transform -1 0 6808 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1354_
timestamp 1649977179
transform 1 0 5336 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1355_
timestamp 1649977179
transform -1 0 7268 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1356_
timestamp 1649977179
transform -1 0 5888 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1357_
timestamp 1649977179
transform -1 0 6900 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1358_
timestamp 1649977179
transform 1 0 5612 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1359_
timestamp 1649977179
transform 1 0 8924 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1360_
timestamp 1649977179
transform 1 0 7452 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1361_
timestamp 1649977179
transform -1 0 7820 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1362_
timestamp 1649977179
transform -1 0 7360 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1363_
timestamp 1649977179
transform -1 0 8004 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1364_
timestamp 1649977179
transform 1 0 6348 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1365_
timestamp 1649977179
transform 1 0 6164 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1366_
timestamp 1649977179
transform -1 0 6072 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1367_
timestamp 1649977179
transform 1 0 5152 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1368_
timestamp 1649977179
transform -1 0 5888 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1369_
timestamp 1649977179
transform 1 0 6348 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1370_
timestamp 1649977179
transform -1 0 8096 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1371_
timestamp 1649977179
transform -1 0 7912 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__nand3_1  _1372_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 10672 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1373_
timestamp 1649977179
transform 1 0 12512 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__nor3_2  _1374_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 20148 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1375_
timestamp 1649977179
transform 1 0 21988 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1376_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 20332 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nor4_2  _1377_
timestamp 1649977179
transform -1 0 22908 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__o21a_1  _1378_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 20056 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a2111oi_2  _1379_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 19780 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__and3b_2  _1380_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 18492 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _1381_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 12788 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1382_
timestamp 1649977179
transform 1 0 27048 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1383_
timestamp 1649977179
transform 1 0 28060 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1384_
timestamp 1649977179
transform 1 0 19228 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1385_
timestamp 1649977179
transform 1 0 20516 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _1386_
timestamp 1649977179
transform 1 0 18124 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1387_
timestamp 1649977179
transform -1 0 21988 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1388_
timestamp 1649977179
transform 1 0 10856 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1389_
timestamp 1649977179
transform 1 0 14352 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1390_
timestamp 1649977179
transform 1 0 19412 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1391_
timestamp 1649977179
transform -1 0 19780 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1392_
timestamp 1649977179
transform -1 0 18492 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__a211o_1  _1393_
timestamp 1649977179
transform -1 0 11684 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1394_
timestamp 1649977179
transform -1 0 20240 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1395_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 11500 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _1396_
timestamp 1649977179
transform 1 0 22816 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1397_
timestamp 1649977179
transform -1 0 23920 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1398_
timestamp 1649977179
transform -1 0 14812 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1399_
timestamp 1649977179
transform 1 0 14076 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1400_
timestamp 1649977179
transform -1 0 16008 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1401_
timestamp 1649977179
transform 1 0 22724 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1402_
timestamp 1649977179
transform -1 0 22448 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1403_
timestamp 1649977179
transform -1 0 29624 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1404_
timestamp 1649977179
transform 1 0 17112 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a2111o_1  _1405_
timestamp 1649977179
transform 1 0 22264 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1406_
timestamp 1649977179
transform -1 0 16008 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1407_
timestamp 1649977179
transform -1 0 12144 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _1408_
timestamp 1649977179
transform 1 0 11776 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1409_
timestamp 1649977179
transform 1 0 12236 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__nand3b_2  _1410_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 18952 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1411_
timestamp 1649977179
transform 1 0 19228 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1412_
timestamp 1649977179
transform -1 0 19320 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1413_
timestamp 1649977179
transform 1 0 18124 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _1414_
timestamp 1649977179
transform 1 0 29992 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1415_
timestamp 1649977179
transform 1 0 30636 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1416_
timestamp 1649977179
transform 1 0 22632 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1417_
timestamp 1649977179
transform 1 0 22540 0 -1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _1418_
timestamp 1649977179
transform 1 0 22816 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1419_
timestamp 1649977179
transform -1 0 23736 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1420_
timestamp 1649977179
transform 1 0 8464 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1421_
timestamp 1649977179
transform 1 0 12512 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a2111o_1  _1422_
timestamp 1649977179
transform 1 0 16652 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1423_
timestamp 1649977179
transform 1 0 14720 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1424_
timestamp 1649977179
transform 1 0 14536 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _1425_
timestamp 1649977179
transform 1 0 16100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1426_
timestamp 1649977179
transform 1 0 14352 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1427_
timestamp 1649977179
transform -1 0 16836 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1428_
timestamp 1649977179
transform -1 0 32016 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1429_
timestamp 1649977179
transform 1 0 15824 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1430_
timestamp 1649977179
transform 1 0 15272 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1431_
timestamp 1649977179
transform -1 0 22264 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1432_
timestamp 1649977179
transform -1 0 21068 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1433_
timestamp 1649977179
transform 1 0 20700 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1434_
timestamp 1649977179
transform -1 0 23828 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1435_
timestamp 1649977179
transform -1 0 21988 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1436_
timestamp 1649977179
transform -1 0 15732 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1437_
timestamp 1649977179
transform 1 0 11592 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _1438_
timestamp 1649977179
transform -1 0 12328 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1439_
timestamp 1649977179
transform -1 0 25024 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1440_
timestamp 1649977179
transform -1 0 24748 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1441_
timestamp 1649977179
transform 1 0 9660 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1442_
timestamp 1649977179
transform 1 0 15548 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1443_
timestamp 1649977179
transform -1 0 23736 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1444_
timestamp 1649977179
transform -1 0 26036 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1445_
timestamp 1649977179
transform -1 0 16192 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _1446_
timestamp 1649977179
transform 1 0 16652 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1447_
timestamp 1649977179
transform -1 0 15640 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1448_
timestamp 1649977179
transform 1 0 14996 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1449_
timestamp 1649977179
transform 1 0 29624 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1450_
timestamp 1649977179
transform -1 0 30452 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1451_
timestamp 1649977179
transform -1 0 26404 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1452_
timestamp 1649977179
transform -1 0 24288 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1453_
timestamp 1649977179
transform 1 0 7820 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1454_
timestamp 1649977179
transform 1 0 14536 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a2111o_1  _1455_
timestamp 1649977179
transform 1 0 16284 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1456_
timestamp 1649977179
transform -1 0 17664 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1457_
timestamp 1649977179
transform -1 0 16744 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1458_
timestamp 1649977179
transform -1 0 25392 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1459_
timestamp 1649977179
transform -1 0 23184 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1460_
timestamp 1649977179
transform 1 0 9844 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1461_
timestamp 1649977179
transform -1 0 17940 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1462_
timestamp 1649977179
transform -1 0 25024 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1463_
timestamp 1649977179
transform -1 0 28152 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1464_
timestamp 1649977179
transform -1 0 17940 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _1465_
timestamp 1649977179
transform 1 0 16008 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1466_
timestamp 1649977179
transform 1 0 14168 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1467_
timestamp 1649977179
transform 1 0 13892 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1468_
timestamp 1649977179
transform -1 0 32752 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a221oi_2  _1469_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 32292 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _1470_
timestamp 1649977179
transform -1 0 20608 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a221oi_1  _1471_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 21804 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1472_
timestamp 1649977179
transform 1 0 8924 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a221oi_1  _1473_
timestamp 1649977179
transform 1 0 13984 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _1474_
timestamp 1649977179
transform 1 0 20976 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _1475_
timestamp 1649977179
transform -1 0 14720 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _1476_
timestamp 1649977179
transform 1 0 14720 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1477_
timestamp 1649977179
transform 1 0 31280 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1478_
timestamp 1649977179
transform 1 0 32200 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1479_
timestamp 1649977179
transform -1 0 26312 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1480_
timestamp 1649977179
transform -1 0 19964 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1481_
timestamp 1649977179
transform 1 0 8924 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1482_
timestamp 1649977179
transform 1 0 12880 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a2111o_1  _1483_
timestamp 1649977179
transform 1 0 14720 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1484_
timestamp 1649977179
transform 1 0 14260 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1485_
timestamp 1649977179
transform 1 0 14260 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1486_
timestamp 1649977179
transform 1 0 29532 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1487_
timestamp 1649977179
transform -1 0 31556 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1488_
timestamp 1649977179
transform -1 0 22080 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1489_
timestamp 1649977179
transform -1 0 20516 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1490_
timestamp 1649977179
transform 1 0 10028 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1491_
timestamp 1649977179
transform 1 0 16836 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a2111o_1  _1492_
timestamp 1649977179
transform -1 0 19504 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1493_
timestamp 1649977179
transform -1 0 18768 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1494_
timestamp 1649977179
transform -1 0 19504 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1495_
timestamp 1649977179
transform 1 0 28428 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1496_
timestamp 1649977179
transform -1 0 29532 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1497_
timestamp 1649977179
transform -1 0 22264 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1498_
timestamp 1649977179
transform -1 0 19964 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1499_
timestamp 1649977179
transform 1 0 9844 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1500_
timestamp 1649977179
transform 1 0 17020 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a2111o_1  _1501_
timestamp 1649977179
transform -1 0 18768 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1502_
timestamp 1649977179
transform -1 0 19780 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1503_
timestamp 1649977179
transform -1 0 19412 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1504_
timestamp 1649977179
transform -1 0 8556 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1505_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 22356 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1506_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 12972 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _1507_
timestamp 1649977179
transform 1 0 10304 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1508_
timestamp 1649977179
transform 1 0 32660 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1509_
timestamp 1649977179
transform -1 0 36340 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1510_
timestamp 1649977179
transform 1 0 39836 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1511_
timestamp 1649977179
transform 1 0 40020 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1512_
timestamp 1649977179
transform 1 0 33948 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1513_
timestamp 1649977179
transform -1 0 37812 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1514_
timestamp 1649977179
transform -1 0 9200 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1515_
timestamp 1649977179
transform -1 0 25116 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1516_
timestamp 1649977179
transform 1 0 26956 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1517_
timestamp 1649977179
transform -1 0 25392 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1518_
timestamp 1649977179
transform 1 0 6992 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1519_
timestamp 1649977179
transform -1 0 5428 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1520_
timestamp 1649977179
transform -1 0 5612 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1521_
timestamp 1649977179
transform -1 0 5152 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1522_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2668 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1523_
timestamp 1649977179
transform 1 0 2944 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1524_
timestamp 1649977179
transform 1 0 2760 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1525_
timestamp 1649977179
transform 1 0 1840 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1526_
timestamp 1649977179
transform 1 0 3772 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1527_
timestamp 1649977179
transform 1 0 13156 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1528_
timestamp 1649977179
transform 1 0 11868 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1529_
timestamp 1649977179
transform 1 0 8740 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1530_
timestamp 1649977179
transform 1 0 13064 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1531_
timestamp 1649977179
transform 1 0 17020 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1532_
timestamp 1649977179
transform -1 0 10672 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1533_
timestamp 1649977179
transform 1 0 6348 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1534_
timestamp 1649977179
transform 1 0 3036 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1535_
timestamp 1649977179
transform 1 0 3588 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1536_
timestamp 1649977179
transform 1 0 3772 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1537_
timestamp 1649977179
transform 1 0 3588 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1538_
timestamp 1649977179
transform -1 0 6716 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1539_
timestamp 1649977179
transform 1 0 12144 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1540_
timestamp 1649977179
transform 1 0 8924 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1541_
timestamp 1649977179
transform 1 0 7728 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1542_
timestamp 1649977179
transform 1 0 10304 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1543_
timestamp 1649977179
transform 1 0 12144 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1544_
timestamp 1649977179
transform 1 0 9752 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1545_
timestamp 1649977179
transform 1 0 5244 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1546_
timestamp 1649977179
transform 1 0 2944 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1547_
timestamp 1649977179
transform 1 0 2852 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1548_
timestamp 1649977179
transform 1 0 4140 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1549_
timestamp 1649977179
transform 1 0 4968 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1550_
timestamp 1649977179
transform -1 0 11500 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1551_
timestamp 1649977179
transform 1 0 6256 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1552_
timestamp 1649977179
transform 1 0 6348 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1553_
timestamp 1649977179
transform 1 0 9568 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1554_
timestamp 1649977179
transform -1 0 11040 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1555_
timestamp 1649977179
transform 1 0 6348 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1556_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3864 0 1 25024
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1557_
timestamp 1649977179
transform 1 0 8648 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1558_
timestamp 1649977179
transform 1 0 11500 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1559_
timestamp 1649977179
transform 1 0 3036 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1560_
timestamp 1649977179
transform -1 0 15548 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1561_
timestamp 1649977179
transform 1 0 17848 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1562_
timestamp 1649977179
transform 1 0 15732 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1563_
timestamp 1649977179
transform 1 0 17296 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1564_
timestamp 1649977179
transform 1 0 18308 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1565_
timestamp 1649977179
transform 1 0 15272 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1566_
timestamp 1649977179
transform 1 0 15456 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1567_
timestamp 1649977179
transform 1 0 11776 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1568_
timestamp 1649977179
transform 1 0 21068 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1569_
timestamp 1649977179
transform 1 0 17664 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1570_
timestamp 1649977179
transform -1 0 23644 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1571_
timestamp 1649977179
transform 1 0 25024 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1572_
timestamp 1649977179
transform -1 0 27968 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1573_
timestamp 1649977179
transform -1 0 23276 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1574_
timestamp 1649977179
transform 1 0 24932 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1575_
timestamp 1649977179
transform -1 0 23552 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1576_
timestamp 1649977179
transform 1 0 19964 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1577_
timestamp 1649977179
transform 1 0 14076 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1578_
timestamp 1649977179
transform 1 0 14076 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1579_
timestamp 1649977179
transform 1 0 11684 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1580_
timestamp 1649977179
transform 1 0 11592 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1581_
timestamp 1649977179
transform 1 0 12144 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1582_
timestamp 1649977179
transform -1 0 15548 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1583_
timestamp 1649977179
transform 1 0 19872 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1584_
timestamp 1649977179
transform -1 0 18676 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1585_
timestamp 1649977179
transform 1 0 16652 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1586_
timestamp 1649977179
transform 1 0 20332 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1587_
timestamp 1649977179
transform 1 0 18860 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1588_
timestamp 1649977179
transform -1 0 24012 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1589_
timestamp 1649977179
transform 1 0 26588 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1590_
timestamp 1649977179
transform 1 0 26312 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1591_
timestamp 1649977179
transform -1 0 24012 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1592_
timestamp 1649977179
transform 1 0 26312 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1593_
timestamp 1649977179
transform 1 0 28336 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1594_
timestamp 1649977179
transform 1 0 26772 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1595_
timestamp 1649977179
transform 1 0 30176 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1596_
timestamp 1649977179
transform 1 0 29808 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1597_
timestamp 1649977179
transform -1 0 32476 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1598_
timestamp 1649977179
transform 1 0 28336 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1599_
timestamp 1649977179
transform 1 0 28520 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1600_
timestamp 1649977179
transform -1 0 25760 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1601_
timestamp 1649977179
transform 1 0 30176 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1602_
timestamp 1649977179
transform -1 0 33580 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1603_
timestamp 1649977179
transform -1 0 27508 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1604_
timestamp 1649977179
transform -1 0 39376 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1605_
timestamp 1649977179
transform -1 0 36156 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1606_
timestamp 1649977179
transform -1 0 33212 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1607_
timestamp 1649977179
transform 1 0 39008 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1608_
timestamp 1649977179
transform 1 0 38640 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1609_
timestamp 1649977179
transform -1 0 33580 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1610_
timestamp 1649977179
transform 1 0 35512 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1611_
timestamp 1649977179
transform 1 0 39100 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1612_
timestamp 1649977179
transform 1 0 39836 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1613_
timestamp 1649977179
transform 1 0 34684 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1614_
timestamp 1649977179
transform 1 0 35328 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1615_
timestamp 1649977179
transform -1 0 39008 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1616_
timestamp 1649977179
transform 1 0 37904 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1617_
timestamp 1649977179
transform 1 0 39836 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1618_
timestamp 1649977179
transform 1 0 38824 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1619_
timestamp 1649977179
transform 1 0 38916 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1620_
timestamp 1649977179
transform 1 0 39008 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1621_
timestamp 1649977179
transform 1 0 37904 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1622_
timestamp 1649977179
transform 1 0 39008 0 -1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1623_
timestamp 1649977179
transform 1 0 38824 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1624_
timestamp 1649977179
transform 1 0 34776 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1625_
timestamp 1649977179
transform 1 0 35052 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1626_
timestamp 1649977179
transform -1 0 32936 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1627_
timestamp 1649977179
transform 1 0 34868 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1628_
timestamp 1649977179
transform 1 0 39836 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1629_
timestamp 1649977179
transform -1 0 38732 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1630_
timestamp 1649977179
transform -1 0 39100 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1631_
timestamp 1649977179
transform 1 0 33304 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1632_
timestamp 1649977179
transform 1 0 24196 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1633_
timestamp 1649977179
transform 1 0 27508 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1634_
timestamp 1649977179
transform 1 0 26220 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1635_
timestamp 1649977179
transform -1 0 24288 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1636_
timestamp 1649977179
transform 1 0 23920 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1637_
timestamp 1649977179
transform -1 0 36064 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1638_
timestamp 1649977179
transform -1 0 36156 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1639_
timestamp 1649977179
transform 1 0 32752 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1640_
timestamp 1649977179
transform -1 0 37444 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1641_
timestamp 1649977179
transform -1 0 33580 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1642_
timestamp 1649977179
transform 1 0 29624 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1643_
timestamp 1649977179
transform 1 0 29992 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1644_
timestamp 1649977179
transform -1 0 33212 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1645_
timestamp 1649977179
transform 1 0 29164 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1646_
timestamp 1649977179
transform 1 0 22632 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1647_
timestamp 1649977179
transform 1 0 22080 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1648_
timestamp 1649977179
transform 1 0 26956 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1649_
timestamp 1649977179
transform 1 0 23368 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1650_
timestamp 1649977179
transform 1 0 26220 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1651_
timestamp 1649977179
transform 1 0 26956 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1652_
timestamp 1649977179
transform 1 0 25668 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1653_
timestamp 1649977179
transform 1 0 21988 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1654_
timestamp 1649977179
transform 1 0 9108 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1655_
timestamp 1649977179
transform 1 0 7268 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1656_
timestamp 1649977179
transform 1 0 6992 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1657_
timestamp 1649977179
transform 1 0 4140 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1658_
timestamp 1649977179
transform 1 0 4048 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1659_
timestamp 1649977179
transform 1 0 3772 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1660_
timestamp 1649977179
transform 1 0 7084 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1661_
timestamp 1649977179
transform 1 0 7728 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1662_
timestamp 1649977179
transform 1 0 4324 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1663_
timestamp 1649977179
transform 1 0 3772 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1664_
timestamp 1649977179
transform -1 0 6624 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1665_
timestamp 1649977179
transform 1 0 7084 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1666_
timestamp 1649977179
transform -1 0 12604 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1667_
timestamp 1649977179
transform -1 0 13524 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1668_
timestamp 1649977179
transform 1 0 16744 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1669_
timestamp 1649977179
transform 1 0 9568 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1670_
timestamp 1649977179
transform -1 0 15548 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1671_
timestamp 1649977179
transform 1 0 16652 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1672_
timestamp 1649977179
transform 1 0 13524 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1673_
timestamp 1649977179
transform -1 0 16008 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1674_
timestamp 1649977179
transform 1 0 12696 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1675_
timestamp 1649977179
transform 1 0 19780 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1676_
timestamp 1649977179
transform 1 0 19964 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1677_
timestamp 1649977179
transform 1 0 9568 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_1  _1678_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 34224 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1679_
timestamp 1649977179
transform 1 0 34960 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dlxtn_1  _1680_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _1681_
timestamp 1649977179
transform 1 0 33488 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_2  _1682_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 38088 0 -1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__dfrtp_1  _1683_
timestamp 1649977179
transform 1 0 39008 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1684_
timestamp 1649977179
transform 1 0 39836 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dlxtn_1  _1685_
timestamp 1649977179
transform -1 0 42872 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _1686_
timestamp 1649977179
transform -1 0 43700 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _1687_
timestamp 1649977179
transform 1 0 42872 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__dfrtp_1  _1688_
timestamp 1649977179
transform 1 0 33028 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1689_
timestamp 1649977179
transform 1 0 36432 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dlxtn_1  _1690_
timestamp 1649977179
transform 1 0 32200 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _1691_
timestamp 1649977179
transform 1 0 35052 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1692_
timestamp 1649977179
transform 1 0 9016 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dlxtn_2  _1693_
timestamp 1649977179
transform -1 0 32200 0 1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__dlxtn_1  _1694_
timestamp 1649977179
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__dfrtp_1  _1695_
timestamp 1649977179
transform -1 0 27784 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1696_
timestamp 1649977179
transform 1 0 24012 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dlxtn_1  _1697_
timestamp 1649977179
transform 1 0 25760 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _1698_
timestamp 1649977179
transform 1 0 21712 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _1699_
timestamp 1649977179
transform 1 0 26128 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__dfrtp_1  _1700_
timestamp 1649977179
transform 1 0 6348 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1701_
timestamp 1649977179
transform 1 0 4140 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dlxtn_1  _1702_
timestamp 1649977179
transform 1 0 4784 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _1703_
timestamp 1649977179
transform -1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_2  _1704_
timestamp 1649977179
transform 1 0 6900 0 -1 30464
box -38 -48 1234 592
use sky130_fd_sc_hd__dfrtp_1  _1705_
timestamp 1649977179
transform -1 0 4968 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1706_
timestamp 1649977179
transform -1 0 4692 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dlxtn_1  _1707_
timestamp 1649977179
transform 1 0 1656 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _1708_
timestamp 1649977179
transform 1 0 1472 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_2  _1709_
timestamp 1649977179
transform 1 0 1564 0 1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wb_clk_i dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 21988 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_0_0_wb_clk_i dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 9200 0 -1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_1_0_wb_clk_i
timestamp 1649977179
transform -1 0 8372 0 1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_2_0_wb_clk_i
timestamp 1649977179
transform -1 0 14352 0 -1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_3_0_wb_clk_i
timestamp 1649977179
transform 1 0 14168 0 -1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_4_0_wb_clk_i
timestamp 1649977179
transform 1 0 7912 0 -1 20672
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_5_0_wb_clk_i
timestamp 1649977179
transform 1 0 8096 0 -1 22848
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_6_0_wb_clk_i
timestamp 1649977179
transform 1 0 14444 0 1 19584
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_7_0_wb_clk_i
timestamp 1649977179
transform 1 0 14444 0 1 22848
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_8_0_wb_clk_i
timestamp 1649977179
transform 1 0 28520 0 -1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_9_0_wb_clk_i
timestamp 1649977179
transform -1 0 29072 0 1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_10_0_wb_clk_i
timestamp 1649977179
transform 1 0 35144 0 1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_11_0_wb_clk_i
timestamp 1649977179
transform 1 0 35696 0 -1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_12_0_wb_clk_i
timestamp 1649977179
transform 1 0 28244 0 -1 20672
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_13_0_wb_clk_i
timestamp 1649977179
transform 1 0 28060 0 1 22848
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_14_0_wb_clk_i
timestamp 1649977179
transform 1 0 35420 0 1 19584
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_15_0_wb_clk_i
timestamp 1649977179
transform 1 0 35420 0 -1 22848
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_2  input1
timestamp 1649977179
transform 1 0 5520 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input2
timestamp 1649977179
transform 1 0 5520 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input3
timestamp 1649977179
transform 1 0 8832 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1649977179
transform -1 0 18584 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1649977179
transform -1 0 19228 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input6
timestamp 1649977179
transform 1 0 6440 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1649977179
transform -1 0 19872 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1649977179
transform -1 0 19412 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input9
timestamp 1649977179
transform 1 0 9568 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input10
timestamp 1649977179
transform 1 0 12696 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input11
timestamp 1649977179
transform 1 0 17388 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input12
timestamp 1649977179
transform 1 0 13248 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input13
timestamp 1649977179
transform 1 0 12512 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1649977179
transform -1 0 5152 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input15
timestamp 1649977179
transform -1 0 6716 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input16
timestamp 1649977179
transform -1 0 15916 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1649977179
transform 1 0 12696 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input18
timestamp 1649977179
transform 1 0 9568 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input19
timestamp 1649977179
transform -1 0 18492 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input20
timestamp 1649977179
transform 1 0 11040 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input21
timestamp 1649977179
transform 1 0 15364 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input22
timestamp 1649977179
transform -1 0 10304 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input23
timestamp 1649977179
transform -1 0 11868 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input24
timestamp 1649977179
transform -1 0 15364 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input25
timestamp 1649977179
transform 1 0 13892 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input26
timestamp 1649977179
transform 1 0 15364 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1649977179
transform -1 0 9200 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1649977179
transform -1 0 7728 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1649977179
transform -1 0 7268 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output30
timestamp 1649977179
transform 1 0 21896 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output31
timestamp 1649977179
transform 1 0 30636 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output32
timestamp 1649977179
transform 1 0 39836 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output33
timestamp 1649977179
transform 1 0 48116 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output34
timestamp 1649977179
transform 1 0 56856 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output35
timestamp 1649977179
transform 1 0 65596 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output36
timestamp 1649977179
transform -1 0 10488 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output37
timestamp 1649977179
transform -1 0 8464 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output38
timestamp 1649977179
transform -1 0 14444 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output39
timestamp 1649977179
transform 1 0 14812 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output40
timestamp 1649977179
transform -1 0 11224 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output41
timestamp 1649977179
transform -1 0 17756 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output42
timestamp 1649977179
transform 1 0 16652 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output43
timestamp 1649977179
transform -1 0 9568 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output44
timestamp 1649977179
transform -1 0 14996 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output45
timestamp 1649977179
transform -1 0 11040 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output46
timestamp 1649977179
transform -1 0 13616 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output47
timestamp 1649977179
transform 1 0 16652 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output48
timestamp 1649977179
transform -1 0 14628 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_49 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 58788 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_50
timestamp 1649977179
transform -1 0 58144 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_51
timestamp 1649977179
transform -1 0 56488 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_52
timestamp 1649977179
transform -1 0 57500 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_53
timestamp 1649977179
transform -1 0 57132 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_54
timestamp 1649977179
transform -1 0 59432 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_55
timestamp 1649977179
transform -1 0 58144 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_56
timestamp 1649977179
transform -1 0 58788 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_57
timestamp 1649977179
transform -1 0 58788 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_58
timestamp 1649977179
transform -1 0 59432 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_59
timestamp 1649977179
transform -1 0 60720 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_60
timestamp 1649977179
transform -1 0 58144 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_61
timestamp 1649977179
transform -1 0 60076 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_62
timestamp 1649977179
transform -1 0 57500 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_63
timestamp 1649977179
transform -1 0 58144 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_64
timestamp 1649977179
transform -1 0 59432 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_65
timestamp 1649977179
transform -1 0 61364 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_66
timestamp 1649977179
transform -1 0 58788 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_67
timestamp 1649977179
transform -1 0 58788 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_68
timestamp 1649977179
transform -1 0 60720 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_69
timestamp 1649977179
transform -1 0 59432 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_70
timestamp 1649977179
transform -1 0 60720 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_71
timestamp 1649977179
transform -1 0 60076 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_72
timestamp 1649977179
transform -1 0 62008 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_73
timestamp 1649977179
transform -1 0 61364 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_74
timestamp 1649977179
transform -1 0 59432 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_75
timestamp 1649977179
transform -1 0 61364 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_76
timestamp 1649977179
transform -1 0 62008 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_77
timestamp 1649977179
transform -1 0 63296 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_78
timestamp 1649977179
transform -1 0 60720 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_79
timestamp 1649977179
transform -1 0 59064 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_80
timestamp 1649977179
transform -1 0 59708 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_81
timestamp 1649977179
transform -1 0 60720 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_82
timestamp 1649977179
transform -1 0 62008 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_83
timestamp 1649977179
transform -1 0 63940 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_84
timestamp 1649977179
transform -1 0 61364 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_85
timestamp 1649977179
transform -1 0 60352 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_86
timestamp 1649977179
transform -1 0 63296 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_87
timestamp 1649977179
transform 1 0 67436 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_88
timestamp 1649977179
transform 1 0 67436 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_89
timestamp 1649977179
transform 1 0 67896 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_90
timestamp 1649977179
transform 1 0 67896 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_91
timestamp 1649977179
transform 1 0 67436 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_92
timestamp 1649977179
transform 1 0 67896 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_93
timestamp 1649977179
transform 1 0 67436 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_94
timestamp 1649977179
transform 1 0 67436 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_95
timestamp 1649977179
transform 1 0 67896 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_96
timestamp 1649977179
transform 1 0 67436 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_97
timestamp 1649977179
transform 1 0 67896 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_98
timestamp 1649977179
transform 1 0 67896 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_99
timestamp 1649977179
transform 1 0 67436 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_100
timestamp 1649977179
transform 1 0 67896 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_101
timestamp 1649977179
transform 1 0 67436 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_102
timestamp 1649977179
transform 1 0 67436 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_103
timestamp 1649977179
transform 1 0 67896 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_104
timestamp 1649977179
transform 1 0 67436 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_105
timestamp 1649977179
transform 1 0 67896 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_106
timestamp 1649977179
transform 1 0 67896 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_107
timestamp 1649977179
transform 1 0 67436 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_108
timestamp 1649977179
transform 1 0 67896 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_109
timestamp 1649977179
transform 1 0 67436 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_110
timestamp 1649977179
transform 1 0 67436 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_111
timestamp 1649977179
transform 1 0 67896 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_112
timestamp 1649977179
transform 1 0 67436 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_113
timestamp 1649977179
transform 1 0 67896 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_114
timestamp 1649977179
transform 1 0 67896 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_115
timestamp 1649977179
transform 1 0 67436 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_116
timestamp 1649977179
transform 1 0 67896 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_117
timestamp 1649977179
transform 1 0 67436 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_118
timestamp 1649977179
transform 1 0 67436 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_119
timestamp 1649977179
transform 1 0 67896 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_120
timestamp 1649977179
transform 1 0 67436 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_121
timestamp 1649977179
transform 1 0 67896 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_122
timestamp 1649977179
transform 1 0 67896 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_123
timestamp 1649977179
transform 1 0 67436 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_124
timestamp 1649977179
transform 1 0 67436 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_125
timestamp 1649977179
transform -1 0 56856 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_126
timestamp 1649977179
transform -1 0 56856 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_127
timestamp 1649977179
transform -1 0 58144 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_128
timestamp 1649977179
transform -1 0 20792 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_129
timestamp 1649977179
transform 1 0 19780 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_130
timestamp 1649977179
transform 1 0 20424 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_131
timestamp 1649977179
transform 1 0 20424 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_132
timestamp 1649977179
transform -1 0 21896 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_133
timestamp 1649977179
transform 1 0 21068 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_134
timestamp 1649977179
transform 1 0 21068 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_135
timestamp 1649977179
transform -1 0 22724 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_136
timestamp 1649977179
transform 1 0 22356 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_137
timestamp 1649977179
transform -1 0 23276 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_138
timestamp 1649977179
transform 1 0 22356 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_139
timestamp 1649977179
transform -1 0 23828 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_140
timestamp 1649977179
transform 1 0 23000 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_141
timestamp 1649977179
transform 1 0 23644 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_142
timestamp 1649977179
transform -1 0 24656 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_143
timestamp 1649977179
transform 1 0 23644 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_144
timestamp 1649977179
transform 1 0 24288 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_145
timestamp 1649977179
transform -1 0 25484 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_146
timestamp 1649977179
transform 1 0 24932 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_147
timestamp 1649977179
transform 1 0 24932 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_148
timestamp 1649977179
transform -1 0 26312 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_149
timestamp 1649977179
transform 1 0 25576 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_150
timestamp 1649977179
transform 1 0 25576 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_151
timestamp 1649977179
transform -1 0 27140 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_152
timestamp 1649977179
transform 1 0 26220 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_153
timestamp 1649977179
transform 1 0 26220 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_154
timestamp 1649977179
transform -1 0 27968 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_155
timestamp 1649977179
transform 1 0 27508 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_156
timestamp 1649977179
transform 1 0 27508 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_157
timestamp 1649977179
transform 1 0 28152 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_158
timestamp 1649977179
transform -1 0 29072 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_159
timestamp 1649977179
transform 1 0 28152 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_160
timestamp 1649977179
transform 1 0 28796 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_161
timestamp 1649977179
transform 1 0 28796 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_162
timestamp 1649977179
transform -1 0 30176 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_163
timestamp 1649977179
transform 1 0 29440 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_164
timestamp 1649977179
transform 1 0 30084 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_165
timestamp 1649977179
transform -1 0 31004 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_166
timestamp 1649977179
transform 1 0 30084 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_167
timestamp 1649977179
transform 1 0 30728 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_168
timestamp 1649977179
transform -1 0 31832 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_169
timestamp 1649977179
transform 1 0 30728 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_170
timestamp 1649977179
transform 1 0 31372 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_171
timestamp 1649977179
transform -1 0 32660 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_172
timestamp 1649977179
transform 1 0 31372 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_173
timestamp 1649977179
transform 1 0 32660 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_174
timestamp 1649977179
transform -1 0 33488 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_175
timestamp 1649977179
transform 1 0 32660 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_176
timestamp 1649977179
transform 1 0 33304 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_177
timestamp 1649977179
transform 1 0 33304 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_178
timestamp 1649977179
transform 1 0 33948 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_179
timestamp 1649977179
transform -1 0 34868 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_180
timestamp 1649977179
transform 1 0 33948 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_181
timestamp 1649977179
transform 1 0 34684 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_182
timestamp 1649977179
transform -1 0 35696 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_183
timestamp 1649977179
transform 1 0 35328 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_184
timestamp 1649977179
transform -1 0 36248 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_185
timestamp 1649977179
transform -1 0 36524 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_186
timestamp 1649977179
transform -1 0 37536 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_187
timestamp 1649977179
transform -1 0 37536 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_188
timestamp 1649977179
transform -1 0 38180 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_189
timestamp 1649977179
transform -1 0 38180 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_190
timestamp 1649977179
transform -1 0 38824 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_191
timestamp 1649977179
transform -1 0 38824 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_192
timestamp 1649977179
transform -1 0 40112 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_193
timestamp 1649977179
transform -1 0 39468 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_194
timestamp 1649977179
transform -1 0 40756 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_195
timestamp 1649977179
transform -1 0 40112 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_196
timestamp 1649977179
transform -1 0 40112 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_197
timestamp 1649977179
transform -1 0 41400 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_198
timestamp 1649977179
transform -1 0 40756 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_199
timestamp 1649977179
transform -1 0 40756 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_200
timestamp 1649977179
transform -1 0 41400 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_201
timestamp 1649977179
transform -1 0 42688 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_202
timestamp 1649977179
transform -1 0 41400 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_203
timestamp 1649977179
transform -1 0 42044 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_204
timestamp 1649977179
transform -1 0 43332 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_205
timestamp 1649977179
transform -1 0 42688 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_206
timestamp 1649977179
transform -1 0 43976 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_207
timestamp 1649977179
transform -1 0 43332 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_208
timestamp 1649977179
transform -1 0 42872 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_209
timestamp 1649977179
transform -1 0 43976 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_210
timestamp 1649977179
transform -1 0 43516 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_211
timestamp 1649977179
transform -1 0 45264 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_212
timestamp 1649977179
transform -1 0 44620 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_213
timestamp 1649977179
transform -1 0 45908 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_214
timestamp 1649977179
transform -1 0 45264 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_215
timestamp 1649977179
transform -1 0 46552 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_216
timestamp 1649977179
transform -1 0 45908 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_217
timestamp 1649977179
transform -1 0 45356 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_218
timestamp 1649977179
transform -1 0 46000 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_219
timestamp 1649977179
transform -1 0 46552 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_220
timestamp 1649977179
transform -1 0 47840 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_221
timestamp 1649977179
transform -1 0 46644 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_222
timestamp 1649977179
transform -1 0 48484 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_223
timestamp 1649977179
transform -1 0 47840 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_224
timestamp 1649977179
transform -1 0 47288 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_225
timestamp 1649977179
transform -1 0 49128 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_226
timestamp 1649977179
transform -1 0 48484 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_227
timestamp 1649977179
transform -1 0 48116 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_228
timestamp 1649977179
transform -1 0 49128 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_229
timestamp 1649977179
transform -1 0 50416 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_230
timestamp 1649977179
transform -1 0 49772 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_231
timestamp 1649977179
transform -1 0 49220 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_232
timestamp 1649977179
transform -1 0 51060 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_233
timestamp 1649977179
transform -1 0 50416 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_234
timestamp 1649977179
transform -1 0 51704 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_235
timestamp 1649977179
transform -1 0 51060 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_236
timestamp 1649977179
transform -1 0 50600 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_237
timestamp 1649977179
transform -1 0 51704 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_238
timestamp 1649977179
transform -1 0 51244 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_239
timestamp 1649977179
transform -1 0 52992 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_240
timestamp 1649977179
transform -1 0 51888 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_241
timestamp 1649977179
transform -1 0 53636 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_242
timestamp 1649977179
transform -1 0 52992 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_243
timestamp 1649977179
transform -1 0 54280 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_244
timestamp 1649977179
transform -1 0 53636 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_245
timestamp 1649977179
transform -1 0 53084 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_246
timestamp 1649977179
transform -1 0 53728 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_247
timestamp 1649977179
transform -1 0 54280 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_248
timestamp 1649977179
transform -1 0 55568 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_249
timestamp 1649977179
transform -1 0 54924 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_250
timestamp 1649977179
transform -1 0 56212 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_251
timestamp 1649977179
transform -1 0 55568 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_252
timestamp 1649977179
transform -1 0 55568 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_253
timestamp 1649977179
transform -1 0 56856 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_254
timestamp 1649977179
transform -1 0 56212 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_255
timestamp 1649977179
transform -1 0 56212 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_256
timestamp 1649977179
transform -1 0 13432 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_257
timestamp 1649977179
transform -1 0 4692 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_258
timestamp 1649977179
transform 1 0 13340 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_259
timestamp 1649977179
transform -1 0 15640 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_260
timestamp 1649977179
transform 1 0 15364 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_261
timestamp 1649977179
transform 1 0 8924 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_262
timestamp 1649977179
transform -1 0 20056 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_263
timestamp 1649977179
transform -1 0 17940 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_264
timestamp 1649977179
transform -1 0 18216 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_265
timestamp 1649977179
transform -1 0 17296 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_266
timestamp 1649977179
transform -1 0 17572 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_267
timestamp 1649977179
transform 1 0 17112 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_268
timestamp 1649977179
transform -1 0 18032 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_269
timestamp 1649977179
transform 1 0 16376 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_270
timestamp 1649977179
transform -1 0 18676 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_271
timestamp 1649977179
transform -1 0 21436 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_272
timestamp 1649977179
transform 1 0 18308 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_273
timestamp 1649977179
transform -1 0 20792 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_274
timestamp 1649977179
transform 1 0 17848 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_275
timestamp 1649977179
transform 1 0 18492 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_276
timestamp 1649977179
transform 1 0 18492 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_277
timestamp 1649977179
transform 1 0 19780 0 -1 3264
box -38 -48 314 592
<< labels >>
flabel metal3 s 0 2184 800 2304 0 FreeSans 480 0 0 0 io_in[0]
port 0 nsew signal input
flabel metal3 s 0 17144 800 17264 0 FreeSans 480 0 0 0 io_in[10]
port 1 nsew signal input
flabel metal3 s 0 18640 800 18760 0 FreeSans 480 0 0 0 io_in[11]
port 2 nsew signal input
flabel metal3 s 0 20136 800 20256 0 FreeSans 480 0 0 0 io_in[12]
port 3 nsew signal input
flabel metal3 s 0 21632 800 21752 0 FreeSans 480 0 0 0 io_in[13]
port 4 nsew signal input
flabel metal3 s 0 23128 800 23248 0 FreeSans 480 0 0 0 io_in[14]
port 5 nsew signal input
flabel metal3 s 0 24624 800 24744 0 FreeSans 480 0 0 0 io_in[15]
port 6 nsew signal input
flabel metal3 s 0 26120 800 26240 0 FreeSans 480 0 0 0 io_in[16]
port 7 nsew signal input
flabel metal3 s 0 27616 800 27736 0 FreeSans 480 0 0 0 io_in[17]
port 8 nsew signal input
flabel metal3 s 0 29112 800 29232 0 FreeSans 480 0 0 0 io_in[18]
port 9 nsew signal input
flabel metal3 s 0 30608 800 30728 0 FreeSans 480 0 0 0 io_in[19]
port 10 nsew signal input
flabel metal3 s 0 3680 800 3800 0 FreeSans 480 0 0 0 io_in[1]
port 11 nsew signal input
flabel metal3 s 0 32104 800 32224 0 FreeSans 480 0 0 0 io_in[20]
port 12 nsew signal input
flabel metal3 s 0 33600 800 33720 0 FreeSans 480 0 0 0 io_in[21]
port 13 nsew signal input
flabel metal3 s 0 35096 800 35216 0 FreeSans 480 0 0 0 io_in[22]
port 14 nsew signal input
flabel metal3 s 0 36592 800 36712 0 FreeSans 480 0 0 0 io_in[23]
port 15 nsew signal input
flabel metal3 s 0 38088 800 38208 0 FreeSans 480 0 0 0 io_in[24]
port 16 nsew signal input
flabel metal3 s 0 39584 800 39704 0 FreeSans 480 0 0 0 io_in[25]
port 17 nsew signal input
flabel metal3 s 0 41080 800 41200 0 FreeSans 480 0 0 0 io_in[26]
port 18 nsew signal input
flabel metal3 s 0 42576 800 42696 0 FreeSans 480 0 0 0 io_in[27]
port 19 nsew signal input
flabel metal3 s 0 44072 800 44192 0 FreeSans 480 0 0 0 io_in[28]
port 20 nsew signal input
flabel metal3 s 0 45568 800 45688 0 FreeSans 480 0 0 0 io_in[29]
port 21 nsew signal input
flabel metal3 s 0 5176 800 5296 0 FreeSans 480 0 0 0 io_in[2]
port 22 nsew signal input
flabel metal3 s 0 47064 800 47184 0 FreeSans 480 0 0 0 io_in[30]
port 23 nsew signal input
flabel metal3 s 0 48560 800 48680 0 FreeSans 480 0 0 0 io_in[31]
port 24 nsew signal input
flabel metal3 s 0 50056 800 50176 0 FreeSans 480 0 0 0 io_in[32]
port 25 nsew signal input
flabel metal3 s 0 51552 800 51672 0 FreeSans 480 0 0 0 io_in[33]
port 26 nsew signal input
flabel metal3 s 0 53048 800 53168 0 FreeSans 480 0 0 0 io_in[34]
port 27 nsew signal input
flabel metal3 s 0 54544 800 54664 0 FreeSans 480 0 0 0 io_in[35]
port 28 nsew signal input
flabel metal3 s 0 56040 800 56160 0 FreeSans 480 0 0 0 io_in[36]
port 29 nsew signal input
flabel metal3 s 0 57536 800 57656 0 FreeSans 480 0 0 0 io_in[37]
port 30 nsew signal input
flabel metal3 s 0 6672 800 6792 0 FreeSans 480 0 0 0 io_in[3]
port 31 nsew signal input
flabel metal3 s 0 8168 800 8288 0 FreeSans 480 0 0 0 io_in[4]
port 32 nsew signal input
flabel metal3 s 0 9664 800 9784 0 FreeSans 480 0 0 0 io_in[5]
port 33 nsew signal input
flabel metal3 s 0 11160 800 11280 0 FreeSans 480 0 0 0 io_in[6]
port 34 nsew signal input
flabel metal3 s 0 12656 800 12776 0 FreeSans 480 0 0 0 io_in[7]
port 35 nsew signal input
flabel metal3 s 0 14152 800 14272 0 FreeSans 480 0 0 0 io_in[8]
port 36 nsew signal input
flabel metal3 s 0 15648 800 15768 0 FreeSans 480 0 0 0 io_in[9]
port 37 nsew signal input
flabel metal2 s 55954 0 56010 800 0 FreeSans 224 90 0 0 io_oeb[0]
port 38 nsew signal tristate
flabel metal2 s 56874 0 56930 800 0 FreeSans 224 90 0 0 io_oeb[10]
port 39 nsew signal tristate
flabel metal2 s 56966 0 57022 800 0 FreeSans 224 90 0 0 io_oeb[11]
port 40 nsew signal tristate
flabel metal2 s 57058 0 57114 800 0 FreeSans 224 90 0 0 io_oeb[12]
port 41 nsew signal tristate
flabel metal2 s 57150 0 57206 800 0 FreeSans 224 90 0 0 io_oeb[13]
port 42 nsew signal tristate
flabel metal2 s 57242 0 57298 800 0 FreeSans 224 90 0 0 io_oeb[14]
port 43 nsew signal tristate
flabel metal2 s 57334 0 57390 800 0 FreeSans 224 90 0 0 io_oeb[15]
port 44 nsew signal tristate
flabel metal2 s 57426 0 57482 800 0 FreeSans 224 90 0 0 io_oeb[16]
port 45 nsew signal tristate
flabel metal2 s 57518 0 57574 800 0 FreeSans 224 90 0 0 io_oeb[17]
port 46 nsew signal tristate
flabel metal2 s 57610 0 57666 800 0 FreeSans 224 90 0 0 io_oeb[18]
port 47 nsew signal tristate
flabel metal2 s 57702 0 57758 800 0 FreeSans 224 90 0 0 io_oeb[19]
port 48 nsew signal tristate
flabel metal2 s 56046 0 56102 800 0 FreeSans 224 90 0 0 io_oeb[1]
port 49 nsew signal tristate
flabel metal2 s 57794 0 57850 800 0 FreeSans 224 90 0 0 io_oeb[20]
port 50 nsew signal tristate
flabel metal2 s 57886 0 57942 800 0 FreeSans 224 90 0 0 io_oeb[21]
port 51 nsew signal tristate
flabel metal2 s 57978 0 58034 800 0 FreeSans 224 90 0 0 io_oeb[22]
port 52 nsew signal tristate
flabel metal2 s 58070 0 58126 800 0 FreeSans 224 90 0 0 io_oeb[23]
port 53 nsew signal tristate
flabel metal2 s 58162 0 58218 800 0 FreeSans 224 90 0 0 io_oeb[24]
port 54 nsew signal tristate
flabel metal2 s 58254 0 58310 800 0 FreeSans 224 90 0 0 io_oeb[25]
port 55 nsew signal tristate
flabel metal2 s 58346 0 58402 800 0 FreeSans 224 90 0 0 io_oeb[26]
port 56 nsew signal tristate
flabel metal2 s 58438 0 58494 800 0 FreeSans 224 90 0 0 io_oeb[27]
port 57 nsew signal tristate
flabel metal2 s 58530 0 58586 800 0 FreeSans 224 90 0 0 io_oeb[28]
port 58 nsew signal tristate
flabel metal2 s 58622 0 58678 800 0 FreeSans 224 90 0 0 io_oeb[29]
port 59 nsew signal tristate
flabel metal2 s 56138 0 56194 800 0 FreeSans 224 90 0 0 io_oeb[2]
port 60 nsew signal tristate
flabel metal2 s 58714 0 58770 800 0 FreeSans 224 90 0 0 io_oeb[30]
port 61 nsew signal tristate
flabel metal2 s 58806 0 58862 800 0 FreeSans 224 90 0 0 io_oeb[31]
port 62 nsew signal tristate
flabel metal2 s 58898 0 58954 800 0 FreeSans 224 90 0 0 io_oeb[32]
port 63 nsew signal tristate
flabel metal2 s 58990 0 59046 800 0 FreeSans 224 90 0 0 io_oeb[33]
port 64 nsew signal tristate
flabel metal2 s 59082 0 59138 800 0 FreeSans 224 90 0 0 io_oeb[34]
port 65 nsew signal tristate
flabel metal2 s 59174 0 59230 800 0 FreeSans 224 90 0 0 io_oeb[35]
port 66 nsew signal tristate
flabel metal2 s 59266 0 59322 800 0 FreeSans 224 90 0 0 io_oeb[36]
port 67 nsew signal tristate
flabel metal2 s 59358 0 59414 800 0 FreeSans 224 90 0 0 io_oeb[37]
port 68 nsew signal tristate
flabel metal2 s 56230 0 56286 800 0 FreeSans 224 90 0 0 io_oeb[3]
port 69 nsew signal tristate
flabel metal2 s 56322 0 56378 800 0 FreeSans 224 90 0 0 io_oeb[4]
port 70 nsew signal tristate
flabel metal2 s 56414 0 56470 800 0 FreeSans 224 90 0 0 io_oeb[5]
port 71 nsew signal tristate
flabel metal2 s 56506 0 56562 800 0 FreeSans 224 90 0 0 io_oeb[6]
port 72 nsew signal tristate
flabel metal2 s 56598 0 56654 800 0 FreeSans 224 90 0 0 io_oeb[7]
port 73 nsew signal tristate
flabel metal2 s 56690 0 56746 800 0 FreeSans 224 90 0 0 io_oeb[8]
port 74 nsew signal tristate
flabel metal2 s 56782 0 56838 800 0 FreeSans 224 90 0 0 io_oeb[9]
port 75 nsew signal tristate
flabel metal3 s 69200 2184 70000 2304 0 FreeSans 480 0 0 0 io_out[0]
port 76 nsew signal tristate
flabel metal3 s 69200 17144 70000 17264 0 FreeSans 480 0 0 0 io_out[10]
port 77 nsew signal tristate
flabel metal3 s 69200 18640 70000 18760 0 FreeSans 480 0 0 0 io_out[11]
port 78 nsew signal tristate
flabel metal3 s 69200 20136 70000 20256 0 FreeSans 480 0 0 0 io_out[12]
port 79 nsew signal tristate
flabel metal3 s 69200 21632 70000 21752 0 FreeSans 480 0 0 0 io_out[13]
port 80 nsew signal tristate
flabel metal3 s 69200 23128 70000 23248 0 FreeSans 480 0 0 0 io_out[14]
port 81 nsew signal tristate
flabel metal3 s 69200 24624 70000 24744 0 FreeSans 480 0 0 0 io_out[15]
port 82 nsew signal tristate
flabel metal3 s 69200 26120 70000 26240 0 FreeSans 480 0 0 0 io_out[16]
port 83 nsew signal tristate
flabel metal3 s 69200 27616 70000 27736 0 FreeSans 480 0 0 0 io_out[17]
port 84 nsew signal tristate
flabel metal3 s 69200 29112 70000 29232 0 FreeSans 480 0 0 0 io_out[18]
port 85 nsew signal tristate
flabel metal3 s 69200 30608 70000 30728 0 FreeSans 480 0 0 0 io_out[19]
port 86 nsew signal tristate
flabel metal3 s 69200 3680 70000 3800 0 FreeSans 480 0 0 0 io_out[1]
port 87 nsew signal tristate
flabel metal3 s 69200 32104 70000 32224 0 FreeSans 480 0 0 0 io_out[20]
port 88 nsew signal tristate
flabel metal3 s 69200 33600 70000 33720 0 FreeSans 480 0 0 0 io_out[21]
port 89 nsew signal tristate
flabel metal3 s 69200 35096 70000 35216 0 FreeSans 480 0 0 0 io_out[22]
port 90 nsew signal tristate
flabel metal3 s 69200 36592 70000 36712 0 FreeSans 480 0 0 0 io_out[23]
port 91 nsew signal tristate
flabel metal3 s 69200 38088 70000 38208 0 FreeSans 480 0 0 0 io_out[24]
port 92 nsew signal tristate
flabel metal3 s 69200 39584 70000 39704 0 FreeSans 480 0 0 0 io_out[25]
port 93 nsew signal tristate
flabel metal3 s 69200 41080 70000 41200 0 FreeSans 480 0 0 0 io_out[26]
port 94 nsew signal tristate
flabel metal3 s 69200 42576 70000 42696 0 FreeSans 480 0 0 0 io_out[27]
port 95 nsew signal tristate
flabel metal3 s 69200 44072 70000 44192 0 FreeSans 480 0 0 0 io_out[28]
port 96 nsew signal tristate
flabel metal3 s 69200 45568 70000 45688 0 FreeSans 480 0 0 0 io_out[29]
port 97 nsew signal tristate
flabel metal3 s 69200 5176 70000 5296 0 FreeSans 480 0 0 0 io_out[2]
port 98 nsew signal tristate
flabel metal3 s 69200 47064 70000 47184 0 FreeSans 480 0 0 0 io_out[30]
port 99 nsew signal tristate
flabel metal3 s 69200 48560 70000 48680 0 FreeSans 480 0 0 0 io_out[31]
port 100 nsew signal tristate
flabel metal3 s 69200 50056 70000 50176 0 FreeSans 480 0 0 0 io_out[32]
port 101 nsew signal tristate
flabel metal3 s 69200 51552 70000 51672 0 FreeSans 480 0 0 0 io_out[33]
port 102 nsew signal tristate
flabel metal3 s 69200 53048 70000 53168 0 FreeSans 480 0 0 0 io_out[34]
port 103 nsew signal tristate
flabel metal3 s 69200 54544 70000 54664 0 FreeSans 480 0 0 0 io_out[35]
port 104 nsew signal tristate
flabel metal3 s 69200 56040 70000 56160 0 FreeSans 480 0 0 0 io_out[36]
port 105 nsew signal tristate
flabel metal3 s 69200 57536 70000 57656 0 FreeSans 480 0 0 0 io_out[37]
port 106 nsew signal tristate
flabel metal3 s 69200 6672 70000 6792 0 FreeSans 480 0 0 0 io_out[3]
port 107 nsew signal tristate
flabel metal3 s 69200 8168 70000 8288 0 FreeSans 480 0 0 0 io_out[4]
port 108 nsew signal tristate
flabel metal3 s 69200 9664 70000 9784 0 FreeSans 480 0 0 0 io_out[5]
port 109 nsew signal tristate
flabel metal3 s 69200 11160 70000 11280 0 FreeSans 480 0 0 0 io_out[6]
port 110 nsew signal tristate
flabel metal3 s 69200 12656 70000 12776 0 FreeSans 480 0 0 0 io_out[7]
port 111 nsew signal tristate
flabel metal3 s 69200 14152 70000 14272 0 FreeSans 480 0 0 0 io_out[8]
port 112 nsew signal tristate
flabel metal3 s 69200 15648 70000 15768 0 FreeSans 480 0 0 0 io_out[9]
port 113 nsew signal tristate
flabel metal2 s 55678 0 55734 800 0 FreeSans 224 90 0 0 irq[0]
port 114 nsew signal tristate
flabel metal2 s 55770 0 55826 800 0 FreeSans 224 90 0 0 irq[1]
port 115 nsew signal tristate
flabel metal2 s 55862 0 55918 800 0 FreeSans 224 90 0 0 irq[2]
port 116 nsew signal tristate
flabel metal2 s 20350 0 20406 800 0 FreeSans 224 90 0 0 la_data_in[0]
port 117 nsew signal input
flabel metal2 s 47950 0 48006 800 0 FreeSans 224 90 0 0 la_data_in[100]
port 118 nsew signal input
flabel metal2 s 48226 0 48282 800 0 FreeSans 224 90 0 0 la_data_in[101]
port 119 nsew signal input
flabel metal2 s 48502 0 48558 800 0 FreeSans 224 90 0 0 la_data_in[102]
port 120 nsew signal input
flabel metal2 s 48778 0 48834 800 0 FreeSans 224 90 0 0 la_data_in[103]
port 121 nsew signal input
flabel metal2 s 49054 0 49110 800 0 FreeSans 224 90 0 0 la_data_in[104]
port 122 nsew signal input
flabel metal2 s 49330 0 49386 800 0 FreeSans 224 90 0 0 la_data_in[105]
port 123 nsew signal input
flabel metal2 s 49606 0 49662 800 0 FreeSans 224 90 0 0 la_data_in[106]
port 124 nsew signal input
flabel metal2 s 49882 0 49938 800 0 FreeSans 224 90 0 0 la_data_in[107]
port 125 nsew signal input
flabel metal2 s 50158 0 50214 800 0 FreeSans 224 90 0 0 la_data_in[108]
port 126 nsew signal input
flabel metal2 s 50434 0 50490 800 0 FreeSans 224 90 0 0 la_data_in[109]
port 127 nsew signal input
flabel metal2 s 23110 0 23166 800 0 FreeSans 224 90 0 0 la_data_in[10]
port 128 nsew signal input
flabel metal2 s 50710 0 50766 800 0 FreeSans 224 90 0 0 la_data_in[110]
port 129 nsew signal input
flabel metal2 s 50986 0 51042 800 0 FreeSans 224 90 0 0 la_data_in[111]
port 130 nsew signal input
flabel metal2 s 51262 0 51318 800 0 FreeSans 224 90 0 0 la_data_in[112]
port 131 nsew signal input
flabel metal2 s 51538 0 51594 800 0 FreeSans 224 90 0 0 la_data_in[113]
port 132 nsew signal input
flabel metal2 s 51814 0 51870 800 0 FreeSans 224 90 0 0 la_data_in[114]
port 133 nsew signal input
flabel metal2 s 52090 0 52146 800 0 FreeSans 224 90 0 0 la_data_in[115]
port 134 nsew signal input
flabel metal2 s 52366 0 52422 800 0 FreeSans 224 90 0 0 la_data_in[116]
port 135 nsew signal input
flabel metal2 s 52642 0 52698 800 0 FreeSans 224 90 0 0 la_data_in[117]
port 136 nsew signal input
flabel metal2 s 52918 0 52974 800 0 FreeSans 224 90 0 0 la_data_in[118]
port 137 nsew signal input
flabel metal2 s 53194 0 53250 800 0 FreeSans 224 90 0 0 la_data_in[119]
port 138 nsew signal input
flabel metal2 s 23386 0 23442 800 0 FreeSans 224 90 0 0 la_data_in[11]
port 139 nsew signal input
flabel metal2 s 53470 0 53526 800 0 FreeSans 224 90 0 0 la_data_in[120]
port 140 nsew signal input
flabel metal2 s 53746 0 53802 800 0 FreeSans 224 90 0 0 la_data_in[121]
port 141 nsew signal input
flabel metal2 s 54022 0 54078 800 0 FreeSans 224 90 0 0 la_data_in[122]
port 142 nsew signal input
flabel metal2 s 54298 0 54354 800 0 FreeSans 224 90 0 0 la_data_in[123]
port 143 nsew signal input
flabel metal2 s 54574 0 54630 800 0 FreeSans 224 90 0 0 la_data_in[124]
port 144 nsew signal input
flabel metal2 s 54850 0 54906 800 0 FreeSans 224 90 0 0 la_data_in[125]
port 145 nsew signal input
flabel metal2 s 55126 0 55182 800 0 FreeSans 224 90 0 0 la_data_in[126]
port 146 nsew signal input
flabel metal2 s 55402 0 55458 800 0 FreeSans 224 90 0 0 la_data_in[127]
port 147 nsew signal input
flabel metal2 s 23662 0 23718 800 0 FreeSans 224 90 0 0 la_data_in[12]
port 148 nsew signal input
flabel metal2 s 23938 0 23994 800 0 FreeSans 224 90 0 0 la_data_in[13]
port 149 nsew signal input
flabel metal2 s 24214 0 24270 800 0 FreeSans 224 90 0 0 la_data_in[14]
port 150 nsew signal input
flabel metal2 s 24490 0 24546 800 0 FreeSans 224 90 0 0 la_data_in[15]
port 151 nsew signal input
flabel metal2 s 24766 0 24822 800 0 FreeSans 224 90 0 0 la_data_in[16]
port 152 nsew signal input
flabel metal2 s 25042 0 25098 800 0 FreeSans 224 90 0 0 la_data_in[17]
port 153 nsew signal input
flabel metal2 s 25318 0 25374 800 0 FreeSans 224 90 0 0 la_data_in[18]
port 154 nsew signal input
flabel metal2 s 25594 0 25650 800 0 FreeSans 224 90 0 0 la_data_in[19]
port 155 nsew signal input
flabel metal2 s 20626 0 20682 800 0 FreeSans 224 90 0 0 la_data_in[1]
port 156 nsew signal input
flabel metal2 s 25870 0 25926 800 0 FreeSans 224 90 0 0 la_data_in[20]
port 157 nsew signal input
flabel metal2 s 26146 0 26202 800 0 FreeSans 224 90 0 0 la_data_in[21]
port 158 nsew signal input
flabel metal2 s 26422 0 26478 800 0 FreeSans 224 90 0 0 la_data_in[22]
port 159 nsew signal input
flabel metal2 s 26698 0 26754 800 0 FreeSans 224 90 0 0 la_data_in[23]
port 160 nsew signal input
flabel metal2 s 26974 0 27030 800 0 FreeSans 224 90 0 0 la_data_in[24]
port 161 nsew signal input
flabel metal2 s 27250 0 27306 800 0 FreeSans 224 90 0 0 la_data_in[25]
port 162 nsew signal input
flabel metal2 s 27526 0 27582 800 0 FreeSans 224 90 0 0 la_data_in[26]
port 163 nsew signal input
flabel metal2 s 27802 0 27858 800 0 FreeSans 224 90 0 0 la_data_in[27]
port 164 nsew signal input
flabel metal2 s 28078 0 28134 800 0 FreeSans 224 90 0 0 la_data_in[28]
port 165 nsew signal input
flabel metal2 s 28354 0 28410 800 0 FreeSans 224 90 0 0 la_data_in[29]
port 166 nsew signal input
flabel metal2 s 20902 0 20958 800 0 FreeSans 224 90 0 0 la_data_in[2]
port 167 nsew signal input
flabel metal2 s 28630 0 28686 800 0 FreeSans 224 90 0 0 la_data_in[30]
port 168 nsew signal input
flabel metal2 s 28906 0 28962 800 0 FreeSans 224 90 0 0 la_data_in[31]
port 169 nsew signal input
flabel metal2 s 29182 0 29238 800 0 FreeSans 224 90 0 0 la_data_in[32]
port 170 nsew signal input
flabel metal2 s 29458 0 29514 800 0 FreeSans 224 90 0 0 la_data_in[33]
port 171 nsew signal input
flabel metal2 s 29734 0 29790 800 0 FreeSans 224 90 0 0 la_data_in[34]
port 172 nsew signal input
flabel metal2 s 30010 0 30066 800 0 FreeSans 224 90 0 0 la_data_in[35]
port 173 nsew signal input
flabel metal2 s 30286 0 30342 800 0 FreeSans 224 90 0 0 la_data_in[36]
port 174 nsew signal input
flabel metal2 s 30562 0 30618 800 0 FreeSans 224 90 0 0 la_data_in[37]
port 175 nsew signal input
flabel metal2 s 30838 0 30894 800 0 FreeSans 224 90 0 0 la_data_in[38]
port 176 nsew signal input
flabel metal2 s 31114 0 31170 800 0 FreeSans 224 90 0 0 la_data_in[39]
port 177 nsew signal input
flabel metal2 s 21178 0 21234 800 0 FreeSans 224 90 0 0 la_data_in[3]
port 178 nsew signal input
flabel metal2 s 31390 0 31446 800 0 FreeSans 224 90 0 0 la_data_in[40]
port 179 nsew signal input
flabel metal2 s 31666 0 31722 800 0 FreeSans 224 90 0 0 la_data_in[41]
port 180 nsew signal input
flabel metal2 s 31942 0 31998 800 0 FreeSans 224 90 0 0 la_data_in[42]
port 181 nsew signal input
flabel metal2 s 32218 0 32274 800 0 FreeSans 224 90 0 0 la_data_in[43]
port 182 nsew signal input
flabel metal2 s 32494 0 32550 800 0 FreeSans 224 90 0 0 la_data_in[44]
port 183 nsew signal input
flabel metal2 s 32770 0 32826 800 0 FreeSans 224 90 0 0 la_data_in[45]
port 184 nsew signal input
flabel metal2 s 33046 0 33102 800 0 FreeSans 224 90 0 0 la_data_in[46]
port 185 nsew signal input
flabel metal2 s 33322 0 33378 800 0 FreeSans 224 90 0 0 la_data_in[47]
port 186 nsew signal input
flabel metal2 s 33598 0 33654 800 0 FreeSans 224 90 0 0 la_data_in[48]
port 187 nsew signal input
flabel metal2 s 33874 0 33930 800 0 FreeSans 224 90 0 0 la_data_in[49]
port 188 nsew signal input
flabel metal2 s 21454 0 21510 800 0 FreeSans 224 90 0 0 la_data_in[4]
port 189 nsew signal input
flabel metal2 s 34150 0 34206 800 0 FreeSans 224 90 0 0 la_data_in[50]
port 190 nsew signal input
flabel metal2 s 34426 0 34482 800 0 FreeSans 224 90 0 0 la_data_in[51]
port 191 nsew signal input
flabel metal2 s 34702 0 34758 800 0 FreeSans 224 90 0 0 la_data_in[52]
port 192 nsew signal input
flabel metal2 s 34978 0 35034 800 0 FreeSans 224 90 0 0 la_data_in[53]
port 193 nsew signal input
flabel metal2 s 35254 0 35310 800 0 FreeSans 224 90 0 0 la_data_in[54]
port 194 nsew signal input
flabel metal2 s 35530 0 35586 800 0 FreeSans 224 90 0 0 la_data_in[55]
port 195 nsew signal input
flabel metal2 s 35806 0 35862 800 0 FreeSans 224 90 0 0 la_data_in[56]
port 196 nsew signal input
flabel metal2 s 36082 0 36138 800 0 FreeSans 224 90 0 0 la_data_in[57]
port 197 nsew signal input
flabel metal2 s 36358 0 36414 800 0 FreeSans 224 90 0 0 la_data_in[58]
port 198 nsew signal input
flabel metal2 s 36634 0 36690 800 0 FreeSans 224 90 0 0 la_data_in[59]
port 199 nsew signal input
flabel metal2 s 21730 0 21786 800 0 FreeSans 224 90 0 0 la_data_in[5]
port 200 nsew signal input
flabel metal2 s 36910 0 36966 800 0 FreeSans 224 90 0 0 la_data_in[60]
port 201 nsew signal input
flabel metal2 s 37186 0 37242 800 0 FreeSans 224 90 0 0 la_data_in[61]
port 202 nsew signal input
flabel metal2 s 37462 0 37518 800 0 FreeSans 224 90 0 0 la_data_in[62]
port 203 nsew signal input
flabel metal2 s 37738 0 37794 800 0 FreeSans 224 90 0 0 la_data_in[63]
port 204 nsew signal input
flabel metal2 s 38014 0 38070 800 0 FreeSans 224 90 0 0 la_data_in[64]
port 205 nsew signal input
flabel metal2 s 38290 0 38346 800 0 FreeSans 224 90 0 0 la_data_in[65]
port 206 nsew signal input
flabel metal2 s 38566 0 38622 800 0 FreeSans 224 90 0 0 la_data_in[66]
port 207 nsew signal input
flabel metal2 s 38842 0 38898 800 0 FreeSans 224 90 0 0 la_data_in[67]
port 208 nsew signal input
flabel metal2 s 39118 0 39174 800 0 FreeSans 224 90 0 0 la_data_in[68]
port 209 nsew signal input
flabel metal2 s 39394 0 39450 800 0 FreeSans 224 90 0 0 la_data_in[69]
port 210 nsew signal input
flabel metal2 s 22006 0 22062 800 0 FreeSans 224 90 0 0 la_data_in[6]
port 211 nsew signal input
flabel metal2 s 39670 0 39726 800 0 FreeSans 224 90 0 0 la_data_in[70]
port 212 nsew signal input
flabel metal2 s 39946 0 40002 800 0 FreeSans 224 90 0 0 la_data_in[71]
port 213 nsew signal input
flabel metal2 s 40222 0 40278 800 0 FreeSans 224 90 0 0 la_data_in[72]
port 214 nsew signal input
flabel metal2 s 40498 0 40554 800 0 FreeSans 224 90 0 0 la_data_in[73]
port 215 nsew signal input
flabel metal2 s 40774 0 40830 800 0 FreeSans 224 90 0 0 la_data_in[74]
port 216 nsew signal input
flabel metal2 s 41050 0 41106 800 0 FreeSans 224 90 0 0 la_data_in[75]
port 217 nsew signal input
flabel metal2 s 41326 0 41382 800 0 FreeSans 224 90 0 0 la_data_in[76]
port 218 nsew signal input
flabel metal2 s 41602 0 41658 800 0 FreeSans 224 90 0 0 la_data_in[77]
port 219 nsew signal input
flabel metal2 s 41878 0 41934 800 0 FreeSans 224 90 0 0 la_data_in[78]
port 220 nsew signal input
flabel metal2 s 42154 0 42210 800 0 FreeSans 224 90 0 0 la_data_in[79]
port 221 nsew signal input
flabel metal2 s 22282 0 22338 800 0 FreeSans 224 90 0 0 la_data_in[7]
port 222 nsew signal input
flabel metal2 s 42430 0 42486 800 0 FreeSans 224 90 0 0 la_data_in[80]
port 223 nsew signal input
flabel metal2 s 42706 0 42762 800 0 FreeSans 224 90 0 0 la_data_in[81]
port 224 nsew signal input
flabel metal2 s 42982 0 43038 800 0 FreeSans 224 90 0 0 la_data_in[82]
port 225 nsew signal input
flabel metal2 s 43258 0 43314 800 0 FreeSans 224 90 0 0 la_data_in[83]
port 226 nsew signal input
flabel metal2 s 43534 0 43590 800 0 FreeSans 224 90 0 0 la_data_in[84]
port 227 nsew signal input
flabel metal2 s 43810 0 43866 800 0 FreeSans 224 90 0 0 la_data_in[85]
port 228 nsew signal input
flabel metal2 s 44086 0 44142 800 0 FreeSans 224 90 0 0 la_data_in[86]
port 229 nsew signal input
flabel metal2 s 44362 0 44418 800 0 FreeSans 224 90 0 0 la_data_in[87]
port 230 nsew signal input
flabel metal2 s 44638 0 44694 800 0 FreeSans 224 90 0 0 la_data_in[88]
port 231 nsew signal input
flabel metal2 s 44914 0 44970 800 0 FreeSans 224 90 0 0 la_data_in[89]
port 232 nsew signal input
flabel metal2 s 22558 0 22614 800 0 FreeSans 224 90 0 0 la_data_in[8]
port 233 nsew signal input
flabel metal2 s 45190 0 45246 800 0 FreeSans 224 90 0 0 la_data_in[90]
port 234 nsew signal input
flabel metal2 s 45466 0 45522 800 0 FreeSans 224 90 0 0 la_data_in[91]
port 235 nsew signal input
flabel metal2 s 45742 0 45798 800 0 FreeSans 224 90 0 0 la_data_in[92]
port 236 nsew signal input
flabel metal2 s 46018 0 46074 800 0 FreeSans 224 90 0 0 la_data_in[93]
port 237 nsew signal input
flabel metal2 s 46294 0 46350 800 0 FreeSans 224 90 0 0 la_data_in[94]
port 238 nsew signal input
flabel metal2 s 46570 0 46626 800 0 FreeSans 224 90 0 0 la_data_in[95]
port 239 nsew signal input
flabel metal2 s 46846 0 46902 800 0 FreeSans 224 90 0 0 la_data_in[96]
port 240 nsew signal input
flabel metal2 s 47122 0 47178 800 0 FreeSans 224 90 0 0 la_data_in[97]
port 241 nsew signal input
flabel metal2 s 47398 0 47454 800 0 FreeSans 224 90 0 0 la_data_in[98]
port 242 nsew signal input
flabel metal2 s 47674 0 47730 800 0 FreeSans 224 90 0 0 la_data_in[99]
port 243 nsew signal input
flabel metal2 s 22834 0 22890 800 0 FreeSans 224 90 0 0 la_data_in[9]
port 244 nsew signal input
flabel metal2 s 20442 0 20498 800 0 FreeSans 224 90 0 0 la_data_out[0]
port 245 nsew signal tristate
flabel metal2 s 48042 0 48098 800 0 FreeSans 224 90 0 0 la_data_out[100]
port 246 nsew signal tristate
flabel metal2 s 48318 0 48374 800 0 FreeSans 224 90 0 0 la_data_out[101]
port 247 nsew signal tristate
flabel metal2 s 48594 0 48650 800 0 FreeSans 224 90 0 0 la_data_out[102]
port 248 nsew signal tristate
flabel metal2 s 48870 0 48926 800 0 FreeSans 224 90 0 0 la_data_out[103]
port 249 nsew signal tristate
flabel metal2 s 49146 0 49202 800 0 FreeSans 224 90 0 0 la_data_out[104]
port 250 nsew signal tristate
flabel metal2 s 49422 0 49478 800 0 FreeSans 224 90 0 0 la_data_out[105]
port 251 nsew signal tristate
flabel metal2 s 49698 0 49754 800 0 FreeSans 224 90 0 0 la_data_out[106]
port 252 nsew signal tristate
flabel metal2 s 49974 0 50030 800 0 FreeSans 224 90 0 0 la_data_out[107]
port 253 nsew signal tristate
flabel metal2 s 50250 0 50306 800 0 FreeSans 224 90 0 0 la_data_out[108]
port 254 nsew signal tristate
flabel metal2 s 50526 0 50582 800 0 FreeSans 224 90 0 0 la_data_out[109]
port 255 nsew signal tristate
flabel metal2 s 23202 0 23258 800 0 FreeSans 224 90 0 0 la_data_out[10]
port 256 nsew signal tristate
flabel metal2 s 50802 0 50858 800 0 FreeSans 224 90 0 0 la_data_out[110]
port 257 nsew signal tristate
flabel metal2 s 51078 0 51134 800 0 FreeSans 224 90 0 0 la_data_out[111]
port 258 nsew signal tristate
flabel metal2 s 51354 0 51410 800 0 FreeSans 224 90 0 0 la_data_out[112]
port 259 nsew signal tristate
flabel metal2 s 51630 0 51686 800 0 FreeSans 224 90 0 0 la_data_out[113]
port 260 nsew signal tristate
flabel metal2 s 51906 0 51962 800 0 FreeSans 224 90 0 0 la_data_out[114]
port 261 nsew signal tristate
flabel metal2 s 52182 0 52238 800 0 FreeSans 224 90 0 0 la_data_out[115]
port 262 nsew signal tristate
flabel metal2 s 52458 0 52514 800 0 FreeSans 224 90 0 0 la_data_out[116]
port 263 nsew signal tristate
flabel metal2 s 52734 0 52790 800 0 FreeSans 224 90 0 0 la_data_out[117]
port 264 nsew signal tristate
flabel metal2 s 53010 0 53066 800 0 FreeSans 224 90 0 0 la_data_out[118]
port 265 nsew signal tristate
flabel metal2 s 53286 0 53342 800 0 FreeSans 224 90 0 0 la_data_out[119]
port 266 nsew signal tristate
flabel metal2 s 23478 0 23534 800 0 FreeSans 224 90 0 0 la_data_out[11]
port 267 nsew signal tristate
flabel metal2 s 53562 0 53618 800 0 FreeSans 224 90 0 0 la_data_out[120]
port 268 nsew signal tristate
flabel metal2 s 53838 0 53894 800 0 FreeSans 224 90 0 0 la_data_out[121]
port 269 nsew signal tristate
flabel metal2 s 54114 0 54170 800 0 FreeSans 224 90 0 0 la_data_out[122]
port 270 nsew signal tristate
flabel metal2 s 54390 0 54446 800 0 FreeSans 224 90 0 0 la_data_out[123]
port 271 nsew signal tristate
flabel metal2 s 54666 0 54722 800 0 FreeSans 224 90 0 0 la_data_out[124]
port 272 nsew signal tristate
flabel metal2 s 54942 0 54998 800 0 FreeSans 224 90 0 0 la_data_out[125]
port 273 nsew signal tristate
flabel metal2 s 55218 0 55274 800 0 FreeSans 224 90 0 0 la_data_out[126]
port 274 nsew signal tristate
flabel metal2 s 55494 0 55550 800 0 FreeSans 224 90 0 0 la_data_out[127]
port 275 nsew signal tristate
flabel metal2 s 23754 0 23810 800 0 FreeSans 224 90 0 0 la_data_out[12]
port 276 nsew signal tristate
flabel metal2 s 24030 0 24086 800 0 FreeSans 224 90 0 0 la_data_out[13]
port 277 nsew signal tristate
flabel metal2 s 24306 0 24362 800 0 FreeSans 224 90 0 0 la_data_out[14]
port 278 nsew signal tristate
flabel metal2 s 24582 0 24638 800 0 FreeSans 224 90 0 0 la_data_out[15]
port 279 nsew signal tristate
flabel metal2 s 24858 0 24914 800 0 FreeSans 224 90 0 0 la_data_out[16]
port 280 nsew signal tristate
flabel metal2 s 25134 0 25190 800 0 FreeSans 224 90 0 0 la_data_out[17]
port 281 nsew signal tristate
flabel metal2 s 25410 0 25466 800 0 FreeSans 224 90 0 0 la_data_out[18]
port 282 nsew signal tristate
flabel metal2 s 25686 0 25742 800 0 FreeSans 224 90 0 0 la_data_out[19]
port 283 nsew signal tristate
flabel metal2 s 20718 0 20774 800 0 FreeSans 224 90 0 0 la_data_out[1]
port 284 nsew signal tristate
flabel metal2 s 25962 0 26018 800 0 FreeSans 224 90 0 0 la_data_out[20]
port 285 nsew signal tristate
flabel metal2 s 26238 0 26294 800 0 FreeSans 224 90 0 0 la_data_out[21]
port 286 nsew signal tristate
flabel metal2 s 26514 0 26570 800 0 FreeSans 224 90 0 0 la_data_out[22]
port 287 nsew signal tristate
flabel metal2 s 26790 0 26846 800 0 FreeSans 224 90 0 0 la_data_out[23]
port 288 nsew signal tristate
flabel metal2 s 27066 0 27122 800 0 FreeSans 224 90 0 0 la_data_out[24]
port 289 nsew signal tristate
flabel metal2 s 27342 0 27398 800 0 FreeSans 224 90 0 0 la_data_out[25]
port 290 nsew signal tristate
flabel metal2 s 27618 0 27674 800 0 FreeSans 224 90 0 0 la_data_out[26]
port 291 nsew signal tristate
flabel metal2 s 27894 0 27950 800 0 FreeSans 224 90 0 0 la_data_out[27]
port 292 nsew signal tristate
flabel metal2 s 28170 0 28226 800 0 FreeSans 224 90 0 0 la_data_out[28]
port 293 nsew signal tristate
flabel metal2 s 28446 0 28502 800 0 FreeSans 224 90 0 0 la_data_out[29]
port 294 nsew signal tristate
flabel metal2 s 20994 0 21050 800 0 FreeSans 224 90 0 0 la_data_out[2]
port 295 nsew signal tristate
flabel metal2 s 28722 0 28778 800 0 FreeSans 224 90 0 0 la_data_out[30]
port 296 nsew signal tristate
flabel metal2 s 28998 0 29054 800 0 FreeSans 224 90 0 0 la_data_out[31]
port 297 nsew signal tristate
flabel metal2 s 29274 0 29330 800 0 FreeSans 224 90 0 0 la_data_out[32]
port 298 nsew signal tristate
flabel metal2 s 29550 0 29606 800 0 FreeSans 224 90 0 0 la_data_out[33]
port 299 nsew signal tristate
flabel metal2 s 29826 0 29882 800 0 FreeSans 224 90 0 0 la_data_out[34]
port 300 nsew signal tristate
flabel metal2 s 30102 0 30158 800 0 FreeSans 224 90 0 0 la_data_out[35]
port 301 nsew signal tristate
flabel metal2 s 30378 0 30434 800 0 FreeSans 224 90 0 0 la_data_out[36]
port 302 nsew signal tristate
flabel metal2 s 30654 0 30710 800 0 FreeSans 224 90 0 0 la_data_out[37]
port 303 nsew signal tristate
flabel metal2 s 30930 0 30986 800 0 FreeSans 224 90 0 0 la_data_out[38]
port 304 nsew signal tristate
flabel metal2 s 31206 0 31262 800 0 FreeSans 224 90 0 0 la_data_out[39]
port 305 nsew signal tristate
flabel metal2 s 21270 0 21326 800 0 FreeSans 224 90 0 0 la_data_out[3]
port 306 nsew signal tristate
flabel metal2 s 31482 0 31538 800 0 FreeSans 224 90 0 0 la_data_out[40]
port 307 nsew signal tristate
flabel metal2 s 31758 0 31814 800 0 FreeSans 224 90 0 0 la_data_out[41]
port 308 nsew signal tristate
flabel metal2 s 32034 0 32090 800 0 FreeSans 224 90 0 0 la_data_out[42]
port 309 nsew signal tristate
flabel metal2 s 32310 0 32366 800 0 FreeSans 224 90 0 0 la_data_out[43]
port 310 nsew signal tristate
flabel metal2 s 32586 0 32642 800 0 FreeSans 224 90 0 0 la_data_out[44]
port 311 nsew signal tristate
flabel metal2 s 32862 0 32918 800 0 FreeSans 224 90 0 0 la_data_out[45]
port 312 nsew signal tristate
flabel metal2 s 33138 0 33194 800 0 FreeSans 224 90 0 0 la_data_out[46]
port 313 nsew signal tristate
flabel metal2 s 33414 0 33470 800 0 FreeSans 224 90 0 0 la_data_out[47]
port 314 nsew signal tristate
flabel metal2 s 33690 0 33746 800 0 FreeSans 224 90 0 0 la_data_out[48]
port 315 nsew signal tristate
flabel metal2 s 33966 0 34022 800 0 FreeSans 224 90 0 0 la_data_out[49]
port 316 nsew signal tristate
flabel metal2 s 21546 0 21602 800 0 FreeSans 224 90 0 0 la_data_out[4]
port 317 nsew signal tristate
flabel metal2 s 34242 0 34298 800 0 FreeSans 224 90 0 0 la_data_out[50]
port 318 nsew signal tristate
flabel metal2 s 34518 0 34574 800 0 FreeSans 224 90 0 0 la_data_out[51]
port 319 nsew signal tristate
flabel metal2 s 34794 0 34850 800 0 FreeSans 224 90 0 0 la_data_out[52]
port 320 nsew signal tristate
flabel metal2 s 35070 0 35126 800 0 FreeSans 224 90 0 0 la_data_out[53]
port 321 nsew signal tristate
flabel metal2 s 35346 0 35402 800 0 FreeSans 224 90 0 0 la_data_out[54]
port 322 nsew signal tristate
flabel metal2 s 35622 0 35678 800 0 FreeSans 224 90 0 0 la_data_out[55]
port 323 nsew signal tristate
flabel metal2 s 35898 0 35954 800 0 FreeSans 224 90 0 0 la_data_out[56]
port 324 nsew signal tristate
flabel metal2 s 36174 0 36230 800 0 FreeSans 224 90 0 0 la_data_out[57]
port 325 nsew signal tristate
flabel metal2 s 36450 0 36506 800 0 FreeSans 224 90 0 0 la_data_out[58]
port 326 nsew signal tristate
flabel metal2 s 36726 0 36782 800 0 FreeSans 224 90 0 0 la_data_out[59]
port 327 nsew signal tristate
flabel metal2 s 21822 0 21878 800 0 FreeSans 224 90 0 0 la_data_out[5]
port 328 nsew signal tristate
flabel metal2 s 37002 0 37058 800 0 FreeSans 224 90 0 0 la_data_out[60]
port 329 nsew signal tristate
flabel metal2 s 37278 0 37334 800 0 FreeSans 224 90 0 0 la_data_out[61]
port 330 nsew signal tristate
flabel metal2 s 37554 0 37610 800 0 FreeSans 224 90 0 0 la_data_out[62]
port 331 nsew signal tristate
flabel metal2 s 37830 0 37886 800 0 FreeSans 224 90 0 0 la_data_out[63]
port 332 nsew signal tristate
flabel metal2 s 38106 0 38162 800 0 FreeSans 224 90 0 0 la_data_out[64]
port 333 nsew signal tristate
flabel metal2 s 38382 0 38438 800 0 FreeSans 224 90 0 0 la_data_out[65]
port 334 nsew signal tristate
flabel metal2 s 38658 0 38714 800 0 FreeSans 224 90 0 0 la_data_out[66]
port 335 nsew signal tristate
flabel metal2 s 38934 0 38990 800 0 FreeSans 224 90 0 0 la_data_out[67]
port 336 nsew signal tristate
flabel metal2 s 39210 0 39266 800 0 FreeSans 224 90 0 0 la_data_out[68]
port 337 nsew signal tristate
flabel metal2 s 39486 0 39542 800 0 FreeSans 224 90 0 0 la_data_out[69]
port 338 nsew signal tristate
flabel metal2 s 22098 0 22154 800 0 FreeSans 224 90 0 0 la_data_out[6]
port 339 nsew signal tristate
flabel metal2 s 39762 0 39818 800 0 FreeSans 224 90 0 0 la_data_out[70]
port 340 nsew signal tristate
flabel metal2 s 40038 0 40094 800 0 FreeSans 224 90 0 0 la_data_out[71]
port 341 nsew signal tristate
flabel metal2 s 40314 0 40370 800 0 FreeSans 224 90 0 0 la_data_out[72]
port 342 nsew signal tristate
flabel metal2 s 40590 0 40646 800 0 FreeSans 224 90 0 0 la_data_out[73]
port 343 nsew signal tristate
flabel metal2 s 40866 0 40922 800 0 FreeSans 224 90 0 0 la_data_out[74]
port 344 nsew signal tristate
flabel metal2 s 41142 0 41198 800 0 FreeSans 224 90 0 0 la_data_out[75]
port 345 nsew signal tristate
flabel metal2 s 41418 0 41474 800 0 FreeSans 224 90 0 0 la_data_out[76]
port 346 nsew signal tristate
flabel metal2 s 41694 0 41750 800 0 FreeSans 224 90 0 0 la_data_out[77]
port 347 nsew signal tristate
flabel metal2 s 41970 0 42026 800 0 FreeSans 224 90 0 0 la_data_out[78]
port 348 nsew signal tristate
flabel metal2 s 42246 0 42302 800 0 FreeSans 224 90 0 0 la_data_out[79]
port 349 nsew signal tristate
flabel metal2 s 22374 0 22430 800 0 FreeSans 224 90 0 0 la_data_out[7]
port 350 nsew signal tristate
flabel metal2 s 42522 0 42578 800 0 FreeSans 224 90 0 0 la_data_out[80]
port 351 nsew signal tristate
flabel metal2 s 42798 0 42854 800 0 FreeSans 224 90 0 0 la_data_out[81]
port 352 nsew signal tristate
flabel metal2 s 43074 0 43130 800 0 FreeSans 224 90 0 0 la_data_out[82]
port 353 nsew signal tristate
flabel metal2 s 43350 0 43406 800 0 FreeSans 224 90 0 0 la_data_out[83]
port 354 nsew signal tristate
flabel metal2 s 43626 0 43682 800 0 FreeSans 224 90 0 0 la_data_out[84]
port 355 nsew signal tristate
flabel metal2 s 43902 0 43958 800 0 FreeSans 224 90 0 0 la_data_out[85]
port 356 nsew signal tristate
flabel metal2 s 44178 0 44234 800 0 FreeSans 224 90 0 0 la_data_out[86]
port 357 nsew signal tristate
flabel metal2 s 44454 0 44510 800 0 FreeSans 224 90 0 0 la_data_out[87]
port 358 nsew signal tristate
flabel metal2 s 44730 0 44786 800 0 FreeSans 224 90 0 0 la_data_out[88]
port 359 nsew signal tristate
flabel metal2 s 45006 0 45062 800 0 FreeSans 224 90 0 0 la_data_out[89]
port 360 nsew signal tristate
flabel metal2 s 22650 0 22706 800 0 FreeSans 224 90 0 0 la_data_out[8]
port 361 nsew signal tristate
flabel metal2 s 45282 0 45338 800 0 FreeSans 224 90 0 0 la_data_out[90]
port 362 nsew signal tristate
flabel metal2 s 45558 0 45614 800 0 FreeSans 224 90 0 0 la_data_out[91]
port 363 nsew signal tristate
flabel metal2 s 45834 0 45890 800 0 FreeSans 224 90 0 0 la_data_out[92]
port 364 nsew signal tristate
flabel metal2 s 46110 0 46166 800 0 FreeSans 224 90 0 0 la_data_out[93]
port 365 nsew signal tristate
flabel metal2 s 46386 0 46442 800 0 FreeSans 224 90 0 0 la_data_out[94]
port 366 nsew signal tristate
flabel metal2 s 46662 0 46718 800 0 FreeSans 224 90 0 0 la_data_out[95]
port 367 nsew signal tristate
flabel metal2 s 46938 0 46994 800 0 FreeSans 224 90 0 0 la_data_out[96]
port 368 nsew signal tristate
flabel metal2 s 47214 0 47270 800 0 FreeSans 224 90 0 0 la_data_out[97]
port 369 nsew signal tristate
flabel metal2 s 47490 0 47546 800 0 FreeSans 224 90 0 0 la_data_out[98]
port 370 nsew signal tristate
flabel metal2 s 47766 0 47822 800 0 FreeSans 224 90 0 0 la_data_out[99]
port 371 nsew signal tristate
flabel metal2 s 22926 0 22982 800 0 FreeSans 224 90 0 0 la_data_out[9]
port 372 nsew signal tristate
flabel metal2 s 20534 0 20590 800 0 FreeSans 224 90 0 0 la_oenb[0]
port 373 nsew signal input
flabel metal2 s 48134 0 48190 800 0 FreeSans 224 90 0 0 la_oenb[100]
port 374 nsew signal input
flabel metal2 s 48410 0 48466 800 0 FreeSans 224 90 0 0 la_oenb[101]
port 375 nsew signal input
flabel metal2 s 48686 0 48742 800 0 FreeSans 224 90 0 0 la_oenb[102]
port 376 nsew signal input
flabel metal2 s 48962 0 49018 800 0 FreeSans 224 90 0 0 la_oenb[103]
port 377 nsew signal input
flabel metal2 s 49238 0 49294 800 0 FreeSans 224 90 0 0 la_oenb[104]
port 378 nsew signal input
flabel metal2 s 49514 0 49570 800 0 FreeSans 224 90 0 0 la_oenb[105]
port 379 nsew signal input
flabel metal2 s 49790 0 49846 800 0 FreeSans 224 90 0 0 la_oenb[106]
port 380 nsew signal input
flabel metal2 s 50066 0 50122 800 0 FreeSans 224 90 0 0 la_oenb[107]
port 381 nsew signal input
flabel metal2 s 50342 0 50398 800 0 FreeSans 224 90 0 0 la_oenb[108]
port 382 nsew signal input
flabel metal2 s 50618 0 50674 800 0 FreeSans 224 90 0 0 la_oenb[109]
port 383 nsew signal input
flabel metal2 s 23294 0 23350 800 0 FreeSans 224 90 0 0 la_oenb[10]
port 384 nsew signal input
flabel metal2 s 50894 0 50950 800 0 FreeSans 224 90 0 0 la_oenb[110]
port 385 nsew signal input
flabel metal2 s 51170 0 51226 800 0 FreeSans 224 90 0 0 la_oenb[111]
port 386 nsew signal input
flabel metal2 s 51446 0 51502 800 0 FreeSans 224 90 0 0 la_oenb[112]
port 387 nsew signal input
flabel metal2 s 51722 0 51778 800 0 FreeSans 224 90 0 0 la_oenb[113]
port 388 nsew signal input
flabel metal2 s 51998 0 52054 800 0 FreeSans 224 90 0 0 la_oenb[114]
port 389 nsew signal input
flabel metal2 s 52274 0 52330 800 0 FreeSans 224 90 0 0 la_oenb[115]
port 390 nsew signal input
flabel metal2 s 52550 0 52606 800 0 FreeSans 224 90 0 0 la_oenb[116]
port 391 nsew signal input
flabel metal2 s 52826 0 52882 800 0 FreeSans 224 90 0 0 la_oenb[117]
port 392 nsew signal input
flabel metal2 s 53102 0 53158 800 0 FreeSans 224 90 0 0 la_oenb[118]
port 393 nsew signal input
flabel metal2 s 53378 0 53434 800 0 FreeSans 224 90 0 0 la_oenb[119]
port 394 nsew signal input
flabel metal2 s 23570 0 23626 800 0 FreeSans 224 90 0 0 la_oenb[11]
port 395 nsew signal input
flabel metal2 s 53654 0 53710 800 0 FreeSans 224 90 0 0 la_oenb[120]
port 396 nsew signal input
flabel metal2 s 53930 0 53986 800 0 FreeSans 224 90 0 0 la_oenb[121]
port 397 nsew signal input
flabel metal2 s 54206 0 54262 800 0 FreeSans 224 90 0 0 la_oenb[122]
port 398 nsew signal input
flabel metal2 s 54482 0 54538 800 0 FreeSans 224 90 0 0 la_oenb[123]
port 399 nsew signal input
flabel metal2 s 54758 0 54814 800 0 FreeSans 224 90 0 0 la_oenb[124]
port 400 nsew signal input
flabel metal2 s 55034 0 55090 800 0 FreeSans 224 90 0 0 la_oenb[125]
port 401 nsew signal input
flabel metal2 s 55310 0 55366 800 0 FreeSans 224 90 0 0 la_oenb[126]
port 402 nsew signal input
flabel metal2 s 55586 0 55642 800 0 FreeSans 224 90 0 0 la_oenb[127]
port 403 nsew signal input
flabel metal2 s 23846 0 23902 800 0 FreeSans 224 90 0 0 la_oenb[12]
port 404 nsew signal input
flabel metal2 s 24122 0 24178 800 0 FreeSans 224 90 0 0 la_oenb[13]
port 405 nsew signal input
flabel metal2 s 24398 0 24454 800 0 FreeSans 224 90 0 0 la_oenb[14]
port 406 nsew signal input
flabel metal2 s 24674 0 24730 800 0 FreeSans 224 90 0 0 la_oenb[15]
port 407 nsew signal input
flabel metal2 s 24950 0 25006 800 0 FreeSans 224 90 0 0 la_oenb[16]
port 408 nsew signal input
flabel metal2 s 25226 0 25282 800 0 FreeSans 224 90 0 0 la_oenb[17]
port 409 nsew signal input
flabel metal2 s 25502 0 25558 800 0 FreeSans 224 90 0 0 la_oenb[18]
port 410 nsew signal input
flabel metal2 s 25778 0 25834 800 0 FreeSans 224 90 0 0 la_oenb[19]
port 411 nsew signal input
flabel metal2 s 20810 0 20866 800 0 FreeSans 224 90 0 0 la_oenb[1]
port 412 nsew signal input
flabel metal2 s 26054 0 26110 800 0 FreeSans 224 90 0 0 la_oenb[20]
port 413 nsew signal input
flabel metal2 s 26330 0 26386 800 0 FreeSans 224 90 0 0 la_oenb[21]
port 414 nsew signal input
flabel metal2 s 26606 0 26662 800 0 FreeSans 224 90 0 0 la_oenb[22]
port 415 nsew signal input
flabel metal2 s 26882 0 26938 800 0 FreeSans 224 90 0 0 la_oenb[23]
port 416 nsew signal input
flabel metal2 s 27158 0 27214 800 0 FreeSans 224 90 0 0 la_oenb[24]
port 417 nsew signal input
flabel metal2 s 27434 0 27490 800 0 FreeSans 224 90 0 0 la_oenb[25]
port 418 nsew signal input
flabel metal2 s 27710 0 27766 800 0 FreeSans 224 90 0 0 la_oenb[26]
port 419 nsew signal input
flabel metal2 s 27986 0 28042 800 0 FreeSans 224 90 0 0 la_oenb[27]
port 420 nsew signal input
flabel metal2 s 28262 0 28318 800 0 FreeSans 224 90 0 0 la_oenb[28]
port 421 nsew signal input
flabel metal2 s 28538 0 28594 800 0 FreeSans 224 90 0 0 la_oenb[29]
port 422 nsew signal input
flabel metal2 s 21086 0 21142 800 0 FreeSans 224 90 0 0 la_oenb[2]
port 423 nsew signal input
flabel metal2 s 28814 0 28870 800 0 FreeSans 224 90 0 0 la_oenb[30]
port 424 nsew signal input
flabel metal2 s 29090 0 29146 800 0 FreeSans 224 90 0 0 la_oenb[31]
port 425 nsew signal input
flabel metal2 s 29366 0 29422 800 0 FreeSans 224 90 0 0 la_oenb[32]
port 426 nsew signal input
flabel metal2 s 29642 0 29698 800 0 FreeSans 224 90 0 0 la_oenb[33]
port 427 nsew signal input
flabel metal2 s 29918 0 29974 800 0 FreeSans 224 90 0 0 la_oenb[34]
port 428 nsew signal input
flabel metal2 s 30194 0 30250 800 0 FreeSans 224 90 0 0 la_oenb[35]
port 429 nsew signal input
flabel metal2 s 30470 0 30526 800 0 FreeSans 224 90 0 0 la_oenb[36]
port 430 nsew signal input
flabel metal2 s 30746 0 30802 800 0 FreeSans 224 90 0 0 la_oenb[37]
port 431 nsew signal input
flabel metal2 s 31022 0 31078 800 0 FreeSans 224 90 0 0 la_oenb[38]
port 432 nsew signal input
flabel metal2 s 31298 0 31354 800 0 FreeSans 224 90 0 0 la_oenb[39]
port 433 nsew signal input
flabel metal2 s 21362 0 21418 800 0 FreeSans 224 90 0 0 la_oenb[3]
port 434 nsew signal input
flabel metal2 s 31574 0 31630 800 0 FreeSans 224 90 0 0 la_oenb[40]
port 435 nsew signal input
flabel metal2 s 31850 0 31906 800 0 FreeSans 224 90 0 0 la_oenb[41]
port 436 nsew signal input
flabel metal2 s 32126 0 32182 800 0 FreeSans 224 90 0 0 la_oenb[42]
port 437 nsew signal input
flabel metal2 s 32402 0 32458 800 0 FreeSans 224 90 0 0 la_oenb[43]
port 438 nsew signal input
flabel metal2 s 32678 0 32734 800 0 FreeSans 224 90 0 0 la_oenb[44]
port 439 nsew signal input
flabel metal2 s 32954 0 33010 800 0 FreeSans 224 90 0 0 la_oenb[45]
port 440 nsew signal input
flabel metal2 s 33230 0 33286 800 0 FreeSans 224 90 0 0 la_oenb[46]
port 441 nsew signal input
flabel metal2 s 33506 0 33562 800 0 FreeSans 224 90 0 0 la_oenb[47]
port 442 nsew signal input
flabel metal2 s 33782 0 33838 800 0 FreeSans 224 90 0 0 la_oenb[48]
port 443 nsew signal input
flabel metal2 s 34058 0 34114 800 0 FreeSans 224 90 0 0 la_oenb[49]
port 444 nsew signal input
flabel metal2 s 21638 0 21694 800 0 FreeSans 224 90 0 0 la_oenb[4]
port 445 nsew signal input
flabel metal2 s 34334 0 34390 800 0 FreeSans 224 90 0 0 la_oenb[50]
port 446 nsew signal input
flabel metal2 s 34610 0 34666 800 0 FreeSans 224 90 0 0 la_oenb[51]
port 447 nsew signal input
flabel metal2 s 34886 0 34942 800 0 FreeSans 224 90 0 0 la_oenb[52]
port 448 nsew signal input
flabel metal2 s 35162 0 35218 800 0 FreeSans 224 90 0 0 la_oenb[53]
port 449 nsew signal input
flabel metal2 s 35438 0 35494 800 0 FreeSans 224 90 0 0 la_oenb[54]
port 450 nsew signal input
flabel metal2 s 35714 0 35770 800 0 FreeSans 224 90 0 0 la_oenb[55]
port 451 nsew signal input
flabel metal2 s 35990 0 36046 800 0 FreeSans 224 90 0 0 la_oenb[56]
port 452 nsew signal input
flabel metal2 s 36266 0 36322 800 0 FreeSans 224 90 0 0 la_oenb[57]
port 453 nsew signal input
flabel metal2 s 36542 0 36598 800 0 FreeSans 224 90 0 0 la_oenb[58]
port 454 nsew signal input
flabel metal2 s 36818 0 36874 800 0 FreeSans 224 90 0 0 la_oenb[59]
port 455 nsew signal input
flabel metal2 s 21914 0 21970 800 0 FreeSans 224 90 0 0 la_oenb[5]
port 456 nsew signal input
flabel metal2 s 37094 0 37150 800 0 FreeSans 224 90 0 0 la_oenb[60]
port 457 nsew signal input
flabel metal2 s 37370 0 37426 800 0 FreeSans 224 90 0 0 la_oenb[61]
port 458 nsew signal input
flabel metal2 s 37646 0 37702 800 0 FreeSans 224 90 0 0 la_oenb[62]
port 459 nsew signal input
flabel metal2 s 37922 0 37978 800 0 FreeSans 224 90 0 0 la_oenb[63]
port 460 nsew signal input
flabel metal2 s 38198 0 38254 800 0 FreeSans 224 90 0 0 la_oenb[64]
port 461 nsew signal input
flabel metal2 s 38474 0 38530 800 0 FreeSans 224 90 0 0 la_oenb[65]
port 462 nsew signal input
flabel metal2 s 38750 0 38806 800 0 FreeSans 224 90 0 0 la_oenb[66]
port 463 nsew signal input
flabel metal2 s 39026 0 39082 800 0 FreeSans 224 90 0 0 la_oenb[67]
port 464 nsew signal input
flabel metal2 s 39302 0 39358 800 0 FreeSans 224 90 0 0 la_oenb[68]
port 465 nsew signal input
flabel metal2 s 39578 0 39634 800 0 FreeSans 224 90 0 0 la_oenb[69]
port 466 nsew signal input
flabel metal2 s 22190 0 22246 800 0 FreeSans 224 90 0 0 la_oenb[6]
port 467 nsew signal input
flabel metal2 s 39854 0 39910 800 0 FreeSans 224 90 0 0 la_oenb[70]
port 468 nsew signal input
flabel metal2 s 40130 0 40186 800 0 FreeSans 224 90 0 0 la_oenb[71]
port 469 nsew signal input
flabel metal2 s 40406 0 40462 800 0 FreeSans 224 90 0 0 la_oenb[72]
port 470 nsew signal input
flabel metal2 s 40682 0 40738 800 0 FreeSans 224 90 0 0 la_oenb[73]
port 471 nsew signal input
flabel metal2 s 40958 0 41014 800 0 FreeSans 224 90 0 0 la_oenb[74]
port 472 nsew signal input
flabel metal2 s 41234 0 41290 800 0 FreeSans 224 90 0 0 la_oenb[75]
port 473 nsew signal input
flabel metal2 s 41510 0 41566 800 0 FreeSans 224 90 0 0 la_oenb[76]
port 474 nsew signal input
flabel metal2 s 41786 0 41842 800 0 FreeSans 224 90 0 0 la_oenb[77]
port 475 nsew signal input
flabel metal2 s 42062 0 42118 800 0 FreeSans 224 90 0 0 la_oenb[78]
port 476 nsew signal input
flabel metal2 s 42338 0 42394 800 0 FreeSans 224 90 0 0 la_oenb[79]
port 477 nsew signal input
flabel metal2 s 22466 0 22522 800 0 FreeSans 224 90 0 0 la_oenb[7]
port 478 nsew signal input
flabel metal2 s 42614 0 42670 800 0 FreeSans 224 90 0 0 la_oenb[80]
port 479 nsew signal input
flabel metal2 s 42890 0 42946 800 0 FreeSans 224 90 0 0 la_oenb[81]
port 480 nsew signal input
flabel metal2 s 43166 0 43222 800 0 FreeSans 224 90 0 0 la_oenb[82]
port 481 nsew signal input
flabel metal2 s 43442 0 43498 800 0 FreeSans 224 90 0 0 la_oenb[83]
port 482 nsew signal input
flabel metal2 s 43718 0 43774 800 0 FreeSans 224 90 0 0 la_oenb[84]
port 483 nsew signal input
flabel metal2 s 43994 0 44050 800 0 FreeSans 224 90 0 0 la_oenb[85]
port 484 nsew signal input
flabel metal2 s 44270 0 44326 800 0 FreeSans 224 90 0 0 la_oenb[86]
port 485 nsew signal input
flabel metal2 s 44546 0 44602 800 0 FreeSans 224 90 0 0 la_oenb[87]
port 486 nsew signal input
flabel metal2 s 44822 0 44878 800 0 FreeSans 224 90 0 0 la_oenb[88]
port 487 nsew signal input
flabel metal2 s 45098 0 45154 800 0 FreeSans 224 90 0 0 la_oenb[89]
port 488 nsew signal input
flabel metal2 s 22742 0 22798 800 0 FreeSans 224 90 0 0 la_oenb[8]
port 489 nsew signal input
flabel metal2 s 45374 0 45430 800 0 FreeSans 224 90 0 0 la_oenb[90]
port 490 nsew signal input
flabel metal2 s 45650 0 45706 800 0 FreeSans 224 90 0 0 la_oenb[91]
port 491 nsew signal input
flabel metal2 s 45926 0 45982 800 0 FreeSans 224 90 0 0 la_oenb[92]
port 492 nsew signal input
flabel metal2 s 46202 0 46258 800 0 FreeSans 224 90 0 0 la_oenb[93]
port 493 nsew signal input
flabel metal2 s 46478 0 46534 800 0 FreeSans 224 90 0 0 la_oenb[94]
port 494 nsew signal input
flabel metal2 s 46754 0 46810 800 0 FreeSans 224 90 0 0 la_oenb[95]
port 495 nsew signal input
flabel metal2 s 47030 0 47086 800 0 FreeSans 224 90 0 0 la_oenb[96]
port 496 nsew signal input
flabel metal2 s 47306 0 47362 800 0 FreeSans 224 90 0 0 la_oenb[97]
port 497 nsew signal input
flabel metal2 s 47582 0 47638 800 0 FreeSans 224 90 0 0 la_oenb[98]
port 498 nsew signal input
flabel metal2 s 47858 0 47914 800 0 FreeSans 224 90 0 0 la_oenb[99]
port 499 nsew signal input
flabel metal2 s 23018 0 23074 800 0 FreeSans 224 90 0 0 la_oenb[9]
port 500 nsew signal input
flabel metal2 s 21822 59200 21878 60000 0 FreeSans 224 90 0 0 out_1
port 501 nsew signal tristate
flabel metal2 s 30562 59200 30618 60000 0 FreeSans 224 90 0 0 out_2
port 502 nsew signal tristate
flabel metal2 s 39302 59200 39358 60000 0 FreeSans 224 90 0 0 out_3
port 503 nsew signal tristate
flabel metal2 s 48042 59200 48098 60000 0 FreeSans 224 90 0 0 out_4
port 504 nsew signal tristate
flabel metal2 s 56782 59200 56838 60000 0 FreeSans 224 90 0 0 out_5
port 505 nsew signal tristate
flabel metal2 s 65522 59200 65578 60000 0 FreeSans 224 90 0 0 out_7
port 506 nsew signal tristate
flabel metal2 s 13082 59200 13138 60000 0 FreeSans 224 90 0 0 rst_o
port 507 nsew signal tristate
flabel metal2 s 4342 59200 4398 60000 0 FreeSans 224 90 0 0 serial_data_rlbp_out
port 508 nsew signal tristate
flabel metal4 s 4208 2128 4528 57712 0 FreeSans 1920 90 0 0 vccd1
port 509 nsew power bidirectional
flabel metal4 s 34928 2128 35248 57712 0 FreeSans 1920 90 0 0 vccd1
port 509 nsew power bidirectional
flabel metal4 s 65648 2128 65968 57712 0 FreeSans 1920 90 0 0 vccd1
port 509 nsew power bidirectional
flabel metal4 s 19568 2128 19888 57712 0 FreeSans 1920 90 0 0 vssd1
port 510 nsew ground bidirectional
flabel metal4 s 50288 2128 50608 57712 0 FreeSans 1920 90 0 0 vssd1
port 510 nsew ground bidirectional
flabel metal2 s 10598 0 10654 800 0 FreeSans 224 90 0 0 wb_clk_i
port 511 nsew signal input
flabel metal2 s 10690 0 10746 800 0 FreeSans 224 90 0 0 wb_rst_i
port 512 nsew signal input
flabel metal2 s 10782 0 10838 800 0 FreeSans 224 90 0 0 wbs_ack_o
port 513 nsew signal tristate
flabel metal2 s 11150 0 11206 800 0 FreeSans 224 90 0 0 wbs_adr_i[0]
port 514 nsew signal input
flabel metal2 s 14278 0 14334 800 0 FreeSans 224 90 0 0 wbs_adr_i[10]
port 515 nsew signal input
flabel metal2 s 14554 0 14610 800 0 FreeSans 224 90 0 0 wbs_adr_i[11]
port 516 nsew signal input
flabel metal2 s 14830 0 14886 800 0 FreeSans 224 90 0 0 wbs_adr_i[12]
port 517 nsew signal input
flabel metal2 s 15106 0 15162 800 0 FreeSans 224 90 0 0 wbs_adr_i[13]
port 518 nsew signal input
flabel metal2 s 15382 0 15438 800 0 FreeSans 224 90 0 0 wbs_adr_i[14]
port 519 nsew signal input
flabel metal2 s 15658 0 15714 800 0 FreeSans 224 90 0 0 wbs_adr_i[15]
port 520 nsew signal input
flabel metal2 s 15934 0 15990 800 0 FreeSans 224 90 0 0 wbs_adr_i[16]
port 521 nsew signal input
flabel metal2 s 16210 0 16266 800 0 FreeSans 224 90 0 0 wbs_adr_i[17]
port 522 nsew signal input
flabel metal2 s 16486 0 16542 800 0 FreeSans 224 90 0 0 wbs_adr_i[18]
port 523 nsew signal input
flabel metal2 s 16762 0 16818 800 0 FreeSans 224 90 0 0 wbs_adr_i[19]
port 524 nsew signal input
flabel metal2 s 11518 0 11574 800 0 FreeSans 224 90 0 0 wbs_adr_i[1]
port 525 nsew signal input
flabel metal2 s 17038 0 17094 800 0 FreeSans 224 90 0 0 wbs_adr_i[20]
port 526 nsew signal input
flabel metal2 s 17314 0 17370 800 0 FreeSans 224 90 0 0 wbs_adr_i[21]
port 527 nsew signal input
flabel metal2 s 17590 0 17646 800 0 FreeSans 224 90 0 0 wbs_adr_i[22]
port 528 nsew signal input
flabel metal2 s 17866 0 17922 800 0 FreeSans 224 90 0 0 wbs_adr_i[23]
port 529 nsew signal input
flabel metal2 s 18142 0 18198 800 0 FreeSans 224 90 0 0 wbs_adr_i[24]
port 530 nsew signal input
flabel metal2 s 18418 0 18474 800 0 FreeSans 224 90 0 0 wbs_adr_i[25]
port 531 nsew signal input
flabel metal2 s 18694 0 18750 800 0 FreeSans 224 90 0 0 wbs_adr_i[26]
port 532 nsew signal input
flabel metal2 s 18970 0 19026 800 0 FreeSans 224 90 0 0 wbs_adr_i[27]
port 533 nsew signal input
flabel metal2 s 19246 0 19302 800 0 FreeSans 224 90 0 0 wbs_adr_i[28]
port 534 nsew signal input
flabel metal2 s 19522 0 19578 800 0 FreeSans 224 90 0 0 wbs_adr_i[29]
port 535 nsew signal input
flabel metal2 s 11886 0 11942 800 0 FreeSans 224 90 0 0 wbs_adr_i[2]
port 536 nsew signal input
flabel metal2 s 19798 0 19854 800 0 FreeSans 224 90 0 0 wbs_adr_i[30]
port 537 nsew signal input
flabel metal2 s 20074 0 20130 800 0 FreeSans 224 90 0 0 wbs_adr_i[31]
port 538 nsew signal input
flabel metal2 s 12254 0 12310 800 0 FreeSans 224 90 0 0 wbs_adr_i[3]
port 539 nsew signal input
flabel metal2 s 12622 0 12678 800 0 FreeSans 224 90 0 0 wbs_adr_i[4]
port 540 nsew signal input
flabel metal2 s 12898 0 12954 800 0 FreeSans 224 90 0 0 wbs_adr_i[5]
port 541 nsew signal input
flabel metal2 s 13174 0 13230 800 0 FreeSans 224 90 0 0 wbs_adr_i[6]
port 542 nsew signal input
flabel metal2 s 13450 0 13506 800 0 FreeSans 224 90 0 0 wbs_adr_i[7]
port 543 nsew signal input
flabel metal2 s 13726 0 13782 800 0 FreeSans 224 90 0 0 wbs_adr_i[8]
port 544 nsew signal input
flabel metal2 s 14002 0 14058 800 0 FreeSans 224 90 0 0 wbs_adr_i[9]
port 545 nsew signal input
flabel metal2 s 10874 0 10930 800 0 FreeSans 224 90 0 0 wbs_cyc_i
port 546 nsew signal input
flabel metal2 s 11242 0 11298 800 0 FreeSans 224 90 0 0 wbs_dat_i[0]
port 547 nsew signal input
flabel metal2 s 14370 0 14426 800 0 FreeSans 224 90 0 0 wbs_dat_i[10]
port 548 nsew signal input
flabel metal2 s 14646 0 14702 800 0 FreeSans 224 90 0 0 wbs_dat_i[11]
port 549 nsew signal input
flabel metal2 s 14922 0 14978 800 0 FreeSans 224 90 0 0 wbs_dat_i[12]
port 550 nsew signal input
flabel metal2 s 15198 0 15254 800 0 FreeSans 224 90 0 0 wbs_dat_i[13]
port 551 nsew signal input
flabel metal2 s 15474 0 15530 800 0 FreeSans 224 90 0 0 wbs_dat_i[14]
port 552 nsew signal input
flabel metal2 s 15750 0 15806 800 0 FreeSans 224 90 0 0 wbs_dat_i[15]
port 553 nsew signal input
flabel metal2 s 16026 0 16082 800 0 FreeSans 224 90 0 0 wbs_dat_i[16]
port 554 nsew signal input
flabel metal2 s 16302 0 16358 800 0 FreeSans 224 90 0 0 wbs_dat_i[17]
port 555 nsew signal input
flabel metal2 s 16578 0 16634 800 0 FreeSans 224 90 0 0 wbs_dat_i[18]
port 556 nsew signal input
flabel metal2 s 16854 0 16910 800 0 FreeSans 224 90 0 0 wbs_dat_i[19]
port 557 nsew signal input
flabel metal2 s 11610 0 11666 800 0 FreeSans 224 90 0 0 wbs_dat_i[1]
port 558 nsew signal input
flabel metal2 s 17130 0 17186 800 0 FreeSans 224 90 0 0 wbs_dat_i[20]
port 559 nsew signal input
flabel metal2 s 17406 0 17462 800 0 FreeSans 224 90 0 0 wbs_dat_i[21]
port 560 nsew signal input
flabel metal2 s 17682 0 17738 800 0 FreeSans 224 90 0 0 wbs_dat_i[22]
port 561 nsew signal input
flabel metal2 s 17958 0 18014 800 0 FreeSans 224 90 0 0 wbs_dat_i[23]
port 562 nsew signal input
flabel metal2 s 18234 0 18290 800 0 FreeSans 224 90 0 0 wbs_dat_i[24]
port 563 nsew signal input
flabel metal2 s 18510 0 18566 800 0 FreeSans 224 90 0 0 wbs_dat_i[25]
port 564 nsew signal input
flabel metal2 s 18786 0 18842 800 0 FreeSans 224 90 0 0 wbs_dat_i[26]
port 565 nsew signal input
flabel metal2 s 19062 0 19118 800 0 FreeSans 224 90 0 0 wbs_dat_i[27]
port 566 nsew signal input
flabel metal2 s 19338 0 19394 800 0 FreeSans 224 90 0 0 wbs_dat_i[28]
port 567 nsew signal input
flabel metal2 s 19614 0 19670 800 0 FreeSans 224 90 0 0 wbs_dat_i[29]
port 568 nsew signal input
flabel metal2 s 11978 0 12034 800 0 FreeSans 224 90 0 0 wbs_dat_i[2]
port 569 nsew signal input
flabel metal2 s 19890 0 19946 800 0 FreeSans 224 90 0 0 wbs_dat_i[30]
port 570 nsew signal input
flabel metal2 s 20166 0 20222 800 0 FreeSans 224 90 0 0 wbs_dat_i[31]
port 571 nsew signal input
flabel metal2 s 12346 0 12402 800 0 FreeSans 224 90 0 0 wbs_dat_i[3]
port 572 nsew signal input
flabel metal2 s 12714 0 12770 800 0 FreeSans 224 90 0 0 wbs_dat_i[4]
port 573 nsew signal input
flabel metal2 s 12990 0 13046 800 0 FreeSans 224 90 0 0 wbs_dat_i[5]
port 574 nsew signal input
flabel metal2 s 13266 0 13322 800 0 FreeSans 224 90 0 0 wbs_dat_i[6]
port 575 nsew signal input
flabel metal2 s 13542 0 13598 800 0 FreeSans 224 90 0 0 wbs_dat_i[7]
port 576 nsew signal input
flabel metal2 s 13818 0 13874 800 0 FreeSans 224 90 0 0 wbs_dat_i[8]
port 577 nsew signal input
flabel metal2 s 14094 0 14150 800 0 FreeSans 224 90 0 0 wbs_dat_i[9]
port 578 nsew signal input
flabel metal2 s 11334 0 11390 800 0 FreeSans 224 90 0 0 wbs_dat_o[0]
port 579 nsew signal tristate
flabel metal2 s 14462 0 14518 800 0 FreeSans 224 90 0 0 wbs_dat_o[10]
port 580 nsew signal tristate
flabel metal2 s 14738 0 14794 800 0 FreeSans 224 90 0 0 wbs_dat_o[11]
port 581 nsew signal tristate
flabel metal2 s 15014 0 15070 800 0 FreeSans 224 90 0 0 wbs_dat_o[12]
port 582 nsew signal tristate
flabel metal2 s 15290 0 15346 800 0 FreeSans 224 90 0 0 wbs_dat_o[13]
port 583 nsew signal tristate
flabel metal2 s 15566 0 15622 800 0 FreeSans 224 90 0 0 wbs_dat_o[14]
port 584 nsew signal tristate
flabel metal2 s 15842 0 15898 800 0 FreeSans 224 90 0 0 wbs_dat_o[15]
port 585 nsew signal tristate
flabel metal2 s 16118 0 16174 800 0 FreeSans 224 90 0 0 wbs_dat_o[16]
port 586 nsew signal tristate
flabel metal2 s 16394 0 16450 800 0 FreeSans 224 90 0 0 wbs_dat_o[17]
port 587 nsew signal tristate
flabel metal2 s 16670 0 16726 800 0 FreeSans 224 90 0 0 wbs_dat_o[18]
port 588 nsew signal tristate
flabel metal2 s 16946 0 17002 800 0 FreeSans 224 90 0 0 wbs_dat_o[19]
port 589 nsew signal tristate
flabel metal2 s 11702 0 11758 800 0 FreeSans 224 90 0 0 wbs_dat_o[1]
port 590 nsew signal tristate
flabel metal2 s 17222 0 17278 800 0 FreeSans 224 90 0 0 wbs_dat_o[20]
port 591 nsew signal tristate
flabel metal2 s 17498 0 17554 800 0 FreeSans 224 90 0 0 wbs_dat_o[21]
port 592 nsew signal tristate
flabel metal2 s 17774 0 17830 800 0 FreeSans 224 90 0 0 wbs_dat_o[22]
port 593 nsew signal tristate
flabel metal2 s 18050 0 18106 800 0 FreeSans 224 90 0 0 wbs_dat_o[23]
port 594 nsew signal tristate
flabel metal2 s 18326 0 18382 800 0 FreeSans 224 90 0 0 wbs_dat_o[24]
port 595 nsew signal tristate
flabel metal2 s 18602 0 18658 800 0 FreeSans 224 90 0 0 wbs_dat_o[25]
port 596 nsew signal tristate
flabel metal2 s 18878 0 18934 800 0 FreeSans 224 90 0 0 wbs_dat_o[26]
port 597 nsew signal tristate
flabel metal2 s 19154 0 19210 800 0 FreeSans 224 90 0 0 wbs_dat_o[27]
port 598 nsew signal tristate
flabel metal2 s 19430 0 19486 800 0 FreeSans 224 90 0 0 wbs_dat_o[28]
port 599 nsew signal tristate
flabel metal2 s 19706 0 19762 800 0 FreeSans 224 90 0 0 wbs_dat_o[29]
port 600 nsew signal tristate
flabel metal2 s 12070 0 12126 800 0 FreeSans 224 90 0 0 wbs_dat_o[2]
port 601 nsew signal tristate
flabel metal2 s 19982 0 20038 800 0 FreeSans 224 90 0 0 wbs_dat_o[30]
port 602 nsew signal tristate
flabel metal2 s 20258 0 20314 800 0 FreeSans 224 90 0 0 wbs_dat_o[31]
port 603 nsew signal tristate
flabel metal2 s 12438 0 12494 800 0 FreeSans 224 90 0 0 wbs_dat_o[3]
port 604 nsew signal tristate
flabel metal2 s 12806 0 12862 800 0 FreeSans 224 90 0 0 wbs_dat_o[4]
port 605 nsew signal tristate
flabel metal2 s 13082 0 13138 800 0 FreeSans 224 90 0 0 wbs_dat_o[5]
port 606 nsew signal tristate
flabel metal2 s 13358 0 13414 800 0 FreeSans 224 90 0 0 wbs_dat_o[6]
port 607 nsew signal tristate
flabel metal2 s 13634 0 13690 800 0 FreeSans 224 90 0 0 wbs_dat_o[7]
port 608 nsew signal tristate
flabel metal2 s 13910 0 13966 800 0 FreeSans 224 90 0 0 wbs_dat_o[8]
port 609 nsew signal tristate
flabel metal2 s 14186 0 14242 800 0 FreeSans 224 90 0 0 wbs_dat_o[9]
port 610 nsew signal tristate
flabel metal2 s 11426 0 11482 800 0 FreeSans 224 90 0 0 wbs_sel_i[0]
port 611 nsew signal input
flabel metal2 s 11794 0 11850 800 0 FreeSans 224 90 0 0 wbs_sel_i[1]
port 612 nsew signal input
flabel metal2 s 12162 0 12218 800 0 FreeSans 224 90 0 0 wbs_sel_i[2]
port 613 nsew signal input
flabel metal2 s 12530 0 12586 800 0 FreeSans 224 90 0 0 wbs_sel_i[3]
port 614 nsew signal input
flabel metal2 s 10966 0 11022 800 0 FreeSans 224 90 0 0 wbs_stb_i
port 615 nsew signal input
flabel metal2 s 11058 0 11114 800 0 FreeSans 224 90 0 0 wbs_we_i
port 616 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 70000 60000
<< end >>
