`default_nettype none

module muler(
    
`ifdef USE_POWER_PINS
    input   VDD,
    input   VSS,
`endif
    
    input  M,
    input  P,
    input  C,
    output OUT

);


endmodule
`default_nettype wire

