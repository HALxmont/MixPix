magic
tech sky130B
magscale 1 2
timestamp 1667828175
<< viali >>
rect 3249 57409 3283 57443
rect 4169 57409 4203 57443
rect 5181 57409 5215 57443
rect 5641 57409 5675 57443
rect 6837 57409 6871 57443
rect 7481 57409 7515 57443
rect 8401 57409 8435 57443
rect 9137 57409 9171 57443
rect 10149 57409 10183 57443
rect 10793 57409 10827 57443
rect 11805 57409 11839 57443
rect 12449 57409 12483 57443
rect 13369 57409 13403 57443
rect 14105 57409 14139 57443
rect 15117 57409 15151 57443
rect 15761 57409 15795 57443
rect 16773 57409 16807 57443
rect 17417 57409 17451 57443
rect 18521 57409 18555 57443
rect 19257 57409 19291 57443
rect 20085 57409 20119 57443
rect 20729 57409 20763 57443
rect 22385 57409 22419 57443
rect 23489 57409 23523 57443
rect 24409 57409 24443 57443
rect 25053 57409 25087 57443
rect 25697 57409 25731 57443
rect 27353 57409 27387 57443
rect 28365 57409 28399 57443
rect 28825 57409 28859 57443
rect 30021 57409 30055 57443
rect 30665 57409 30699 57443
rect 31585 57409 31619 57443
rect 32321 57409 32355 57443
rect 33333 57409 33367 57443
rect 33977 57409 34011 57443
rect 34989 57409 35023 57443
rect 35633 57409 35667 57443
rect 37289 57409 37323 57443
rect 38577 57409 38611 57443
rect 40049 57409 40083 57443
rect 40693 57409 40727 57443
rect 41705 57409 41739 57443
rect 42441 57409 42475 57443
rect 43361 57409 43395 57443
rect 44005 57409 44039 57443
rect 45017 57409 45051 57443
rect 46673 57409 46707 57443
rect 47593 57409 47627 57443
rect 48329 57409 48363 57443
rect 48973 57409 49007 57443
rect 50169 57409 50203 57443
rect 50813 57409 50847 57443
rect 51641 57409 51675 57443
rect 52745 57409 52779 57443
rect 53389 57409 53423 57443
rect 54033 57409 54067 57443
rect 55321 57409 55355 57443
rect 55965 57409 55999 57443
rect 56609 57409 56643 57443
rect 57897 57409 57931 57443
rect 58541 57409 58575 57443
rect 59185 57409 59219 57443
rect 60473 57409 60507 57443
rect 61117 57409 61151 57443
rect 61761 57409 61795 57443
rect 63233 57409 63267 57443
rect 63877 57409 63911 57443
rect 65625 57409 65659 57443
rect 67097 57409 67131 57443
rect 45661 57341 45695 57375
rect 64889 57341 64923 57375
rect 37933 57273 37967 57307
rect 21833 57001 21867 57035
rect 26801 57001 26835 57035
rect 38945 57001 38979 57035
rect 62129 57001 62163 57035
rect 11897 14365 11931 14399
rect 11989 14365 12023 14399
rect 12102 14359 12136 14393
rect 12265 14365 12299 14399
rect 15301 14365 15335 14399
rect 15390 14365 15424 14399
rect 15506 14365 15540 14399
rect 15669 14365 15703 14399
rect 11621 14229 11655 14263
rect 15025 14229 15059 14263
rect 4353 14025 4387 14059
rect 8401 14025 8435 14059
rect 14197 14025 14231 14059
rect 4261 13889 4295 13923
rect 4445 13889 4479 13923
rect 7297 13889 7331 13923
rect 8033 13889 8067 13923
rect 8861 13889 8895 13923
rect 10609 13889 10643 13923
rect 10698 13889 10732 13923
rect 10793 13892 10827 13926
rect 10977 13889 11011 13923
rect 12081 13889 12115 13923
rect 13093 13889 13127 13923
rect 13256 13889 13290 13923
rect 13369 13889 13403 13923
rect 13461 13889 13495 13923
rect 15025 13889 15059 13923
rect 4997 13821 5031 13855
rect 8125 13821 8159 13855
rect 8953 13821 8987 13855
rect 10333 13821 10367 13855
rect 12357 13821 12391 13855
rect 13737 13821 13771 13855
rect 14749 13821 14783 13855
rect 7481 13685 7515 13719
rect 8217 13685 8251 13719
rect 9045 13685 9079 13719
rect 9229 13685 9263 13719
rect 8125 13481 8159 13515
rect 9045 13481 9079 13515
rect 11529 13481 11563 13515
rect 8309 13413 8343 13447
rect 9321 13413 9355 13447
rect 7297 13277 7331 13311
rect 7941 13277 7975 13311
rect 8125 13277 8159 13311
rect 8953 13277 8987 13311
rect 9137 13277 9171 13311
rect 10563 13277 10597 13311
rect 10714 13271 10748 13305
rect 10814 13271 10848 13305
rect 10977 13277 11011 13311
rect 12817 13277 12851 13311
rect 12906 13277 12940 13311
rect 13006 13271 13040 13305
rect 13197 13277 13231 13311
rect 15393 13277 15427 13311
rect 15482 13277 15516 13311
rect 15577 13277 15611 13311
rect 15773 13277 15807 13311
rect 16451 13277 16485 13311
rect 16586 13274 16620 13308
rect 16686 13277 16720 13311
rect 16865 13277 16899 13311
rect 7481 13141 7515 13175
rect 10333 13141 10367 13175
rect 12541 13141 12575 13175
rect 15117 13141 15151 13175
rect 16221 13141 16255 13175
rect 9413 12937 9447 12971
rect 13728 12869 13762 12903
rect 4721 12801 4755 12835
rect 4900 12801 4934 12835
rect 4997 12801 5031 12835
rect 5135 12801 5169 12835
rect 9045 12801 9079 12835
rect 13461 12801 13495 12835
rect 15853 12801 15887 12835
rect 9137 12733 9171 12767
rect 16129 12733 16163 12767
rect 5365 12665 5399 12699
rect 7665 12597 7699 12631
rect 9045 12597 9079 12631
rect 14841 12597 14875 12631
rect 22845 12393 22879 12427
rect 20637 12325 20671 12359
rect 5273 12257 5307 12291
rect 5549 12189 5583 12223
rect 7021 12189 7055 12223
rect 10149 12189 10183 12223
rect 11989 12189 12023 12223
rect 12256 12189 12290 12223
rect 15485 12189 15519 12223
rect 17325 12189 17359 12223
rect 19257 12189 19291 12223
rect 21327 12189 21361 12223
rect 21462 12189 21496 12223
rect 21562 12189 21596 12223
rect 21741 12189 21775 12223
rect 22201 12189 22235 12223
rect 22380 12189 22414 12223
rect 22480 12189 22514 12223
rect 22569 12189 22603 12223
rect 7266 12121 7300 12155
rect 10416 12121 10450 12155
rect 15752 12121 15786 12155
rect 17592 12121 17626 12155
rect 19524 12121 19558 12155
rect 21097 12121 21131 12155
rect 8401 12053 8435 12087
rect 11529 12053 11563 12087
rect 13369 12053 13403 12087
rect 16865 12053 16899 12087
rect 18705 12053 18739 12087
rect 5365 11849 5399 11883
rect 9045 11849 9079 11883
rect 20637 11849 20671 11883
rect 10158 11781 10192 11815
rect 14924 11781 14958 11815
rect 4721 11713 4755 11747
rect 4884 11713 4918 11747
rect 4984 11713 5018 11747
rect 5089 11713 5123 11747
rect 7461 11713 7495 11747
rect 14657 11713 14691 11747
rect 18429 11713 18463 11747
rect 18696 11713 18730 11747
rect 20913 11713 20947 11747
rect 21005 11713 21039 11747
rect 21097 11713 21131 11747
rect 21281 11713 21315 11747
rect 7205 11645 7239 11679
rect 10425 11645 10459 11679
rect 8585 11509 8619 11543
rect 16037 11509 16071 11543
rect 19809 11509 19843 11543
rect 4445 11305 4479 11339
rect 4629 11305 4663 11339
rect 6377 11305 6411 11339
rect 10333 11305 10367 11339
rect 12173 11305 12207 11339
rect 22385 11305 22419 11339
rect 23213 11305 23247 11339
rect 22753 11237 22787 11271
rect 11713 11169 11747 11203
rect 13553 11169 13587 11203
rect 22477 11169 22511 11203
rect 4353 11101 4387 11135
rect 4445 11101 4479 11135
rect 5733 11101 5767 11135
rect 5912 11101 5946 11135
rect 6009 11101 6043 11135
rect 6101 11101 6135 11135
rect 11457 11101 11491 11135
rect 13297 11101 13331 11135
rect 22385 11101 22419 11135
rect 23397 11101 23431 11135
rect 23489 11101 23523 11135
rect 4169 11033 4203 11067
rect 23213 11033 23247 11067
rect 23673 10965 23707 10999
rect 4629 10761 4663 10795
rect 5825 10761 5859 10795
rect 10977 10761 11011 10795
rect 14381 10761 14415 10795
rect 20453 10761 20487 10795
rect 4169 10693 4203 10727
rect 9864 10693 9898 10727
rect 16681 10693 16715 10727
rect 24225 10693 24259 10727
rect 4445 10625 4479 10659
rect 5365 10625 5399 10659
rect 5641 10625 5675 10659
rect 6377 10625 6411 10659
rect 6561 10631 6595 10665
rect 6653 10625 6687 10659
rect 6745 10625 6779 10659
rect 7757 10625 7791 10659
rect 8013 10625 8047 10659
rect 9597 10625 9631 10659
rect 13001 10625 13035 10659
rect 13268 10625 13302 10659
rect 16937 10625 16971 10659
rect 17046 10625 17080 10659
rect 17141 10628 17175 10662
rect 17325 10625 17359 10659
rect 18153 10625 18187 10659
rect 18420 10625 18454 10659
rect 20683 10625 20717 10659
rect 20821 10625 20855 10659
rect 20913 10628 20947 10662
rect 21097 10625 21131 10659
rect 22017 10625 22051 10659
rect 22201 10625 22235 10659
rect 23029 10625 23063 10659
rect 23857 10625 23891 10659
rect 4353 10557 4387 10591
rect 5457 10557 5491 10591
rect 7021 10557 7055 10591
rect 23121 10557 23155 10591
rect 23949 10557 23983 10591
rect 24041 10489 24075 10523
rect 4445 10421 4479 10455
rect 5457 10421 5491 10455
rect 9137 10421 9171 10455
rect 19533 10421 19567 10455
rect 21833 10421 21867 10455
rect 22109 10421 22143 10455
rect 23029 10421 23063 10455
rect 23397 10421 23431 10455
rect 24225 10421 24259 10455
rect 4353 10217 4387 10251
rect 5273 10217 5307 10251
rect 5457 10217 5491 10251
rect 8401 10217 8435 10251
rect 16773 10217 16807 10251
rect 20177 10217 20211 10251
rect 22661 10217 22695 10251
rect 23489 10217 23523 10251
rect 18705 10149 18739 10183
rect 22753 10081 22787 10115
rect 3249 10013 3283 10047
rect 4169 10013 4203 10047
rect 5181 10013 5215 10047
rect 5273 10013 5307 10047
rect 5917 10013 5951 10047
rect 6080 10007 6114 10041
rect 6193 10013 6227 10047
rect 6331 10013 6365 10047
rect 7021 10013 7055 10047
rect 15393 10013 15427 10047
rect 17325 10013 17359 10047
rect 20453 10013 20487 10047
rect 20545 10013 20579 10047
rect 20637 10013 20671 10047
rect 20821 10013 20855 10047
rect 22661 10013 22695 10047
rect 23489 10013 23523 10047
rect 23581 10013 23615 10047
rect 4997 9945 5031 9979
rect 6561 9945 6595 9979
rect 7266 9945 7300 9979
rect 15660 9945 15694 9979
rect 17592 9945 17626 9979
rect 11161 9877 11195 9911
rect 11989 9877 12023 9911
rect 13093 9877 13127 9911
rect 14197 9877 14231 9911
rect 14749 9877 14783 9911
rect 21741 9877 21775 9911
rect 23029 9877 23063 9911
rect 23857 9877 23891 9911
rect 3525 9673 3559 9707
rect 6837 9673 6871 9707
rect 6377 9605 6411 9639
rect 22753 9605 22787 9639
rect 3341 9537 3375 9571
rect 5457 9537 5491 9571
rect 6653 9537 6687 9571
rect 12817 9537 12851 9571
rect 20545 9537 20579 9571
rect 21097 9537 21131 9571
rect 21833 9537 21867 9571
rect 23029 9537 23063 9571
rect 23121 9537 23155 9571
rect 23213 9537 23247 9571
rect 23397 9537 23431 9571
rect 4537 9469 4571 9503
rect 4813 9469 4847 9503
rect 6469 9469 6503 9503
rect 12541 9469 12575 9503
rect 15577 9469 15611 9503
rect 15853 9469 15887 9503
rect 16681 9469 16715 9503
rect 16957 9469 16991 9503
rect 5273 9401 5307 9435
rect 7389 9401 7423 9435
rect 18061 9401 18095 9435
rect 22017 9401 22051 9435
rect 6377 9333 6411 9367
rect 7849 9333 7883 9367
rect 8585 9333 8619 9367
rect 9321 9333 9355 9367
rect 10977 9333 11011 9367
rect 13461 9333 13495 9367
rect 14565 9333 14599 9367
rect 18521 9333 18555 9367
rect 21281 9333 21315 9367
rect 17325 9061 17359 9095
rect 3249 8993 3283 9027
rect 5273 8993 5307 9027
rect 6561 8993 6595 9027
rect 10333 8993 10367 9027
rect 13001 8993 13035 9027
rect 21649 8993 21683 9027
rect 2697 8925 2731 8959
rect 2973 8925 3007 8959
rect 3065 8925 3099 8959
rect 4997 8925 5031 8959
rect 6285 8925 6319 8959
rect 7021 8925 7055 8959
rect 9413 8925 9447 8959
rect 12725 8925 12759 8959
rect 14105 8925 14139 8959
rect 15945 8925 15979 8959
rect 20545 8925 20579 8959
rect 20637 8925 20671 8959
rect 20729 8925 20763 8959
rect 20913 8925 20947 8959
rect 21373 8925 21407 8959
rect 23029 8925 23063 8959
rect 23121 8925 23155 8959
rect 23213 8925 23247 8959
rect 23397 8925 23431 8959
rect 7288 8857 7322 8891
rect 10578 8857 10612 8891
rect 14350 8857 14384 8891
rect 16212 8857 16246 8891
rect 20269 8857 20303 8891
rect 3801 8789 3835 8823
rect 8401 8789 8435 8823
rect 9597 8789 9631 8823
rect 11713 8789 11747 8823
rect 12265 8789 12299 8823
rect 15485 8789 15519 8823
rect 17877 8789 17911 8823
rect 18429 8789 18463 8823
rect 19349 8789 19383 8823
rect 22753 8789 22787 8823
rect 7021 8585 7055 8619
rect 8401 8585 8435 8619
rect 10149 8585 10183 8619
rect 13185 8585 13219 8619
rect 19533 8585 19567 8619
rect 20453 8585 20487 8619
rect 7481 8517 7515 8551
rect 15402 8517 15436 8551
rect 18420 8517 18454 8551
rect 5089 8449 5123 8483
rect 5549 8449 5583 8483
rect 6377 8449 6411 8483
rect 6540 8449 6574 8483
rect 6656 8449 6690 8483
rect 6791 8449 6825 8483
rect 7665 8449 7699 8483
rect 8309 8449 8343 8483
rect 9045 8449 9079 8483
rect 9505 8449 9539 8483
rect 10425 8449 10459 8483
rect 10530 8449 10564 8483
rect 10630 8449 10664 8483
rect 10793 8449 10827 8483
rect 11621 8449 11655 8483
rect 11897 8449 11931 8483
rect 12541 8449 12575 8483
rect 12725 8449 12759 8483
rect 12817 8449 12851 8483
rect 12909 8449 12943 8483
rect 13829 8449 13863 8483
rect 18153 8449 18187 8483
rect 19993 8449 20027 8483
rect 20269 8449 20303 8483
rect 21833 8449 21867 8483
rect 22109 8449 22143 8483
rect 23213 8449 23247 8483
rect 23397 8449 23431 8483
rect 23489 8449 23523 8483
rect 23581 8449 23615 8483
rect 24317 8449 24351 8483
rect 4813 8381 4847 8415
rect 11805 8381 11839 8415
rect 15669 8381 15703 8415
rect 16681 8381 16715 8415
rect 16957 8381 16991 8415
rect 20085 8381 20119 8415
rect 21281 8381 21315 8415
rect 12081 8313 12115 8347
rect 13645 8313 13679 8347
rect 14289 8313 14323 8347
rect 23857 8313 23891 8347
rect 5733 8245 5767 8279
rect 9689 8245 9723 8279
rect 11621 8245 11655 8279
rect 20085 8245 20119 8279
rect 4997 8041 5031 8075
rect 8401 8041 8435 8075
rect 9597 8041 9631 8075
rect 10149 8041 10183 8075
rect 10609 8041 10643 8075
rect 11069 8041 11103 8075
rect 11989 8041 12023 8075
rect 13553 8041 13587 8075
rect 16957 8041 16991 8075
rect 21557 8041 21591 8075
rect 25053 8041 25087 8075
rect 9597 7905 9631 7939
rect 10333 7905 10367 7939
rect 11253 7905 11287 7939
rect 12081 7905 12115 7939
rect 21557 7905 21591 7939
rect 5457 7837 5491 7871
rect 5641 7837 5675 7871
rect 5733 7837 5767 7871
rect 5825 7837 5859 7871
rect 7021 7837 7055 7871
rect 9413 7837 9447 7871
rect 10425 7837 10459 7871
rect 11345 7837 11379 7871
rect 12265 7837 12299 7871
rect 12909 7837 12943 7871
rect 13093 7837 13127 7871
rect 13185 7837 13219 7871
rect 13277 7837 13311 7871
rect 14565 7837 14599 7871
rect 15209 7837 15243 7871
rect 18061 7837 18095 7871
rect 19257 7837 19291 7871
rect 21465 7837 21499 7871
rect 22937 7837 22971 7871
rect 23029 7837 23063 7871
rect 23121 7837 23155 7871
rect 23305 7837 23339 7871
rect 24593 7837 24627 7871
rect 4261 7769 4295 7803
rect 6101 7769 6135 7803
rect 7266 7769 7300 7803
rect 9689 7769 9723 7803
rect 10149 7769 10183 7803
rect 11069 7769 11103 7803
rect 11989 7769 12023 7803
rect 15669 7769 15703 7803
rect 19524 7769 19558 7803
rect 22661 7769 22695 7803
rect 4353 7701 4387 7735
rect 9229 7701 9263 7735
rect 11529 7701 11563 7735
rect 12449 7701 12483 7735
rect 14381 7701 14415 7735
rect 15025 7701 15059 7735
rect 17877 7701 17911 7735
rect 18705 7701 18739 7735
rect 20637 7701 20671 7735
rect 21833 7701 21867 7735
rect 24409 7701 24443 7735
rect 4261 7497 4295 7531
rect 5181 7497 5215 7531
rect 6837 7497 6871 7531
rect 19533 7497 19567 7531
rect 21833 7497 21867 7531
rect 22845 7497 22879 7531
rect 4721 7429 4755 7463
rect 6377 7429 6411 7463
rect 7849 7429 7883 7463
rect 18420 7429 18454 7463
rect 4077 7361 4111 7395
rect 4997 7361 5031 7395
rect 5641 7361 5675 7395
rect 6653 7361 6687 7395
rect 9597 7361 9631 7395
rect 10057 7361 10091 7395
rect 10236 7361 10270 7395
rect 10336 7367 10370 7401
rect 10425 7361 10459 7395
rect 11621 7345 11655 7379
rect 12265 7361 12299 7395
rect 12428 7361 12462 7395
rect 12528 7364 12562 7398
rect 12633 7361 12667 7395
rect 13369 7361 13403 7395
rect 15945 7361 15979 7395
rect 16911 7361 16945 7395
rect 17049 7367 17083 7401
rect 17141 7361 17175 7395
rect 17325 7361 17359 7395
rect 18153 7361 18187 7395
rect 20821 7361 20855 7395
rect 21005 7361 21039 7395
rect 22017 7361 22051 7395
rect 22477 7361 22511 7395
rect 23305 7361 23339 7395
rect 4905 7293 4939 7327
rect 6469 7293 6503 7327
rect 22569 7293 22603 7327
rect 23397 7293 23431 7327
rect 5825 7225 5859 7259
rect 16129 7225 16163 7259
rect 20637 7225 20671 7259
rect 4997 7157 5031 7191
rect 6377 7157 6411 7191
rect 7389 7157 7423 7191
rect 10701 7157 10735 7191
rect 11805 7157 11839 7191
rect 12909 7157 12943 7191
rect 14657 7157 14691 7191
rect 16681 7157 16715 7191
rect 20177 7157 20211 7191
rect 21005 7157 21039 7191
rect 22661 7157 22695 7191
rect 23489 7157 23523 7191
rect 23673 7157 23707 7191
rect 5457 6953 5491 6987
rect 9229 6953 9263 6987
rect 10333 6953 10367 6987
rect 13369 6953 13403 6987
rect 14933 6953 14967 6987
rect 15485 6953 15519 6987
rect 17509 6953 17543 6987
rect 20361 6953 20395 6987
rect 24409 6953 24443 6987
rect 12725 6885 12759 6919
rect 14197 6885 14231 6919
rect 18705 6885 18739 6919
rect 22109 6885 22143 6919
rect 4629 6817 4663 6851
rect 6561 6817 6595 6851
rect 16129 6817 16163 6851
rect 24501 6817 24535 6851
rect 4353 6749 4387 6783
rect 5917 6749 5951 6783
rect 6101 6749 6135 6783
rect 6193 6749 6227 6783
rect 6285 6749 6319 6783
rect 7021 6749 7055 6783
rect 9229 6749 9263 6783
rect 9413 6749 9447 6783
rect 9505 6749 9539 6783
rect 10149 6749 10183 6783
rect 10977 6749 11011 6783
rect 11621 6749 11655 6783
rect 12265 6749 12299 6783
rect 12909 6749 12943 6783
rect 13553 6749 13587 6783
rect 14841 6749 14875 6783
rect 15025 6749 15059 6783
rect 15669 6749 15703 6783
rect 16396 6749 16430 6783
rect 18521 6749 18555 6783
rect 19257 6749 19291 6783
rect 21281 6749 21315 6783
rect 21373 6749 21407 6783
rect 21465 6749 21499 6783
rect 21649 6749 21683 6783
rect 23397 6749 23431 6783
rect 23489 6749 23523 6783
rect 23581 6749 23615 6783
rect 23765 6749 23799 6783
rect 24409 6749 24443 6783
rect 7266 6681 7300 6715
rect 18061 6681 18095 6715
rect 20453 6681 20487 6715
rect 8401 6613 8435 6647
rect 9689 6613 9723 6647
rect 10793 6613 10827 6647
rect 11437 6613 11471 6647
rect 12081 6613 12115 6647
rect 14657 6613 14691 6647
rect 19441 6613 19475 6647
rect 21005 6613 21039 6647
rect 23121 6613 23155 6647
rect 24777 6613 24811 6647
rect 4905 6409 4939 6443
rect 8861 6409 8895 6443
rect 10241 6409 10275 6443
rect 14289 6409 14323 6443
rect 18153 6409 18187 6443
rect 5365 6341 5399 6375
rect 13154 6341 13188 6375
rect 19288 6341 19322 6375
rect 21833 6341 21867 6375
rect 2697 6273 2731 6307
rect 3341 6273 3375 6307
rect 3985 6273 4019 6307
rect 4077 6273 4111 6307
rect 5549 6273 5583 6307
rect 5641 6273 5675 6307
rect 9321 6273 9355 6307
rect 10057 6273 10091 6307
rect 10333 6273 10367 6307
rect 10517 6273 10551 6307
rect 10793 6273 10827 6307
rect 11621 6273 11655 6307
rect 12449 6273 12483 6307
rect 15025 6273 15059 6307
rect 15117 6273 15151 6307
rect 16129 6273 16163 6307
rect 16865 6273 16899 6307
rect 17693 6273 17727 6307
rect 20637 6273 20671 6307
rect 21097 6273 21131 6307
rect 22109 6273 22143 6307
rect 22201 6273 22235 6307
rect 22293 6273 22327 6307
rect 22477 6273 22511 6307
rect 23213 6273 23247 6307
rect 12909 6205 12943 6239
rect 19533 6205 19567 6239
rect 22937 6205 22971 6239
rect 2881 6137 2915 6171
rect 4353 6137 4387 6171
rect 7205 6137 7239 6171
rect 12265 6137 12299 6171
rect 15393 6137 15427 6171
rect 17509 6137 17543 6171
rect 3525 6069 3559 6103
rect 3985 6069 4019 6103
rect 5457 6069 5491 6103
rect 5825 6069 5859 6103
rect 6653 6069 6687 6103
rect 7757 6069 7791 6103
rect 8309 6069 8343 6103
rect 9505 6069 9539 6103
rect 11805 6069 11839 6103
rect 15025 6069 15059 6103
rect 15945 6069 15979 6103
rect 17049 6069 17083 6103
rect 20453 6069 20487 6103
rect 21281 6069 21315 6103
rect 3985 5865 4019 5899
rect 5457 5865 5491 5899
rect 7757 5865 7791 5899
rect 9045 5865 9079 5899
rect 9505 5865 9539 5899
rect 14933 5865 14967 5899
rect 16957 5865 16991 5899
rect 20637 5865 20671 5899
rect 23857 5865 23891 5899
rect 4169 5797 4203 5831
rect 12725 5797 12759 5831
rect 5457 5729 5491 5763
rect 14933 5729 14967 5763
rect 19257 5729 19291 5763
rect 21925 5729 21959 5763
rect 22201 5729 22235 5763
rect 3801 5661 3835 5695
rect 3985 5661 4019 5695
rect 5273 5661 5307 5695
rect 5549 5661 5583 5695
rect 6193 5661 6227 5695
rect 6377 5661 6411 5695
rect 6469 5661 6503 5695
rect 6561 5661 6595 5695
rect 7941 5661 7975 5695
rect 9689 5661 9723 5695
rect 10149 5661 10183 5695
rect 10793 5661 10827 5695
rect 13185 5661 13219 5695
rect 14197 5661 14231 5695
rect 14841 5661 14875 5695
rect 15669 5661 15703 5695
rect 17877 5661 17911 5695
rect 18521 5661 18555 5695
rect 21281 5661 21315 5695
rect 11060 5593 11094 5627
rect 19524 5593 19558 5627
rect 5733 5525 5767 5559
rect 6837 5525 6871 5559
rect 10333 5525 10367 5559
rect 12173 5525 12207 5559
rect 13369 5525 13403 5559
rect 14381 5525 14415 5559
rect 15209 5525 15243 5559
rect 18061 5525 18095 5559
rect 18705 5525 18739 5559
rect 23213 5525 23247 5559
rect 4537 5321 4571 5355
rect 10517 5321 10551 5355
rect 15761 5321 15795 5355
rect 16681 5321 16715 5355
rect 19625 5321 19659 5355
rect 21005 5321 21039 5355
rect 9597 5253 9631 5287
rect 15301 5253 15335 5287
rect 17816 5253 17850 5287
rect 3525 5185 3559 5219
rect 5825 5185 5859 5219
rect 6377 5185 6411 5219
rect 6561 5185 6595 5219
rect 6653 5185 6687 5219
rect 6745 5185 6779 5219
rect 10057 5185 10091 5219
rect 10333 5185 10367 5219
rect 11713 5185 11747 5219
rect 12817 5185 12851 5219
rect 12909 5185 12943 5219
rect 13001 5185 13035 5219
rect 13185 5185 13219 5219
rect 13645 5185 13679 5219
rect 15577 5185 15611 5219
rect 18061 5185 18095 5219
rect 19809 5185 19843 5219
rect 20085 5185 20119 5219
rect 20545 5185 20579 5219
rect 20821 5185 20855 5219
rect 22017 5185 22051 5219
rect 23581 5185 23615 5219
rect 23673 5185 23707 5219
rect 23765 5185 23799 5219
rect 23949 5185 23983 5219
rect 3617 5117 3651 5151
rect 5549 5117 5583 5151
rect 10149 5117 10183 5151
rect 11805 5117 11839 5151
rect 13921 5117 13955 5151
rect 15485 5117 15519 5151
rect 19993 5117 20027 5151
rect 20637 5117 20671 5151
rect 24409 5117 24443 5151
rect 3893 5049 3927 5083
rect 19165 5049 19199 5083
rect 23305 5049 23339 5083
rect 3709 4981 3743 5015
rect 7021 4981 7055 5015
rect 8309 4981 8343 5015
rect 10333 4981 10367 5015
rect 11713 4981 11747 5015
rect 12081 4981 12115 5015
rect 12541 4981 12575 5015
rect 15301 4981 15335 5015
rect 20085 4981 20119 5015
rect 20821 4981 20855 5015
rect 21833 4981 21867 5015
rect 22477 4981 22511 5015
rect 3985 4777 4019 4811
rect 4905 4777 4939 4811
rect 5733 4777 5767 4811
rect 5917 4777 5951 4811
rect 8401 4777 8435 4811
rect 9689 4777 9723 4811
rect 12357 4777 12391 4811
rect 12725 4777 12759 4811
rect 14565 4777 14599 4811
rect 15485 4777 15519 4811
rect 15945 4777 15979 4811
rect 16405 4777 16439 4811
rect 16865 4777 16899 4811
rect 17325 4777 17359 4811
rect 17785 4777 17819 4811
rect 20269 4777 20303 4811
rect 20913 4777 20947 4811
rect 21281 4777 21315 4811
rect 21925 4777 21959 4811
rect 19809 4709 19843 4743
rect 22293 4709 22327 4743
rect 3893 4641 3927 4675
rect 5549 4641 5583 4675
rect 12449 4641 12483 4675
rect 14749 4641 14783 4675
rect 15669 4641 15703 4675
rect 17509 4641 17543 4675
rect 21189 4641 21223 4675
rect 21925 4641 21959 4675
rect 3801 4573 3835 4607
rect 4813 4573 4847 4607
rect 5457 4573 5491 4607
rect 5733 4573 5767 4607
rect 6561 4573 6595 4607
rect 7021 4573 7055 4607
rect 9505 4573 9539 4607
rect 10149 4573 10183 4607
rect 12357 4573 12391 4607
rect 13277 4573 13311 4607
rect 14565 4573 14599 4607
rect 14841 4573 14875 4607
rect 15761 4573 15795 4607
rect 16589 4573 16623 4607
rect 16697 4573 16731 4607
rect 17601 4573 17635 4607
rect 18521 4573 18555 4607
rect 19625 4573 19659 4607
rect 20453 4573 20487 4607
rect 21097 4573 21131 4607
rect 22109 4573 22143 4607
rect 23305 4573 23339 4607
rect 23394 4573 23428 4607
rect 23489 4573 23523 4607
rect 23673 4573 23707 4607
rect 24409 4573 24443 4607
rect 7288 4505 7322 4539
rect 10416 4505 10450 4539
rect 15485 4505 15519 4539
rect 16405 4505 16439 4539
rect 17325 4505 17359 4539
rect 21373 4505 21407 4539
rect 21833 4505 21867 4539
rect 4169 4437 4203 4471
rect 9045 4437 9079 4471
rect 11529 4437 11563 4471
rect 13461 4437 13495 4471
rect 15025 4437 15059 4471
rect 18337 4437 18371 4471
rect 23029 4437 23063 4471
rect 7941 4233 7975 4267
rect 11621 4233 11655 4267
rect 20453 4233 20487 4267
rect 10885 4165 10919 4199
rect 21833 4165 21867 4199
rect 2881 4097 2915 4131
rect 3341 4097 3375 4131
rect 5641 4097 5675 4131
rect 5825 4097 5859 4131
rect 6561 4097 6595 4131
rect 6828 4097 6862 4131
rect 8401 4097 8435 4131
rect 8657 4097 8691 4131
rect 12081 4097 12115 4131
rect 12265 4097 12299 4131
rect 12357 4097 12391 4131
rect 12449 4097 12483 4131
rect 13185 4097 13219 4131
rect 13441 4097 13475 4131
rect 15117 4097 15151 4131
rect 15853 4097 15887 4131
rect 17233 4097 17267 4131
rect 17969 4097 18003 4131
rect 18236 4097 18270 4131
rect 20637 4097 20671 4131
rect 21097 4097 21131 4131
rect 22109 4097 22143 4131
rect 3433 4029 3467 4063
rect 4997 4029 5031 4063
rect 10701 4029 10735 4063
rect 12725 4029 12759 4063
rect 21925 4029 21959 4063
rect 23397 4029 23431 4063
rect 16773 3961 16807 3995
rect 19993 3961 20027 3995
rect 22293 3961 22327 3995
rect 3525 3893 3559 3927
rect 3709 3893 3743 3927
rect 4767 3893 4801 3927
rect 5733 3893 5767 3927
rect 9781 3893 9815 3927
rect 14565 3893 14599 3927
rect 15301 3893 15335 3927
rect 16037 3893 16071 3927
rect 17417 3893 17451 3927
rect 19349 3893 19383 3927
rect 21281 3893 21315 3927
rect 21925 3893 21959 3927
rect 22753 3893 22787 3927
rect 24041 3893 24075 3927
rect 24685 3893 24719 3927
rect 5917 3689 5951 3723
rect 21741 3689 21775 3723
rect 4261 3621 4295 3655
rect 14473 3621 14507 3655
rect 17233 3621 17267 3655
rect 20085 3621 20119 3655
rect 21925 3621 21959 3655
rect 52101 3621 52135 3655
rect 10333 3553 10367 3587
rect 13277 3553 13311 3587
rect 24409 3553 24443 3587
rect 5273 3485 5307 3519
rect 5436 3482 5470 3516
rect 5536 3479 5570 3513
rect 5687 3485 5721 3519
rect 6377 3485 6411 3519
rect 6561 3485 6595 3519
rect 6653 3485 6687 3519
rect 6745 3485 6779 3519
rect 7757 3485 7791 3519
rect 8217 3485 8251 3519
rect 8953 3485 8987 3519
rect 9505 3485 9539 3519
rect 13001 3485 13035 3519
rect 14289 3485 14323 3519
rect 15301 3485 15335 3519
rect 15749 3485 15783 3519
rect 15945 3485 15979 3519
rect 16037 3485 16071 3519
rect 16175 3485 16209 3519
rect 18613 3485 18647 3519
rect 19533 3485 19567 3519
rect 20269 3485 20303 3519
rect 21281 3485 21315 3519
rect 21373 3485 21407 3519
rect 21741 3485 21775 3519
rect 22845 3485 22879 3519
rect 23673 3485 23707 3519
rect 26157 3485 26191 3519
rect 27261 3485 27295 3519
rect 27721 3485 27755 3519
rect 28365 3485 28399 3519
rect 29561 3485 29595 3519
rect 30297 3485 30331 3519
rect 31401 3485 31435 3519
rect 32229 3485 32263 3519
rect 33057 3485 33091 3519
rect 39957 3485 39991 3519
rect 40601 3485 40635 3519
rect 41245 3485 41279 3519
rect 41889 3485 41923 3519
rect 42717 3485 42751 3519
rect 43821 3485 43855 3519
rect 45201 3485 45235 3519
rect 45845 3485 45879 3519
rect 46489 3485 46523 3519
rect 47685 3485 47719 3519
rect 48329 3485 48363 3519
rect 50169 3485 50203 3519
rect 50813 3485 50847 3519
rect 51457 3485 51491 3519
rect 52929 3485 52963 3519
rect 53573 3485 53607 3519
rect 55413 3485 55447 3519
rect 56057 3485 56091 3519
rect 56701 3485 56735 3519
rect 57345 3485 57379 3519
rect 57989 3485 58023 3519
rect 10578 3417 10612 3451
rect 16405 3417 16439 3451
rect 18346 3417 18380 3451
rect 4813 3349 4847 3383
rect 7021 3349 7055 3383
rect 7573 3349 7607 3383
rect 8401 3349 8435 3383
rect 9689 3349 9723 3383
rect 11713 3349 11747 3383
rect 15117 3349 15151 3383
rect 19349 3349 19383 3383
rect 25053 3349 25087 3383
rect 3065 3145 3099 3179
rect 4721 3145 4755 3179
rect 10701 3145 10735 3179
rect 17969 3145 18003 3179
rect 14197 3077 14231 3111
rect 15770 3077 15804 3111
rect 18696 3077 18730 3111
rect 4077 3009 4111 3043
rect 4240 3009 4274 3043
rect 4340 3009 4374 3043
rect 4445 3009 4479 3043
rect 5181 3009 5215 3043
rect 5344 3009 5378 3043
rect 5457 3009 5491 3043
rect 5595 3009 5629 3043
rect 6745 3009 6779 3043
rect 7205 3009 7239 3043
rect 7461 3009 7495 3043
rect 9321 3009 9355 3043
rect 9577 3009 9611 3043
rect 11989 3009 12023 3043
rect 12725 3009 12759 3043
rect 12909 3009 12943 3043
rect 13541 3009 13575 3043
rect 13737 3009 13771 3043
rect 13829 3009 13863 3043
rect 13921 3009 13955 3043
rect 16681 3009 16715 3043
rect 16865 3009 16899 3043
rect 16957 3009 16991 3043
rect 17049 3009 17083 3043
rect 17785 3009 17819 3043
rect 20545 3009 20579 3043
rect 16037 2941 16071 2975
rect 18429 2941 18463 2975
rect 21281 2941 21315 2975
rect 25145 2941 25179 2975
rect 38577 2941 38611 2975
rect 40509 2941 40543 2975
rect 44373 2941 44407 2975
rect 48237 2941 48271 2975
rect 50169 2941 50203 2975
rect 55965 2941 55999 2975
rect 5825 2873 5859 2907
rect 20361 2873 20395 2907
rect 39221 2873 39255 2907
rect 41153 2873 41187 2907
rect 43085 2873 43119 2907
rect 45017 2873 45051 2907
rect 46305 2873 46339 2907
rect 48881 2873 48915 2907
rect 50813 2873 50847 2907
rect 53389 2873 53423 2907
rect 54677 2873 54711 2907
rect 58541 2873 58575 2907
rect 3525 2805 3559 2839
rect 6561 2805 6595 2839
rect 8585 2805 8619 2839
rect 12173 2805 12207 2839
rect 12817 2805 12851 2839
rect 14657 2805 14691 2839
rect 17325 2805 17359 2839
rect 19809 2805 19843 2839
rect 21833 2805 21867 2839
rect 22569 2805 22603 2839
rect 23213 2805 23247 2839
rect 23857 2805 23891 2839
rect 24501 2805 24535 2839
rect 25789 2805 25823 2839
rect 26249 2805 26283 2839
rect 26985 2805 27019 2839
rect 27721 2805 27755 2839
rect 28365 2805 28399 2839
rect 29009 2805 29043 2839
rect 29653 2805 29687 2839
rect 30297 2805 30331 2839
rect 30941 2805 30975 2839
rect 31585 2805 31619 2839
rect 32505 2805 32539 2839
rect 33149 2805 33183 2839
rect 33793 2805 33827 2839
rect 34253 2805 34287 2839
rect 34897 2805 34931 2839
rect 35541 2805 35575 2839
rect 36369 2805 36403 2839
rect 37289 2805 37323 2839
rect 37933 2805 37967 2839
rect 39865 2805 39899 2839
rect 42441 2805 42475 2839
rect 43729 2805 43763 2839
rect 45661 2805 45695 2839
rect 47593 2805 47627 2839
rect 49525 2805 49559 2839
rect 51457 2805 51491 2839
rect 52745 2805 52779 2839
rect 54033 2805 54067 2839
rect 55321 2805 55355 2839
rect 56609 2805 56643 2839
rect 57897 2805 57931 2839
rect 4537 2601 4571 2635
rect 6377 2601 6411 2635
rect 9321 2601 9355 2635
rect 14565 2601 14599 2635
rect 17049 2601 17083 2635
rect 4077 2533 4111 2567
rect 8401 2533 8435 2567
rect 11989 2533 12023 2567
rect 12725 2533 12759 2567
rect 19533 2533 19567 2567
rect 21925 2533 21959 2567
rect 23213 2533 23247 2567
rect 30941 2533 30975 2567
rect 32873 2533 32907 2567
rect 41153 2533 41187 2567
rect 45017 2533 45051 2567
rect 48881 2533 48915 2567
rect 52745 2533 52779 2567
rect 56609 2533 56643 2567
rect 58541 2533 58575 2567
rect 7021 2465 7055 2499
rect 18429 2465 18463 2499
rect 25697 2465 25731 2499
rect 37933 2465 37967 2499
rect 39865 2465 39899 2499
rect 42441 2465 42475 2499
rect 45661 2465 45695 2499
rect 47593 2465 47627 2499
rect 50169 2465 50203 2499
rect 53389 2465 53423 2499
rect 55321 2465 55355 2499
rect 59185 2465 59219 2499
rect 3893 2397 3927 2431
rect 4721 2397 4755 2431
rect 5181 2397 5215 2431
rect 5365 2397 5399 2431
rect 5457 2397 5491 2431
rect 5595 2397 5629 2431
rect 6561 2397 6595 2431
rect 9505 2397 9539 2431
rect 10241 2397 10275 2431
rect 10977 2397 11011 2431
rect 11805 2397 11839 2431
rect 12541 2397 12575 2431
rect 13277 2397 13311 2431
rect 14381 2397 14415 2431
rect 15393 2397 15427 2431
rect 16129 2397 16163 2431
rect 18162 2397 18196 2431
rect 19717 2397 19751 2431
rect 20453 2397 20487 2431
rect 21189 2397 21223 2431
rect 22109 2397 22143 2431
rect 23857 2397 23891 2431
rect 26157 2397 26191 2431
rect 26985 2397 27019 2431
rect 28365 2397 28399 2431
rect 29009 2397 29043 2431
rect 30297 2397 30331 2431
rect 31585 2397 31619 2431
rect 33517 2397 33551 2431
rect 34161 2397 34195 2431
rect 34989 2397 35023 2431
rect 35633 2397 35667 2431
rect 36093 2397 36127 2431
rect 37289 2397 37323 2431
rect 38577 2397 38611 2431
rect 40509 2397 40543 2431
rect 43085 2397 43119 2431
rect 43729 2397 43763 2431
rect 46305 2397 46339 2431
rect 48237 2397 48271 2431
rect 50813 2397 50847 2431
rect 51457 2397 51491 2431
rect 54033 2397 54067 2431
rect 55965 2397 55999 2431
rect 57897 2397 57931 2431
rect 2697 2329 2731 2363
rect 5825 2329 5859 2363
rect 7266 2329 7300 2363
rect 3249 2261 3283 2295
rect 10057 2261 10091 2295
rect 10793 2261 10827 2295
rect 13461 2261 13495 2295
rect 15209 2261 15243 2295
rect 15945 2261 15979 2295
rect 20269 2261 20303 2295
rect 21005 2261 21039 2295
rect 25053 2261 25087 2295
rect 26341 2261 26375 2295
rect 27169 2261 27203 2295
<< metal1 >>
rect 1104 57690 68816 57712
rect 1104 57638 19574 57690
rect 19626 57638 19638 57690
rect 19690 57638 19702 57690
rect 19754 57638 19766 57690
rect 19818 57638 19830 57690
rect 19882 57638 50294 57690
rect 50346 57638 50358 57690
rect 50410 57638 50422 57690
rect 50474 57638 50486 57690
rect 50538 57638 50550 57690
rect 50602 57638 68816 57690
rect 1104 57616 68816 57638
rect 3237 57443 3295 57449
rect 3237 57409 3249 57443
rect 3283 57440 3295 57443
rect 3510 57440 3516 57452
rect 3283 57412 3516 57440
rect 3283 57409 3295 57412
rect 3237 57403 3295 57409
rect 3510 57400 3516 57412
rect 3568 57400 3574 57452
rect 4154 57440 4160 57452
rect 4115 57412 4160 57440
rect 4154 57400 4160 57412
rect 4212 57400 4218 57452
rect 5166 57440 5172 57452
rect 5127 57412 5172 57440
rect 5166 57400 5172 57412
rect 5224 57400 5230 57452
rect 5629 57443 5687 57449
rect 5629 57409 5641 57443
rect 5675 57440 5687 57443
rect 5718 57440 5724 57452
rect 5675 57412 5724 57440
rect 5675 57409 5687 57412
rect 5629 57403 5687 57409
rect 5718 57400 5724 57412
rect 5776 57400 5782 57452
rect 6822 57440 6828 57452
rect 6783 57412 6828 57440
rect 6822 57400 6828 57412
rect 6880 57400 6886 57452
rect 7374 57400 7380 57452
rect 7432 57440 7438 57452
rect 7469 57443 7527 57449
rect 7469 57440 7481 57443
rect 7432 57412 7481 57440
rect 7432 57400 7438 57412
rect 7469 57409 7481 57412
rect 7515 57409 7527 57443
rect 7469 57403 7527 57409
rect 8389 57443 8447 57449
rect 8389 57409 8401 57443
rect 8435 57440 8447 57443
rect 8478 57440 8484 57452
rect 8435 57412 8484 57440
rect 8435 57409 8447 57412
rect 8389 57403 8447 57409
rect 8478 57400 8484 57412
rect 8536 57400 8542 57452
rect 9030 57400 9036 57452
rect 9088 57440 9094 57452
rect 9125 57443 9183 57449
rect 9125 57440 9137 57443
rect 9088 57412 9137 57440
rect 9088 57400 9094 57412
rect 9125 57409 9137 57412
rect 9171 57409 9183 57443
rect 10134 57440 10140 57452
rect 10095 57412 10140 57440
rect 9125 57403 9183 57409
rect 10134 57400 10140 57412
rect 10192 57400 10198 57452
rect 10686 57400 10692 57452
rect 10744 57440 10750 57452
rect 10781 57443 10839 57449
rect 10781 57440 10793 57443
rect 10744 57412 10793 57440
rect 10744 57400 10750 57412
rect 10781 57409 10793 57412
rect 10827 57409 10839 57443
rect 11790 57440 11796 57452
rect 11751 57412 11796 57440
rect 10781 57403 10839 57409
rect 11790 57400 11796 57412
rect 11848 57400 11854 57452
rect 12434 57440 12440 57452
rect 12395 57412 12440 57440
rect 12434 57400 12440 57412
rect 12492 57400 12498 57452
rect 13357 57443 13415 57449
rect 13357 57409 13369 57443
rect 13403 57440 13415 57443
rect 13446 57440 13452 57452
rect 13403 57412 13452 57440
rect 13403 57409 13415 57412
rect 13357 57403 13415 57409
rect 13446 57400 13452 57412
rect 13504 57400 13510 57452
rect 13998 57400 14004 57452
rect 14056 57440 14062 57452
rect 14093 57443 14151 57449
rect 14093 57440 14105 57443
rect 14056 57412 14105 57440
rect 14056 57400 14062 57412
rect 14093 57409 14105 57412
rect 14139 57409 14151 57443
rect 15102 57440 15108 57452
rect 15063 57412 15108 57440
rect 14093 57403 14151 57409
rect 15102 57400 15108 57412
rect 15160 57400 15166 57452
rect 15654 57400 15660 57452
rect 15712 57440 15718 57452
rect 15749 57443 15807 57449
rect 15749 57440 15761 57443
rect 15712 57412 15761 57440
rect 15712 57400 15718 57412
rect 15749 57409 15761 57412
rect 15795 57409 15807 57443
rect 16758 57440 16764 57452
rect 16719 57412 16764 57440
rect 15749 57403 15807 57409
rect 16758 57400 16764 57412
rect 16816 57400 16822 57452
rect 17310 57400 17316 57452
rect 17368 57440 17374 57452
rect 17405 57443 17463 57449
rect 17405 57440 17417 57443
rect 17368 57412 17417 57440
rect 17368 57400 17374 57412
rect 17405 57409 17417 57412
rect 17451 57409 17463 57443
rect 17405 57403 17463 57409
rect 18414 57400 18420 57452
rect 18472 57440 18478 57452
rect 18509 57443 18567 57449
rect 18509 57440 18521 57443
rect 18472 57412 18521 57440
rect 18472 57400 18478 57412
rect 18509 57409 18521 57412
rect 18555 57409 18567 57443
rect 18509 57403 18567 57409
rect 18966 57400 18972 57452
rect 19024 57440 19030 57452
rect 19245 57443 19303 57449
rect 19245 57440 19257 57443
rect 19024 57412 19257 57440
rect 19024 57400 19030 57412
rect 19245 57409 19257 57412
rect 19291 57409 19303 57443
rect 20070 57440 20076 57452
rect 20031 57412 20076 57440
rect 19245 57403 19303 57409
rect 20070 57400 20076 57412
rect 20128 57400 20134 57452
rect 20714 57440 20720 57452
rect 20675 57412 20720 57440
rect 20714 57400 20720 57412
rect 20772 57400 20778 57452
rect 22278 57400 22284 57452
rect 22336 57440 22342 57452
rect 22373 57443 22431 57449
rect 22373 57440 22385 57443
rect 22336 57412 22385 57440
rect 22336 57400 22342 57412
rect 22373 57409 22385 57412
rect 22419 57409 22431 57443
rect 23474 57440 23480 57452
rect 23435 57412 23480 57440
rect 22373 57403 22431 57409
rect 23474 57400 23480 57412
rect 23532 57400 23538 57452
rect 23934 57400 23940 57452
rect 23992 57440 23998 57452
rect 24397 57443 24455 57449
rect 24397 57440 24409 57443
rect 23992 57412 24409 57440
rect 23992 57400 23998 57412
rect 24397 57409 24409 57412
rect 24443 57409 24455 57443
rect 25038 57440 25044 57452
rect 24999 57412 25044 57440
rect 24397 57403 24455 57409
rect 25038 57400 25044 57412
rect 25096 57400 25102 57452
rect 25590 57400 25596 57452
rect 25648 57440 25654 57452
rect 25685 57443 25743 57449
rect 25685 57440 25697 57443
rect 25648 57412 25697 57440
rect 25648 57400 25654 57412
rect 25685 57409 25697 57412
rect 25731 57409 25743 57443
rect 25685 57403 25743 57409
rect 27246 57400 27252 57452
rect 27304 57440 27310 57452
rect 27341 57443 27399 57449
rect 27341 57440 27353 57443
rect 27304 57412 27353 57440
rect 27304 57400 27310 57412
rect 27341 57409 27353 57412
rect 27387 57409 27399 57443
rect 28350 57440 28356 57452
rect 28311 57412 28356 57440
rect 27341 57403 27399 57409
rect 28350 57400 28356 57412
rect 28408 57400 28414 57452
rect 28813 57443 28871 57449
rect 28813 57409 28825 57443
rect 28859 57440 28871 57443
rect 28902 57440 28908 57452
rect 28859 57412 28908 57440
rect 28859 57409 28871 57412
rect 28813 57403 28871 57409
rect 28902 57400 28908 57412
rect 28960 57400 28966 57452
rect 30006 57440 30012 57452
rect 29967 57412 30012 57440
rect 30006 57400 30012 57412
rect 30064 57400 30070 57452
rect 30558 57400 30564 57452
rect 30616 57440 30622 57452
rect 30653 57443 30711 57449
rect 30653 57440 30665 57443
rect 30616 57412 30665 57440
rect 30616 57400 30622 57412
rect 30653 57409 30665 57412
rect 30699 57409 30711 57443
rect 30653 57403 30711 57409
rect 31573 57443 31631 57449
rect 31573 57409 31585 57443
rect 31619 57440 31631 57443
rect 31662 57440 31668 57452
rect 31619 57412 31668 57440
rect 31619 57409 31631 57412
rect 31573 57403 31631 57409
rect 31662 57400 31668 57412
rect 31720 57400 31726 57452
rect 32214 57400 32220 57452
rect 32272 57440 32278 57452
rect 32309 57443 32367 57449
rect 32309 57440 32321 57443
rect 32272 57412 32321 57440
rect 32272 57400 32278 57412
rect 32309 57409 32321 57412
rect 32355 57409 32367 57443
rect 33318 57440 33324 57452
rect 33279 57412 33324 57440
rect 32309 57403 32367 57409
rect 33318 57400 33324 57412
rect 33376 57400 33382 57452
rect 33870 57400 33876 57452
rect 33928 57440 33934 57452
rect 33965 57443 34023 57449
rect 33965 57440 33977 57443
rect 33928 57412 33977 57440
rect 33928 57400 33934 57412
rect 33965 57409 33977 57412
rect 34011 57409 34023 57443
rect 34974 57440 34980 57452
rect 34935 57412 34980 57440
rect 33965 57403 34023 57409
rect 34974 57400 34980 57412
rect 35032 57400 35038 57452
rect 35526 57400 35532 57452
rect 35584 57440 35590 57452
rect 35621 57443 35679 57449
rect 35621 57440 35633 57443
rect 35584 57412 35633 57440
rect 35584 57400 35590 57412
rect 35621 57409 35633 57412
rect 35667 57409 35679 57443
rect 35621 57403 35679 57409
rect 36630 57400 36636 57452
rect 36688 57440 36694 57452
rect 37277 57443 37335 57449
rect 37277 57440 37289 57443
rect 36688 57412 37289 57440
rect 36688 57400 36694 57412
rect 37277 57409 37289 57412
rect 37323 57409 37335 57443
rect 37277 57403 37335 57409
rect 38286 57400 38292 57452
rect 38344 57440 38350 57452
rect 38565 57443 38623 57449
rect 38565 57440 38577 57443
rect 38344 57412 38577 57440
rect 38344 57400 38350 57412
rect 38565 57409 38577 57412
rect 38611 57409 38623 57443
rect 40034 57440 40040 57452
rect 39995 57412 40040 57440
rect 38565 57403 38623 57409
rect 40034 57400 40040 57412
rect 40092 57400 40098 57452
rect 40494 57400 40500 57452
rect 40552 57440 40558 57452
rect 40681 57443 40739 57449
rect 40681 57440 40693 57443
rect 40552 57412 40693 57440
rect 40552 57400 40558 57412
rect 40681 57409 40693 57412
rect 40727 57409 40739 57443
rect 40681 57403 40739 57409
rect 41598 57400 41604 57452
rect 41656 57440 41662 57452
rect 41693 57443 41751 57449
rect 41693 57440 41705 57443
rect 41656 57412 41705 57440
rect 41656 57400 41662 57412
rect 41693 57409 41705 57412
rect 41739 57409 41751 57443
rect 41693 57403 41751 57409
rect 42150 57400 42156 57452
rect 42208 57440 42214 57452
rect 42429 57443 42487 57449
rect 42429 57440 42441 57443
rect 42208 57412 42441 57440
rect 42208 57400 42214 57412
rect 42429 57409 42441 57412
rect 42475 57409 42487 57443
rect 42429 57403 42487 57409
rect 43254 57400 43260 57452
rect 43312 57440 43318 57452
rect 43349 57443 43407 57449
rect 43349 57440 43361 57443
rect 43312 57412 43361 57440
rect 43312 57400 43318 57412
rect 43349 57409 43361 57412
rect 43395 57409 43407 57443
rect 43349 57403 43407 57409
rect 43806 57400 43812 57452
rect 43864 57440 43870 57452
rect 43993 57443 44051 57449
rect 43993 57440 44005 57443
rect 43864 57412 44005 57440
rect 43864 57400 43870 57412
rect 43993 57409 44005 57412
rect 44039 57409 44051 57443
rect 43993 57403 44051 57409
rect 44910 57400 44916 57452
rect 44968 57440 44974 57452
rect 45005 57443 45063 57449
rect 45005 57440 45017 57443
rect 44968 57412 45017 57440
rect 44968 57400 44974 57412
rect 45005 57409 45017 57412
rect 45051 57409 45063 57443
rect 45005 57403 45063 57409
rect 46566 57400 46572 57452
rect 46624 57440 46630 57452
rect 46661 57443 46719 57449
rect 46661 57440 46673 57443
rect 46624 57412 46673 57440
rect 46624 57400 46630 57412
rect 46661 57409 46673 57412
rect 46707 57409 46719 57443
rect 46661 57403 46719 57409
rect 47118 57400 47124 57452
rect 47176 57440 47182 57452
rect 47581 57443 47639 57449
rect 47581 57440 47593 57443
rect 47176 57412 47593 57440
rect 47176 57400 47182 57412
rect 47581 57409 47593 57412
rect 47627 57409 47639 57443
rect 48314 57440 48320 57452
rect 48275 57412 48320 57440
rect 47581 57403 47639 57409
rect 48314 57400 48320 57412
rect 48372 57400 48378 57452
rect 48774 57400 48780 57452
rect 48832 57440 48838 57452
rect 48961 57443 49019 57449
rect 48961 57440 48973 57443
rect 48832 57412 48973 57440
rect 48832 57400 48838 57412
rect 48961 57409 48973 57412
rect 49007 57409 49019 57443
rect 48961 57403 49019 57409
rect 49878 57400 49884 57452
rect 49936 57440 49942 57452
rect 50157 57443 50215 57449
rect 50157 57440 50169 57443
rect 49936 57412 50169 57440
rect 49936 57400 49942 57412
rect 50157 57409 50169 57412
rect 50203 57409 50215 57443
rect 50157 57403 50215 57409
rect 50614 57400 50620 57452
rect 50672 57440 50678 57452
rect 50801 57443 50859 57449
rect 50801 57440 50813 57443
rect 50672 57412 50813 57440
rect 50672 57400 50678 57412
rect 50801 57409 50813 57412
rect 50847 57409 50859 57443
rect 50801 57403 50859 57409
rect 51534 57400 51540 57452
rect 51592 57440 51598 57452
rect 51629 57443 51687 57449
rect 51629 57440 51641 57443
rect 51592 57412 51641 57440
rect 51592 57400 51598 57412
rect 51629 57409 51641 57412
rect 51675 57409 51687 57443
rect 51629 57403 51687 57409
rect 52454 57400 52460 57452
rect 52512 57440 52518 57452
rect 52733 57443 52791 57449
rect 52733 57440 52745 57443
rect 52512 57412 52745 57440
rect 52512 57400 52518 57412
rect 52733 57409 52745 57412
rect 52779 57409 52791 57443
rect 52733 57403 52791 57409
rect 53190 57400 53196 57452
rect 53248 57440 53254 57452
rect 53377 57443 53435 57449
rect 53377 57440 53389 57443
rect 53248 57412 53389 57440
rect 53248 57400 53254 57412
rect 53377 57409 53389 57412
rect 53423 57409 53435 57443
rect 53377 57403 53435 57409
rect 53834 57400 53840 57452
rect 53892 57440 53898 57452
rect 54021 57443 54079 57449
rect 54021 57440 54033 57443
rect 53892 57412 54033 57440
rect 53892 57400 53898 57412
rect 54021 57409 54033 57412
rect 54067 57409 54079 57443
rect 54021 57403 54079 57409
rect 54846 57400 54852 57452
rect 54904 57440 54910 57452
rect 55309 57443 55367 57449
rect 55309 57440 55321 57443
rect 54904 57412 55321 57440
rect 54904 57400 54910 57412
rect 55309 57409 55321 57412
rect 55355 57409 55367 57443
rect 55309 57403 55367 57409
rect 55398 57400 55404 57452
rect 55456 57440 55462 57452
rect 55953 57443 56011 57449
rect 55953 57440 55965 57443
rect 55456 57412 55965 57440
rect 55456 57400 55462 57412
rect 55953 57409 55965 57412
rect 55999 57409 56011 57443
rect 56594 57440 56600 57452
rect 56555 57412 56600 57440
rect 55953 57403 56011 57409
rect 56594 57400 56600 57412
rect 56652 57400 56658 57452
rect 57054 57400 57060 57452
rect 57112 57440 57118 57452
rect 57885 57443 57943 57449
rect 57885 57440 57897 57443
rect 57112 57412 57897 57440
rect 57112 57400 57118 57412
rect 57885 57409 57897 57412
rect 57931 57409 57943 57443
rect 57885 57403 57943 57409
rect 58158 57400 58164 57452
rect 58216 57440 58222 57452
rect 58529 57443 58587 57449
rect 58529 57440 58541 57443
rect 58216 57412 58541 57440
rect 58216 57400 58222 57412
rect 58529 57409 58541 57412
rect 58575 57409 58587 57443
rect 58529 57403 58587 57409
rect 58710 57400 58716 57452
rect 58768 57440 58774 57452
rect 59173 57443 59231 57449
rect 59173 57440 59185 57443
rect 58768 57412 59185 57440
rect 58768 57400 58774 57412
rect 59173 57409 59185 57412
rect 59219 57409 59231 57443
rect 59173 57403 59231 57409
rect 59814 57400 59820 57452
rect 59872 57440 59878 57452
rect 60461 57443 60519 57449
rect 60461 57440 60473 57443
rect 59872 57412 60473 57440
rect 59872 57400 59878 57412
rect 60461 57409 60473 57412
rect 60507 57409 60519 57443
rect 60461 57403 60519 57409
rect 60734 57400 60740 57452
rect 60792 57440 60798 57452
rect 61105 57443 61163 57449
rect 61105 57440 61117 57443
rect 60792 57412 61117 57440
rect 60792 57400 60798 57412
rect 61105 57409 61117 57412
rect 61151 57409 61163 57443
rect 61105 57403 61163 57409
rect 61470 57400 61476 57452
rect 61528 57440 61534 57452
rect 61749 57443 61807 57449
rect 61749 57440 61761 57443
rect 61528 57412 61761 57440
rect 61528 57400 61534 57412
rect 61749 57409 61761 57412
rect 61795 57409 61807 57443
rect 61749 57403 61807 57409
rect 63126 57400 63132 57452
rect 63184 57440 63190 57452
rect 63221 57443 63279 57449
rect 63221 57440 63233 57443
rect 63184 57412 63233 57440
rect 63184 57400 63190 57412
rect 63221 57409 63233 57412
rect 63267 57409 63279 57443
rect 63221 57403 63279 57409
rect 63678 57400 63684 57452
rect 63736 57440 63742 57452
rect 63865 57443 63923 57449
rect 63865 57440 63877 57443
rect 63736 57412 63877 57440
rect 63736 57400 63742 57412
rect 63865 57409 63877 57412
rect 63911 57409 63923 57443
rect 63865 57403 63923 57409
rect 65334 57400 65340 57452
rect 65392 57440 65398 57452
rect 65613 57443 65671 57449
rect 65613 57440 65625 57443
rect 65392 57412 65625 57440
rect 65392 57400 65398 57412
rect 65613 57409 65625 57412
rect 65659 57409 65671 57443
rect 65613 57403 65671 57409
rect 66990 57400 66996 57452
rect 67048 57440 67054 57452
rect 67085 57443 67143 57449
rect 67085 57440 67097 57443
rect 67048 57412 67097 57440
rect 67048 57400 67054 57412
rect 67085 57409 67097 57412
rect 67131 57409 67143 57443
rect 67085 57403 67143 57409
rect 45462 57332 45468 57384
rect 45520 57372 45526 57384
rect 45649 57375 45707 57381
rect 45649 57372 45661 57375
rect 45520 57344 45661 57372
rect 45520 57332 45526 57344
rect 45649 57341 45661 57344
rect 45695 57341 45707 57375
rect 45649 57335 45707 57341
rect 64782 57332 64788 57384
rect 64840 57372 64846 57384
rect 64877 57375 64935 57381
rect 64877 57372 64889 57375
rect 64840 57344 64889 57372
rect 64840 57332 64846 57344
rect 64877 57341 64889 57344
rect 64923 57341 64935 57375
rect 64877 57335 64935 57341
rect 37274 57264 37280 57316
rect 37332 57304 37338 57316
rect 37921 57307 37979 57313
rect 37921 57304 37933 57307
rect 37332 57276 37933 57304
rect 37332 57264 37338 57276
rect 37921 57273 37933 57276
rect 37967 57273 37979 57307
rect 37921 57267 37979 57273
rect 1104 57146 68816 57168
rect 1104 57094 4214 57146
rect 4266 57094 4278 57146
rect 4330 57094 4342 57146
rect 4394 57094 4406 57146
rect 4458 57094 4470 57146
rect 4522 57094 34934 57146
rect 34986 57094 34998 57146
rect 35050 57094 35062 57146
rect 35114 57094 35126 57146
rect 35178 57094 35190 57146
rect 35242 57094 65654 57146
rect 65706 57094 65718 57146
rect 65770 57094 65782 57146
rect 65834 57094 65846 57146
rect 65898 57094 65910 57146
rect 65962 57094 68816 57146
rect 1104 57072 68816 57094
rect 21726 56992 21732 57044
rect 21784 57032 21790 57044
rect 21821 57035 21879 57041
rect 21821 57032 21833 57035
rect 21784 57004 21833 57032
rect 21784 56992 21790 57004
rect 21821 57001 21833 57004
rect 21867 57001 21879 57035
rect 21821 56995 21879 57001
rect 26694 56992 26700 57044
rect 26752 57032 26758 57044
rect 26789 57035 26847 57041
rect 26789 57032 26801 57035
rect 26752 57004 26801 57032
rect 26752 56992 26758 57004
rect 26789 57001 26801 57004
rect 26835 57001 26847 57035
rect 26789 56995 26847 57001
rect 38838 56992 38844 57044
rect 38896 57032 38902 57044
rect 38933 57035 38991 57041
rect 38933 57032 38945 57035
rect 38896 57004 38945 57032
rect 38896 56992 38902 57004
rect 38933 57001 38945 57004
rect 38979 57001 38991 57035
rect 62114 57032 62120 57044
rect 62075 57004 62120 57032
rect 38933 56995 38991 57001
rect 62114 56992 62120 57004
rect 62172 56992 62178 57044
rect 1104 56602 68816 56624
rect 1104 56550 19574 56602
rect 19626 56550 19638 56602
rect 19690 56550 19702 56602
rect 19754 56550 19766 56602
rect 19818 56550 19830 56602
rect 19882 56550 50294 56602
rect 50346 56550 50358 56602
rect 50410 56550 50422 56602
rect 50474 56550 50486 56602
rect 50538 56550 50550 56602
rect 50602 56550 68816 56602
rect 1104 56528 68816 56550
rect 1104 56058 68816 56080
rect 1104 56006 4214 56058
rect 4266 56006 4278 56058
rect 4330 56006 4342 56058
rect 4394 56006 4406 56058
rect 4458 56006 4470 56058
rect 4522 56006 34934 56058
rect 34986 56006 34998 56058
rect 35050 56006 35062 56058
rect 35114 56006 35126 56058
rect 35178 56006 35190 56058
rect 35242 56006 65654 56058
rect 65706 56006 65718 56058
rect 65770 56006 65782 56058
rect 65834 56006 65846 56058
rect 65898 56006 65910 56058
rect 65962 56006 68816 56058
rect 1104 55984 68816 56006
rect 1104 55514 68816 55536
rect 1104 55462 19574 55514
rect 19626 55462 19638 55514
rect 19690 55462 19702 55514
rect 19754 55462 19766 55514
rect 19818 55462 19830 55514
rect 19882 55462 50294 55514
rect 50346 55462 50358 55514
rect 50410 55462 50422 55514
rect 50474 55462 50486 55514
rect 50538 55462 50550 55514
rect 50602 55462 68816 55514
rect 1104 55440 68816 55462
rect 1104 54970 68816 54992
rect 1104 54918 4214 54970
rect 4266 54918 4278 54970
rect 4330 54918 4342 54970
rect 4394 54918 4406 54970
rect 4458 54918 4470 54970
rect 4522 54918 34934 54970
rect 34986 54918 34998 54970
rect 35050 54918 35062 54970
rect 35114 54918 35126 54970
rect 35178 54918 35190 54970
rect 35242 54918 65654 54970
rect 65706 54918 65718 54970
rect 65770 54918 65782 54970
rect 65834 54918 65846 54970
rect 65898 54918 65910 54970
rect 65962 54918 68816 54970
rect 1104 54896 68816 54918
rect 1104 54426 68816 54448
rect 1104 54374 19574 54426
rect 19626 54374 19638 54426
rect 19690 54374 19702 54426
rect 19754 54374 19766 54426
rect 19818 54374 19830 54426
rect 19882 54374 50294 54426
rect 50346 54374 50358 54426
rect 50410 54374 50422 54426
rect 50474 54374 50486 54426
rect 50538 54374 50550 54426
rect 50602 54374 68816 54426
rect 1104 54352 68816 54374
rect 1104 53882 68816 53904
rect 1104 53830 4214 53882
rect 4266 53830 4278 53882
rect 4330 53830 4342 53882
rect 4394 53830 4406 53882
rect 4458 53830 4470 53882
rect 4522 53830 34934 53882
rect 34986 53830 34998 53882
rect 35050 53830 35062 53882
rect 35114 53830 35126 53882
rect 35178 53830 35190 53882
rect 35242 53830 65654 53882
rect 65706 53830 65718 53882
rect 65770 53830 65782 53882
rect 65834 53830 65846 53882
rect 65898 53830 65910 53882
rect 65962 53830 68816 53882
rect 1104 53808 68816 53830
rect 1104 53338 68816 53360
rect 1104 53286 19574 53338
rect 19626 53286 19638 53338
rect 19690 53286 19702 53338
rect 19754 53286 19766 53338
rect 19818 53286 19830 53338
rect 19882 53286 50294 53338
rect 50346 53286 50358 53338
rect 50410 53286 50422 53338
rect 50474 53286 50486 53338
rect 50538 53286 50550 53338
rect 50602 53286 68816 53338
rect 1104 53264 68816 53286
rect 1104 52794 68816 52816
rect 1104 52742 4214 52794
rect 4266 52742 4278 52794
rect 4330 52742 4342 52794
rect 4394 52742 4406 52794
rect 4458 52742 4470 52794
rect 4522 52742 34934 52794
rect 34986 52742 34998 52794
rect 35050 52742 35062 52794
rect 35114 52742 35126 52794
rect 35178 52742 35190 52794
rect 35242 52742 65654 52794
rect 65706 52742 65718 52794
rect 65770 52742 65782 52794
rect 65834 52742 65846 52794
rect 65898 52742 65910 52794
rect 65962 52742 68816 52794
rect 1104 52720 68816 52742
rect 1104 52250 68816 52272
rect 1104 52198 19574 52250
rect 19626 52198 19638 52250
rect 19690 52198 19702 52250
rect 19754 52198 19766 52250
rect 19818 52198 19830 52250
rect 19882 52198 50294 52250
rect 50346 52198 50358 52250
rect 50410 52198 50422 52250
rect 50474 52198 50486 52250
rect 50538 52198 50550 52250
rect 50602 52198 68816 52250
rect 1104 52176 68816 52198
rect 1104 51706 68816 51728
rect 1104 51654 4214 51706
rect 4266 51654 4278 51706
rect 4330 51654 4342 51706
rect 4394 51654 4406 51706
rect 4458 51654 4470 51706
rect 4522 51654 34934 51706
rect 34986 51654 34998 51706
rect 35050 51654 35062 51706
rect 35114 51654 35126 51706
rect 35178 51654 35190 51706
rect 35242 51654 65654 51706
rect 65706 51654 65718 51706
rect 65770 51654 65782 51706
rect 65834 51654 65846 51706
rect 65898 51654 65910 51706
rect 65962 51654 68816 51706
rect 1104 51632 68816 51654
rect 1104 51162 68816 51184
rect 1104 51110 19574 51162
rect 19626 51110 19638 51162
rect 19690 51110 19702 51162
rect 19754 51110 19766 51162
rect 19818 51110 19830 51162
rect 19882 51110 50294 51162
rect 50346 51110 50358 51162
rect 50410 51110 50422 51162
rect 50474 51110 50486 51162
rect 50538 51110 50550 51162
rect 50602 51110 68816 51162
rect 1104 51088 68816 51110
rect 1104 50618 68816 50640
rect 1104 50566 4214 50618
rect 4266 50566 4278 50618
rect 4330 50566 4342 50618
rect 4394 50566 4406 50618
rect 4458 50566 4470 50618
rect 4522 50566 34934 50618
rect 34986 50566 34998 50618
rect 35050 50566 35062 50618
rect 35114 50566 35126 50618
rect 35178 50566 35190 50618
rect 35242 50566 65654 50618
rect 65706 50566 65718 50618
rect 65770 50566 65782 50618
rect 65834 50566 65846 50618
rect 65898 50566 65910 50618
rect 65962 50566 68816 50618
rect 1104 50544 68816 50566
rect 1104 50074 68816 50096
rect 1104 50022 19574 50074
rect 19626 50022 19638 50074
rect 19690 50022 19702 50074
rect 19754 50022 19766 50074
rect 19818 50022 19830 50074
rect 19882 50022 50294 50074
rect 50346 50022 50358 50074
rect 50410 50022 50422 50074
rect 50474 50022 50486 50074
rect 50538 50022 50550 50074
rect 50602 50022 68816 50074
rect 1104 50000 68816 50022
rect 1104 49530 68816 49552
rect 1104 49478 4214 49530
rect 4266 49478 4278 49530
rect 4330 49478 4342 49530
rect 4394 49478 4406 49530
rect 4458 49478 4470 49530
rect 4522 49478 34934 49530
rect 34986 49478 34998 49530
rect 35050 49478 35062 49530
rect 35114 49478 35126 49530
rect 35178 49478 35190 49530
rect 35242 49478 65654 49530
rect 65706 49478 65718 49530
rect 65770 49478 65782 49530
rect 65834 49478 65846 49530
rect 65898 49478 65910 49530
rect 65962 49478 68816 49530
rect 1104 49456 68816 49478
rect 1104 48986 68816 49008
rect 1104 48934 19574 48986
rect 19626 48934 19638 48986
rect 19690 48934 19702 48986
rect 19754 48934 19766 48986
rect 19818 48934 19830 48986
rect 19882 48934 50294 48986
rect 50346 48934 50358 48986
rect 50410 48934 50422 48986
rect 50474 48934 50486 48986
rect 50538 48934 50550 48986
rect 50602 48934 68816 48986
rect 1104 48912 68816 48934
rect 1104 48442 68816 48464
rect 1104 48390 4214 48442
rect 4266 48390 4278 48442
rect 4330 48390 4342 48442
rect 4394 48390 4406 48442
rect 4458 48390 4470 48442
rect 4522 48390 34934 48442
rect 34986 48390 34998 48442
rect 35050 48390 35062 48442
rect 35114 48390 35126 48442
rect 35178 48390 35190 48442
rect 35242 48390 65654 48442
rect 65706 48390 65718 48442
rect 65770 48390 65782 48442
rect 65834 48390 65846 48442
rect 65898 48390 65910 48442
rect 65962 48390 68816 48442
rect 1104 48368 68816 48390
rect 1104 47898 68816 47920
rect 1104 47846 19574 47898
rect 19626 47846 19638 47898
rect 19690 47846 19702 47898
rect 19754 47846 19766 47898
rect 19818 47846 19830 47898
rect 19882 47846 50294 47898
rect 50346 47846 50358 47898
rect 50410 47846 50422 47898
rect 50474 47846 50486 47898
rect 50538 47846 50550 47898
rect 50602 47846 68816 47898
rect 1104 47824 68816 47846
rect 1104 47354 68816 47376
rect 1104 47302 4214 47354
rect 4266 47302 4278 47354
rect 4330 47302 4342 47354
rect 4394 47302 4406 47354
rect 4458 47302 4470 47354
rect 4522 47302 34934 47354
rect 34986 47302 34998 47354
rect 35050 47302 35062 47354
rect 35114 47302 35126 47354
rect 35178 47302 35190 47354
rect 35242 47302 65654 47354
rect 65706 47302 65718 47354
rect 65770 47302 65782 47354
rect 65834 47302 65846 47354
rect 65898 47302 65910 47354
rect 65962 47302 68816 47354
rect 1104 47280 68816 47302
rect 1104 46810 68816 46832
rect 1104 46758 19574 46810
rect 19626 46758 19638 46810
rect 19690 46758 19702 46810
rect 19754 46758 19766 46810
rect 19818 46758 19830 46810
rect 19882 46758 50294 46810
rect 50346 46758 50358 46810
rect 50410 46758 50422 46810
rect 50474 46758 50486 46810
rect 50538 46758 50550 46810
rect 50602 46758 68816 46810
rect 1104 46736 68816 46758
rect 1104 46266 68816 46288
rect 1104 46214 4214 46266
rect 4266 46214 4278 46266
rect 4330 46214 4342 46266
rect 4394 46214 4406 46266
rect 4458 46214 4470 46266
rect 4522 46214 34934 46266
rect 34986 46214 34998 46266
rect 35050 46214 35062 46266
rect 35114 46214 35126 46266
rect 35178 46214 35190 46266
rect 35242 46214 65654 46266
rect 65706 46214 65718 46266
rect 65770 46214 65782 46266
rect 65834 46214 65846 46266
rect 65898 46214 65910 46266
rect 65962 46214 68816 46266
rect 1104 46192 68816 46214
rect 1104 45722 68816 45744
rect 1104 45670 19574 45722
rect 19626 45670 19638 45722
rect 19690 45670 19702 45722
rect 19754 45670 19766 45722
rect 19818 45670 19830 45722
rect 19882 45670 50294 45722
rect 50346 45670 50358 45722
rect 50410 45670 50422 45722
rect 50474 45670 50486 45722
rect 50538 45670 50550 45722
rect 50602 45670 68816 45722
rect 1104 45648 68816 45670
rect 1104 45178 68816 45200
rect 1104 45126 4214 45178
rect 4266 45126 4278 45178
rect 4330 45126 4342 45178
rect 4394 45126 4406 45178
rect 4458 45126 4470 45178
rect 4522 45126 34934 45178
rect 34986 45126 34998 45178
rect 35050 45126 35062 45178
rect 35114 45126 35126 45178
rect 35178 45126 35190 45178
rect 35242 45126 65654 45178
rect 65706 45126 65718 45178
rect 65770 45126 65782 45178
rect 65834 45126 65846 45178
rect 65898 45126 65910 45178
rect 65962 45126 68816 45178
rect 1104 45104 68816 45126
rect 1104 44634 68816 44656
rect 1104 44582 19574 44634
rect 19626 44582 19638 44634
rect 19690 44582 19702 44634
rect 19754 44582 19766 44634
rect 19818 44582 19830 44634
rect 19882 44582 50294 44634
rect 50346 44582 50358 44634
rect 50410 44582 50422 44634
rect 50474 44582 50486 44634
rect 50538 44582 50550 44634
rect 50602 44582 68816 44634
rect 1104 44560 68816 44582
rect 1104 44090 68816 44112
rect 1104 44038 4214 44090
rect 4266 44038 4278 44090
rect 4330 44038 4342 44090
rect 4394 44038 4406 44090
rect 4458 44038 4470 44090
rect 4522 44038 34934 44090
rect 34986 44038 34998 44090
rect 35050 44038 35062 44090
rect 35114 44038 35126 44090
rect 35178 44038 35190 44090
rect 35242 44038 65654 44090
rect 65706 44038 65718 44090
rect 65770 44038 65782 44090
rect 65834 44038 65846 44090
rect 65898 44038 65910 44090
rect 65962 44038 68816 44090
rect 1104 44016 68816 44038
rect 1104 43546 68816 43568
rect 1104 43494 19574 43546
rect 19626 43494 19638 43546
rect 19690 43494 19702 43546
rect 19754 43494 19766 43546
rect 19818 43494 19830 43546
rect 19882 43494 50294 43546
rect 50346 43494 50358 43546
rect 50410 43494 50422 43546
rect 50474 43494 50486 43546
rect 50538 43494 50550 43546
rect 50602 43494 68816 43546
rect 1104 43472 68816 43494
rect 1104 43002 68816 43024
rect 1104 42950 4214 43002
rect 4266 42950 4278 43002
rect 4330 42950 4342 43002
rect 4394 42950 4406 43002
rect 4458 42950 4470 43002
rect 4522 42950 34934 43002
rect 34986 42950 34998 43002
rect 35050 42950 35062 43002
rect 35114 42950 35126 43002
rect 35178 42950 35190 43002
rect 35242 42950 65654 43002
rect 65706 42950 65718 43002
rect 65770 42950 65782 43002
rect 65834 42950 65846 43002
rect 65898 42950 65910 43002
rect 65962 42950 68816 43002
rect 1104 42928 68816 42950
rect 1104 42458 68816 42480
rect 1104 42406 19574 42458
rect 19626 42406 19638 42458
rect 19690 42406 19702 42458
rect 19754 42406 19766 42458
rect 19818 42406 19830 42458
rect 19882 42406 50294 42458
rect 50346 42406 50358 42458
rect 50410 42406 50422 42458
rect 50474 42406 50486 42458
rect 50538 42406 50550 42458
rect 50602 42406 68816 42458
rect 1104 42384 68816 42406
rect 1104 41914 68816 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 34934 41914
rect 34986 41862 34998 41914
rect 35050 41862 35062 41914
rect 35114 41862 35126 41914
rect 35178 41862 35190 41914
rect 35242 41862 65654 41914
rect 65706 41862 65718 41914
rect 65770 41862 65782 41914
rect 65834 41862 65846 41914
rect 65898 41862 65910 41914
rect 65962 41862 68816 41914
rect 1104 41840 68816 41862
rect 1104 41370 68816 41392
rect 1104 41318 19574 41370
rect 19626 41318 19638 41370
rect 19690 41318 19702 41370
rect 19754 41318 19766 41370
rect 19818 41318 19830 41370
rect 19882 41318 50294 41370
rect 50346 41318 50358 41370
rect 50410 41318 50422 41370
rect 50474 41318 50486 41370
rect 50538 41318 50550 41370
rect 50602 41318 68816 41370
rect 1104 41296 68816 41318
rect 1104 40826 68816 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 34934 40826
rect 34986 40774 34998 40826
rect 35050 40774 35062 40826
rect 35114 40774 35126 40826
rect 35178 40774 35190 40826
rect 35242 40774 65654 40826
rect 65706 40774 65718 40826
rect 65770 40774 65782 40826
rect 65834 40774 65846 40826
rect 65898 40774 65910 40826
rect 65962 40774 68816 40826
rect 1104 40752 68816 40774
rect 1104 40282 68816 40304
rect 1104 40230 19574 40282
rect 19626 40230 19638 40282
rect 19690 40230 19702 40282
rect 19754 40230 19766 40282
rect 19818 40230 19830 40282
rect 19882 40230 50294 40282
rect 50346 40230 50358 40282
rect 50410 40230 50422 40282
rect 50474 40230 50486 40282
rect 50538 40230 50550 40282
rect 50602 40230 68816 40282
rect 1104 40208 68816 40230
rect 1104 39738 68816 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 65654 39738
rect 65706 39686 65718 39738
rect 65770 39686 65782 39738
rect 65834 39686 65846 39738
rect 65898 39686 65910 39738
rect 65962 39686 68816 39738
rect 1104 39664 68816 39686
rect 1104 39194 68816 39216
rect 1104 39142 19574 39194
rect 19626 39142 19638 39194
rect 19690 39142 19702 39194
rect 19754 39142 19766 39194
rect 19818 39142 19830 39194
rect 19882 39142 50294 39194
rect 50346 39142 50358 39194
rect 50410 39142 50422 39194
rect 50474 39142 50486 39194
rect 50538 39142 50550 39194
rect 50602 39142 68816 39194
rect 1104 39120 68816 39142
rect 1104 38650 68816 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 65654 38650
rect 65706 38598 65718 38650
rect 65770 38598 65782 38650
rect 65834 38598 65846 38650
rect 65898 38598 65910 38650
rect 65962 38598 68816 38650
rect 1104 38576 68816 38598
rect 1104 38106 68816 38128
rect 1104 38054 19574 38106
rect 19626 38054 19638 38106
rect 19690 38054 19702 38106
rect 19754 38054 19766 38106
rect 19818 38054 19830 38106
rect 19882 38054 50294 38106
rect 50346 38054 50358 38106
rect 50410 38054 50422 38106
rect 50474 38054 50486 38106
rect 50538 38054 50550 38106
rect 50602 38054 68816 38106
rect 1104 38032 68816 38054
rect 1104 37562 68816 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 65654 37562
rect 65706 37510 65718 37562
rect 65770 37510 65782 37562
rect 65834 37510 65846 37562
rect 65898 37510 65910 37562
rect 65962 37510 68816 37562
rect 1104 37488 68816 37510
rect 1104 37018 68816 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 50294 37018
rect 50346 36966 50358 37018
rect 50410 36966 50422 37018
rect 50474 36966 50486 37018
rect 50538 36966 50550 37018
rect 50602 36966 68816 37018
rect 1104 36944 68816 36966
rect 1104 36474 68816 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 65654 36474
rect 65706 36422 65718 36474
rect 65770 36422 65782 36474
rect 65834 36422 65846 36474
rect 65898 36422 65910 36474
rect 65962 36422 68816 36474
rect 1104 36400 68816 36422
rect 1104 35930 68816 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 50294 35930
rect 50346 35878 50358 35930
rect 50410 35878 50422 35930
rect 50474 35878 50486 35930
rect 50538 35878 50550 35930
rect 50602 35878 68816 35930
rect 1104 35856 68816 35878
rect 1104 35386 68816 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 65654 35386
rect 65706 35334 65718 35386
rect 65770 35334 65782 35386
rect 65834 35334 65846 35386
rect 65898 35334 65910 35386
rect 65962 35334 68816 35386
rect 1104 35312 68816 35334
rect 1104 34842 68816 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 50294 34842
rect 50346 34790 50358 34842
rect 50410 34790 50422 34842
rect 50474 34790 50486 34842
rect 50538 34790 50550 34842
rect 50602 34790 68816 34842
rect 1104 34768 68816 34790
rect 1104 34298 68816 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 65654 34298
rect 65706 34246 65718 34298
rect 65770 34246 65782 34298
rect 65834 34246 65846 34298
rect 65898 34246 65910 34298
rect 65962 34246 68816 34298
rect 1104 34224 68816 34246
rect 1104 33754 68816 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 50294 33754
rect 50346 33702 50358 33754
rect 50410 33702 50422 33754
rect 50474 33702 50486 33754
rect 50538 33702 50550 33754
rect 50602 33702 68816 33754
rect 1104 33680 68816 33702
rect 1104 33210 68816 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 65654 33210
rect 65706 33158 65718 33210
rect 65770 33158 65782 33210
rect 65834 33158 65846 33210
rect 65898 33158 65910 33210
rect 65962 33158 68816 33210
rect 1104 33136 68816 33158
rect 1104 32666 68816 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 50294 32666
rect 50346 32614 50358 32666
rect 50410 32614 50422 32666
rect 50474 32614 50486 32666
rect 50538 32614 50550 32666
rect 50602 32614 68816 32666
rect 1104 32592 68816 32614
rect 1104 32122 68816 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 65654 32122
rect 65706 32070 65718 32122
rect 65770 32070 65782 32122
rect 65834 32070 65846 32122
rect 65898 32070 65910 32122
rect 65962 32070 68816 32122
rect 1104 32048 68816 32070
rect 1104 31578 68816 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 50294 31578
rect 50346 31526 50358 31578
rect 50410 31526 50422 31578
rect 50474 31526 50486 31578
rect 50538 31526 50550 31578
rect 50602 31526 68816 31578
rect 1104 31504 68816 31526
rect 1104 31034 68816 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 65654 31034
rect 65706 30982 65718 31034
rect 65770 30982 65782 31034
rect 65834 30982 65846 31034
rect 65898 30982 65910 31034
rect 65962 30982 68816 31034
rect 1104 30960 68816 30982
rect 1104 30490 68816 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 50294 30490
rect 50346 30438 50358 30490
rect 50410 30438 50422 30490
rect 50474 30438 50486 30490
rect 50538 30438 50550 30490
rect 50602 30438 68816 30490
rect 1104 30416 68816 30438
rect 1104 29946 68816 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 65654 29946
rect 65706 29894 65718 29946
rect 65770 29894 65782 29946
rect 65834 29894 65846 29946
rect 65898 29894 65910 29946
rect 65962 29894 68816 29946
rect 1104 29872 68816 29894
rect 1104 29402 68816 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 50294 29402
rect 50346 29350 50358 29402
rect 50410 29350 50422 29402
rect 50474 29350 50486 29402
rect 50538 29350 50550 29402
rect 50602 29350 68816 29402
rect 1104 29328 68816 29350
rect 1104 28858 68816 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 65654 28858
rect 65706 28806 65718 28858
rect 65770 28806 65782 28858
rect 65834 28806 65846 28858
rect 65898 28806 65910 28858
rect 65962 28806 68816 28858
rect 1104 28784 68816 28806
rect 1104 28314 68816 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 50294 28314
rect 50346 28262 50358 28314
rect 50410 28262 50422 28314
rect 50474 28262 50486 28314
rect 50538 28262 50550 28314
rect 50602 28262 68816 28314
rect 1104 28240 68816 28262
rect 1104 27770 68816 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 65654 27770
rect 65706 27718 65718 27770
rect 65770 27718 65782 27770
rect 65834 27718 65846 27770
rect 65898 27718 65910 27770
rect 65962 27718 68816 27770
rect 1104 27696 68816 27718
rect 1104 27226 68816 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 50294 27226
rect 50346 27174 50358 27226
rect 50410 27174 50422 27226
rect 50474 27174 50486 27226
rect 50538 27174 50550 27226
rect 50602 27174 68816 27226
rect 1104 27152 68816 27174
rect 1104 26682 68816 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 65654 26682
rect 65706 26630 65718 26682
rect 65770 26630 65782 26682
rect 65834 26630 65846 26682
rect 65898 26630 65910 26682
rect 65962 26630 68816 26682
rect 1104 26608 68816 26630
rect 1104 26138 68816 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 50294 26138
rect 50346 26086 50358 26138
rect 50410 26086 50422 26138
rect 50474 26086 50486 26138
rect 50538 26086 50550 26138
rect 50602 26086 68816 26138
rect 1104 26064 68816 26086
rect 1104 25594 68816 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 65654 25594
rect 65706 25542 65718 25594
rect 65770 25542 65782 25594
rect 65834 25542 65846 25594
rect 65898 25542 65910 25594
rect 65962 25542 68816 25594
rect 1104 25520 68816 25542
rect 1104 25050 68816 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 50294 25050
rect 50346 24998 50358 25050
rect 50410 24998 50422 25050
rect 50474 24998 50486 25050
rect 50538 24998 50550 25050
rect 50602 24998 68816 25050
rect 1104 24976 68816 24998
rect 1104 24506 68816 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 65654 24506
rect 65706 24454 65718 24506
rect 65770 24454 65782 24506
rect 65834 24454 65846 24506
rect 65898 24454 65910 24506
rect 65962 24454 68816 24506
rect 1104 24432 68816 24454
rect 1104 23962 68816 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 50294 23962
rect 50346 23910 50358 23962
rect 50410 23910 50422 23962
rect 50474 23910 50486 23962
rect 50538 23910 50550 23962
rect 50602 23910 68816 23962
rect 1104 23888 68816 23910
rect 1104 23418 68816 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 65654 23418
rect 65706 23366 65718 23418
rect 65770 23366 65782 23418
rect 65834 23366 65846 23418
rect 65898 23366 65910 23418
rect 65962 23366 68816 23418
rect 1104 23344 68816 23366
rect 1104 22874 68816 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 50294 22874
rect 50346 22822 50358 22874
rect 50410 22822 50422 22874
rect 50474 22822 50486 22874
rect 50538 22822 50550 22874
rect 50602 22822 68816 22874
rect 1104 22800 68816 22822
rect 1104 22330 68816 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 65654 22330
rect 65706 22278 65718 22330
rect 65770 22278 65782 22330
rect 65834 22278 65846 22330
rect 65898 22278 65910 22330
rect 65962 22278 68816 22330
rect 1104 22256 68816 22278
rect 1104 21786 68816 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 50294 21786
rect 50346 21734 50358 21786
rect 50410 21734 50422 21786
rect 50474 21734 50486 21786
rect 50538 21734 50550 21786
rect 50602 21734 68816 21786
rect 1104 21712 68816 21734
rect 1104 21242 68816 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 65654 21242
rect 65706 21190 65718 21242
rect 65770 21190 65782 21242
rect 65834 21190 65846 21242
rect 65898 21190 65910 21242
rect 65962 21190 68816 21242
rect 1104 21168 68816 21190
rect 1104 20698 68816 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 50294 20698
rect 50346 20646 50358 20698
rect 50410 20646 50422 20698
rect 50474 20646 50486 20698
rect 50538 20646 50550 20698
rect 50602 20646 68816 20698
rect 1104 20624 68816 20646
rect 1104 20154 68816 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 65654 20154
rect 65706 20102 65718 20154
rect 65770 20102 65782 20154
rect 65834 20102 65846 20154
rect 65898 20102 65910 20154
rect 65962 20102 68816 20154
rect 1104 20080 68816 20102
rect 1104 19610 68816 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 50294 19610
rect 50346 19558 50358 19610
rect 50410 19558 50422 19610
rect 50474 19558 50486 19610
rect 50538 19558 50550 19610
rect 50602 19558 68816 19610
rect 1104 19536 68816 19558
rect 1104 19066 68816 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 65654 19066
rect 65706 19014 65718 19066
rect 65770 19014 65782 19066
rect 65834 19014 65846 19066
rect 65898 19014 65910 19066
rect 65962 19014 68816 19066
rect 1104 18992 68816 19014
rect 1104 18522 68816 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 50294 18522
rect 50346 18470 50358 18522
rect 50410 18470 50422 18522
rect 50474 18470 50486 18522
rect 50538 18470 50550 18522
rect 50602 18470 68816 18522
rect 1104 18448 68816 18470
rect 1104 17978 68816 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 65654 17978
rect 65706 17926 65718 17978
rect 65770 17926 65782 17978
rect 65834 17926 65846 17978
rect 65898 17926 65910 17978
rect 65962 17926 68816 17978
rect 1104 17904 68816 17926
rect 1104 17434 68816 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 50294 17434
rect 50346 17382 50358 17434
rect 50410 17382 50422 17434
rect 50474 17382 50486 17434
rect 50538 17382 50550 17434
rect 50602 17382 68816 17434
rect 1104 17360 68816 17382
rect 1104 16890 68816 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 65654 16890
rect 65706 16838 65718 16890
rect 65770 16838 65782 16890
rect 65834 16838 65846 16890
rect 65898 16838 65910 16890
rect 65962 16838 68816 16890
rect 1104 16816 68816 16838
rect 1104 16346 68816 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 50294 16346
rect 50346 16294 50358 16346
rect 50410 16294 50422 16346
rect 50474 16294 50486 16346
rect 50538 16294 50550 16346
rect 50602 16294 68816 16346
rect 1104 16272 68816 16294
rect 1104 15802 68816 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 65654 15802
rect 65706 15750 65718 15802
rect 65770 15750 65782 15802
rect 65834 15750 65846 15802
rect 65898 15750 65910 15802
rect 65962 15750 68816 15802
rect 1104 15728 68816 15750
rect 1104 15258 68816 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 50294 15258
rect 50346 15206 50358 15258
rect 50410 15206 50422 15258
rect 50474 15206 50486 15258
rect 50538 15206 50550 15258
rect 50602 15206 68816 15258
rect 1104 15184 68816 15206
rect 1104 14714 68816 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 65654 14714
rect 65706 14662 65718 14714
rect 65770 14662 65782 14714
rect 65834 14662 65846 14714
rect 65898 14662 65910 14714
rect 65962 14662 68816 14714
rect 1104 14640 68816 14662
rect 11698 14424 11704 14476
rect 11756 14464 11762 14476
rect 11756 14436 12020 14464
rect 11756 14424 11762 14436
rect 10502 14356 10508 14408
rect 10560 14396 10566 14408
rect 11992 14405 12020 14436
rect 11885 14399 11943 14405
rect 10560 14390 11744 14396
rect 11885 14390 11897 14399
rect 10560 14368 11897 14390
rect 10560 14356 10566 14368
rect 11716 14365 11897 14368
rect 11931 14365 11943 14399
rect 11716 14362 11943 14365
rect 11885 14359 11943 14362
rect 11977 14399 12035 14405
rect 12253 14399 12311 14405
rect 11977 14365 11989 14399
rect 12023 14365 12035 14399
rect 11977 14359 12035 14365
rect 12090 14393 12148 14399
rect 12090 14359 12102 14393
rect 12136 14390 12148 14393
rect 12136 14362 12204 14390
rect 12136 14359 12148 14362
rect 12090 14353 12148 14359
rect 10410 14288 10416 14340
rect 10468 14328 10474 14340
rect 10468 14300 11744 14328
rect 10468 14288 10474 14300
rect 4338 14220 4344 14272
rect 4396 14260 4402 14272
rect 5074 14260 5080 14272
rect 4396 14232 5080 14260
rect 4396 14220 4402 14232
rect 5074 14220 5080 14232
rect 5132 14260 5138 14272
rect 11422 14260 11428 14272
rect 5132 14232 11428 14260
rect 5132 14220 5138 14232
rect 11422 14220 11428 14232
rect 11480 14220 11486 14272
rect 11606 14260 11612 14272
rect 11567 14232 11612 14260
rect 11606 14220 11612 14232
rect 11664 14220 11670 14272
rect 11716 14260 11744 14300
rect 12176 14260 12204 14362
rect 12253 14365 12265 14399
rect 12299 14396 12311 14399
rect 12434 14396 12440 14408
rect 12299 14368 12440 14396
rect 12299 14365 12311 14368
rect 12253 14359 12311 14365
rect 12434 14356 12440 14368
rect 12492 14356 12498 14408
rect 15194 14356 15200 14408
rect 15252 14396 15258 14408
rect 15289 14399 15347 14405
rect 15289 14396 15301 14399
rect 15252 14368 15301 14396
rect 15252 14356 15258 14368
rect 15289 14365 15301 14368
rect 15335 14365 15347 14399
rect 15289 14359 15347 14365
rect 15378 14399 15436 14405
rect 15378 14365 15390 14399
rect 15424 14365 15436 14399
rect 15378 14359 15436 14365
rect 15494 14399 15552 14405
rect 15494 14365 15506 14399
rect 15540 14396 15552 14399
rect 15657 14399 15715 14405
rect 15540 14368 15608 14396
rect 15540 14365 15552 14368
rect 15494 14359 15552 14365
rect 15010 14260 15016 14272
rect 11716 14232 12204 14260
rect 14971 14232 15016 14260
rect 15010 14220 15016 14232
rect 15068 14220 15074 14272
rect 15396 14260 15424 14359
rect 15580 14328 15608 14368
rect 15657 14365 15669 14399
rect 15703 14396 15715 14399
rect 16850 14396 16856 14408
rect 15703 14368 16856 14396
rect 15703 14365 15715 14368
rect 15657 14359 15715 14365
rect 16850 14356 16856 14368
rect 16908 14356 16914 14408
rect 16298 14328 16304 14340
rect 15580 14300 16304 14328
rect 16298 14288 16304 14300
rect 16356 14288 16362 14340
rect 15654 14260 15660 14272
rect 15396 14232 15660 14260
rect 15654 14220 15660 14232
rect 15712 14220 15718 14272
rect 1104 14170 68816 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 50294 14170
rect 50346 14118 50358 14170
rect 50410 14118 50422 14170
rect 50474 14118 50486 14170
rect 50538 14118 50550 14170
rect 50602 14118 68816 14170
rect 1104 14096 68816 14118
rect 4338 14056 4344 14068
rect 4299 14028 4344 14056
rect 4338 14016 4344 14028
rect 4396 14016 4402 14068
rect 8389 14059 8447 14065
rect 8389 14025 8401 14059
rect 8435 14025 8447 14059
rect 8389 14019 8447 14025
rect 8404 13988 8432 14019
rect 11422 14016 11428 14068
rect 11480 14056 11486 14068
rect 14185 14059 14243 14065
rect 14185 14056 14197 14059
rect 11480 14028 14197 14056
rect 11480 14016 11486 14028
rect 14185 14025 14197 14028
rect 14231 14056 14243 14059
rect 14734 14056 14740 14068
rect 14231 14028 14740 14056
rect 14231 14025 14243 14028
rect 14185 14019 14243 14025
rect 14734 14016 14740 14028
rect 14792 14016 14798 14068
rect 8404 13960 10824 13988
rect 10796 13932 10824 13960
rect 12894 13948 12900 14000
rect 12952 13988 12958 14000
rect 12952 13960 15056 13988
rect 12952 13948 12958 13960
rect 4249 13923 4307 13929
rect 4249 13889 4261 13923
rect 4295 13889 4307 13923
rect 4249 13883 4307 13889
rect 4433 13923 4491 13929
rect 4433 13889 4445 13923
rect 4479 13920 4491 13923
rect 5810 13920 5816 13932
rect 4479 13892 5816 13920
rect 4479 13889 4491 13892
rect 4433 13883 4491 13889
rect 4264 13852 4292 13883
rect 5810 13880 5816 13892
rect 5868 13920 5874 13932
rect 7285 13923 7343 13929
rect 7285 13920 7297 13923
rect 5868 13892 7297 13920
rect 5868 13880 5874 13892
rect 7285 13889 7297 13892
rect 7331 13889 7343 13923
rect 7285 13883 7343 13889
rect 8021 13923 8079 13929
rect 8021 13889 8033 13923
rect 8067 13920 8079 13923
rect 8846 13920 8852 13932
rect 8067 13892 8852 13920
rect 8067 13889 8079 13892
rect 8021 13883 8079 13889
rect 8846 13880 8852 13892
rect 8904 13880 8910 13932
rect 10594 13920 10600 13932
rect 10555 13892 10600 13920
rect 10594 13880 10600 13892
rect 10652 13880 10658 13932
rect 10686 13923 10744 13929
rect 10686 13889 10698 13923
rect 10732 13889 10744 13923
rect 10686 13883 10744 13889
rect 10781 13926 10839 13932
rect 10781 13892 10793 13926
rect 10827 13892 10839 13926
rect 10781 13886 10839 13892
rect 10965 13923 11023 13929
rect 10965 13889 10977 13923
rect 11011 13920 11023 13923
rect 11146 13920 11152 13932
rect 11011 13892 11152 13920
rect 11011 13889 11023 13892
rect 10965 13883 11023 13889
rect 4985 13855 5043 13861
rect 4985 13852 4997 13855
rect 4264 13824 4997 13852
rect 4985 13821 4997 13824
rect 5031 13852 5043 13855
rect 8110 13852 8116 13864
rect 5031 13824 7328 13852
rect 8071 13824 8116 13852
rect 5031 13821 5043 13824
rect 4985 13815 5043 13821
rect 7300 13796 7328 13824
rect 8110 13812 8116 13824
rect 8168 13812 8174 13864
rect 8754 13812 8760 13864
rect 8812 13852 8818 13864
rect 8941 13855 8999 13861
rect 8941 13852 8953 13855
rect 8812 13824 8953 13852
rect 8812 13812 8818 13824
rect 8941 13821 8953 13824
rect 8987 13821 8999 13855
rect 8941 13815 8999 13821
rect 9858 13812 9864 13864
rect 9916 13852 9922 13864
rect 10321 13855 10379 13861
rect 10321 13852 10333 13855
rect 9916 13824 10333 13852
rect 9916 13812 9922 13824
rect 10321 13821 10333 13824
rect 10367 13821 10379 13855
rect 10704 13852 10732 13883
rect 11146 13880 11152 13892
rect 11204 13920 11210 13932
rect 12069 13923 12127 13929
rect 12069 13920 12081 13923
rect 11204 13892 12081 13920
rect 11204 13880 11210 13892
rect 12069 13889 12081 13892
rect 12115 13920 12127 13923
rect 12434 13920 12440 13932
rect 12115 13892 12440 13920
rect 12115 13889 12127 13892
rect 12069 13883 12127 13889
rect 12434 13880 12440 13892
rect 12492 13920 12498 13932
rect 13078 13920 13084 13932
rect 12492 13892 13084 13920
rect 12492 13880 12498 13892
rect 13078 13880 13084 13892
rect 13136 13880 13142 13932
rect 13372 13929 13400 13960
rect 15028 13929 15056 13960
rect 13244 13923 13302 13929
rect 13244 13920 13256 13923
rect 13188 13892 13256 13920
rect 10870 13852 10876 13864
rect 10704 13824 10876 13852
rect 10321 13815 10379 13821
rect 10870 13812 10876 13824
rect 10928 13812 10934 13864
rect 11514 13812 11520 13864
rect 11572 13852 11578 13864
rect 12345 13855 12403 13861
rect 12345 13852 12357 13855
rect 11572 13824 12357 13852
rect 11572 13812 11578 13824
rect 12345 13821 12357 13824
rect 12391 13821 12403 13855
rect 12345 13815 12403 13821
rect 12710 13812 12716 13864
rect 12768 13852 12774 13864
rect 13188 13852 13216 13892
rect 13244 13889 13256 13892
rect 13290 13889 13302 13923
rect 13244 13883 13302 13889
rect 13357 13923 13415 13929
rect 13357 13889 13369 13923
rect 13403 13889 13415 13923
rect 13357 13883 13415 13889
rect 13449 13923 13507 13929
rect 13449 13889 13461 13923
rect 13495 13889 13507 13923
rect 13449 13883 13507 13889
rect 15013 13923 15071 13929
rect 15013 13889 15025 13923
rect 15059 13889 15071 13923
rect 15013 13883 15071 13889
rect 12768 13824 13216 13852
rect 12768 13812 12774 13824
rect 7282 13744 7288 13796
rect 7340 13744 7346 13796
rect 10778 13744 10784 13796
rect 10836 13784 10842 13796
rect 11698 13784 11704 13796
rect 10836 13756 11704 13784
rect 10836 13744 10842 13756
rect 11698 13744 11704 13756
rect 11756 13744 11762 13796
rect 12158 13744 12164 13796
rect 12216 13784 12222 13796
rect 13464 13784 13492 13883
rect 13722 13852 13728 13864
rect 13683 13824 13728 13852
rect 13722 13812 13728 13824
rect 13780 13812 13786 13864
rect 14734 13852 14740 13864
rect 14695 13824 14740 13852
rect 14734 13812 14740 13824
rect 14792 13852 14798 13864
rect 21542 13852 21548 13864
rect 14792 13824 21548 13852
rect 14792 13812 14798 13824
rect 21542 13812 21548 13824
rect 21600 13812 21606 13864
rect 12216 13756 13492 13784
rect 12216 13744 12222 13756
rect 7469 13719 7527 13725
rect 7469 13685 7481 13719
rect 7515 13716 7527 13719
rect 8205 13719 8263 13725
rect 8205 13716 8217 13719
rect 7515 13688 8217 13716
rect 7515 13685 7527 13688
rect 7469 13679 7527 13685
rect 8205 13685 8217 13688
rect 8251 13716 8263 13719
rect 9030 13716 9036 13728
rect 8251 13688 9036 13716
rect 8251 13685 8263 13688
rect 8205 13679 8263 13685
rect 9030 13676 9036 13688
rect 9088 13676 9094 13728
rect 9217 13719 9275 13725
rect 9217 13685 9229 13719
rect 9263 13716 9275 13719
rect 13078 13716 13084 13728
rect 9263 13688 13084 13716
rect 9263 13685 9275 13688
rect 9217 13679 9275 13685
rect 13078 13676 13084 13688
rect 13136 13676 13142 13728
rect 1104 13626 68816 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 65654 13626
rect 65706 13574 65718 13626
rect 65770 13574 65782 13626
rect 65834 13574 65846 13626
rect 65898 13574 65910 13626
rect 65962 13574 68816 13626
rect 1104 13552 68816 13574
rect 8113 13515 8171 13521
rect 8113 13481 8125 13515
rect 8159 13512 8171 13515
rect 9030 13512 9036 13524
rect 8159 13484 9036 13512
rect 8159 13481 8171 13484
rect 8113 13475 8171 13481
rect 9030 13472 9036 13484
rect 9088 13472 9094 13524
rect 10410 13512 10416 13524
rect 9232 13484 10416 13512
rect 8297 13447 8355 13453
rect 8297 13413 8309 13447
rect 8343 13444 8355 13447
rect 9232 13444 9260 13484
rect 10410 13472 10416 13484
rect 10468 13472 10474 13524
rect 10520 13484 11468 13512
rect 8343 13416 9260 13444
rect 9309 13447 9367 13453
rect 8343 13413 8355 13416
rect 8297 13407 8355 13413
rect 9309 13413 9321 13447
rect 9355 13444 9367 13447
rect 10520 13444 10548 13484
rect 10778 13444 10784 13456
rect 9355 13416 10548 13444
rect 10717 13416 10784 13444
rect 9355 13413 9367 13416
rect 9309 13407 9367 13413
rect 7282 13308 7288 13320
rect 7243 13280 7288 13308
rect 7282 13268 7288 13280
rect 7340 13268 7346 13320
rect 7929 13311 7987 13317
rect 7929 13277 7941 13311
rect 7975 13277 7987 13311
rect 7929 13271 7987 13277
rect 8113 13311 8171 13317
rect 8113 13277 8125 13311
rect 8159 13308 8171 13311
rect 8570 13308 8576 13320
rect 8159 13280 8576 13308
rect 8159 13277 8171 13280
rect 8113 13271 8171 13277
rect 7944 13240 7972 13271
rect 8570 13268 8576 13280
rect 8628 13268 8634 13320
rect 8938 13308 8944 13320
rect 8899 13280 8944 13308
rect 8938 13268 8944 13280
rect 8996 13268 9002 13320
rect 9125 13311 9183 13317
rect 9125 13277 9137 13311
rect 9171 13308 9183 13311
rect 9214 13308 9220 13320
rect 9171 13280 9220 13308
rect 9171 13277 9183 13280
rect 9125 13271 9183 13277
rect 9214 13268 9220 13280
rect 9272 13268 9278 13320
rect 10551 13311 10609 13317
rect 10717 13311 10745 13416
rect 10778 13404 10784 13416
rect 10836 13404 10842 13456
rect 11440 13444 11468 13484
rect 11514 13472 11520 13524
rect 11572 13512 11578 13524
rect 12710 13512 12716 13524
rect 11572 13484 11617 13512
rect 12176 13484 12716 13512
rect 11572 13472 11578 13484
rect 12176 13444 12204 13484
rect 12710 13472 12716 13484
rect 12768 13472 12774 13524
rect 11440 13416 12204 13444
rect 12894 13404 12900 13456
rect 12952 13404 12958 13456
rect 16850 13444 16856 13456
rect 15764 13416 16856 13444
rect 10551 13277 10563 13311
rect 10597 13277 10609 13311
rect 10551 13271 10609 13277
rect 8956 13240 8984 13268
rect 7944 13212 8984 13240
rect 10581 13240 10609 13271
rect 10702 13305 10760 13311
rect 10702 13271 10714 13305
rect 10748 13271 10760 13305
rect 10702 13265 10760 13271
rect 10799 13262 10805 13314
rect 10857 13302 10863 13314
rect 10965 13311 11023 13317
rect 10857 13274 10902 13302
rect 10965 13277 10977 13311
rect 11011 13308 11023 13311
rect 11146 13308 11152 13320
rect 11011 13280 11152 13308
rect 11011 13277 11023 13280
rect 10857 13262 10863 13274
rect 10965 13271 11023 13277
rect 11146 13268 11152 13280
rect 11204 13268 11210 13320
rect 12909 13317 12937 13404
rect 13078 13336 13084 13388
rect 13136 13336 13142 13388
rect 15654 13376 15660 13388
rect 15488 13348 15660 13376
rect 12805 13311 12863 13317
rect 12805 13277 12817 13311
rect 12851 13277 12863 13311
rect 12805 13271 12863 13277
rect 12894 13311 12952 13317
rect 12894 13277 12906 13311
rect 12940 13277 12952 13311
rect 12894 13271 12952 13277
rect 12994 13305 13052 13311
rect 12994 13271 13006 13305
rect 13040 13284 13052 13305
rect 13096 13284 13124 13336
rect 13040 13271 13124 13284
rect 10581 13212 10640 13240
rect 7469 13175 7527 13181
rect 7469 13141 7481 13175
rect 7515 13172 7527 13175
rect 7944 13172 7972 13212
rect 10318 13172 10324 13184
rect 7515 13144 7972 13172
rect 10279 13144 10324 13172
rect 7515 13141 7527 13144
rect 7469 13135 7527 13141
rect 10318 13132 10324 13144
rect 10376 13132 10382 13184
rect 10612 13172 10640 13212
rect 11422 13172 11428 13184
rect 10612 13144 11428 13172
rect 11422 13132 11428 13144
rect 11480 13132 11486 13184
rect 12526 13172 12532 13184
rect 12487 13144 12532 13172
rect 12526 13132 12532 13144
rect 12584 13132 12590 13184
rect 12820 13172 12848 13271
rect 12994 13265 13124 13271
rect 13170 13268 13176 13320
rect 13228 13317 13234 13320
rect 13228 13311 13243 13317
rect 13231 13277 13243 13311
rect 13228 13271 13243 13277
rect 13228 13268 13234 13271
rect 15286 13268 15292 13320
rect 15344 13308 15350 13320
rect 15488 13317 15516 13348
rect 15654 13336 15660 13348
rect 15712 13336 15718 13388
rect 15764 13317 15792 13416
rect 16850 13404 16856 13416
rect 16908 13404 16914 13456
rect 15381 13311 15439 13317
rect 15381 13308 15393 13311
rect 15344 13280 15393 13308
rect 15344 13268 15350 13280
rect 15381 13277 15393 13280
rect 15427 13277 15439 13311
rect 15381 13271 15439 13277
rect 15470 13311 15528 13317
rect 15470 13277 15482 13311
rect 15516 13277 15528 13311
rect 15470 13271 15528 13277
rect 15565 13311 15623 13317
rect 15565 13277 15577 13311
rect 15611 13308 15623 13311
rect 15761 13311 15819 13317
rect 15611 13280 15691 13308
rect 15611 13277 15623 13280
rect 15565 13271 15623 13277
rect 13004 13256 13124 13265
rect 15663 13240 15691 13280
rect 15761 13277 15773 13311
rect 15807 13277 15819 13311
rect 15761 13271 15819 13277
rect 16390 13268 16396 13320
rect 16448 13317 16454 13320
rect 16448 13311 16497 13317
rect 16448 13277 16451 13311
rect 16485 13277 16497 13311
rect 16448 13271 16497 13277
rect 16574 13308 16632 13314
rect 16574 13274 16586 13308
rect 16620 13274 16632 13308
rect 16448 13268 16454 13271
rect 16574 13268 16632 13274
rect 16666 13268 16672 13320
rect 16724 13317 16730 13320
rect 16724 13308 16732 13317
rect 16724 13280 16769 13308
rect 16724 13271 16732 13280
rect 16724 13268 16730 13271
rect 16850 13268 16856 13320
rect 16908 13308 16914 13320
rect 17310 13308 17316 13320
rect 16908 13280 17316 13308
rect 16908 13268 16914 13280
rect 17310 13268 17316 13280
rect 17368 13268 17374 13320
rect 16592 13240 16620 13268
rect 15663 13212 16436 13240
rect 16592 13212 16712 13240
rect 16408 13184 16436 13212
rect 13262 13172 13268 13184
rect 12820 13144 13268 13172
rect 13262 13132 13268 13144
rect 13320 13132 13326 13184
rect 14918 13132 14924 13184
rect 14976 13172 14982 13184
rect 15105 13175 15163 13181
rect 15105 13172 15117 13175
rect 14976 13144 15117 13172
rect 14976 13132 14982 13144
rect 15105 13141 15117 13144
rect 15151 13141 15163 13175
rect 16206 13172 16212 13184
rect 16167 13144 16212 13172
rect 15105 13135 15163 13141
rect 16206 13132 16212 13144
rect 16264 13132 16270 13184
rect 16390 13132 16396 13184
rect 16448 13132 16454 13184
rect 16574 13132 16580 13184
rect 16632 13172 16638 13184
rect 16684 13172 16712 13212
rect 16632 13144 16712 13172
rect 16632 13132 16638 13144
rect 1104 13082 68816 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 50294 13082
rect 50346 13030 50358 13082
rect 50410 13030 50422 13082
rect 50474 13030 50486 13082
rect 50538 13030 50550 13082
rect 50602 13030 68816 13082
rect 1104 13008 68816 13030
rect 9401 12971 9459 12977
rect 9401 12937 9413 12971
rect 9447 12968 9459 12971
rect 10778 12968 10784 12980
rect 9447 12940 10784 12968
rect 9447 12937 9459 12940
rect 9401 12931 9459 12937
rect 10778 12928 10784 12940
rect 10836 12928 10842 12980
rect 15654 12928 15660 12980
rect 15712 12968 15718 12980
rect 16574 12968 16580 12980
rect 15712 12940 16580 12968
rect 15712 12928 15718 12940
rect 16574 12928 16580 12940
rect 16632 12928 16638 12980
rect 13716 12903 13774 12909
rect 13716 12869 13728 12903
rect 13762 12900 13774 12903
rect 15010 12900 15016 12912
rect 13762 12872 15016 12900
rect 13762 12869 13774 12872
rect 13716 12863 13774 12869
rect 15010 12860 15016 12872
rect 15068 12860 15074 12912
rect 4706 12832 4712 12844
rect 4667 12804 4712 12832
rect 4706 12792 4712 12804
rect 4764 12792 4770 12844
rect 4888 12835 4946 12841
rect 4888 12801 4900 12835
rect 4934 12801 4946 12835
rect 4888 12795 4946 12801
rect 4985 12835 5043 12841
rect 4985 12801 4997 12835
rect 5031 12801 5043 12835
rect 4985 12795 5043 12801
rect 5123 12835 5181 12841
rect 5123 12801 5135 12835
rect 5169 12832 5181 12835
rect 8754 12832 8760 12844
rect 5169 12804 8760 12832
rect 5169 12801 5181 12804
rect 5123 12795 5181 12801
rect 4614 12724 4620 12776
rect 4672 12764 4678 12776
rect 4903 12764 4931 12795
rect 4672 12736 4931 12764
rect 5000 12764 5028 12795
rect 8754 12792 8760 12804
rect 8812 12792 8818 12844
rect 8938 12792 8944 12844
rect 8996 12832 9002 12844
rect 9033 12835 9091 12841
rect 9033 12832 9045 12835
rect 8996 12804 9045 12832
rect 8996 12792 9002 12804
rect 9033 12801 9045 12804
rect 9079 12801 9091 12835
rect 9033 12795 9091 12801
rect 13449 12835 13507 12841
rect 13449 12801 13461 12835
rect 13495 12832 13507 12835
rect 13538 12832 13544 12844
rect 13495 12804 13544 12832
rect 13495 12801 13507 12804
rect 13449 12795 13507 12801
rect 13538 12792 13544 12804
rect 13596 12792 13602 12844
rect 15841 12835 15899 12841
rect 15841 12801 15853 12835
rect 15887 12832 15899 12835
rect 21726 12832 21732 12844
rect 15887 12804 21732 12832
rect 15887 12801 15899 12804
rect 15841 12795 15899 12801
rect 21726 12792 21732 12804
rect 21784 12792 21790 12844
rect 6178 12764 6184 12776
rect 5000 12736 6184 12764
rect 4672 12724 4678 12736
rect 6178 12724 6184 12736
rect 6236 12724 6242 12776
rect 8386 12724 8392 12776
rect 8444 12764 8450 12776
rect 9125 12767 9183 12773
rect 9125 12764 9137 12767
rect 8444 12736 9137 12764
rect 8444 12724 8450 12736
rect 9125 12733 9137 12736
rect 9171 12733 9183 12767
rect 16114 12764 16120 12776
rect 16075 12736 16120 12764
rect 9125 12727 9183 12733
rect 16114 12724 16120 12736
rect 16172 12724 16178 12776
rect 5353 12699 5411 12705
rect 5353 12665 5365 12699
rect 5399 12696 5411 12699
rect 10134 12696 10140 12708
rect 5399 12668 10140 12696
rect 5399 12665 5411 12668
rect 5353 12659 5411 12665
rect 10134 12656 10140 12668
rect 10192 12656 10198 12708
rect 7282 12588 7288 12640
rect 7340 12628 7346 12640
rect 7653 12631 7711 12637
rect 7653 12628 7665 12631
rect 7340 12600 7665 12628
rect 7340 12588 7346 12600
rect 7653 12597 7665 12600
rect 7699 12628 7711 12631
rect 8846 12628 8852 12640
rect 7699 12600 8852 12628
rect 7699 12597 7711 12600
rect 7653 12591 7711 12597
rect 8846 12588 8852 12600
rect 8904 12588 8910 12640
rect 9030 12628 9036 12640
rect 8991 12600 9036 12628
rect 9030 12588 9036 12600
rect 9088 12588 9094 12640
rect 14829 12631 14887 12637
rect 14829 12597 14841 12631
rect 14875 12628 14887 12631
rect 15194 12628 15200 12640
rect 14875 12600 15200 12628
rect 14875 12597 14887 12600
rect 14829 12591 14887 12597
rect 15194 12588 15200 12600
rect 15252 12628 15258 12640
rect 20070 12628 20076 12640
rect 15252 12600 20076 12628
rect 15252 12588 15258 12600
rect 20070 12588 20076 12600
rect 20128 12588 20134 12640
rect 1104 12538 68816 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 65654 12538
rect 65706 12486 65718 12538
rect 65770 12486 65782 12538
rect 65834 12486 65846 12538
rect 65898 12486 65910 12538
rect 65962 12486 68816 12538
rect 1104 12464 68816 12486
rect 22833 12427 22891 12433
rect 22833 12424 22845 12427
rect 17236 12396 22845 12424
rect 4706 12248 4712 12300
rect 4764 12288 4770 12300
rect 5261 12291 5319 12297
rect 5261 12288 5273 12291
rect 4764 12260 5273 12288
rect 4764 12248 4770 12260
rect 5261 12257 5273 12260
rect 5307 12257 5319 12291
rect 5261 12251 5319 12257
rect 5534 12220 5540 12232
rect 5495 12192 5540 12220
rect 5534 12180 5540 12192
rect 5592 12180 5598 12232
rect 7009 12223 7067 12229
rect 7009 12189 7021 12223
rect 7055 12220 7067 12223
rect 7098 12220 7104 12232
rect 7055 12192 7104 12220
rect 7055 12189 7067 12192
rect 7009 12183 7067 12189
rect 7098 12180 7104 12192
rect 7156 12180 7162 12232
rect 10137 12223 10195 12229
rect 10137 12189 10149 12223
rect 10183 12220 10195 12223
rect 11698 12220 11704 12232
rect 10183 12192 11704 12220
rect 10183 12189 10195 12192
rect 10137 12183 10195 12189
rect 11698 12180 11704 12192
rect 11756 12220 11762 12232
rect 11977 12223 12035 12229
rect 11977 12220 11989 12223
rect 11756 12192 11989 12220
rect 11756 12180 11762 12192
rect 11977 12189 11989 12192
rect 12023 12189 12035 12223
rect 11977 12183 12035 12189
rect 12244 12223 12302 12229
rect 12244 12189 12256 12223
rect 12290 12220 12302 12223
rect 12526 12220 12532 12232
rect 12290 12192 12532 12220
rect 12290 12189 12302 12192
rect 12244 12183 12302 12189
rect 12526 12180 12532 12192
rect 12584 12180 12590 12232
rect 14642 12180 14648 12232
rect 14700 12220 14706 12232
rect 15473 12223 15531 12229
rect 15473 12220 15485 12223
rect 14700 12192 15485 12220
rect 14700 12180 14706 12192
rect 15473 12189 15485 12192
rect 15519 12220 15531 12223
rect 16942 12220 16948 12232
rect 15519 12192 16948 12220
rect 15519 12189 15531 12192
rect 15473 12183 15531 12189
rect 16942 12180 16948 12192
rect 17000 12180 17006 12232
rect 5350 12112 5356 12164
rect 5408 12152 5414 12164
rect 10410 12161 10416 12164
rect 7254 12155 7312 12161
rect 7254 12152 7266 12155
rect 5408 12124 7266 12152
rect 5408 12112 5414 12124
rect 7254 12121 7266 12124
rect 7300 12121 7312 12155
rect 7254 12115 7312 12121
rect 10404 12115 10416 12161
rect 10468 12152 10474 12164
rect 15740 12155 15798 12161
rect 10468 12124 10504 12152
rect 10410 12112 10416 12115
rect 10468 12112 10474 12124
rect 15740 12121 15752 12155
rect 15786 12152 15798 12155
rect 17236 12152 17264 12396
rect 22833 12393 22845 12396
rect 22879 12393 22891 12427
rect 22833 12387 22891 12393
rect 20625 12359 20683 12365
rect 20625 12325 20637 12359
rect 20671 12356 20683 12359
rect 20898 12356 20904 12368
rect 20671 12328 20904 12356
rect 20671 12325 20683 12328
rect 20625 12319 20683 12325
rect 20898 12316 20904 12328
rect 20956 12316 20962 12368
rect 21465 12328 22508 12356
rect 20806 12248 20812 12300
rect 20864 12288 20870 12300
rect 21465 12288 21493 12328
rect 20864 12260 21493 12288
rect 20864 12248 20870 12260
rect 17313 12223 17371 12229
rect 17313 12189 17325 12223
rect 17359 12220 17371 12223
rect 17862 12220 17868 12232
rect 17359 12192 17868 12220
rect 17359 12189 17371 12192
rect 17313 12183 17371 12189
rect 15786 12124 17264 12152
rect 15786 12121 15798 12124
rect 15740 12115 15798 12121
rect 8386 12084 8392 12096
rect 8347 12056 8392 12084
rect 8386 12044 8392 12056
rect 8444 12044 8450 12096
rect 11422 12044 11428 12096
rect 11480 12084 11486 12096
rect 11517 12087 11575 12093
rect 11517 12084 11529 12087
rect 11480 12056 11529 12084
rect 11480 12044 11486 12056
rect 11517 12053 11529 12056
rect 11563 12053 11575 12087
rect 11517 12047 11575 12053
rect 13262 12044 13268 12096
rect 13320 12084 13326 12096
rect 13357 12087 13415 12093
rect 13357 12084 13369 12087
rect 13320 12056 13369 12084
rect 13320 12044 13326 12056
rect 13357 12053 13369 12056
rect 13403 12053 13415 12087
rect 16850 12084 16856 12096
rect 16811 12056 16856 12084
rect 13357 12047 13415 12053
rect 16850 12044 16856 12056
rect 16908 12044 16914 12096
rect 16942 12044 16948 12096
rect 17000 12084 17006 12096
rect 17328 12084 17356 12183
rect 17862 12180 17868 12192
rect 17920 12220 17926 12232
rect 18414 12220 18420 12232
rect 17920 12192 18420 12220
rect 17920 12180 17926 12192
rect 18414 12180 18420 12192
rect 18472 12220 18478 12232
rect 19245 12223 19303 12229
rect 19245 12220 19257 12223
rect 18472 12192 19257 12220
rect 18472 12180 18478 12192
rect 19245 12189 19257 12192
rect 19291 12189 19303 12223
rect 19245 12183 19303 12189
rect 19352 12192 21128 12220
rect 17580 12155 17638 12161
rect 17580 12121 17592 12155
rect 17626 12152 17638 12155
rect 19352 12152 19380 12192
rect 17626 12124 19380 12152
rect 19512 12155 19570 12161
rect 17626 12121 17638 12124
rect 17580 12115 17638 12121
rect 19512 12121 19524 12155
rect 19558 12152 19570 12155
rect 20530 12152 20536 12164
rect 19558 12124 20536 12152
rect 19558 12121 19570 12124
rect 19512 12115 19570 12121
rect 20530 12112 20536 12124
rect 20588 12112 20594 12164
rect 21100 12161 21128 12192
rect 21266 12180 21272 12232
rect 21324 12229 21330 12232
rect 21465 12229 21493 12260
rect 21324 12223 21373 12229
rect 21324 12189 21327 12223
rect 21361 12189 21373 12223
rect 21324 12183 21373 12189
rect 21450 12223 21508 12229
rect 21450 12189 21462 12223
rect 21496 12189 21508 12223
rect 21450 12183 21508 12189
rect 21550 12223 21608 12229
rect 21550 12189 21562 12223
rect 21596 12220 21608 12223
rect 21596 12192 21680 12220
rect 21596 12189 21608 12192
rect 21550 12183 21608 12189
rect 21324 12180 21330 12183
rect 21085 12155 21143 12161
rect 21085 12121 21097 12155
rect 21131 12121 21143 12155
rect 21085 12115 21143 12121
rect 21652 12096 21680 12192
rect 21726 12180 21732 12232
rect 21784 12220 21790 12232
rect 22370 12229 22376 12232
rect 22189 12223 22247 12229
rect 22189 12220 22201 12223
rect 21784 12192 22201 12220
rect 21784 12180 21790 12192
rect 22189 12189 22201 12192
rect 22235 12189 22247 12223
rect 22368 12220 22376 12229
rect 22331 12192 22376 12220
rect 22189 12183 22247 12189
rect 22368 12183 22376 12192
rect 22370 12180 22376 12183
rect 22428 12180 22434 12232
rect 22480 12229 22508 12328
rect 22468 12223 22526 12229
rect 22468 12189 22480 12223
rect 22514 12189 22526 12223
rect 22468 12183 22526 12189
rect 22557 12223 22615 12229
rect 22557 12189 22569 12223
rect 22603 12189 22615 12223
rect 22557 12183 22615 12189
rect 22572 12152 22600 12183
rect 22572 12124 22692 12152
rect 18690 12084 18696 12096
rect 17000 12056 17356 12084
rect 18651 12056 18696 12084
rect 17000 12044 17006 12056
rect 18690 12044 18696 12056
rect 18748 12044 18754 12096
rect 21634 12044 21640 12096
rect 21692 12044 21698 12096
rect 22554 12044 22560 12096
rect 22612 12084 22618 12096
rect 22664 12084 22692 12124
rect 22612 12056 22692 12084
rect 22612 12044 22618 12056
rect 1104 11994 68816 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 50294 11994
rect 50346 11942 50358 11994
rect 50410 11942 50422 11994
rect 50474 11942 50486 11994
rect 50538 11942 50550 11994
rect 50602 11942 68816 11994
rect 1104 11920 68816 11942
rect 5350 11880 5356 11892
rect 5311 11852 5356 11880
rect 5350 11840 5356 11852
rect 5408 11840 5414 11892
rect 5534 11840 5540 11892
rect 5592 11880 5598 11892
rect 5592 11852 8524 11880
rect 5592 11840 5598 11852
rect 8386 11812 8392 11824
rect 5092 11784 8392 11812
rect 4706 11744 4712 11756
rect 4667 11716 4712 11744
rect 4706 11704 4712 11716
rect 4764 11704 4770 11756
rect 5092 11753 5120 11784
rect 8386 11772 8392 11784
rect 8444 11772 8450 11824
rect 8496 11812 8524 11852
rect 8754 11840 8760 11892
rect 8812 11880 8818 11892
rect 9033 11883 9091 11889
rect 9033 11880 9045 11883
rect 8812 11852 9045 11880
rect 8812 11840 8818 11852
rect 9033 11849 9045 11852
rect 9079 11849 9091 11883
rect 12710 11880 12716 11892
rect 9033 11843 9091 11849
rect 9232 11852 12716 11880
rect 9232 11812 9260 11852
rect 12710 11840 12716 11852
rect 12768 11880 12774 11892
rect 16114 11880 16120 11892
rect 12768 11852 16120 11880
rect 12768 11840 12774 11852
rect 16114 11840 16120 11852
rect 16172 11840 16178 11892
rect 20530 11840 20536 11892
rect 20588 11880 20594 11892
rect 20625 11883 20683 11889
rect 20625 11880 20637 11883
rect 20588 11852 20637 11880
rect 20588 11840 20594 11852
rect 20625 11849 20637 11852
rect 20671 11849 20683 11883
rect 20625 11843 20683 11849
rect 8496 11784 9260 11812
rect 10134 11772 10140 11824
rect 10192 11821 10198 11824
rect 14918 11821 14924 11824
rect 10192 11812 10204 11821
rect 14912 11812 14924 11821
rect 10192 11784 10237 11812
rect 14879 11784 14924 11812
rect 10192 11775 10204 11784
rect 14912 11775 14924 11784
rect 10192 11772 10198 11775
rect 14918 11772 14924 11775
rect 14976 11772 14982 11824
rect 16850 11772 16856 11824
rect 16908 11812 16914 11824
rect 22554 11812 22560 11824
rect 16908 11784 22560 11812
rect 16908 11772 16914 11784
rect 22554 11772 22560 11784
rect 22612 11772 22618 11824
rect 4872 11747 4930 11753
rect 4872 11744 4884 11747
rect 4816 11716 4884 11744
rect 4816 11620 4844 11716
rect 4872 11713 4884 11716
rect 4918 11713 4930 11747
rect 4872 11707 4930 11713
rect 4972 11747 5030 11753
rect 4972 11713 4984 11747
rect 5018 11713 5030 11747
rect 4972 11707 5030 11713
rect 5077 11747 5135 11753
rect 5077 11713 5089 11747
rect 5123 11713 5135 11747
rect 5077 11707 5135 11713
rect 4987 11676 5015 11707
rect 6362 11704 6368 11756
rect 6420 11744 6426 11756
rect 7449 11747 7507 11753
rect 7449 11744 7461 11747
rect 6420 11716 7461 11744
rect 6420 11704 6426 11716
rect 7449 11713 7461 11716
rect 7495 11713 7507 11747
rect 7449 11707 7507 11713
rect 13538 11704 13544 11756
rect 13596 11744 13602 11756
rect 14642 11744 14648 11756
rect 13596 11716 14648 11744
rect 13596 11704 13602 11716
rect 14642 11704 14648 11716
rect 14700 11704 14706 11756
rect 18414 11744 18420 11756
rect 18375 11716 18420 11744
rect 18414 11704 18420 11716
rect 18472 11704 18478 11756
rect 18684 11747 18742 11753
rect 18684 11713 18696 11747
rect 18730 11744 18742 11747
rect 20438 11744 20444 11756
rect 18730 11716 20444 11744
rect 18730 11713 18742 11716
rect 18684 11707 18742 11713
rect 20438 11704 20444 11716
rect 20496 11704 20502 11756
rect 20898 11744 20904 11756
rect 20859 11716 20904 11744
rect 20898 11704 20904 11716
rect 20956 11704 20962 11756
rect 20993 11747 21051 11753
rect 20993 11713 21005 11747
rect 21039 11713 21051 11747
rect 20993 11707 21051 11713
rect 6178 11676 6184 11688
rect 4987 11648 6184 11676
rect 6178 11636 6184 11648
rect 6236 11636 6242 11688
rect 7190 11676 7196 11688
rect 7151 11648 7196 11676
rect 7190 11636 7196 11648
rect 7248 11636 7254 11688
rect 10413 11679 10471 11685
rect 10413 11645 10425 11679
rect 10459 11676 10471 11679
rect 11698 11676 11704 11688
rect 10459 11648 11704 11676
rect 10459 11645 10471 11648
rect 10413 11639 10471 11645
rect 4798 11568 4804 11620
rect 4856 11568 4862 11620
rect 8570 11540 8576 11552
rect 8531 11512 8576 11540
rect 8570 11500 8576 11512
rect 8628 11500 8634 11552
rect 9490 11500 9496 11552
rect 9548 11540 9554 11552
rect 10428 11540 10456 11639
rect 11698 11636 11704 11648
rect 11756 11636 11762 11688
rect 20806 11636 20812 11688
rect 20864 11676 20870 11688
rect 21008 11676 21036 11707
rect 21082 11704 21088 11756
rect 21140 11744 21146 11756
rect 21140 11716 21185 11744
rect 21140 11704 21146 11716
rect 21266 11704 21272 11756
rect 21324 11744 21330 11756
rect 21726 11744 21732 11756
rect 21324 11716 21732 11744
rect 21324 11704 21330 11716
rect 21726 11704 21732 11716
rect 21784 11704 21790 11756
rect 20864 11648 21036 11676
rect 20864 11636 20870 11648
rect 9548 11512 10456 11540
rect 9548 11500 9554 11512
rect 15286 11500 15292 11552
rect 15344 11540 15350 11552
rect 16022 11540 16028 11552
rect 15344 11512 16028 11540
rect 15344 11500 15350 11512
rect 16022 11500 16028 11512
rect 16080 11500 16086 11552
rect 19794 11540 19800 11552
rect 19755 11512 19800 11540
rect 19794 11500 19800 11512
rect 19852 11500 19858 11552
rect 1104 11450 68816 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 65654 11450
rect 65706 11398 65718 11450
rect 65770 11398 65782 11450
rect 65834 11398 65846 11450
rect 65898 11398 65910 11450
rect 65962 11398 68816 11450
rect 1104 11376 68816 11398
rect 4430 11336 4436 11348
rect 4391 11308 4436 11336
rect 4430 11296 4436 11308
rect 4488 11296 4494 11348
rect 4614 11336 4620 11348
rect 4575 11308 4620 11336
rect 4614 11296 4620 11308
rect 4672 11296 4678 11348
rect 6362 11336 6368 11348
rect 6323 11308 6368 11336
rect 6362 11296 6368 11308
rect 6420 11296 6426 11348
rect 9950 11296 9956 11348
rect 10008 11336 10014 11348
rect 10321 11339 10379 11345
rect 10321 11336 10333 11339
rect 10008 11308 10333 11336
rect 10008 11296 10014 11308
rect 10321 11305 10333 11308
rect 10367 11336 10379 11339
rect 10502 11336 10508 11348
rect 10367 11308 10508 11336
rect 10367 11305 10379 11308
rect 10321 11299 10379 11305
rect 10502 11296 10508 11308
rect 10560 11296 10566 11348
rect 12158 11336 12164 11348
rect 12119 11308 12164 11336
rect 12158 11296 12164 11308
rect 12216 11296 12222 11348
rect 22094 11296 22100 11348
rect 22152 11336 22158 11348
rect 22373 11339 22431 11345
rect 22373 11336 22385 11339
rect 22152 11308 22385 11336
rect 22152 11296 22158 11308
rect 22373 11305 22385 11308
rect 22419 11305 22431 11339
rect 23198 11336 23204 11348
rect 22373 11299 22431 11305
rect 22480 11308 23204 11336
rect 4448 11240 9674 11268
rect 4338 11132 4344 11144
rect 4299 11104 4344 11132
rect 4338 11092 4344 11104
rect 4396 11092 4402 11144
rect 4448 11141 4476 11240
rect 5442 11160 5448 11212
rect 5500 11200 5506 11212
rect 6178 11200 6184 11212
rect 5500 11172 5856 11200
rect 5500 11160 5506 11172
rect 4433 11135 4491 11141
rect 4433 11101 4445 11135
rect 4479 11101 4491 11135
rect 4433 11095 4491 11101
rect 4706 11092 4712 11144
rect 4764 11132 4770 11144
rect 5718 11132 5724 11144
rect 4764 11104 5724 11132
rect 4764 11092 4770 11104
rect 5718 11092 5724 11104
rect 5776 11092 5782 11144
rect 5828 11132 5856 11172
rect 6012 11172 6184 11200
rect 6012 11141 6040 11172
rect 6178 11160 6184 11172
rect 6236 11160 6242 11212
rect 5900 11135 5958 11141
rect 5900 11132 5912 11135
rect 5828 11104 5912 11132
rect 5900 11101 5912 11104
rect 5946 11101 5958 11135
rect 5900 11095 5958 11101
rect 5997 11135 6055 11141
rect 5997 11101 6009 11135
rect 6043 11101 6055 11135
rect 5997 11095 6055 11101
rect 6089 11135 6147 11141
rect 6089 11101 6101 11135
rect 6135 11126 6147 11135
rect 8570 11132 8576 11144
rect 6288 11126 8576 11132
rect 6135 11104 8576 11126
rect 6135 11101 6316 11104
rect 6089 11098 6316 11101
rect 6089 11095 6147 11098
rect 8570 11092 8576 11104
rect 8628 11092 8634 11144
rect 4154 11064 4160 11076
rect 4115 11036 4160 11064
rect 4154 11024 4160 11036
rect 4212 11024 4218 11076
rect 9646 11064 9674 11240
rect 19794 11228 19800 11280
rect 19852 11268 19858 11280
rect 20622 11268 20628 11280
rect 19852 11240 20628 11268
rect 19852 11228 19858 11240
rect 20622 11228 20628 11240
rect 20680 11268 20686 11280
rect 22480 11268 22508 11308
rect 23198 11296 23204 11308
rect 23256 11296 23262 11348
rect 20680 11240 22508 11268
rect 22741 11271 22799 11277
rect 20680 11228 20686 11240
rect 22741 11237 22753 11271
rect 22787 11268 22799 11271
rect 23106 11268 23112 11280
rect 22787 11240 23112 11268
rect 22787 11237 22799 11240
rect 22741 11231 22799 11237
rect 23106 11228 23112 11240
rect 23164 11228 23170 11280
rect 23842 11268 23848 11280
rect 23216 11240 23848 11268
rect 11698 11200 11704 11212
rect 11659 11172 11704 11200
rect 11698 11160 11704 11172
rect 11756 11160 11762 11212
rect 13538 11200 13544 11212
rect 13499 11172 13544 11200
rect 13538 11160 13544 11172
rect 13596 11160 13602 11212
rect 18690 11160 18696 11212
rect 18748 11200 18754 11212
rect 21358 11200 21364 11212
rect 18748 11172 21364 11200
rect 18748 11160 18754 11172
rect 21358 11160 21364 11172
rect 21416 11200 21422 11212
rect 22465 11203 22523 11209
rect 22465 11200 22477 11203
rect 21416 11172 22477 11200
rect 21416 11160 21422 11172
rect 22465 11169 22477 11172
rect 22511 11200 22523 11203
rect 23216 11200 23244 11240
rect 23842 11228 23848 11240
rect 23900 11228 23906 11280
rect 22511 11172 23244 11200
rect 22511 11169 22523 11172
rect 22465 11163 22523 11169
rect 11445 11135 11503 11141
rect 11445 11101 11457 11135
rect 11491 11132 11503 11135
rect 11606 11132 11612 11144
rect 11491 11104 11612 11132
rect 11491 11101 11503 11104
rect 11445 11095 11503 11101
rect 11606 11092 11612 11104
rect 11664 11092 11670 11144
rect 13285 11135 13343 11141
rect 13285 11101 13297 11135
rect 13331 11132 13343 11135
rect 13722 11132 13728 11144
rect 13331 11104 13728 11132
rect 13331 11101 13343 11104
rect 13285 11095 13343 11101
rect 13722 11092 13728 11104
rect 13780 11092 13786 11144
rect 22370 11132 22376 11144
rect 22331 11104 22376 11132
rect 22370 11092 22376 11104
rect 22428 11092 22434 11144
rect 23014 11092 23020 11144
rect 23072 11132 23078 11144
rect 23385 11135 23443 11141
rect 23385 11132 23397 11135
rect 23072 11104 23397 11132
rect 23072 11092 23078 11104
rect 23385 11101 23397 11104
rect 23431 11101 23443 11135
rect 23385 11095 23443 11101
rect 23477 11135 23535 11141
rect 23477 11101 23489 11135
rect 23523 11132 23535 11135
rect 23566 11132 23572 11144
rect 23523 11104 23572 11132
rect 23523 11101 23535 11104
rect 23477 11095 23535 11101
rect 23566 11092 23572 11104
rect 23624 11092 23630 11144
rect 10686 11064 10692 11076
rect 9646 11036 10692 11064
rect 10686 11024 10692 11036
rect 10744 11024 10750 11076
rect 16022 11024 16028 11076
rect 16080 11064 16086 11076
rect 23201 11067 23259 11073
rect 23201 11064 23213 11067
rect 16080 11036 23213 11064
rect 16080 11024 16086 11036
rect 23201 11033 23213 11036
rect 23247 11064 23259 11067
rect 24486 11064 24492 11076
rect 23247 11036 24492 11064
rect 23247 11033 23259 11036
rect 23201 11027 23259 11033
rect 24486 11024 24492 11036
rect 24544 11024 24550 11076
rect 23658 10996 23664 11008
rect 23619 10968 23664 10996
rect 23658 10956 23664 10968
rect 23716 10956 23722 11008
rect 1104 10906 68816 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 50294 10906
rect 50346 10854 50358 10906
rect 50410 10854 50422 10906
rect 50474 10854 50486 10906
rect 50538 10854 50550 10906
rect 50602 10854 68816 10906
rect 1104 10832 68816 10854
rect 4617 10795 4675 10801
rect 4617 10761 4629 10795
rect 4663 10792 4675 10795
rect 4798 10792 4804 10804
rect 4663 10764 4804 10792
rect 4663 10761 4675 10764
rect 4617 10755 4675 10761
rect 4798 10752 4804 10764
rect 4856 10752 4862 10804
rect 5813 10795 5871 10801
rect 5813 10761 5825 10795
rect 5859 10792 5871 10795
rect 5859 10764 6592 10792
rect 5859 10761 5871 10764
rect 5813 10755 5871 10761
rect 4154 10724 4160 10736
rect 4067 10696 4160 10724
rect 4154 10684 4160 10696
rect 4212 10724 4218 10736
rect 5994 10724 6000 10736
rect 4212 10696 5028 10724
rect 4212 10684 4218 10696
rect 5000 10668 5028 10696
rect 5644 10696 6000 10724
rect 4433 10659 4491 10665
rect 4433 10625 4445 10659
rect 4479 10656 4491 10659
rect 4706 10656 4712 10668
rect 4479 10628 4712 10656
rect 4479 10625 4491 10628
rect 4433 10619 4491 10625
rect 4706 10616 4712 10628
rect 4764 10616 4770 10668
rect 4982 10616 4988 10668
rect 5040 10656 5046 10668
rect 5644 10665 5672 10696
rect 5994 10684 6000 10696
rect 6052 10684 6058 10736
rect 6564 10671 6592 10764
rect 10594 10752 10600 10804
rect 10652 10792 10658 10804
rect 10965 10795 11023 10801
rect 10965 10792 10977 10795
rect 10652 10764 10977 10792
rect 10652 10752 10658 10764
rect 10965 10761 10977 10764
rect 11011 10792 11023 10795
rect 14369 10795 14427 10801
rect 11011 10764 12434 10792
rect 11011 10761 11023 10764
rect 10965 10755 11023 10761
rect 7190 10684 7196 10736
rect 7248 10724 7254 10736
rect 9858 10733 9864 10736
rect 9852 10724 9864 10733
rect 7248 10696 9536 10724
rect 9819 10696 9864 10724
rect 7248 10684 7254 10696
rect 5353 10659 5411 10665
rect 5353 10656 5365 10659
rect 5040 10628 5365 10656
rect 5040 10616 5046 10628
rect 5353 10625 5365 10628
rect 5399 10625 5411 10659
rect 5353 10619 5411 10625
rect 5629 10659 5687 10665
rect 5629 10625 5641 10659
rect 5675 10625 5687 10659
rect 5629 10619 5687 10625
rect 5718 10616 5724 10668
rect 5776 10656 5782 10668
rect 6549 10665 6607 10671
rect 7760 10665 7788 10696
rect 9508 10668 9536 10696
rect 9852 10687 9864 10696
rect 9858 10684 9864 10687
rect 9916 10684 9922 10736
rect 6365 10659 6423 10665
rect 6365 10656 6377 10659
rect 5776 10628 6377 10656
rect 5776 10616 5782 10628
rect 6365 10625 6377 10628
rect 6411 10625 6423 10659
rect 6549 10631 6561 10665
rect 6595 10631 6607 10665
rect 6549 10625 6607 10631
rect 6641 10659 6699 10665
rect 6641 10625 6653 10659
rect 6687 10625 6699 10659
rect 6365 10619 6423 10625
rect 6641 10619 6699 10625
rect 6733 10659 6791 10665
rect 6733 10625 6745 10659
rect 6779 10625 6791 10659
rect 6733 10619 6791 10625
rect 7745 10659 7803 10665
rect 7745 10625 7757 10659
rect 7791 10625 7803 10659
rect 8001 10659 8059 10665
rect 8001 10656 8013 10659
rect 7745 10619 7803 10625
rect 7852 10628 8013 10656
rect 4338 10588 4344 10600
rect 4251 10560 4344 10588
rect 4338 10548 4344 10560
rect 4396 10588 4402 10600
rect 5166 10588 5172 10600
rect 4396 10560 5172 10588
rect 4396 10548 4402 10560
rect 5166 10548 5172 10560
rect 5224 10588 5230 10600
rect 5445 10591 5503 10597
rect 5445 10588 5457 10591
rect 5224 10560 5457 10588
rect 5224 10548 5230 10560
rect 5445 10557 5457 10560
rect 5491 10557 5503 10591
rect 5445 10551 5503 10557
rect 6178 10548 6184 10600
rect 6236 10588 6242 10600
rect 6656 10588 6684 10619
rect 6236 10560 6684 10588
rect 6236 10548 6242 10560
rect 4430 10452 4436 10464
rect 4343 10424 4436 10452
rect 4430 10412 4436 10424
rect 4488 10452 4494 10464
rect 5258 10452 5264 10464
rect 4488 10424 5264 10452
rect 4488 10412 4494 10424
rect 5258 10412 5264 10424
rect 5316 10452 5322 10464
rect 5445 10455 5503 10461
rect 5445 10452 5457 10455
rect 5316 10424 5457 10452
rect 5316 10412 5322 10424
rect 5445 10421 5457 10424
rect 5491 10452 5503 10455
rect 6362 10452 6368 10464
rect 5491 10424 6368 10452
rect 5491 10421 5503 10424
rect 5445 10415 5503 10421
rect 6362 10412 6368 10424
rect 6420 10412 6426 10464
rect 6748 10452 6776 10619
rect 7009 10591 7067 10597
rect 7009 10557 7021 10591
rect 7055 10588 7067 10591
rect 7852 10588 7880 10628
rect 8001 10625 8013 10628
rect 8047 10625 8059 10659
rect 8001 10619 8059 10625
rect 9490 10616 9496 10668
rect 9548 10656 9554 10668
rect 9585 10659 9643 10665
rect 9585 10656 9597 10659
rect 9548 10628 9597 10656
rect 9548 10616 9554 10628
rect 9585 10625 9597 10628
rect 9631 10625 9643 10659
rect 9585 10619 9643 10625
rect 7055 10560 7880 10588
rect 7055 10557 7067 10560
rect 7009 10551 7067 10557
rect 9125 10455 9183 10461
rect 9125 10452 9137 10455
rect 6748 10424 9137 10452
rect 9125 10421 9137 10424
rect 9171 10452 9183 10455
rect 9214 10452 9220 10464
rect 9171 10424 9220 10452
rect 9171 10421 9183 10424
rect 9125 10415 9183 10421
rect 9214 10412 9220 10424
rect 9272 10412 9278 10464
rect 12406 10452 12434 10764
rect 14369 10761 14381 10795
rect 14415 10792 14427 10795
rect 20438 10792 20444 10804
rect 14415 10764 16988 10792
rect 20399 10764 20444 10792
rect 14415 10761 14427 10764
rect 14369 10755 14427 10761
rect 13538 10724 13544 10736
rect 13004 10696 13544 10724
rect 13004 10665 13032 10696
rect 13538 10684 13544 10696
rect 13596 10684 13602 10736
rect 16669 10727 16727 10733
rect 16669 10693 16681 10727
rect 16715 10693 16727 10727
rect 16669 10687 16727 10693
rect 16960 10724 16988 10764
rect 20438 10752 20444 10764
rect 20496 10752 20502 10804
rect 20806 10792 20812 10804
rect 20732 10764 20812 10792
rect 19150 10724 19156 10736
rect 16960 10696 19156 10724
rect 12989 10659 13047 10665
rect 12989 10625 13001 10659
rect 13035 10625 13047 10659
rect 12989 10619 13047 10625
rect 13256 10659 13314 10665
rect 13256 10625 13268 10659
rect 13302 10656 13314 10659
rect 16684 10656 16712 10687
rect 16960 10665 16988 10696
rect 19150 10684 19156 10696
rect 19208 10684 19214 10736
rect 20732 10724 20760 10764
rect 20806 10752 20812 10764
rect 20864 10752 20870 10804
rect 20898 10752 20904 10804
rect 20956 10792 20962 10804
rect 20956 10764 22048 10792
rect 20956 10752 20962 10764
rect 20732 10696 20852 10724
rect 13302 10628 16712 10656
rect 16925 10659 16988 10665
rect 13302 10625 13314 10628
rect 13256 10619 13314 10625
rect 16925 10625 16937 10659
rect 16971 10628 16988 10659
rect 17034 10659 17092 10665
rect 16971 10625 16983 10628
rect 16925 10619 16983 10625
rect 17034 10625 17046 10659
rect 17080 10625 17092 10659
rect 17034 10619 17092 10625
rect 17129 10662 17187 10668
rect 17129 10628 17141 10662
rect 17175 10628 17187 10662
rect 17310 10656 17316 10668
rect 17271 10628 17316 10656
rect 17129 10622 17187 10628
rect 15654 10480 15660 10532
rect 15712 10520 15718 10532
rect 16942 10520 16948 10532
rect 15712 10492 16948 10520
rect 15712 10480 15718 10492
rect 16942 10480 16948 10492
rect 17000 10520 17006 10532
rect 17052 10520 17080 10619
rect 17144 10588 17172 10622
rect 17310 10616 17316 10628
rect 17368 10616 17374 10668
rect 17862 10616 17868 10668
rect 17920 10656 17926 10668
rect 18141 10659 18199 10665
rect 18141 10656 18153 10659
rect 17920 10628 18153 10656
rect 17920 10616 17926 10628
rect 18141 10625 18153 10628
rect 18187 10625 18199 10659
rect 18141 10619 18199 10625
rect 18408 10659 18466 10665
rect 18408 10625 18420 10659
rect 18454 10656 18466 10659
rect 20162 10656 20168 10668
rect 18454 10628 20168 10656
rect 18454 10625 18466 10628
rect 18408 10619 18466 10625
rect 20162 10616 20168 10628
rect 20220 10616 20226 10668
rect 20622 10616 20628 10668
rect 20680 10665 20686 10668
rect 20824 10665 20852 10696
rect 20680 10659 20729 10665
rect 20680 10625 20683 10659
rect 20717 10625 20729 10659
rect 20680 10619 20729 10625
rect 20809 10659 20867 10665
rect 20809 10625 20821 10659
rect 20855 10625 20867 10659
rect 20809 10619 20867 10625
rect 20898 10619 20904 10671
rect 20956 10659 20962 10671
rect 21085 10659 21143 10665
rect 20956 10631 21001 10659
rect 20956 10619 20962 10631
rect 21085 10625 21097 10659
rect 21131 10656 21143 10659
rect 21266 10656 21272 10668
rect 21131 10628 21272 10656
rect 21131 10625 21143 10628
rect 21085 10619 21143 10625
rect 20680 10616 20686 10619
rect 17770 10588 17776 10600
rect 17144 10560 17776 10588
rect 17770 10548 17776 10560
rect 17828 10548 17834 10600
rect 20990 10548 20996 10600
rect 21048 10588 21054 10600
rect 21100 10588 21128 10619
rect 21266 10616 21272 10628
rect 21324 10616 21330 10668
rect 22020 10665 22048 10764
rect 23658 10684 23664 10736
rect 23716 10724 23722 10736
rect 24213 10727 24271 10733
rect 24213 10724 24225 10727
rect 23716 10696 24225 10724
rect 23716 10684 23722 10696
rect 24213 10693 24225 10696
rect 24259 10693 24271 10727
rect 24213 10687 24271 10693
rect 22005 10659 22063 10665
rect 22005 10625 22017 10659
rect 22051 10625 22063 10659
rect 22005 10619 22063 10625
rect 22189 10659 22247 10665
rect 22189 10625 22201 10659
rect 22235 10656 22247 10659
rect 22370 10656 22376 10668
rect 22235 10628 22376 10656
rect 22235 10625 22247 10628
rect 22189 10619 22247 10625
rect 22370 10616 22376 10628
rect 22428 10656 22434 10668
rect 22646 10656 22652 10668
rect 22428 10628 22652 10656
rect 22428 10616 22434 10628
rect 22646 10616 22652 10628
rect 22704 10656 22710 10668
rect 23017 10659 23075 10665
rect 23017 10656 23029 10659
rect 22704 10628 23029 10656
rect 22704 10616 22710 10628
rect 23017 10625 23029 10628
rect 23063 10625 23075 10659
rect 23842 10656 23848 10668
rect 23803 10628 23848 10656
rect 23017 10619 23075 10625
rect 23842 10616 23848 10628
rect 23900 10616 23906 10668
rect 21048 10560 21128 10588
rect 21048 10548 21054 10560
rect 22554 10548 22560 10600
rect 22612 10588 22618 10600
rect 23109 10591 23167 10597
rect 23109 10588 23121 10591
rect 22612 10560 23121 10588
rect 22612 10548 22618 10560
rect 23109 10557 23121 10560
rect 23155 10588 23167 10591
rect 23937 10591 23995 10597
rect 23937 10588 23949 10591
rect 23155 10560 23949 10588
rect 23155 10557 23167 10560
rect 23109 10551 23167 10557
rect 23937 10557 23949 10560
rect 23983 10557 23995 10591
rect 23937 10551 23995 10557
rect 17000 10492 17080 10520
rect 17000 10480 17006 10492
rect 20530 10480 20536 10532
rect 20588 10520 20594 10532
rect 24029 10523 24087 10529
rect 24029 10520 24041 10523
rect 20588 10492 24041 10520
rect 20588 10480 20594 10492
rect 24029 10489 24041 10492
rect 24075 10489 24087 10523
rect 24029 10483 24087 10489
rect 12986 10452 12992 10464
rect 12406 10424 12992 10452
rect 12986 10412 12992 10424
rect 13044 10412 13050 10464
rect 19521 10455 19579 10461
rect 19521 10421 19533 10455
rect 19567 10452 19579 10455
rect 20438 10452 20444 10464
rect 19567 10424 20444 10452
rect 19567 10421 19579 10424
rect 19521 10415 19579 10421
rect 20438 10412 20444 10424
rect 20496 10412 20502 10464
rect 20714 10412 20720 10464
rect 20772 10452 20778 10464
rect 21821 10455 21879 10461
rect 21821 10452 21833 10455
rect 20772 10424 21833 10452
rect 20772 10412 20778 10424
rect 21821 10421 21833 10424
rect 21867 10421 21879 10455
rect 22094 10452 22100 10464
rect 22055 10424 22100 10452
rect 21821 10415 21879 10421
rect 22094 10412 22100 10424
rect 22152 10452 22158 10464
rect 23017 10455 23075 10461
rect 23017 10452 23029 10455
rect 22152 10424 23029 10452
rect 22152 10412 22158 10424
rect 23017 10421 23029 10424
rect 23063 10421 23075 10455
rect 23382 10452 23388 10464
rect 23343 10424 23388 10452
rect 23017 10415 23075 10421
rect 23382 10412 23388 10424
rect 23440 10412 23446 10464
rect 24213 10455 24271 10461
rect 24213 10421 24225 10455
rect 24259 10452 24271 10455
rect 26970 10452 26976 10464
rect 24259 10424 26976 10452
rect 24259 10421 24271 10424
rect 24213 10415 24271 10421
rect 26970 10412 26976 10424
rect 27028 10412 27034 10464
rect 1104 10362 68816 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 65654 10362
rect 65706 10310 65718 10362
rect 65770 10310 65782 10362
rect 65834 10310 65846 10362
rect 65898 10310 65910 10362
rect 65962 10310 68816 10362
rect 1104 10288 68816 10310
rect 4341 10251 4399 10257
rect 4341 10217 4353 10251
rect 4387 10248 4399 10251
rect 5258 10248 5264 10260
rect 4387 10220 5264 10248
rect 4387 10217 4399 10220
rect 4341 10211 4399 10217
rect 5258 10208 5264 10220
rect 5316 10208 5322 10260
rect 5442 10248 5448 10260
rect 5403 10220 5448 10248
rect 5442 10208 5448 10220
rect 5500 10208 5506 10260
rect 8110 10248 8116 10260
rect 6932 10220 8116 10248
rect 5442 10112 5448 10124
rect 4172 10084 5448 10112
rect 4172 10053 4200 10084
rect 5442 10072 5448 10084
rect 5500 10072 5506 10124
rect 3237 10047 3295 10053
rect 3237 10013 3249 10047
rect 3283 10044 3295 10047
rect 4157 10047 4215 10053
rect 4157 10044 4169 10047
rect 3283 10016 4169 10044
rect 3283 10013 3295 10016
rect 3237 10007 3295 10013
rect 4157 10013 4169 10016
rect 4203 10013 4215 10047
rect 5166 10044 5172 10056
rect 5127 10016 5172 10044
rect 4157 10007 4215 10013
rect 5166 10004 5172 10016
rect 5224 10004 5230 10056
rect 5258 10004 5264 10056
rect 5316 10044 5322 10056
rect 5316 10016 5361 10044
rect 5316 10004 5322 10016
rect 5718 10004 5724 10056
rect 5776 10044 5782 10056
rect 5905 10047 5963 10053
rect 6181 10047 6239 10053
rect 5905 10044 5917 10047
rect 5776 10016 5917 10044
rect 5776 10004 5782 10016
rect 5905 10013 5917 10016
rect 5951 10013 5963 10047
rect 6068 10041 6126 10047
rect 6068 10038 6080 10041
rect 5905 10007 5963 10013
rect 6012 10010 6080 10038
rect 4982 9976 4988 9988
rect 4943 9948 4988 9976
rect 4982 9936 4988 9948
rect 5040 9936 5046 9988
rect 6012 9908 6040 10010
rect 6068 10007 6080 10010
rect 6114 10007 6126 10041
rect 6181 10013 6193 10047
rect 6227 10013 6239 10047
rect 6181 10007 6239 10013
rect 6319 10047 6377 10053
rect 6319 10013 6331 10047
rect 6365 10044 6377 10047
rect 6932 10044 6960 10220
rect 8110 10208 8116 10220
rect 8168 10248 8174 10260
rect 8389 10251 8447 10257
rect 8389 10248 8401 10251
rect 8168 10220 8401 10248
rect 8168 10208 8174 10220
rect 8389 10217 8401 10220
rect 8435 10217 8447 10251
rect 8389 10211 8447 10217
rect 16482 10208 16488 10260
rect 16540 10248 16546 10260
rect 16761 10251 16819 10257
rect 16761 10248 16773 10251
rect 16540 10220 16773 10248
rect 16540 10208 16546 10220
rect 16761 10217 16773 10220
rect 16807 10217 16819 10251
rect 20162 10248 20168 10260
rect 20123 10220 20168 10248
rect 16761 10211 16819 10217
rect 20162 10208 20168 10220
rect 20220 10208 20226 10260
rect 22094 10208 22100 10260
rect 22152 10248 22158 10260
rect 22649 10251 22707 10257
rect 22649 10248 22661 10251
rect 22152 10220 22661 10248
rect 22152 10208 22158 10220
rect 22649 10217 22661 10220
rect 22695 10248 22707 10251
rect 23477 10251 23535 10257
rect 23477 10248 23489 10251
rect 22695 10220 23489 10248
rect 22695 10217 22707 10220
rect 22649 10211 22707 10217
rect 23477 10217 23489 10220
rect 23523 10217 23535 10251
rect 23477 10211 23535 10217
rect 18693 10183 18751 10189
rect 18693 10149 18705 10183
rect 18739 10180 18751 10183
rect 22554 10180 22560 10192
rect 18739 10152 22560 10180
rect 18739 10149 18751 10152
rect 18693 10143 18751 10149
rect 22554 10140 22560 10152
rect 22612 10140 22618 10192
rect 23566 10180 23572 10192
rect 22756 10152 23572 10180
rect 22756 10121 22784 10152
rect 23566 10140 23572 10152
rect 23624 10140 23630 10192
rect 22741 10115 22799 10121
rect 22741 10112 22753 10115
rect 20456 10084 22753 10112
rect 20456 10056 20484 10084
rect 22741 10081 22753 10084
rect 22787 10081 22799 10115
rect 22741 10075 22799 10081
rect 23198 10072 23204 10124
rect 23256 10112 23262 10124
rect 23256 10084 23612 10112
rect 23256 10072 23262 10084
rect 6365 10016 6960 10044
rect 7009 10047 7067 10053
rect 6365 10013 6377 10016
rect 6319 10007 6377 10013
rect 7009 10013 7021 10047
rect 7055 10044 7067 10047
rect 7098 10044 7104 10056
rect 7055 10016 7104 10044
rect 7055 10013 7067 10016
rect 7009 10007 7067 10013
rect 6068 10001 6126 10007
rect 6183 9920 6211 10007
rect 7098 10004 7104 10016
rect 7156 10004 7162 10056
rect 15381 10047 15439 10053
rect 15381 10013 15393 10047
rect 15427 10044 15439 10047
rect 16574 10044 16580 10056
rect 15427 10016 16580 10044
rect 15427 10013 15439 10016
rect 15381 10007 15439 10013
rect 16574 10004 16580 10016
rect 16632 10044 16638 10056
rect 17313 10047 17371 10053
rect 17313 10044 17325 10047
rect 16632 10016 17325 10044
rect 16632 10004 16638 10016
rect 17313 10013 17325 10016
rect 17359 10044 17371 10047
rect 17862 10044 17868 10056
rect 17359 10016 17868 10044
rect 17359 10013 17371 10016
rect 17313 10007 17371 10013
rect 17862 10004 17868 10016
rect 17920 10004 17926 10056
rect 20438 10044 20444 10056
rect 20399 10016 20444 10044
rect 20438 10004 20444 10016
rect 20496 10004 20502 10056
rect 20533 10047 20591 10053
rect 20533 10013 20545 10047
rect 20579 10013 20591 10047
rect 20533 10007 20591 10013
rect 6549 9979 6607 9985
rect 6549 9945 6561 9979
rect 6595 9976 6607 9979
rect 7254 9979 7312 9985
rect 7254 9976 7266 9979
rect 6595 9948 7266 9976
rect 6595 9945 6607 9948
rect 6549 9939 6607 9945
rect 7254 9945 7266 9948
rect 7300 9945 7312 9979
rect 7254 9939 7312 9945
rect 15648 9979 15706 9985
rect 15648 9945 15660 9979
rect 15694 9976 15706 9979
rect 16206 9976 16212 9988
rect 15694 9948 16212 9976
rect 15694 9945 15706 9948
rect 15648 9939 15706 9945
rect 16206 9936 16212 9948
rect 16264 9936 16270 9988
rect 17580 9979 17638 9985
rect 17580 9945 17592 9979
rect 17626 9976 17638 9979
rect 19242 9976 19248 9988
rect 17626 9948 19248 9976
rect 17626 9945 17638 9948
rect 17580 9939 17638 9945
rect 19242 9936 19248 9948
rect 19300 9936 19306 9988
rect 6086 9908 6092 9920
rect 6012 9880 6092 9908
rect 6086 9868 6092 9880
rect 6144 9868 6150 9920
rect 6178 9868 6184 9920
rect 6236 9868 6242 9920
rect 11149 9911 11207 9917
rect 11149 9877 11161 9911
rect 11195 9908 11207 9911
rect 11238 9908 11244 9920
rect 11195 9880 11244 9908
rect 11195 9877 11207 9880
rect 11149 9871 11207 9877
rect 11238 9868 11244 9880
rect 11296 9868 11302 9920
rect 11977 9911 12035 9917
rect 11977 9877 11989 9911
rect 12023 9908 12035 9911
rect 12434 9908 12440 9920
rect 12023 9880 12440 9908
rect 12023 9877 12035 9880
rect 11977 9871 12035 9877
rect 12434 9868 12440 9880
rect 12492 9868 12498 9920
rect 13078 9908 13084 9920
rect 13039 9880 13084 9908
rect 13078 9868 13084 9880
rect 13136 9868 13142 9920
rect 14182 9908 14188 9920
rect 14143 9880 14188 9908
rect 14182 9868 14188 9880
rect 14240 9868 14246 9920
rect 14734 9908 14740 9920
rect 14695 9880 14740 9908
rect 14734 9868 14740 9880
rect 14792 9868 14798 9920
rect 15562 9868 15568 9920
rect 15620 9908 15626 9920
rect 20548 9908 20576 10007
rect 20622 10004 20628 10056
rect 20680 10044 20686 10056
rect 20809 10047 20867 10053
rect 20680 10016 20725 10044
rect 20680 10004 20686 10016
rect 20809 10013 20821 10047
rect 20855 10044 20867 10047
rect 20990 10044 20996 10056
rect 20855 10016 20996 10044
rect 20855 10013 20867 10016
rect 20809 10007 20867 10013
rect 20990 10004 20996 10016
rect 21048 10004 21054 10056
rect 22646 10044 22652 10056
rect 22607 10016 22652 10044
rect 22646 10004 22652 10016
rect 22704 10004 22710 10056
rect 23584 10053 23612 10084
rect 23477 10047 23535 10053
rect 23477 10013 23489 10047
rect 23523 10013 23535 10047
rect 23477 10007 23535 10013
rect 23569 10047 23627 10053
rect 23569 10013 23581 10047
rect 23615 10013 23627 10047
rect 23569 10007 23627 10013
rect 22664 9976 22692 10004
rect 23492 9976 23520 10007
rect 22664 9948 23520 9976
rect 20806 9908 20812 9920
rect 15620 9880 20812 9908
rect 15620 9868 15626 9880
rect 20806 9868 20812 9880
rect 20864 9868 20870 9920
rect 21726 9908 21732 9920
rect 21687 9880 21732 9908
rect 21726 9868 21732 9880
rect 21784 9868 21790 9920
rect 23017 9911 23075 9917
rect 23017 9877 23029 9911
rect 23063 9908 23075 9911
rect 23198 9908 23204 9920
rect 23063 9880 23204 9908
rect 23063 9877 23075 9880
rect 23017 9871 23075 9877
rect 23198 9868 23204 9880
rect 23256 9868 23262 9920
rect 23290 9868 23296 9920
rect 23348 9908 23354 9920
rect 23845 9911 23903 9917
rect 23845 9908 23857 9911
rect 23348 9880 23857 9908
rect 23348 9868 23354 9880
rect 23845 9877 23857 9880
rect 23891 9877 23903 9911
rect 23845 9871 23903 9877
rect 1104 9818 68816 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 50294 9818
rect 50346 9766 50358 9818
rect 50410 9766 50422 9818
rect 50474 9766 50486 9818
rect 50538 9766 50550 9818
rect 50602 9766 68816 9818
rect 1104 9744 68816 9766
rect 3513 9707 3571 9713
rect 3513 9673 3525 9707
rect 3559 9673 3571 9707
rect 3513 9667 3571 9673
rect 3528 9636 3556 9667
rect 6086 9664 6092 9716
rect 6144 9704 6150 9716
rect 6825 9707 6883 9713
rect 6825 9704 6837 9707
rect 6144 9676 6837 9704
rect 6144 9664 6150 9676
rect 6825 9673 6837 9676
rect 6871 9673 6883 9707
rect 6825 9667 6883 9673
rect 16482 9664 16488 9716
rect 16540 9704 16546 9716
rect 23014 9704 23020 9716
rect 16540 9676 23020 9704
rect 16540 9664 16546 9676
rect 23014 9664 23020 9676
rect 23072 9664 23078 9716
rect 4982 9636 4988 9648
rect 3528 9608 4988 9636
rect 4982 9596 4988 9608
rect 5040 9636 5046 9648
rect 6365 9639 6423 9645
rect 6365 9636 6377 9639
rect 5040 9608 6377 9636
rect 5040 9596 5046 9608
rect 6365 9605 6377 9608
rect 6411 9605 6423 9639
rect 6365 9599 6423 9605
rect 12894 9596 12900 9648
rect 12952 9636 12958 9648
rect 12952 9608 19196 9636
rect 12952 9596 12958 9608
rect 3326 9568 3332 9580
rect 3287 9540 3332 9568
rect 3326 9528 3332 9540
rect 3384 9528 3390 9580
rect 5445 9571 5503 9577
rect 5445 9537 5457 9571
rect 5491 9568 5503 9571
rect 6086 9568 6092 9580
rect 5491 9540 6092 9568
rect 5491 9537 5503 9540
rect 5445 9531 5503 9537
rect 6086 9528 6092 9540
rect 6144 9568 6150 9580
rect 6641 9571 6699 9577
rect 6144 9540 6592 9568
rect 6144 9528 6150 9540
rect 4525 9503 4583 9509
rect 4525 9469 4537 9503
rect 4571 9469 4583 9503
rect 4525 9463 4583 9469
rect 4540 9432 4568 9463
rect 4614 9460 4620 9512
rect 4672 9500 4678 9512
rect 4801 9503 4859 9509
rect 4801 9500 4813 9503
rect 4672 9472 4813 9500
rect 4672 9460 4678 9472
rect 4801 9469 4813 9472
rect 4847 9469 4859 9503
rect 4801 9463 4859 9469
rect 5166 9460 5172 9512
rect 5224 9500 5230 9512
rect 6457 9503 6515 9509
rect 6457 9500 6469 9503
rect 5224 9472 6469 9500
rect 5224 9460 5230 9472
rect 5276 9441 5304 9472
rect 6457 9469 6469 9472
rect 6503 9469 6515 9503
rect 6564 9500 6592 9540
rect 6641 9537 6653 9571
rect 6687 9568 6699 9571
rect 7742 9568 7748 9580
rect 6687 9540 7748 9568
rect 6687 9537 6699 9540
rect 6641 9531 6699 9537
rect 7742 9528 7748 9540
rect 7800 9528 7806 9580
rect 12802 9568 12808 9580
rect 12715 9540 12808 9568
rect 12802 9528 12808 9540
rect 12860 9568 12866 9580
rect 19168 9568 19196 9608
rect 19242 9596 19248 9648
rect 19300 9636 19306 9648
rect 22741 9639 22799 9645
rect 22741 9636 22753 9639
rect 19300 9608 22753 9636
rect 19300 9596 19306 9608
rect 22741 9605 22753 9608
rect 22787 9605 22799 9639
rect 22741 9599 22799 9605
rect 20533 9571 20591 9577
rect 20533 9568 20545 9571
rect 12860 9540 15884 9568
rect 19168 9540 20545 9568
rect 12860 9528 12866 9540
rect 12529 9503 12587 9509
rect 6564 9472 7420 9500
rect 6457 9463 6515 9469
rect 7392 9441 7420 9472
rect 12529 9469 12541 9503
rect 12575 9500 12587 9503
rect 12618 9500 12624 9512
rect 12575 9472 12624 9500
rect 12575 9469 12587 9472
rect 12529 9463 12587 9469
rect 12618 9460 12624 9472
rect 12676 9460 12682 9512
rect 15562 9500 15568 9512
rect 15523 9472 15568 9500
rect 15562 9460 15568 9472
rect 15620 9460 15626 9512
rect 15856 9509 15884 9540
rect 20533 9537 20545 9540
rect 20579 9568 20591 9571
rect 20806 9568 20812 9580
rect 20579 9540 20812 9568
rect 20579 9537 20591 9540
rect 20533 9531 20591 9537
rect 20806 9528 20812 9540
rect 20864 9568 20870 9580
rect 21085 9571 21143 9577
rect 21085 9568 21097 9571
rect 20864 9540 21097 9568
rect 20864 9528 20870 9540
rect 21085 9537 21097 9540
rect 21131 9537 21143 9571
rect 21085 9531 21143 9537
rect 21821 9571 21879 9577
rect 21821 9537 21833 9571
rect 21867 9537 21879 9571
rect 21821 9531 21879 9537
rect 15841 9503 15899 9509
rect 15841 9469 15853 9503
rect 15887 9500 15899 9503
rect 16669 9503 16727 9509
rect 16669 9500 16681 9503
rect 15887 9472 16681 9500
rect 15887 9469 15899 9472
rect 15841 9463 15899 9469
rect 16669 9469 16681 9472
rect 16715 9469 16727 9503
rect 16942 9500 16948 9512
rect 16903 9472 16948 9500
rect 16669 9463 16727 9469
rect 16942 9460 16948 9472
rect 17000 9460 17006 9512
rect 20438 9460 20444 9512
rect 20496 9500 20502 9512
rect 21726 9500 21732 9512
rect 20496 9472 21732 9500
rect 20496 9460 20502 9472
rect 21726 9460 21732 9472
rect 21784 9500 21790 9512
rect 21836 9500 21864 9531
rect 22554 9528 22560 9580
rect 22612 9568 22618 9580
rect 23017 9571 23075 9577
rect 23017 9568 23029 9571
rect 22612 9540 23029 9568
rect 22612 9528 22618 9540
rect 23017 9537 23029 9540
rect 23063 9537 23075 9571
rect 23017 9531 23075 9537
rect 23109 9571 23167 9577
rect 23109 9537 23121 9571
rect 23155 9537 23167 9571
rect 23109 9531 23167 9537
rect 21784 9472 21864 9500
rect 21784 9460 21790 9472
rect 22922 9460 22928 9512
rect 22980 9500 22986 9512
rect 23124 9500 23152 9531
rect 23198 9528 23204 9580
rect 23256 9568 23262 9580
rect 23385 9571 23443 9577
rect 23256 9540 23301 9568
rect 23256 9528 23262 9540
rect 23385 9537 23397 9571
rect 23431 9537 23443 9571
rect 23385 9531 23443 9537
rect 23400 9500 23428 9531
rect 22980 9472 23152 9500
rect 23216 9472 23428 9500
rect 22980 9460 22986 9472
rect 23216 9444 23244 9472
rect 5261 9435 5319 9441
rect 4540 9404 5212 9432
rect 5184 9364 5212 9404
rect 5261 9401 5273 9435
rect 5307 9401 5319 9435
rect 5261 9395 5319 9401
rect 7377 9435 7435 9441
rect 7377 9401 7389 9435
rect 7423 9432 7435 9435
rect 9030 9432 9036 9444
rect 7423 9404 9036 9432
rect 7423 9401 7435 9404
rect 7377 9395 7435 9401
rect 9030 9392 9036 9404
rect 9088 9392 9094 9444
rect 18049 9435 18107 9441
rect 18049 9401 18061 9435
rect 18095 9432 18107 9435
rect 19978 9432 19984 9444
rect 18095 9404 19984 9432
rect 18095 9401 18107 9404
rect 18049 9395 18107 9401
rect 19978 9392 19984 9404
rect 20036 9392 20042 9444
rect 22005 9435 22063 9441
rect 22005 9401 22017 9435
rect 22051 9432 22063 9435
rect 22094 9432 22100 9444
rect 22051 9404 22100 9432
rect 22051 9401 22063 9404
rect 22005 9395 22063 9401
rect 22094 9392 22100 9404
rect 22152 9392 22158 9444
rect 23198 9392 23204 9444
rect 23256 9392 23262 9444
rect 5626 9364 5632 9376
rect 5184 9336 5632 9364
rect 5626 9324 5632 9336
rect 5684 9324 5690 9376
rect 6362 9364 6368 9376
rect 6323 9336 6368 9364
rect 6362 9324 6368 9336
rect 6420 9324 6426 9376
rect 7834 9364 7840 9376
rect 7795 9336 7840 9364
rect 7834 9324 7840 9336
rect 7892 9364 7898 9376
rect 8573 9367 8631 9373
rect 8573 9364 8585 9367
rect 7892 9336 8585 9364
rect 7892 9324 7898 9336
rect 8573 9333 8585 9336
rect 8619 9333 8631 9367
rect 9306 9364 9312 9376
rect 9267 9336 9312 9364
rect 8573 9327 8631 9333
rect 9306 9324 9312 9336
rect 9364 9324 9370 9376
rect 10965 9367 11023 9373
rect 10965 9333 10977 9367
rect 11011 9364 11023 9367
rect 11514 9364 11520 9376
rect 11011 9336 11520 9364
rect 11011 9333 11023 9336
rect 10965 9327 11023 9333
rect 11514 9324 11520 9336
rect 11572 9324 11578 9376
rect 13446 9364 13452 9376
rect 13407 9336 13452 9364
rect 13446 9324 13452 9336
rect 13504 9324 13510 9376
rect 14553 9367 14611 9373
rect 14553 9333 14565 9367
rect 14599 9364 14611 9367
rect 15194 9364 15200 9376
rect 14599 9336 15200 9364
rect 14599 9333 14611 9336
rect 14553 9327 14611 9333
rect 15194 9324 15200 9336
rect 15252 9324 15258 9376
rect 18230 9324 18236 9376
rect 18288 9364 18294 9376
rect 18509 9367 18567 9373
rect 18509 9364 18521 9367
rect 18288 9336 18521 9364
rect 18288 9324 18294 9336
rect 18509 9333 18521 9336
rect 18555 9333 18567 9367
rect 18509 9327 18567 9333
rect 21269 9367 21327 9373
rect 21269 9333 21281 9367
rect 21315 9364 21327 9367
rect 22646 9364 22652 9376
rect 21315 9336 22652 9364
rect 21315 9333 21327 9336
rect 21269 9327 21327 9333
rect 22646 9324 22652 9336
rect 22704 9324 22710 9376
rect 1104 9274 68816 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 65654 9274
rect 65706 9222 65718 9274
rect 65770 9222 65782 9274
rect 65834 9222 65846 9274
rect 65898 9222 65910 9274
rect 65962 9222 68816 9274
rect 1104 9200 68816 9222
rect 12802 9160 12808 9172
rect 6564 9132 12808 9160
rect 6564 9033 6592 9132
rect 12802 9120 12808 9132
rect 12860 9120 12866 9172
rect 20438 9160 20444 9172
rect 14108 9132 20444 9160
rect 14108 9092 14136 9132
rect 20438 9120 20444 9132
rect 20496 9120 20502 9172
rect 22094 9160 22100 9172
rect 20640 9132 22100 9160
rect 12406 9064 14136 9092
rect 17313 9095 17371 9101
rect 3237 9027 3295 9033
rect 3237 8993 3249 9027
rect 3283 9024 3295 9027
rect 5261 9027 5319 9033
rect 5261 9024 5273 9027
rect 3283 8996 5273 9024
rect 3283 8993 3295 8996
rect 3237 8987 3295 8993
rect 5261 8993 5273 8996
rect 5307 9024 5319 9027
rect 6549 9027 6607 9033
rect 6549 9024 6561 9027
rect 5307 8996 6561 9024
rect 5307 8993 5319 8996
rect 5261 8987 5319 8993
rect 6549 8993 6561 8996
rect 6595 8993 6607 9027
rect 6549 8987 6607 8993
rect 9490 8984 9496 9036
rect 9548 9024 9554 9036
rect 10321 9027 10379 9033
rect 10321 9024 10333 9027
rect 9548 8996 10333 9024
rect 9548 8984 9554 8996
rect 10321 8993 10333 8996
rect 10367 8993 10379 9027
rect 10321 8987 10379 8993
rect 2682 8956 2688 8968
rect 2643 8928 2688 8956
rect 2682 8916 2688 8928
rect 2740 8916 2746 8968
rect 2961 8959 3019 8965
rect 2961 8925 2973 8959
rect 3007 8925 3019 8959
rect 2961 8919 3019 8925
rect 3053 8959 3111 8965
rect 3053 8925 3065 8959
rect 3099 8956 3111 8959
rect 3326 8956 3332 8968
rect 3099 8928 3332 8956
rect 3099 8925 3111 8928
rect 3053 8919 3111 8925
rect 2976 8888 3004 8919
rect 3326 8916 3332 8928
rect 3384 8956 3390 8968
rect 3878 8956 3884 8968
rect 3384 8928 3884 8956
rect 3384 8916 3390 8928
rect 3878 8916 3884 8928
rect 3936 8916 3942 8968
rect 4985 8959 5043 8965
rect 4985 8925 4997 8959
rect 5031 8956 5043 8959
rect 6178 8956 6184 8968
rect 5031 8928 6184 8956
rect 5031 8925 5043 8928
rect 4985 8919 5043 8925
rect 6178 8916 6184 8928
rect 6236 8916 6242 8968
rect 6273 8959 6331 8965
rect 6273 8925 6285 8959
rect 6319 8956 6331 8959
rect 6638 8956 6644 8968
rect 6319 8928 6644 8956
rect 6319 8925 6331 8928
rect 6273 8919 6331 8925
rect 6638 8916 6644 8928
rect 6696 8916 6702 8968
rect 7009 8959 7067 8965
rect 7009 8925 7021 8959
rect 7055 8956 7067 8959
rect 7098 8956 7104 8968
rect 7055 8928 7104 8956
rect 7055 8925 7067 8928
rect 7009 8919 7067 8925
rect 7098 8916 7104 8928
rect 7156 8916 7162 8968
rect 9306 8916 9312 8968
rect 9364 8956 9370 8968
rect 9401 8959 9459 8965
rect 9401 8956 9413 8959
rect 9364 8928 9413 8956
rect 9364 8916 9370 8928
rect 9401 8925 9413 8928
rect 9447 8956 9459 8959
rect 12406 8956 12434 9064
rect 17313 9061 17325 9095
rect 17359 9092 17371 9095
rect 17359 9064 20208 9092
rect 17359 9061 17371 9064
rect 17313 9055 17371 9061
rect 12526 8984 12532 9036
rect 12584 9024 12590 9036
rect 12989 9027 13047 9033
rect 12989 9024 13001 9027
rect 12584 8996 13001 9024
rect 12584 8984 12590 8996
rect 12989 8993 13001 8996
rect 13035 8993 13047 9027
rect 12989 8987 13047 8993
rect 20180 8968 20208 9064
rect 12710 8956 12716 8968
rect 9447 8928 12434 8956
rect 12623 8928 12716 8956
rect 9447 8925 9459 8928
rect 9401 8919 9459 8925
rect 12710 8916 12716 8928
rect 12768 8916 12774 8968
rect 14093 8959 14151 8965
rect 14093 8925 14105 8959
rect 14139 8956 14151 8959
rect 15933 8959 15991 8965
rect 15933 8956 15945 8959
rect 14139 8928 15945 8956
rect 14139 8925 14151 8928
rect 14093 8919 14151 8925
rect 15933 8925 15945 8928
rect 15979 8956 15991 8959
rect 16574 8956 16580 8968
rect 15979 8928 16580 8956
rect 15979 8925 15991 8928
rect 15933 8919 15991 8925
rect 16574 8916 16580 8928
rect 16632 8916 16638 8968
rect 20162 8916 20168 8968
rect 20220 8956 20226 8968
rect 20640 8965 20668 9132
rect 22094 9120 22100 9132
rect 22152 9120 22158 9172
rect 23198 9052 23204 9104
rect 23256 9052 23262 9104
rect 21637 9027 21695 9033
rect 21637 9024 21649 9027
rect 20916 8996 21649 9024
rect 20533 8959 20591 8965
rect 20533 8956 20545 8959
rect 20220 8928 20545 8956
rect 20220 8916 20226 8928
rect 20533 8925 20545 8928
rect 20579 8925 20591 8959
rect 20533 8919 20591 8925
rect 20625 8959 20683 8965
rect 20625 8925 20637 8959
rect 20671 8925 20683 8959
rect 20625 8919 20683 8925
rect 20714 8916 20720 8968
rect 20772 8956 20778 8968
rect 20916 8965 20944 8996
rect 21637 8993 21649 8996
rect 21683 9024 21695 9027
rect 23216 9024 23244 9052
rect 21683 8996 23428 9024
rect 21683 8993 21695 8996
rect 21637 8987 21695 8993
rect 20901 8959 20959 8965
rect 20772 8928 20817 8956
rect 20772 8916 20778 8928
rect 20901 8925 20913 8959
rect 20947 8925 20959 8959
rect 20901 8919 20959 8925
rect 21266 8916 21272 8968
rect 21324 8956 21330 8968
rect 21361 8959 21419 8965
rect 21361 8956 21373 8959
rect 21324 8928 21373 8956
rect 21324 8916 21330 8928
rect 21361 8925 21373 8928
rect 21407 8925 21419 8959
rect 23017 8959 23075 8965
rect 23017 8956 23029 8959
rect 21361 8919 21419 8925
rect 21468 8928 23029 8956
rect 7282 8897 7288 8900
rect 2976 8860 3740 8888
rect 3712 8832 3740 8860
rect 6288 8860 6914 8888
rect 6288 8832 6316 8860
rect 6886 8832 6914 8860
rect 7276 8851 7288 8897
rect 7340 8888 7346 8900
rect 7340 8860 7376 8888
rect 7282 8848 7288 8851
rect 7340 8848 7346 8860
rect 10134 8848 10140 8900
rect 10192 8888 10198 8900
rect 10566 8891 10624 8897
rect 10566 8888 10578 8891
rect 10192 8860 10578 8888
rect 10192 8848 10198 8860
rect 10566 8857 10578 8860
rect 10612 8857 10624 8891
rect 10566 8851 10624 8857
rect 3694 8780 3700 8832
rect 3752 8820 3758 8832
rect 3789 8823 3847 8829
rect 3789 8820 3801 8823
rect 3752 8792 3801 8820
rect 3752 8780 3758 8792
rect 3789 8789 3801 8792
rect 3835 8789 3847 8823
rect 3789 8783 3847 8789
rect 6270 8780 6276 8832
rect 6328 8780 6334 8832
rect 6886 8820 6920 8832
rect 6827 8792 6920 8820
rect 6914 8780 6920 8792
rect 6972 8820 6978 8832
rect 8389 8823 8447 8829
rect 8389 8820 8401 8823
rect 6972 8792 8401 8820
rect 6972 8780 6978 8792
rect 8389 8789 8401 8792
rect 8435 8789 8447 8823
rect 9582 8820 9588 8832
rect 9543 8792 9588 8820
rect 8389 8783 8447 8789
rect 9582 8780 9588 8792
rect 9640 8780 9646 8832
rect 10410 8780 10416 8832
rect 10468 8820 10474 8832
rect 11701 8823 11759 8829
rect 11701 8820 11713 8823
rect 10468 8792 11713 8820
rect 10468 8780 10474 8792
rect 11701 8789 11713 8792
rect 11747 8789 11759 8823
rect 11701 8783 11759 8789
rect 12253 8823 12311 8829
rect 12253 8789 12265 8823
rect 12299 8820 12311 8823
rect 12342 8820 12348 8832
rect 12299 8792 12348 8820
rect 12299 8789 12311 8792
rect 12253 8783 12311 8789
rect 12342 8780 12348 8792
rect 12400 8780 12406 8832
rect 12728 8820 12756 8916
rect 13170 8848 13176 8900
rect 13228 8888 13234 8900
rect 14338 8891 14396 8897
rect 14338 8888 14350 8891
rect 13228 8860 14350 8888
rect 13228 8848 13234 8860
rect 14338 8857 14350 8860
rect 14384 8857 14396 8891
rect 16200 8891 16258 8897
rect 14338 8851 14396 8857
rect 14476 8860 15608 8888
rect 14476 8820 14504 8860
rect 15470 8820 15476 8832
rect 12728 8792 14504 8820
rect 15431 8792 15476 8820
rect 15470 8780 15476 8792
rect 15528 8780 15534 8832
rect 15580 8820 15608 8860
rect 16200 8857 16212 8891
rect 16246 8888 16258 8891
rect 20257 8891 20315 8897
rect 20257 8888 20269 8891
rect 16246 8860 20269 8888
rect 16246 8857 16258 8860
rect 16200 8851 16258 8857
rect 20257 8857 20269 8860
rect 20303 8857 20315 8891
rect 20257 8851 20315 8857
rect 20346 8848 20352 8900
rect 20404 8888 20410 8900
rect 21468 8888 21496 8928
rect 23017 8925 23029 8928
rect 23063 8925 23075 8959
rect 23017 8919 23075 8925
rect 23109 8959 23167 8965
rect 23109 8925 23121 8959
rect 23155 8925 23167 8959
rect 23109 8919 23167 8925
rect 23201 8959 23259 8965
rect 23201 8925 23213 8959
rect 23247 8956 23259 8959
rect 23290 8956 23296 8968
rect 23247 8928 23296 8956
rect 23247 8925 23259 8928
rect 23201 8919 23259 8925
rect 20404 8860 21496 8888
rect 20404 8848 20410 8860
rect 22094 8848 22100 8900
rect 22152 8888 22158 8900
rect 22922 8888 22928 8900
rect 22152 8860 22928 8888
rect 22152 8848 22158 8860
rect 22922 8848 22928 8860
rect 22980 8888 22986 8900
rect 23124 8888 23152 8919
rect 23290 8916 23296 8928
rect 23348 8916 23354 8968
rect 23400 8965 23428 8996
rect 23385 8959 23443 8965
rect 23385 8925 23397 8959
rect 23431 8925 23443 8959
rect 23385 8919 23443 8925
rect 22980 8860 23152 8888
rect 22980 8848 22986 8860
rect 16666 8820 16672 8832
rect 15580 8792 16672 8820
rect 16666 8780 16672 8792
rect 16724 8780 16730 8832
rect 17862 8820 17868 8832
rect 17823 8792 17868 8820
rect 17862 8780 17868 8792
rect 17920 8780 17926 8832
rect 18417 8823 18475 8829
rect 18417 8789 18429 8823
rect 18463 8820 18475 8823
rect 18506 8820 18512 8832
rect 18463 8792 18512 8820
rect 18463 8789 18475 8792
rect 18417 8783 18475 8789
rect 18506 8780 18512 8792
rect 18564 8780 18570 8832
rect 19337 8823 19395 8829
rect 19337 8789 19349 8823
rect 19383 8820 19395 8823
rect 19426 8820 19432 8832
rect 19383 8792 19432 8820
rect 19383 8789 19395 8792
rect 19337 8783 19395 8789
rect 19426 8780 19432 8792
rect 19484 8780 19490 8832
rect 22738 8820 22744 8832
rect 22699 8792 22744 8820
rect 22738 8780 22744 8792
rect 22796 8780 22802 8832
rect 23124 8820 23152 8860
rect 23290 8820 23296 8832
rect 23124 8792 23296 8820
rect 23290 8780 23296 8792
rect 23348 8780 23354 8832
rect 1104 8730 68816 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 50294 8730
rect 50346 8678 50358 8730
rect 50410 8678 50422 8730
rect 50474 8678 50486 8730
rect 50538 8678 50550 8730
rect 50602 8678 68816 8730
rect 1104 8656 68816 8678
rect 5902 8616 5908 8628
rect 4724 8588 5908 8616
rect 2682 8304 2688 8356
rect 2740 8344 2746 8356
rect 4724 8344 4752 8588
rect 5902 8576 5908 8588
rect 5960 8616 5966 8628
rect 7009 8619 7067 8625
rect 5960 8588 6868 8616
rect 5960 8576 5966 8588
rect 5626 8548 5632 8560
rect 5092 8520 5632 8548
rect 5092 8489 5120 8520
rect 5626 8508 5632 8520
rect 5684 8508 5690 8560
rect 6840 8548 6868 8588
rect 7009 8585 7021 8619
rect 7055 8616 7067 8619
rect 7282 8616 7288 8628
rect 7055 8588 7288 8616
rect 7055 8585 7067 8588
rect 7009 8579 7067 8585
rect 7282 8576 7288 8588
rect 7340 8576 7346 8628
rect 8389 8619 8447 8625
rect 8389 8585 8401 8619
rect 8435 8616 8447 8619
rect 9306 8616 9312 8628
rect 8435 8588 9312 8616
rect 8435 8585 8447 8588
rect 8389 8579 8447 8585
rect 7469 8551 7527 8557
rect 7469 8548 7481 8551
rect 6840 8520 7481 8548
rect 7469 8517 7481 8520
rect 7515 8517 7527 8551
rect 7469 8511 7527 8517
rect 5077 8483 5135 8489
rect 5077 8449 5089 8483
rect 5123 8449 5135 8483
rect 5077 8443 5135 8449
rect 5442 8440 5448 8492
rect 5500 8480 5506 8492
rect 5537 8483 5595 8489
rect 5537 8480 5549 8483
rect 5500 8452 5549 8480
rect 5500 8440 5506 8452
rect 5537 8449 5549 8452
rect 5583 8449 5595 8483
rect 6365 8483 6423 8489
rect 6365 8480 6377 8483
rect 5537 8443 5595 8449
rect 5644 8452 6377 8480
rect 4801 8415 4859 8421
rect 4801 8381 4813 8415
rect 4847 8381 4859 8415
rect 5644 8412 5672 8452
rect 6365 8449 6377 8452
rect 6411 8449 6423 8483
rect 6528 8483 6586 8489
rect 6528 8480 6540 8483
rect 6365 8443 6423 8449
rect 6472 8452 6540 8480
rect 4801 8375 4859 8381
rect 5552 8384 5672 8412
rect 2740 8316 4752 8344
rect 4816 8344 4844 8375
rect 5552 8356 5580 8384
rect 6178 8372 6184 8424
rect 6236 8412 6242 8424
rect 6472 8412 6500 8452
rect 6528 8449 6540 8452
rect 6574 8449 6586 8483
rect 6528 8443 6586 8449
rect 6641 8440 6647 8492
rect 6699 8480 6705 8492
rect 6779 8483 6837 8489
rect 6699 8452 6744 8480
rect 6699 8440 6705 8452
rect 6779 8449 6791 8483
rect 6825 8480 6837 8483
rect 6914 8480 6920 8492
rect 6825 8452 6920 8480
rect 6825 8449 6837 8452
rect 6779 8443 6837 8449
rect 6886 8440 6920 8452
rect 6972 8440 6978 8492
rect 7653 8483 7711 8489
rect 7653 8449 7665 8483
rect 7699 8480 7711 8483
rect 7834 8480 7840 8492
rect 7699 8452 7840 8480
rect 7699 8449 7711 8452
rect 7653 8443 7711 8449
rect 7834 8440 7840 8452
rect 7892 8480 7898 8492
rect 8297 8483 8355 8489
rect 8297 8480 8309 8483
rect 7892 8452 8309 8480
rect 7892 8440 7898 8452
rect 8297 8449 8309 8452
rect 8343 8449 8355 8483
rect 8297 8443 8355 8449
rect 6886 8436 6960 8440
rect 6236 8384 6500 8412
rect 6236 8372 6242 8384
rect 5534 8344 5540 8356
rect 4816 8316 5540 8344
rect 2740 8304 2746 8316
rect 5534 8304 5540 8316
rect 5592 8304 5598 8356
rect 8404 8344 8432 8579
rect 9306 8576 9312 8588
rect 9364 8576 9370 8628
rect 10134 8616 10140 8628
rect 10095 8588 10140 8616
rect 10134 8576 10140 8588
rect 10192 8576 10198 8628
rect 12894 8616 12900 8628
rect 10244 8588 12900 8616
rect 9030 8480 9036 8492
rect 8943 8452 9036 8480
rect 9030 8440 9036 8452
rect 9088 8480 9094 8492
rect 9493 8483 9551 8489
rect 9493 8480 9505 8483
rect 9088 8452 9505 8480
rect 9088 8440 9094 8452
rect 9493 8449 9505 8452
rect 9539 8480 9551 8483
rect 10244 8480 10272 8588
rect 12894 8576 12900 8588
rect 12952 8576 12958 8628
rect 13170 8616 13176 8628
rect 13131 8588 13176 8616
rect 13170 8576 13176 8588
rect 13228 8576 13234 8628
rect 15102 8616 15108 8628
rect 13280 8588 15108 8616
rect 13280 8548 13308 8588
rect 15102 8576 15108 8588
rect 15160 8616 15166 8628
rect 15470 8616 15476 8628
rect 15160 8588 15476 8616
rect 15160 8576 15166 8588
rect 15470 8576 15476 8588
rect 15528 8616 15534 8628
rect 15528 8588 18276 8616
rect 15528 8576 15534 8588
rect 10796 8520 12388 8548
rect 10796 8492 10824 8520
rect 10410 8480 10416 8492
rect 9539 8452 10272 8480
rect 10371 8452 10416 8480
rect 9539 8449 9551 8452
rect 9493 8443 9551 8449
rect 10410 8440 10416 8452
rect 10468 8440 10474 8492
rect 10518 8483 10576 8489
rect 10518 8449 10530 8483
rect 10564 8449 10576 8483
rect 10518 8443 10576 8449
rect 10618 8483 10676 8489
rect 10618 8449 10630 8483
rect 10664 8480 10676 8483
rect 10664 8452 10732 8480
rect 10664 8449 10676 8452
rect 10618 8443 10676 8449
rect 10318 8372 10324 8424
rect 10376 8412 10382 8424
rect 10520 8412 10548 8443
rect 10376 8384 10548 8412
rect 10704 8412 10732 8452
rect 10778 8440 10784 8492
rect 10836 8480 10842 8492
rect 11606 8480 11612 8492
rect 10836 8452 10881 8480
rect 11567 8452 11612 8480
rect 10836 8440 10842 8452
rect 11606 8440 11612 8452
rect 11664 8440 11670 8492
rect 11885 8483 11943 8489
rect 11885 8449 11897 8483
rect 11931 8480 11943 8483
rect 12250 8480 12256 8492
rect 11931 8452 12256 8480
rect 11931 8449 11943 8452
rect 11885 8443 11943 8449
rect 12250 8440 12256 8452
rect 12308 8440 12314 8492
rect 12360 8480 12388 8520
rect 12912 8520 13308 8548
rect 12526 8480 12532 8492
rect 12360 8452 12532 8480
rect 12526 8440 12532 8452
rect 12584 8440 12590 8492
rect 12912 8489 12940 8520
rect 13538 8508 13544 8560
rect 13596 8548 13602 8560
rect 15390 8551 15448 8557
rect 15390 8548 15402 8551
rect 13596 8520 15402 8548
rect 13596 8508 13602 8520
rect 15390 8517 15402 8520
rect 15436 8517 15448 8551
rect 15390 8511 15448 8517
rect 12713 8483 12771 8489
rect 12713 8449 12725 8483
rect 12759 8449 12771 8483
rect 12713 8443 12771 8449
rect 12805 8483 12863 8489
rect 12805 8449 12817 8483
rect 12851 8449 12863 8483
rect 12805 8443 12863 8449
rect 12897 8483 12955 8489
rect 12897 8449 12909 8483
rect 12943 8449 12955 8483
rect 12897 8443 12955 8449
rect 10870 8412 10876 8424
rect 10704 8384 10876 8412
rect 10376 8372 10382 8384
rect 5644 8316 8432 8344
rect 10520 8344 10548 8384
rect 10870 8372 10876 8384
rect 10928 8372 10934 8424
rect 11790 8412 11796 8424
rect 11751 8384 11796 8412
rect 11790 8372 11796 8384
rect 11848 8372 11854 8424
rect 12728 8412 12756 8443
rect 12084 8384 12756 8412
rect 12084 8353 12112 8384
rect 12069 8347 12127 8353
rect 10520 8316 12020 8344
rect 5442 8236 5448 8288
rect 5500 8276 5506 8288
rect 5644 8276 5672 8316
rect 5500 8248 5672 8276
rect 5500 8236 5506 8248
rect 5718 8236 5724 8288
rect 5776 8276 5782 8288
rect 9674 8276 9680 8288
rect 5776 8248 5821 8276
rect 9635 8248 9680 8276
rect 5776 8236 5782 8248
rect 9674 8236 9680 8248
rect 9732 8236 9738 8288
rect 10042 8236 10048 8288
rect 10100 8276 10106 8288
rect 10778 8276 10784 8288
rect 10100 8248 10784 8276
rect 10100 8236 10106 8248
rect 10778 8236 10784 8248
rect 10836 8236 10842 8288
rect 11606 8276 11612 8288
rect 11567 8248 11612 8276
rect 11606 8236 11612 8248
rect 11664 8236 11670 8288
rect 11992 8276 12020 8316
rect 12069 8313 12081 8347
rect 12115 8313 12127 8347
rect 12069 8307 12127 8313
rect 12820 8288 12848 8443
rect 13170 8440 13176 8492
rect 13228 8480 13234 8492
rect 13446 8480 13452 8492
rect 13228 8452 13452 8480
rect 13228 8440 13234 8452
rect 13446 8440 13452 8452
rect 13504 8480 13510 8492
rect 13817 8483 13875 8489
rect 13817 8480 13829 8483
rect 13504 8452 13829 8480
rect 13504 8440 13510 8452
rect 13817 8449 13829 8452
rect 13863 8449 13875 8483
rect 18138 8480 18144 8492
rect 13817 8443 13875 8449
rect 16132 8452 18144 8480
rect 16132 8424 16160 8452
rect 18138 8440 18144 8452
rect 18196 8440 18202 8492
rect 18248 8480 18276 8588
rect 18966 8576 18972 8628
rect 19024 8616 19030 8628
rect 19521 8619 19579 8625
rect 19521 8616 19533 8619
rect 19024 8588 19533 8616
rect 19024 8576 19030 8588
rect 19521 8585 19533 8588
rect 19567 8616 19579 8619
rect 20346 8616 20352 8628
rect 19567 8588 20352 8616
rect 19567 8585 19579 8588
rect 19521 8579 19579 8585
rect 20346 8576 20352 8588
rect 20404 8576 20410 8628
rect 20441 8619 20499 8625
rect 20441 8585 20453 8619
rect 20487 8616 20499 8619
rect 20530 8616 20536 8628
rect 20487 8588 20536 8616
rect 20487 8585 20499 8588
rect 20441 8579 20499 8585
rect 20530 8576 20536 8588
rect 20588 8576 20594 8628
rect 18408 8551 18466 8557
rect 18408 8517 18420 8551
rect 18454 8548 18466 8551
rect 22738 8548 22744 8560
rect 18454 8520 22744 8548
rect 18454 8517 18466 8520
rect 18408 8511 18466 8517
rect 22738 8508 22744 8520
rect 22796 8508 22802 8560
rect 23290 8508 23296 8560
rect 23348 8548 23354 8560
rect 23348 8520 23520 8548
rect 23348 8508 23354 8520
rect 19981 8483 20039 8489
rect 19981 8480 19993 8483
rect 18248 8452 19993 8480
rect 19981 8449 19993 8452
rect 20027 8449 20039 8483
rect 20254 8480 20260 8492
rect 20215 8452 20260 8480
rect 19981 8443 20039 8449
rect 20254 8440 20260 8452
rect 20312 8440 20318 8492
rect 20438 8440 20444 8492
rect 20496 8480 20502 8492
rect 20496 8452 21404 8480
rect 20496 8440 20502 8452
rect 15657 8415 15715 8421
rect 15657 8381 15669 8415
rect 15703 8412 15715 8415
rect 16114 8412 16120 8424
rect 15703 8384 16120 8412
rect 15703 8381 15715 8384
rect 15657 8375 15715 8381
rect 16114 8372 16120 8384
rect 16172 8372 16178 8424
rect 16666 8412 16672 8424
rect 16627 8384 16672 8412
rect 16666 8372 16672 8384
rect 16724 8372 16730 8424
rect 16945 8415 17003 8421
rect 16945 8381 16957 8415
rect 16991 8412 17003 8415
rect 17310 8412 17316 8424
rect 16991 8384 17316 8412
rect 16991 8381 17003 8384
rect 16945 8375 17003 8381
rect 17310 8372 17316 8384
rect 17368 8372 17374 8424
rect 19150 8372 19156 8424
rect 19208 8412 19214 8424
rect 20073 8415 20131 8421
rect 20073 8412 20085 8415
rect 19208 8384 20085 8412
rect 19208 8372 19214 8384
rect 20073 8381 20085 8384
rect 20119 8381 20131 8415
rect 21266 8412 21272 8424
rect 21227 8384 21272 8412
rect 20073 8375 20131 8381
rect 21266 8372 21272 8384
rect 21324 8372 21330 8424
rect 21376 8412 21404 8452
rect 21542 8440 21548 8492
rect 21600 8480 21606 8492
rect 21821 8483 21879 8489
rect 21821 8480 21833 8483
rect 21600 8452 21833 8480
rect 21600 8440 21606 8452
rect 21821 8449 21833 8452
rect 21867 8480 21879 8483
rect 21910 8480 21916 8492
rect 21867 8452 21916 8480
rect 21867 8449 21879 8452
rect 21821 8443 21879 8449
rect 21910 8440 21916 8452
rect 21968 8440 21974 8492
rect 22094 8480 22100 8492
rect 22055 8452 22100 8480
rect 22094 8440 22100 8452
rect 22152 8440 22158 8492
rect 23198 8480 23204 8492
rect 23159 8452 23204 8480
rect 23198 8440 23204 8452
rect 23256 8440 23262 8492
rect 23382 8480 23388 8492
rect 23343 8452 23388 8480
rect 23382 8440 23388 8452
rect 23440 8440 23446 8492
rect 23492 8489 23520 8520
rect 23477 8483 23535 8489
rect 23477 8449 23489 8483
rect 23523 8449 23535 8483
rect 23477 8443 23535 8449
rect 23569 8483 23627 8489
rect 23569 8449 23581 8483
rect 23615 8449 23627 8483
rect 24302 8480 24308 8492
rect 24263 8452 24308 8480
rect 23569 8443 23627 8449
rect 23584 8412 23612 8443
rect 24302 8440 24308 8452
rect 24360 8440 24366 8492
rect 21376 8384 23612 8412
rect 13630 8344 13636 8356
rect 13591 8316 13636 8344
rect 13630 8304 13636 8316
rect 13688 8304 13694 8356
rect 14274 8344 14280 8356
rect 14235 8316 14280 8344
rect 14274 8304 14280 8316
rect 14332 8304 14338 8356
rect 19334 8304 19340 8356
rect 19392 8344 19398 8356
rect 23845 8347 23903 8353
rect 23845 8344 23857 8347
rect 19392 8316 23857 8344
rect 19392 8304 19398 8316
rect 23845 8313 23857 8316
rect 23891 8313 23903 8347
rect 23845 8307 23903 8313
rect 12618 8276 12624 8288
rect 11992 8248 12624 8276
rect 12618 8236 12624 8248
rect 12676 8276 12682 8288
rect 12802 8276 12808 8288
rect 12676 8248 12808 8276
rect 12676 8236 12682 8248
rect 12802 8236 12808 8248
rect 12860 8236 12866 8288
rect 20070 8276 20076 8288
rect 20031 8248 20076 8276
rect 20070 8236 20076 8248
rect 20128 8236 20134 8288
rect 1104 8186 68816 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 65654 8186
rect 65706 8134 65718 8186
rect 65770 8134 65782 8186
rect 65834 8134 65846 8186
rect 65898 8134 65910 8186
rect 65962 8134 68816 8186
rect 1104 8112 68816 8134
rect 4985 8075 5043 8081
rect 4985 8041 4997 8075
rect 5031 8072 5043 8075
rect 5442 8072 5448 8084
rect 5031 8044 5448 8072
rect 5031 8041 5043 8044
rect 4985 8035 5043 8041
rect 5442 8032 5448 8044
rect 5500 8032 5506 8084
rect 8386 8072 8392 8084
rect 5920 8044 8392 8072
rect 4062 7964 4068 8016
rect 4120 8004 4126 8016
rect 5920 8004 5948 8044
rect 8386 8032 8392 8044
rect 8444 8032 8450 8084
rect 9582 8072 9588 8084
rect 9543 8044 9588 8072
rect 9582 8032 9588 8044
rect 9640 8072 9646 8084
rect 10137 8075 10195 8081
rect 10137 8072 10149 8075
rect 9640 8044 10149 8072
rect 9640 8032 9646 8044
rect 10137 8041 10149 8044
rect 10183 8041 10195 8075
rect 10137 8035 10195 8041
rect 10597 8075 10655 8081
rect 10597 8041 10609 8075
rect 10643 8072 10655 8075
rect 10870 8072 10876 8084
rect 10643 8044 10876 8072
rect 10643 8041 10655 8044
rect 10597 8035 10655 8041
rect 4120 7976 5948 8004
rect 10152 8004 10180 8035
rect 10870 8032 10876 8044
rect 10928 8032 10934 8084
rect 11057 8075 11115 8081
rect 11057 8041 11069 8075
rect 11103 8072 11115 8075
rect 11606 8072 11612 8084
rect 11103 8044 11612 8072
rect 11103 8041 11115 8044
rect 11057 8035 11115 8041
rect 11072 8004 11100 8035
rect 11606 8032 11612 8044
rect 11664 8072 11670 8084
rect 11977 8075 12035 8081
rect 11977 8072 11989 8075
rect 11664 8044 11989 8072
rect 11664 8032 11670 8044
rect 11977 8041 11989 8044
rect 12023 8041 12035 8075
rect 13354 8072 13360 8084
rect 11977 8035 12035 8041
rect 12176 8044 13360 8072
rect 10152 7976 11100 8004
rect 4120 7964 4126 7976
rect 5534 7936 5540 7948
rect 5460 7908 5540 7936
rect 5460 7877 5488 7908
rect 5534 7896 5540 7908
rect 5592 7896 5598 7948
rect 5445 7871 5503 7877
rect 5445 7837 5457 7871
rect 5491 7837 5503 7871
rect 5626 7868 5632 7880
rect 5587 7840 5632 7868
rect 5445 7831 5503 7837
rect 5626 7828 5632 7840
rect 5684 7828 5690 7880
rect 5721 7871 5779 7877
rect 5721 7837 5733 7871
rect 5767 7837 5779 7871
rect 5721 7831 5779 7837
rect 5813 7871 5871 7877
rect 5813 7837 5825 7871
rect 5859 7868 5871 7871
rect 5920 7868 5948 7976
rect 9585 7939 9643 7945
rect 9585 7905 9597 7939
rect 9631 7936 9643 7939
rect 9674 7936 9680 7948
rect 9631 7908 9680 7936
rect 9631 7905 9643 7908
rect 9585 7899 9643 7905
rect 9674 7896 9680 7908
rect 9732 7936 9738 7948
rect 10321 7939 10379 7945
rect 10321 7936 10333 7939
rect 9732 7908 10333 7936
rect 9732 7896 9738 7908
rect 10321 7905 10333 7908
rect 10367 7936 10379 7939
rect 11241 7939 11299 7945
rect 11241 7936 11253 7939
rect 10367 7908 11253 7936
rect 10367 7905 10379 7908
rect 10321 7899 10379 7905
rect 11241 7905 11253 7908
rect 11287 7936 11299 7939
rect 11790 7936 11796 7948
rect 11287 7908 11796 7936
rect 11287 7905 11299 7908
rect 11241 7899 11299 7905
rect 11790 7896 11796 7908
rect 11848 7936 11854 7948
rect 12069 7939 12127 7945
rect 12069 7936 12081 7939
rect 11848 7908 12081 7936
rect 11848 7896 11854 7908
rect 12069 7905 12081 7908
rect 12115 7905 12127 7939
rect 12069 7899 12127 7905
rect 5859 7840 5948 7868
rect 7009 7871 7067 7877
rect 5859 7837 5871 7840
rect 5813 7831 5871 7837
rect 7009 7837 7021 7871
rect 7055 7868 7067 7871
rect 7098 7868 7104 7880
rect 7055 7840 7104 7868
rect 7055 7837 7067 7840
rect 7009 7831 7067 7837
rect 4249 7803 4307 7809
rect 4249 7769 4261 7803
rect 4295 7800 4307 7803
rect 4614 7800 4620 7812
rect 4295 7772 4620 7800
rect 4295 7769 4307 7772
rect 4249 7763 4307 7769
rect 4614 7760 4620 7772
rect 4672 7760 4678 7812
rect 4341 7735 4399 7741
rect 4341 7701 4353 7735
rect 4387 7732 4399 7735
rect 4798 7732 4804 7744
rect 4387 7704 4804 7732
rect 4387 7701 4399 7704
rect 4341 7695 4399 7701
rect 4798 7692 4804 7704
rect 4856 7692 4862 7744
rect 5736 7732 5764 7831
rect 7098 7828 7104 7840
rect 7156 7828 7162 7880
rect 9398 7868 9404 7880
rect 9359 7840 9404 7868
rect 9398 7828 9404 7840
rect 9456 7828 9462 7880
rect 10413 7871 10471 7877
rect 10413 7868 10425 7871
rect 9508 7840 10425 7868
rect 6089 7803 6147 7809
rect 6089 7769 6101 7803
rect 6135 7800 6147 7803
rect 7254 7803 7312 7809
rect 7254 7800 7266 7803
rect 6135 7772 7266 7800
rect 6135 7769 6147 7772
rect 6089 7763 6147 7769
rect 7254 7769 7266 7772
rect 7300 7769 7312 7803
rect 7254 7763 7312 7769
rect 8754 7760 8760 7812
rect 8812 7800 8818 7812
rect 9508 7800 9536 7840
rect 10413 7837 10425 7840
rect 10459 7837 10471 7871
rect 10413 7831 10471 7837
rect 11333 7871 11391 7877
rect 11333 7837 11345 7871
rect 11379 7868 11391 7871
rect 12176 7868 12204 8044
rect 13354 8032 13360 8044
rect 13412 8032 13418 8084
rect 13538 8072 13544 8084
rect 13499 8044 13544 8072
rect 13538 8032 13544 8044
rect 13596 8032 13602 8084
rect 16574 8032 16580 8084
rect 16632 8072 16638 8084
rect 16945 8075 17003 8081
rect 16945 8072 16957 8075
rect 16632 8044 16957 8072
rect 16632 8032 16638 8044
rect 16945 8041 16957 8044
rect 16991 8041 17003 8075
rect 21542 8072 21548 8084
rect 21503 8044 21548 8072
rect 16945 8035 17003 8041
rect 21542 8032 21548 8044
rect 21600 8032 21606 8084
rect 21726 8032 21732 8084
rect 21784 8072 21790 8084
rect 25041 8075 25099 8081
rect 25041 8072 25053 8075
rect 21784 8044 25053 8072
rect 21784 8032 21790 8044
rect 15470 8004 15476 8016
rect 12268 7976 15476 8004
rect 12268 7877 12296 7976
rect 15470 7964 15476 7976
rect 15528 7964 15534 8016
rect 20346 7964 20352 8016
rect 20404 8004 20410 8016
rect 23290 8004 23296 8016
rect 20404 7976 22968 8004
rect 20404 7964 20410 7976
rect 12802 7896 12808 7948
rect 12860 7936 12866 7948
rect 21545 7939 21603 7945
rect 21545 7936 21557 7939
rect 12860 7908 13216 7936
rect 12860 7896 12866 7908
rect 11379 7840 12204 7868
rect 12253 7871 12311 7877
rect 11379 7837 11391 7840
rect 11333 7831 11391 7837
rect 12253 7837 12265 7871
rect 12299 7837 12311 7871
rect 12253 7831 12311 7837
rect 12526 7828 12532 7880
rect 12584 7868 12590 7880
rect 13188 7877 13216 7908
rect 20548 7908 21557 7936
rect 12897 7871 12955 7877
rect 12897 7868 12909 7871
rect 12584 7840 12909 7868
rect 12584 7828 12590 7840
rect 12897 7837 12909 7840
rect 12943 7837 12955 7871
rect 12897 7831 12955 7837
rect 13081 7871 13139 7877
rect 13081 7837 13093 7871
rect 13127 7837 13139 7871
rect 13081 7831 13139 7837
rect 13173 7871 13231 7877
rect 13173 7837 13185 7871
rect 13219 7837 13231 7871
rect 13173 7831 13231 7837
rect 13265 7871 13323 7877
rect 13265 7837 13277 7871
rect 13311 7868 13323 7871
rect 14274 7868 14280 7880
rect 13311 7840 14280 7868
rect 13311 7837 13323 7840
rect 13265 7831 13323 7837
rect 8812 7772 9536 7800
rect 9677 7803 9735 7809
rect 8812 7760 8818 7772
rect 9677 7769 9689 7803
rect 9723 7800 9735 7803
rect 10137 7803 10195 7809
rect 10137 7800 10149 7803
rect 9723 7772 10149 7800
rect 9723 7769 9735 7772
rect 9677 7763 9735 7769
rect 10137 7769 10149 7772
rect 10183 7800 10195 7803
rect 10502 7800 10508 7812
rect 10183 7772 10508 7800
rect 10183 7769 10195 7772
rect 10137 7763 10195 7769
rect 10502 7760 10508 7772
rect 10560 7800 10566 7812
rect 11057 7803 11115 7809
rect 11057 7800 11069 7803
rect 10560 7772 11069 7800
rect 10560 7760 10566 7772
rect 11057 7769 11069 7772
rect 11103 7800 11115 7803
rect 11698 7800 11704 7812
rect 11103 7772 11704 7800
rect 11103 7769 11115 7772
rect 11057 7763 11115 7769
rect 11698 7760 11704 7772
rect 11756 7800 11762 7812
rect 11977 7803 12035 7809
rect 11977 7800 11989 7803
rect 11756 7772 11989 7800
rect 11756 7760 11762 7772
rect 11977 7769 11989 7772
rect 12023 7769 12035 7803
rect 13096 7800 13124 7831
rect 14274 7828 14280 7840
rect 14332 7828 14338 7880
rect 14553 7871 14611 7877
rect 14553 7837 14565 7871
rect 14599 7837 14611 7871
rect 15194 7868 15200 7880
rect 15107 7840 15200 7868
rect 14553 7831 14611 7837
rect 11977 7763 12035 7769
rect 12452 7772 13124 7800
rect 14568 7800 14596 7831
rect 15194 7828 15200 7840
rect 15252 7868 15258 7880
rect 16022 7868 16028 7880
rect 15252 7840 16028 7868
rect 15252 7828 15258 7840
rect 16022 7828 16028 7840
rect 16080 7828 16086 7880
rect 17862 7828 17868 7880
rect 17920 7868 17926 7880
rect 18049 7871 18107 7877
rect 18049 7868 18061 7871
rect 17920 7840 18061 7868
rect 17920 7828 17926 7840
rect 18049 7837 18061 7840
rect 18095 7837 18107 7871
rect 18049 7831 18107 7837
rect 18138 7828 18144 7880
rect 18196 7868 18202 7880
rect 19245 7871 19303 7877
rect 19245 7868 19257 7871
rect 18196 7840 19257 7868
rect 18196 7828 18202 7840
rect 19245 7837 19257 7840
rect 19291 7837 19303 7871
rect 19245 7831 19303 7837
rect 20070 7828 20076 7880
rect 20128 7868 20134 7880
rect 20548 7868 20576 7908
rect 21545 7905 21557 7908
rect 21591 7905 21603 7939
rect 21545 7899 21603 7905
rect 21450 7868 21456 7880
rect 20128 7840 20576 7868
rect 21411 7840 21456 7868
rect 20128 7828 20134 7840
rect 21450 7828 21456 7840
rect 21508 7828 21514 7880
rect 22940 7877 22968 7976
rect 23032 7976 23296 8004
rect 23032 7877 23060 7976
rect 23290 7964 23296 7976
rect 23348 7964 23354 8016
rect 23198 7896 23204 7948
rect 23256 7936 23262 7948
rect 23256 7908 23336 7936
rect 23256 7896 23262 7908
rect 22925 7871 22983 7877
rect 22925 7837 22937 7871
rect 22971 7837 22983 7871
rect 22925 7831 22983 7837
rect 23017 7871 23075 7877
rect 23017 7837 23029 7871
rect 23063 7837 23075 7871
rect 23017 7831 23075 7837
rect 23106 7828 23112 7880
rect 23164 7868 23170 7880
rect 23308 7877 23336 7908
rect 24596 7877 24624 8044
rect 25041 8041 25053 8044
rect 25087 8041 25099 8075
rect 25041 8035 25099 8041
rect 23293 7871 23351 7877
rect 23164 7840 23209 7868
rect 23164 7828 23170 7840
rect 23293 7837 23305 7871
rect 23339 7837 23351 7871
rect 23293 7831 23351 7837
rect 24581 7871 24639 7877
rect 24581 7837 24593 7871
rect 24627 7837 24639 7871
rect 24581 7831 24639 7837
rect 14734 7800 14740 7812
rect 14568 7772 14740 7800
rect 6638 7732 6644 7744
rect 5736 7704 6644 7732
rect 6638 7692 6644 7704
rect 6696 7692 6702 7744
rect 9217 7735 9275 7741
rect 9217 7701 9229 7735
rect 9263 7732 9275 7735
rect 10226 7732 10232 7744
rect 9263 7704 10232 7732
rect 9263 7701 9275 7704
rect 9217 7695 9275 7701
rect 10226 7692 10232 7704
rect 10284 7692 10290 7744
rect 11517 7735 11575 7741
rect 11517 7701 11529 7735
rect 11563 7732 11575 7735
rect 11882 7732 11888 7744
rect 11563 7704 11888 7732
rect 11563 7701 11575 7704
rect 11517 7695 11575 7701
rect 11882 7692 11888 7704
rect 11940 7692 11946 7744
rect 12452 7741 12480 7772
rect 14734 7760 14740 7772
rect 14792 7800 14798 7812
rect 15378 7800 15384 7812
rect 14792 7772 15384 7800
rect 14792 7760 14798 7772
rect 15378 7760 15384 7772
rect 15436 7760 15442 7812
rect 15654 7800 15660 7812
rect 15615 7772 15660 7800
rect 15654 7760 15660 7772
rect 15712 7760 15718 7812
rect 19512 7803 19570 7809
rect 19512 7769 19524 7803
rect 19558 7800 19570 7803
rect 22649 7803 22707 7809
rect 22649 7800 22661 7803
rect 19558 7772 22661 7800
rect 19558 7769 19570 7772
rect 19512 7763 19570 7769
rect 22649 7769 22661 7772
rect 22695 7769 22707 7803
rect 22649 7763 22707 7769
rect 12437 7735 12495 7741
rect 12437 7701 12449 7735
rect 12483 7701 12495 7735
rect 14366 7732 14372 7744
rect 14327 7704 14372 7732
rect 12437 7695 12495 7701
rect 14366 7692 14372 7704
rect 14424 7692 14430 7744
rect 15010 7732 15016 7744
rect 14971 7704 15016 7732
rect 15010 7692 15016 7704
rect 15068 7692 15074 7744
rect 15194 7692 15200 7744
rect 15252 7732 15258 7744
rect 17865 7735 17923 7741
rect 17865 7732 17877 7735
rect 15252 7704 17877 7732
rect 15252 7692 15258 7704
rect 17865 7701 17877 7704
rect 17911 7701 17923 7735
rect 17865 7695 17923 7701
rect 18693 7735 18751 7741
rect 18693 7701 18705 7735
rect 18739 7732 18751 7735
rect 18874 7732 18880 7744
rect 18739 7704 18880 7732
rect 18739 7701 18751 7704
rect 18693 7695 18751 7701
rect 18874 7692 18880 7704
rect 18932 7692 18938 7744
rect 20346 7692 20352 7744
rect 20404 7732 20410 7744
rect 20625 7735 20683 7741
rect 20625 7732 20637 7735
rect 20404 7704 20637 7732
rect 20404 7692 20410 7704
rect 20625 7701 20637 7704
rect 20671 7701 20683 7735
rect 20625 7695 20683 7701
rect 21821 7735 21879 7741
rect 21821 7701 21833 7735
rect 21867 7732 21879 7735
rect 22278 7732 22284 7744
rect 21867 7704 22284 7732
rect 21867 7701 21879 7704
rect 21821 7695 21879 7701
rect 22278 7692 22284 7704
rect 22336 7692 22342 7744
rect 24394 7732 24400 7744
rect 24355 7704 24400 7732
rect 24394 7692 24400 7704
rect 24452 7692 24458 7744
rect 1104 7642 68816 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 50294 7642
rect 50346 7590 50358 7642
rect 50410 7590 50422 7642
rect 50474 7590 50486 7642
rect 50538 7590 50550 7642
rect 50602 7590 68816 7642
rect 1104 7568 68816 7590
rect 4249 7531 4307 7537
rect 4249 7497 4261 7531
rect 4295 7497 4307 7531
rect 4249 7491 4307 7497
rect 5169 7531 5227 7537
rect 5169 7497 5181 7531
rect 5215 7528 5227 7531
rect 5626 7528 5632 7540
rect 5215 7500 5632 7528
rect 5215 7497 5227 7500
rect 5169 7491 5227 7497
rect 4264 7460 4292 7491
rect 5626 7488 5632 7500
rect 5684 7488 5690 7540
rect 6178 7488 6184 7540
rect 6236 7528 6242 7540
rect 6825 7531 6883 7537
rect 6825 7528 6837 7531
rect 6236 7500 6837 7528
rect 6236 7488 6242 7500
rect 6825 7497 6837 7500
rect 6871 7497 6883 7531
rect 6825 7491 6883 7497
rect 10318 7488 10324 7540
rect 10376 7488 10382 7540
rect 11698 7488 11704 7540
rect 11756 7528 11762 7540
rect 12434 7528 12440 7540
rect 11756 7500 12440 7528
rect 11756 7488 11762 7500
rect 12434 7488 12440 7500
rect 12492 7488 12498 7540
rect 16942 7488 16948 7540
rect 17000 7528 17006 7540
rect 19521 7531 19579 7537
rect 17000 7500 17080 7528
rect 17000 7488 17006 7500
rect 4709 7463 4767 7469
rect 4709 7460 4721 7463
rect 4264 7432 4721 7460
rect 4709 7429 4721 7432
rect 4755 7460 4767 7463
rect 5350 7460 5356 7472
rect 4755 7432 5356 7460
rect 4755 7429 4767 7432
rect 4709 7423 4767 7429
rect 5350 7420 5356 7432
rect 5408 7460 5414 7472
rect 6365 7463 6423 7469
rect 6365 7460 6377 7463
rect 5408 7432 6377 7460
rect 5408 7420 5414 7432
rect 6365 7429 6377 7432
rect 6411 7429 6423 7463
rect 6365 7423 6423 7429
rect 7098 7420 7104 7472
rect 7156 7460 7162 7472
rect 7837 7463 7895 7469
rect 7837 7460 7849 7463
rect 7156 7432 7849 7460
rect 7156 7420 7162 7432
rect 7837 7429 7849 7432
rect 7883 7429 7895 7463
rect 7837 7423 7895 7429
rect 10336 7407 10364 7488
rect 10778 7420 10784 7472
rect 10836 7460 10842 7472
rect 10836 7432 11836 7460
rect 10836 7420 10842 7432
rect 3878 7352 3884 7404
rect 3936 7392 3942 7404
rect 4065 7395 4123 7401
rect 4065 7392 4077 7395
rect 3936 7364 4077 7392
rect 3936 7352 3942 7364
rect 4065 7361 4077 7364
rect 4111 7361 4123 7395
rect 4982 7392 4988 7404
rect 4943 7364 4988 7392
rect 4065 7355 4123 7361
rect 4982 7352 4988 7364
rect 5040 7352 5046 7404
rect 5629 7395 5687 7401
rect 5629 7361 5641 7395
rect 5675 7392 5687 7395
rect 6086 7392 6092 7404
rect 5675 7364 6092 7392
rect 5675 7361 5687 7364
rect 5629 7355 5687 7361
rect 6086 7352 6092 7364
rect 6144 7352 6150 7404
rect 6641 7395 6699 7401
rect 6641 7361 6653 7395
rect 6687 7392 6699 7395
rect 9490 7392 9496 7404
rect 6687 7364 9496 7392
rect 6687 7361 6699 7364
rect 6641 7355 6699 7361
rect 9490 7352 9496 7364
rect 9548 7352 9554 7404
rect 9582 7352 9588 7404
rect 9640 7392 9646 7404
rect 10042 7392 10048 7404
rect 9640 7364 9685 7392
rect 10003 7364 10048 7392
rect 9640 7352 9646 7364
rect 10042 7352 10048 7364
rect 10100 7352 10106 7404
rect 10226 7401 10232 7404
rect 10224 7392 10232 7401
rect 10187 7364 10232 7392
rect 10224 7355 10232 7364
rect 10226 7352 10232 7355
rect 10284 7352 10290 7404
rect 10324 7401 10382 7407
rect 10324 7367 10336 7401
rect 10370 7367 10382 7401
rect 10324 7361 10382 7367
rect 10413 7395 10471 7401
rect 10413 7361 10425 7395
rect 10459 7361 10471 7395
rect 11808 7392 11836 7432
rect 11882 7420 11888 7472
rect 11940 7460 11946 7472
rect 12802 7460 12808 7472
rect 11940 7432 12434 7460
rect 11940 7420 11946 7432
rect 12406 7401 12434 7432
rect 12531 7432 12808 7460
rect 12531 7404 12559 7432
rect 12802 7420 12808 7432
rect 12860 7420 12866 7472
rect 17052 7407 17080 7500
rect 19521 7497 19533 7531
rect 19567 7528 19579 7531
rect 20438 7528 20444 7540
rect 19567 7500 20444 7528
rect 19567 7497 19579 7500
rect 19521 7491 19579 7497
rect 20438 7488 20444 7500
rect 20496 7488 20502 7540
rect 21450 7528 21456 7540
rect 21008 7500 21456 7528
rect 18408 7463 18466 7469
rect 18408 7429 18420 7463
rect 18454 7460 18466 7463
rect 19334 7460 19340 7472
rect 18454 7432 19340 7460
rect 18454 7429 18466 7432
rect 18408 7423 18466 7429
rect 19334 7420 19340 7432
rect 19392 7420 19398 7472
rect 12253 7395 12311 7401
rect 12253 7392 12265 7395
rect 10413 7355 10471 7361
rect 11609 7379 11667 7385
rect 4893 7327 4951 7333
rect 4893 7293 4905 7327
rect 4939 7324 4951 7327
rect 5534 7324 5540 7336
rect 4939 7296 5540 7324
rect 4939 7293 4951 7296
rect 4893 7287 4951 7293
rect 5534 7284 5540 7296
rect 5592 7324 5598 7336
rect 6457 7327 6515 7333
rect 6457 7324 6469 7327
rect 5592 7296 6469 7324
rect 5592 7284 5598 7296
rect 5828 7265 5856 7296
rect 6457 7293 6469 7296
rect 6503 7293 6515 7327
rect 6457 7287 6515 7293
rect 5813 7259 5871 7265
rect 5813 7225 5825 7259
rect 5859 7225 5871 7259
rect 5813 7219 5871 7225
rect 10318 7216 10324 7268
rect 10376 7256 10382 7268
rect 10428 7256 10456 7355
rect 11609 7345 11621 7379
rect 11655 7345 11667 7379
rect 11808 7364 12265 7392
rect 12253 7361 12265 7364
rect 12299 7361 12311 7395
rect 12406 7395 12474 7401
rect 12406 7364 12428 7395
rect 12253 7355 12311 7361
rect 12416 7361 12428 7364
rect 12462 7361 12474 7395
rect 12416 7355 12474 7361
rect 12516 7398 12574 7404
rect 12516 7364 12528 7398
rect 12562 7364 12574 7398
rect 12516 7358 12574 7364
rect 12621 7395 12679 7401
rect 12710 7395 12716 7404
rect 12621 7361 12633 7395
rect 12667 7367 12716 7395
rect 12667 7361 12679 7367
rect 12621 7355 12679 7361
rect 12710 7352 12716 7367
rect 12768 7352 12774 7404
rect 13357 7395 13415 7401
rect 13357 7361 13369 7395
rect 13403 7361 13415 7395
rect 15930 7392 15936 7404
rect 15843 7364 15936 7392
rect 13357 7355 13415 7361
rect 11609 7339 11667 7345
rect 10376 7228 10456 7256
rect 11624 7256 11652 7339
rect 11698 7256 11704 7268
rect 11624 7228 11704 7256
rect 10376 7216 10382 7228
rect 11698 7216 11704 7228
rect 11756 7216 11762 7268
rect 12158 7216 12164 7268
rect 12216 7256 12222 7268
rect 12710 7256 12716 7268
rect 12216 7228 12716 7256
rect 12216 7216 12222 7228
rect 12710 7216 12716 7228
rect 12768 7216 12774 7268
rect 13372 7256 13400 7355
rect 15930 7352 15936 7364
rect 15988 7392 15994 7404
rect 15988 7364 16068 7392
rect 15988 7352 15994 7364
rect 16040 7324 16068 7364
rect 16850 7352 16856 7404
rect 16908 7401 16914 7404
rect 17037 7401 17095 7407
rect 16908 7395 16957 7401
rect 16908 7361 16911 7395
rect 16945 7361 16957 7395
rect 17037 7367 17049 7401
rect 17083 7367 17095 7401
rect 17037 7361 17095 7367
rect 16908 7355 16957 7361
rect 16908 7352 16914 7355
rect 17126 7352 17132 7404
rect 17184 7392 17190 7404
rect 17184 7364 17229 7392
rect 17184 7352 17190 7364
rect 17310 7352 17316 7404
rect 17368 7392 17374 7404
rect 18138 7392 18144 7404
rect 17368 7364 17413 7392
rect 18099 7364 18144 7392
rect 17368 7352 17374 7364
rect 18138 7352 18144 7364
rect 18196 7352 18202 7404
rect 19150 7352 19156 7404
rect 19208 7392 19214 7404
rect 21008 7401 21036 7500
rect 21450 7488 21456 7500
rect 21508 7528 21514 7540
rect 21821 7531 21879 7537
rect 21821 7528 21833 7531
rect 21508 7500 21833 7528
rect 21508 7488 21514 7500
rect 21821 7497 21833 7500
rect 21867 7528 21879 7531
rect 22833 7531 22891 7537
rect 21867 7500 22508 7528
rect 21867 7497 21879 7500
rect 21821 7491 21879 7497
rect 20809 7395 20867 7401
rect 20809 7392 20821 7395
rect 19208 7364 20821 7392
rect 19208 7352 19214 7364
rect 20809 7361 20821 7364
rect 20855 7361 20867 7395
rect 20809 7355 20867 7361
rect 20993 7395 21051 7401
rect 20993 7361 21005 7395
rect 21039 7361 21051 7395
rect 22002 7392 22008 7404
rect 21963 7364 22008 7392
rect 20993 7355 21051 7361
rect 22002 7352 22008 7364
rect 22060 7352 22066 7404
rect 22480 7401 22508 7500
rect 22833 7497 22845 7531
rect 22879 7528 22891 7531
rect 23750 7528 23756 7540
rect 22879 7500 23756 7528
rect 22879 7497 22891 7500
rect 22833 7491 22891 7497
rect 23750 7488 23756 7500
rect 23808 7488 23814 7540
rect 22465 7395 22523 7401
rect 22465 7361 22477 7395
rect 22511 7392 22523 7395
rect 23290 7392 23296 7404
rect 22511 7364 23296 7392
rect 22511 7361 22523 7364
rect 22465 7355 22523 7361
rect 23290 7352 23296 7364
rect 23348 7352 23354 7404
rect 17494 7324 17500 7336
rect 16040 7296 17500 7324
rect 17494 7284 17500 7296
rect 17552 7284 17558 7336
rect 22554 7324 22560 7336
rect 22515 7296 22560 7324
rect 22554 7284 22560 7296
rect 22612 7284 22618 7336
rect 23014 7284 23020 7336
rect 23072 7324 23078 7336
rect 23385 7327 23443 7333
rect 23385 7324 23397 7327
rect 23072 7296 23397 7324
rect 23072 7284 23078 7296
rect 23385 7293 23397 7296
rect 23431 7293 23443 7327
rect 24394 7324 24400 7336
rect 23385 7287 23443 7293
rect 23492 7296 24400 7324
rect 12820 7228 13400 7256
rect 16117 7259 16175 7265
rect 4985 7191 5043 7197
rect 4985 7157 4997 7191
rect 5031 7188 5043 7191
rect 5718 7188 5724 7200
rect 5031 7160 5724 7188
rect 5031 7157 5043 7160
rect 4985 7151 5043 7157
rect 5718 7148 5724 7160
rect 5776 7188 5782 7200
rect 6365 7191 6423 7197
rect 6365 7188 6377 7191
rect 5776 7160 6377 7188
rect 5776 7148 5782 7160
rect 6365 7157 6377 7160
rect 6411 7157 6423 7191
rect 6365 7151 6423 7157
rect 7377 7191 7435 7197
rect 7377 7157 7389 7191
rect 7423 7188 7435 7191
rect 7926 7188 7932 7200
rect 7423 7160 7932 7188
rect 7423 7157 7435 7160
rect 7377 7151 7435 7157
rect 7926 7148 7932 7160
rect 7984 7148 7990 7200
rect 10689 7191 10747 7197
rect 10689 7157 10701 7191
rect 10735 7188 10747 7191
rect 11054 7188 11060 7200
rect 10735 7160 11060 7188
rect 10735 7157 10747 7160
rect 10689 7151 10747 7157
rect 11054 7148 11060 7160
rect 11112 7148 11118 7200
rect 11793 7191 11851 7197
rect 11793 7157 11805 7191
rect 11839 7188 11851 7191
rect 11882 7188 11888 7200
rect 11839 7160 11888 7188
rect 11839 7157 11851 7160
rect 11793 7151 11851 7157
rect 11882 7148 11888 7160
rect 11940 7148 11946 7200
rect 12342 7148 12348 7200
rect 12400 7188 12406 7200
rect 12820 7188 12848 7228
rect 16117 7225 16129 7259
rect 16163 7256 16175 7259
rect 17586 7256 17592 7268
rect 16163 7228 17592 7256
rect 16163 7225 16175 7228
rect 16117 7219 16175 7225
rect 17586 7216 17592 7228
rect 17644 7216 17650 7268
rect 20625 7259 20683 7265
rect 20625 7225 20637 7259
rect 20671 7256 20683 7259
rect 21450 7256 21456 7268
rect 20671 7228 21456 7256
rect 20671 7225 20683 7228
rect 20625 7219 20683 7225
rect 21450 7216 21456 7228
rect 21508 7216 21514 7268
rect 22066 7228 22692 7256
rect 12400 7160 12848 7188
rect 12400 7148 12406 7160
rect 12894 7148 12900 7200
rect 12952 7188 12958 7200
rect 14642 7188 14648 7200
rect 12952 7160 12997 7188
rect 14603 7160 14648 7188
rect 12952 7148 12958 7160
rect 14642 7148 14648 7160
rect 14700 7188 14706 7200
rect 15654 7188 15660 7200
rect 14700 7160 15660 7188
rect 14700 7148 14706 7160
rect 15654 7148 15660 7160
rect 15712 7148 15718 7200
rect 16666 7188 16672 7200
rect 16627 7160 16672 7188
rect 16666 7148 16672 7160
rect 16724 7148 16730 7200
rect 20165 7191 20223 7197
rect 20165 7157 20177 7191
rect 20211 7188 20223 7191
rect 20714 7188 20720 7200
rect 20211 7160 20720 7188
rect 20211 7157 20223 7160
rect 20165 7151 20223 7157
rect 20714 7148 20720 7160
rect 20772 7148 20778 7200
rect 20993 7191 21051 7197
rect 20993 7157 21005 7191
rect 21039 7188 21051 7191
rect 21542 7188 21548 7200
rect 21039 7160 21548 7188
rect 21039 7157 21051 7160
rect 20993 7151 21051 7157
rect 21542 7148 21548 7160
rect 21600 7188 21606 7200
rect 22066 7188 22094 7228
rect 22664 7197 22692 7228
rect 23492 7197 23520 7296
rect 24394 7284 24400 7296
rect 24452 7284 24458 7336
rect 21600 7160 22094 7188
rect 22649 7191 22707 7197
rect 21600 7148 21606 7160
rect 22649 7157 22661 7191
rect 22695 7188 22707 7191
rect 23477 7191 23535 7197
rect 23477 7188 23489 7191
rect 22695 7160 23489 7188
rect 22695 7157 22707 7160
rect 22649 7151 22707 7157
rect 23477 7157 23489 7160
rect 23523 7157 23535 7191
rect 23477 7151 23535 7157
rect 23566 7148 23572 7200
rect 23624 7188 23630 7200
rect 23661 7191 23719 7197
rect 23661 7188 23673 7191
rect 23624 7160 23673 7188
rect 23624 7148 23630 7160
rect 23661 7157 23673 7160
rect 23707 7157 23719 7191
rect 23661 7151 23719 7157
rect 1104 7098 68816 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 65654 7098
rect 65706 7046 65718 7098
rect 65770 7046 65782 7098
rect 65834 7046 65846 7098
rect 65898 7046 65910 7098
rect 65962 7046 68816 7098
rect 1104 7024 68816 7046
rect 5445 6987 5503 6993
rect 5445 6953 5457 6987
rect 5491 6984 5503 6987
rect 6086 6984 6092 6996
rect 5491 6956 6092 6984
rect 5491 6953 5503 6956
rect 5445 6947 5503 6953
rect 6086 6944 6092 6956
rect 6144 6944 6150 6996
rect 8386 6944 8392 6996
rect 8444 6984 8450 6996
rect 9217 6987 9275 6993
rect 9217 6984 9229 6987
rect 8444 6956 9229 6984
rect 8444 6944 8450 6956
rect 9217 6953 9229 6956
rect 9263 6953 9275 6987
rect 9217 6947 9275 6953
rect 10321 6987 10379 6993
rect 10321 6953 10333 6987
rect 10367 6984 10379 6987
rect 10502 6984 10508 6996
rect 10367 6956 10508 6984
rect 10367 6953 10379 6956
rect 10321 6947 10379 6953
rect 10502 6944 10508 6956
rect 10560 6944 10566 6996
rect 13354 6984 13360 6996
rect 13315 6956 13360 6984
rect 13354 6944 13360 6956
rect 13412 6944 13418 6996
rect 14918 6984 14924 6996
rect 14879 6956 14924 6984
rect 14918 6944 14924 6956
rect 14976 6944 14982 6996
rect 15470 6984 15476 6996
rect 15431 6956 15476 6984
rect 15470 6944 15476 6956
rect 15528 6944 15534 6996
rect 16850 6944 16856 6996
rect 16908 6984 16914 6996
rect 17497 6987 17555 6993
rect 17497 6984 17509 6987
rect 16908 6956 17509 6984
rect 16908 6944 16914 6956
rect 17497 6953 17509 6956
rect 17543 6984 17555 6987
rect 20254 6984 20260 6996
rect 17543 6956 20260 6984
rect 17543 6953 17555 6956
rect 17497 6947 17555 6953
rect 20254 6944 20260 6956
rect 20312 6944 20318 6996
rect 20349 6987 20407 6993
rect 20349 6953 20361 6987
rect 20395 6984 20407 6987
rect 20806 6984 20812 6996
rect 20395 6956 20812 6984
rect 20395 6953 20407 6956
rect 20349 6947 20407 6953
rect 20806 6944 20812 6956
rect 20864 6944 20870 6996
rect 24394 6984 24400 6996
rect 24355 6956 24400 6984
rect 24394 6944 24400 6956
rect 24452 6944 24458 6996
rect 12526 6876 12532 6928
rect 12584 6916 12590 6928
rect 12713 6919 12771 6925
rect 12713 6916 12725 6919
rect 12584 6888 12725 6916
rect 12584 6876 12590 6888
rect 12713 6885 12725 6888
rect 12759 6885 12771 6919
rect 12713 6879 12771 6885
rect 14185 6919 14243 6925
rect 14185 6885 14197 6919
rect 14231 6916 14243 6919
rect 18693 6919 18751 6925
rect 14231 6888 14412 6916
rect 14231 6885 14243 6888
rect 14185 6879 14243 6885
rect 2682 6808 2688 6860
rect 2740 6848 2746 6860
rect 4617 6851 4675 6857
rect 4617 6848 4629 6851
rect 2740 6820 4629 6848
rect 2740 6808 2746 6820
rect 4617 6817 4629 6820
rect 4663 6817 4675 6851
rect 4617 6811 4675 6817
rect 5166 6808 5172 6860
rect 5224 6848 5230 6860
rect 6549 6851 6607 6857
rect 5224 6820 6316 6848
rect 5224 6808 5230 6820
rect 4341 6783 4399 6789
rect 4341 6749 4353 6783
rect 4387 6780 4399 6783
rect 5442 6780 5448 6792
rect 4387 6752 5448 6780
rect 4387 6749 4399 6752
rect 4341 6743 4399 6749
rect 5442 6740 5448 6752
rect 5500 6740 5506 6792
rect 5626 6740 5632 6792
rect 5684 6780 5690 6792
rect 5905 6783 5963 6789
rect 5905 6780 5917 6783
rect 5684 6752 5917 6780
rect 5684 6740 5690 6752
rect 5905 6749 5917 6752
rect 5951 6749 5963 6783
rect 6086 6780 6092 6792
rect 6047 6752 6092 6780
rect 5905 6743 5963 6749
rect 6086 6740 6092 6752
rect 6144 6740 6150 6792
rect 6288 6789 6316 6820
rect 6549 6817 6561 6851
rect 6595 6848 6607 6851
rect 6595 6820 6960 6848
rect 6595 6817 6607 6820
rect 6549 6811 6607 6817
rect 6181 6783 6239 6789
rect 6181 6749 6193 6783
rect 6227 6749 6239 6783
rect 6181 6743 6239 6749
rect 6273 6783 6331 6789
rect 6273 6749 6285 6783
rect 6319 6780 6331 6783
rect 6319 6752 6776 6780
rect 6319 6749 6331 6752
rect 6273 6743 6331 6749
rect 6196 6712 6224 6743
rect 6638 6712 6644 6724
rect 6196 6684 6644 6712
rect 6638 6672 6644 6684
rect 6696 6672 6702 6724
rect 6748 6644 6776 6752
rect 6932 6712 6960 6820
rect 10778 6808 10784 6860
rect 10836 6848 10842 6860
rect 14274 6848 14280 6860
rect 10836 6820 14280 6848
rect 10836 6808 10842 6820
rect 14274 6808 14280 6820
rect 14332 6808 14338 6860
rect 14384 6848 14412 6888
rect 18693 6885 18705 6919
rect 18739 6885 18751 6919
rect 20824 6916 20852 6944
rect 22002 6916 22008 6928
rect 20824 6888 22008 6916
rect 18693 6879 18751 6885
rect 15930 6848 15936 6860
rect 14384 6820 15936 6848
rect 15930 6808 15936 6820
rect 15988 6808 15994 6860
rect 16114 6848 16120 6860
rect 16075 6820 16120 6848
rect 16114 6808 16120 6820
rect 16172 6808 16178 6860
rect 18708 6848 18736 6879
rect 22002 6876 22008 6888
rect 22060 6916 22066 6928
rect 22097 6919 22155 6925
rect 22097 6916 22109 6919
rect 22060 6888 22109 6916
rect 22060 6876 22066 6888
rect 22097 6885 22109 6888
rect 22143 6885 22155 6919
rect 22097 6879 22155 6885
rect 20990 6848 20996 6860
rect 18708 6820 20996 6848
rect 20990 6808 20996 6820
rect 21048 6808 21054 6860
rect 23290 6808 23296 6860
rect 23348 6848 23354 6860
rect 24486 6848 24492 6860
rect 23348 6820 23888 6848
rect 24447 6820 24492 6848
rect 23348 6808 23354 6820
rect 7009 6783 7067 6789
rect 7009 6749 7021 6783
rect 7055 6780 7067 6783
rect 8294 6780 8300 6792
rect 7055 6752 8300 6780
rect 7055 6749 7067 6752
rect 7009 6743 7067 6749
rect 8294 6740 8300 6752
rect 8352 6740 8358 6792
rect 9214 6780 9220 6792
rect 9175 6752 9220 6780
rect 9214 6740 9220 6752
rect 9272 6740 9278 6792
rect 9401 6783 9459 6789
rect 9401 6749 9413 6783
rect 9447 6749 9459 6783
rect 9401 6743 9459 6749
rect 9493 6783 9551 6789
rect 9493 6749 9505 6783
rect 9539 6749 9551 6783
rect 10134 6780 10140 6792
rect 10095 6752 10140 6780
rect 9493 6743 9551 6749
rect 7254 6715 7312 6721
rect 7254 6712 7266 6715
rect 6932 6684 7266 6712
rect 7254 6681 7266 6684
rect 7300 6681 7312 6715
rect 9416 6712 9444 6743
rect 7254 6675 7312 6681
rect 8404 6684 9444 6712
rect 8404 6653 8432 6684
rect 8389 6647 8447 6653
rect 8389 6644 8401 6647
rect 6748 6616 8401 6644
rect 8389 6613 8401 6616
rect 8435 6613 8447 6647
rect 8389 6607 8447 6613
rect 9214 6604 9220 6656
rect 9272 6644 9278 6656
rect 9508 6644 9536 6743
rect 10134 6740 10140 6752
rect 10192 6740 10198 6792
rect 10965 6783 11023 6789
rect 10965 6749 10977 6783
rect 11011 6780 11023 6783
rect 11238 6780 11244 6792
rect 11011 6752 11244 6780
rect 11011 6749 11023 6752
rect 10965 6743 11023 6749
rect 11238 6740 11244 6752
rect 11296 6740 11302 6792
rect 11514 6740 11520 6792
rect 11572 6780 11578 6792
rect 11609 6783 11667 6789
rect 11609 6780 11621 6783
rect 11572 6752 11621 6780
rect 11572 6740 11578 6752
rect 11609 6749 11621 6752
rect 11655 6749 11667 6783
rect 11609 6743 11667 6749
rect 12253 6783 12311 6789
rect 12253 6749 12265 6783
rect 12299 6780 12311 6783
rect 12897 6783 12955 6789
rect 12299 6752 12848 6780
rect 12299 6749 12311 6752
rect 12253 6743 12311 6749
rect 10042 6672 10048 6724
rect 10100 6712 10106 6724
rect 12268 6712 12296 6743
rect 10100 6684 12296 6712
rect 10100 6672 10106 6684
rect 9272 6616 9536 6644
rect 9677 6647 9735 6653
rect 9272 6604 9278 6616
rect 9677 6613 9689 6647
rect 9723 6644 9735 6647
rect 10594 6644 10600 6656
rect 9723 6616 10600 6644
rect 9723 6613 9735 6616
rect 9677 6607 9735 6613
rect 10594 6604 10600 6616
rect 10652 6604 10658 6656
rect 10686 6604 10692 6656
rect 10744 6644 10750 6656
rect 10781 6647 10839 6653
rect 10781 6644 10793 6647
rect 10744 6616 10793 6644
rect 10744 6604 10750 6616
rect 10781 6613 10793 6616
rect 10827 6613 10839 6647
rect 10781 6607 10839 6613
rect 11330 6604 11336 6656
rect 11388 6644 11394 6656
rect 11425 6647 11483 6653
rect 11425 6644 11437 6647
rect 11388 6616 11437 6644
rect 11388 6604 11394 6616
rect 11425 6613 11437 6616
rect 11471 6613 11483 6647
rect 12066 6644 12072 6656
rect 12027 6616 12072 6644
rect 11425 6607 11483 6613
rect 12066 6604 12072 6616
rect 12124 6604 12130 6656
rect 12820 6644 12848 6752
rect 12897 6749 12909 6783
rect 12943 6749 12955 6783
rect 13538 6780 13544 6792
rect 13499 6752 13544 6780
rect 12897 6743 12955 6749
rect 12912 6712 12940 6743
rect 13538 6740 13544 6752
rect 13596 6740 13602 6792
rect 14090 6740 14096 6792
rect 14148 6780 14154 6792
rect 14829 6783 14887 6789
rect 14829 6780 14841 6783
rect 14148 6752 14841 6780
rect 14148 6740 14154 6752
rect 14829 6749 14841 6752
rect 14875 6749 14887 6783
rect 15010 6780 15016 6792
rect 14971 6752 15016 6780
rect 14829 6743 14887 6749
rect 15010 6740 15016 6752
rect 15068 6740 15074 6792
rect 15657 6783 15715 6789
rect 15657 6749 15669 6783
rect 15703 6780 15715 6783
rect 15746 6780 15752 6792
rect 15703 6752 15752 6780
rect 15703 6749 15715 6752
rect 15657 6743 15715 6749
rect 15746 6740 15752 6752
rect 15804 6740 15810 6792
rect 16384 6783 16442 6789
rect 16384 6749 16396 6783
rect 16430 6780 16442 6783
rect 16666 6780 16672 6792
rect 16430 6752 16672 6780
rect 16430 6749 16442 6752
rect 16384 6743 16442 6749
rect 16666 6740 16672 6752
rect 16724 6740 16730 6792
rect 18509 6783 18567 6789
rect 18509 6749 18521 6783
rect 18555 6780 18567 6783
rect 18874 6780 18880 6792
rect 18555 6752 18880 6780
rect 18555 6749 18567 6752
rect 18509 6743 18567 6749
rect 18874 6740 18880 6752
rect 18932 6740 18938 6792
rect 19245 6783 19303 6789
rect 19245 6780 19257 6783
rect 18984 6752 19257 6780
rect 13078 6712 13084 6724
rect 12912 6684 13084 6712
rect 13078 6672 13084 6684
rect 13136 6712 13142 6724
rect 14734 6712 14740 6724
rect 13136 6684 14740 6712
rect 13136 6672 13142 6684
rect 14734 6672 14740 6684
rect 14792 6672 14798 6724
rect 18049 6715 18107 6721
rect 18049 6681 18061 6715
rect 18095 6712 18107 6715
rect 18782 6712 18788 6724
rect 18095 6684 18788 6712
rect 18095 6681 18107 6684
rect 18049 6675 18107 6681
rect 18782 6672 18788 6684
rect 18840 6712 18846 6724
rect 18984 6712 19012 6752
rect 19245 6749 19257 6752
rect 19291 6749 19303 6783
rect 21269 6783 21327 6789
rect 21269 6780 21281 6783
rect 19245 6743 19303 6749
rect 19352 6752 21281 6780
rect 19352 6712 19380 6752
rect 21269 6749 21281 6752
rect 21315 6749 21327 6783
rect 21269 6743 21327 6749
rect 21361 6783 21419 6789
rect 21361 6749 21373 6783
rect 21407 6749 21419 6783
rect 21361 6743 21419 6749
rect 18840 6684 19012 6712
rect 19260 6684 19380 6712
rect 20441 6715 20499 6721
rect 18840 6672 18846 6684
rect 13814 6644 13820 6656
rect 12820 6616 13820 6644
rect 13814 6604 13820 6616
rect 13872 6604 13878 6656
rect 13906 6604 13912 6656
rect 13964 6644 13970 6656
rect 14645 6647 14703 6653
rect 14645 6644 14657 6647
rect 13964 6616 14657 6644
rect 13964 6604 13970 6616
rect 14645 6613 14657 6616
rect 14691 6613 14703 6647
rect 14645 6607 14703 6613
rect 16666 6604 16672 6656
rect 16724 6644 16730 6656
rect 19260 6644 19288 6684
rect 20441 6681 20453 6715
rect 20487 6712 20499 6715
rect 20530 6712 20536 6724
rect 20487 6684 20536 6712
rect 20487 6681 20499 6684
rect 20441 6675 20499 6681
rect 20530 6672 20536 6684
rect 20588 6672 20594 6724
rect 21376 6712 21404 6743
rect 21450 6740 21456 6792
rect 21508 6780 21514 6792
rect 21637 6783 21695 6789
rect 21508 6752 21553 6780
rect 21508 6740 21514 6752
rect 21637 6749 21649 6783
rect 21683 6780 21695 6783
rect 22462 6780 22468 6792
rect 21683 6752 22468 6780
rect 21683 6749 21695 6752
rect 21637 6743 21695 6749
rect 22462 6740 22468 6752
rect 22520 6740 22526 6792
rect 23382 6780 23388 6792
rect 23343 6752 23388 6780
rect 23382 6740 23388 6752
rect 23440 6740 23446 6792
rect 23477 6783 23535 6789
rect 23477 6749 23489 6783
rect 23523 6749 23535 6783
rect 23477 6743 23535 6749
rect 23569 6783 23627 6789
rect 23569 6749 23581 6783
rect 23615 6749 23627 6783
rect 23569 6743 23627 6749
rect 22094 6712 22100 6724
rect 21376 6684 22100 6712
rect 22094 6672 22100 6684
rect 22152 6712 22158 6724
rect 23290 6712 23296 6724
rect 22152 6684 23296 6712
rect 22152 6672 22158 6684
rect 23290 6672 23296 6684
rect 23348 6712 23354 6724
rect 23492 6712 23520 6743
rect 23348 6684 23520 6712
rect 23348 6672 23354 6684
rect 19426 6644 19432 6656
rect 16724 6616 19288 6644
rect 19387 6616 19432 6644
rect 16724 6604 16730 6616
rect 19426 6604 19432 6616
rect 19484 6604 19490 6656
rect 20714 6604 20720 6656
rect 20772 6644 20778 6656
rect 20993 6647 21051 6653
rect 20993 6644 21005 6647
rect 20772 6616 21005 6644
rect 20772 6604 20778 6616
rect 20993 6613 21005 6616
rect 21039 6613 21051 6647
rect 20993 6607 21051 6613
rect 21174 6604 21180 6656
rect 21232 6644 21238 6656
rect 23109 6647 23167 6653
rect 23109 6644 23121 6647
rect 21232 6616 23121 6644
rect 21232 6604 21238 6616
rect 23109 6613 23121 6616
rect 23155 6613 23167 6647
rect 23584 6644 23612 6743
rect 23658 6740 23664 6792
rect 23716 6780 23722 6792
rect 23753 6783 23811 6789
rect 23753 6780 23765 6783
rect 23716 6752 23765 6780
rect 23716 6740 23722 6752
rect 23753 6749 23765 6752
rect 23799 6749 23811 6783
rect 23860 6780 23888 6820
rect 24486 6808 24492 6820
rect 24544 6808 24550 6860
rect 24397 6783 24455 6789
rect 24397 6780 24409 6783
rect 23860 6752 24409 6780
rect 23753 6743 23811 6749
rect 24397 6749 24409 6752
rect 24443 6749 24455 6783
rect 24397 6743 24455 6749
rect 24765 6647 24823 6653
rect 24765 6644 24777 6647
rect 23584 6616 24777 6644
rect 23109 6607 23167 6613
rect 24765 6613 24777 6616
rect 24811 6613 24823 6647
rect 24765 6607 24823 6613
rect 1104 6554 68816 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 50294 6554
rect 50346 6502 50358 6554
rect 50410 6502 50422 6554
rect 50474 6502 50486 6554
rect 50538 6502 50550 6554
rect 50602 6502 68816 6554
rect 1104 6480 68816 6502
rect 4893 6443 4951 6449
rect 4893 6409 4905 6443
rect 4939 6440 4951 6443
rect 8386 6440 8392 6452
rect 4939 6412 8392 6440
rect 4939 6409 4951 6412
rect 4893 6403 4951 6409
rect 3694 6372 3700 6384
rect 3344 6344 3700 6372
rect 2682 6304 2688 6316
rect 2643 6276 2688 6304
rect 2682 6264 2688 6276
rect 2740 6264 2746 6316
rect 3344 6313 3372 6344
rect 3694 6332 3700 6344
rect 3752 6372 3758 6384
rect 4908 6372 4936 6403
rect 8386 6400 8392 6412
rect 8444 6400 8450 6452
rect 8849 6443 8907 6449
rect 8849 6409 8861 6443
rect 8895 6440 8907 6443
rect 10042 6440 10048 6452
rect 8895 6412 10048 6440
rect 8895 6409 8907 6412
rect 8849 6403 8907 6409
rect 10042 6400 10048 6412
rect 10100 6400 10106 6452
rect 10226 6440 10232 6452
rect 10187 6412 10232 6440
rect 10226 6400 10232 6412
rect 10284 6400 10290 6452
rect 12526 6440 12532 6452
rect 10336 6412 12532 6440
rect 5350 6372 5356 6384
rect 3752 6344 4936 6372
rect 5311 6344 5356 6372
rect 3752 6332 3758 6344
rect 5350 6332 5356 6344
rect 5408 6332 5414 6384
rect 10336 6372 10364 6412
rect 12526 6400 12532 6412
rect 12584 6400 12590 6452
rect 12802 6400 12808 6452
rect 12860 6440 12866 6452
rect 14090 6440 14096 6452
rect 12860 6412 14096 6440
rect 12860 6400 12866 6412
rect 14090 6400 14096 6412
rect 14148 6440 14154 6452
rect 14277 6443 14335 6449
rect 14277 6440 14289 6443
rect 14148 6412 14289 6440
rect 14148 6400 14154 6412
rect 14277 6409 14289 6412
rect 14323 6409 14335 6443
rect 16942 6440 16948 6452
rect 14277 6403 14335 6409
rect 14384 6412 16948 6440
rect 10594 6372 10600 6384
rect 5644 6344 10364 6372
rect 10428 6344 10600 6372
rect 3329 6307 3387 6313
rect 3329 6273 3341 6307
rect 3375 6273 3387 6307
rect 3329 6267 3387 6273
rect 3786 6264 3792 6316
rect 3844 6304 3850 6316
rect 3973 6307 4031 6313
rect 3973 6304 3985 6307
rect 3844 6276 3985 6304
rect 3844 6264 3850 6276
rect 3973 6273 3985 6276
rect 4019 6273 4031 6307
rect 3973 6267 4031 6273
rect 4062 6264 4068 6316
rect 4120 6304 4126 6316
rect 5534 6304 5540 6316
rect 4120 6276 4165 6304
rect 5495 6276 5540 6304
rect 4120 6264 4126 6276
rect 5534 6264 5540 6276
rect 5592 6264 5598 6316
rect 5644 6313 5672 6344
rect 5629 6307 5687 6313
rect 5629 6273 5641 6307
rect 5675 6273 5687 6307
rect 5629 6267 5687 6273
rect 6270 6264 6276 6316
rect 6328 6304 6334 6316
rect 9214 6304 9220 6316
rect 6328 6276 9220 6304
rect 6328 6264 6334 6276
rect 9214 6264 9220 6276
rect 9272 6264 9278 6316
rect 9309 6307 9367 6313
rect 9309 6273 9321 6307
rect 9355 6304 9367 6307
rect 9355 6276 9996 6304
rect 9355 6273 9367 6276
rect 9309 6267 9367 6273
rect 3878 6196 3884 6248
rect 3936 6236 3942 6248
rect 3936 6208 5396 6236
rect 3936 6196 3942 6208
rect 2869 6171 2927 6177
rect 2869 6137 2881 6171
rect 2915 6168 2927 6171
rect 4341 6171 4399 6177
rect 2915 6140 4016 6168
rect 2915 6137 2927 6140
rect 2869 6131 2927 6137
rect 3988 6112 4016 6140
rect 4341 6137 4353 6171
rect 4387 6168 4399 6171
rect 5258 6168 5264 6180
rect 4387 6140 5264 6168
rect 4387 6137 4399 6140
rect 4341 6131 4399 6137
rect 5258 6128 5264 6140
rect 5316 6128 5322 6180
rect 5368 6168 5396 6208
rect 5442 6196 5448 6248
rect 5500 6236 5506 6248
rect 9858 6236 9864 6248
rect 5500 6208 9864 6236
rect 5500 6196 5506 6208
rect 9858 6196 9864 6208
rect 9916 6196 9922 6248
rect 6546 6168 6552 6180
rect 5368 6140 6552 6168
rect 6546 6128 6552 6140
rect 6604 6128 6610 6180
rect 7193 6171 7251 6177
rect 7193 6137 7205 6171
rect 7239 6168 7251 6171
rect 9968 6168 9996 6276
rect 10042 6264 10048 6316
rect 10100 6304 10106 6316
rect 10321 6307 10379 6313
rect 10100 6276 10145 6304
rect 10100 6264 10106 6276
rect 10321 6273 10333 6307
rect 10367 6304 10379 6307
rect 10428 6304 10456 6344
rect 10594 6332 10600 6344
rect 10652 6332 10658 6384
rect 12158 6372 12164 6384
rect 10796 6344 12164 6372
rect 10367 6276 10456 6304
rect 10505 6307 10563 6313
rect 10367 6273 10379 6276
rect 10321 6267 10379 6273
rect 10505 6273 10517 6307
rect 10551 6304 10563 6307
rect 10686 6304 10692 6316
rect 10551 6276 10692 6304
rect 10551 6273 10563 6276
rect 10505 6267 10563 6273
rect 10686 6264 10692 6276
rect 10744 6264 10750 6316
rect 10796 6313 10824 6344
rect 12158 6332 12164 6344
rect 12216 6332 12222 6384
rect 12710 6372 12716 6384
rect 12268 6344 12716 6372
rect 10781 6307 10839 6313
rect 10781 6273 10793 6307
rect 10827 6273 10839 6307
rect 11606 6304 11612 6316
rect 11567 6276 11612 6304
rect 10781 6267 10839 6273
rect 11606 6264 11612 6276
rect 11664 6264 11670 6316
rect 11698 6264 11704 6316
rect 11756 6304 11762 6316
rect 12268 6304 12296 6344
rect 12710 6332 12716 6344
rect 12768 6332 12774 6384
rect 12894 6332 12900 6384
rect 12952 6372 12958 6384
rect 13142 6375 13200 6381
rect 13142 6372 13154 6375
rect 12952 6344 13154 6372
rect 12952 6332 12958 6344
rect 13142 6341 13154 6344
rect 13188 6341 13200 6375
rect 13142 6335 13200 6341
rect 13538 6332 13544 6384
rect 13596 6372 13602 6384
rect 14182 6372 14188 6384
rect 13596 6344 14188 6372
rect 13596 6332 13602 6344
rect 14182 6332 14188 6344
rect 14240 6372 14246 6384
rect 14384 6372 14412 6412
rect 16942 6400 16948 6412
rect 17000 6400 17006 6452
rect 18141 6443 18199 6449
rect 18141 6409 18153 6443
rect 18187 6440 18199 6443
rect 18414 6440 18420 6452
rect 18187 6412 18420 6440
rect 18187 6409 18199 6412
rect 18141 6403 18199 6409
rect 18414 6400 18420 6412
rect 18472 6440 18478 6452
rect 18472 6412 21956 6440
rect 18472 6400 18478 6412
rect 14240 6344 14412 6372
rect 16868 6344 18644 6372
rect 14240 6332 14246 6344
rect 11756 6276 12296 6304
rect 12437 6307 12495 6313
rect 11756 6264 11762 6276
rect 12437 6273 12449 6307
rect 12483 6304 12495 6307
rect 12802 6304 12808 6316
rect 12483 6276 12808 6304
rect 12483 6273 12495 6276
rect 12437 6267 12495 6273
rect 12802 6264 12808 6276
rect 12860 6264 12866 6316
rect 13722 6264 13728 6316
rect 13780 6304 13786 6316
rect 15010 6304 15016 6316
rect 13780 6276 15016 6304
rect 13780 6264 13786 6276
rect 15010 6264 15016 6276
rect 15068 6264 15074 6316
rect 15102 6264 15108 6316
rect 15160 6304 15166 6316
rect 16868 6313 16896 6344
rect 16117 6307 16175 6313
rect 15160 6276 15205 6304
rect 15160 6264 15166 6276
rect 16117 6273 16129 6307
rect 16163 6273 16175 6307
rect 16117 6267 16175 6273
rect 16853 6307 16911 6313
rect 16853 6273 16865 6307
rect 16899 6273 16911 6307
rect 16853 6267 16911 6273
rect 17681 6307 17739 6313
rect 17681 6273 17693 6307
rect 17727 6304 17739 6307
rect 18506 6304 18512 6316
rect 17727 6276 18512 6304
rect 17727 6273 17739 6276
rect 17681 6267 17739 6273
rect 12894 6236 12900 6248
rect 10612 6208 12664 6236
rect 12855 6208 12900 6236
rect 10612 6168 10640 6208
rect 12636 6180 12664 6208
rect 12894 6196 12900 6208
rect 12952 6196 12958 6248
rect 16132 6236 16160 6267
rect 18506 6264 18512 6276
rect 18564 6264 18570 6316
rect 18616 6304 18644 6344
rect 19058 6332 19064 6384
rect 19116 6332 19122 6384
rect 19276 6375 19334 6381
rect 19276 6341 19288 6375
rect 19322 6372 19334 6375
rect 21821 6375 21879 6381
rect 21821 6372 21833 6375
rect 19322 6344 21833 6372
rect 19322 6341 19334 6344
rect 19276 6335 19334 6341
rect 21821 6341 21833 6344
rect 21867 6341 21879 6375
rect 21821 6335 21879 6341
rect 19076 6304 19104 6332
rect 19978 6304 19984 6316
rect 18616 6276 19984 6304
rect 19978 6264 19984 6276
rect 20036 6264 20042 6316
rect 20530 6264 20536 6316
rect 20588 6304 20594 6316
rect 20625 6307 20683 6313
rect 20625 6304 20637 6307
rect 20588 6276 20637 6304
rect 20588 6264 20594 6276
rect 20625 6273 20637 6276
rect 20671 6273 20683 6307
rect 20625 6267 20683 6273
rect 20806 6264 20812 6316
rect 20864 6304 20870 6316
rect 21085 6307 21143 6313
rect 21085 6304 21097 6307
rect 20864 6276 21097 6304
rect 20864 6264 20870 6276
rect 21085 6273 21097 6276
rect 21131 6273 21143 6307
rect 21928 6304 21956 6412
rect 22094 6400 22100 6452
rect 22152 6400 22158 6452
rect 22112 6372 22140 6400
rect 22112 6344 22232 6372
rect 22204 6313 22232 6344
rect 22097 6307 22155 6313
rect 22097 6304 22109 6307
rect 21928 6276 22109 6304
rect 21085 6267 21143 6273
rect 22097 6273 22109 6276
rect 22143 6273 22155 6307
rect 22097 6267 22155 6273
rect 22189 6307 22247 6313
rect 22189 6273 22201 6307
rect 22235 6273 22247 6307
rect 22189 6267 22247 6273
rect 22278 6264 22284 6316
rect 22336 6304 22342 6316
rect 22336 6276 22381 6304
rect 22336 6264 22342 6276
rect 22462 6264 22468 6316
rect 22520 6304 22526 6316
rect 23201 6307 23259 6313
rect 23201 6304 23213 6307
rect 22520 6276 23213 6304
rect 22520 6264 22526 6276
rect 23201 6273 23213 6276
rect 23247 6304 23259 6307
rect 23658 6304 23664 6316
rect 23247 6276 23664 6304
rect 23247 6273 23259 6276
rect 23201 6267 23259 6273
rect 23658 6264 23664 6276
rect 23716 6264 23722 6316
rect 18230 6236 18236 6248
rect 16132 6208 18236 6236
rect 18230 6196 18236 6208
rect 18288 6196 18294 6248
rect 19521 6239 19579 6245
rect 19521 6205 19533 6239
rect 19567 6205 19579 6239
rect 22922 6236 22928 6248
rect 22835 6208 22928 6236
rect 19521 6199 19579 6205
rect 7239 6140 10640 6168
rect 7239 6137 7251 6140
rect 7193 6131 7251 6137
rect 12250 6128 12256 6180
rect 12308 6168 12314 6180
rect 12308 6140 12353 6168
rect 12308 6128 12314 6140
rect 12618 6128 12624 6180
rect 12676 6128 12682 6180
rect 15286 6168 15292 6180
rect 13832 6140 15292 6168
rect 3513 6103 3571 6109
rect 3513 6069 3525 6103
rect 3559 6100 3571 6103
rect 3786 6100 3792 6112
rect 3559 6072 3792 6100
rect 3559 6069 3571 6072
rect 3513 6063 3571 6069
rect 3786 6060 3792 6072
rect 3844 6060 3850 6112
rect 3970 6060 3976 6112
rect 4028 6100 4034 6112
rect 5445 6103 5503 6109
rect 4028 6072 4121 6100
rect 4028 6060 4034 6072
rect 5445 6069 5457 6103
rect 5491 6100 5503 6103
rect 5718 6100 5724 6112
rect 5491 6072 5724 6100
rect 5491 6069 5503 6072
rect 5445 6063 5503 6069
rect 5718 6060 5724 6072
rect 5776 6060 5782 6112
rect 5813 6103 5871 6109
rect 5813 6069 5825 6103
rect 5859 6100 5871 6103
rect 6086 6100 6092 6112
rect 5859 6072 6092 6100
rect 5859 6069 5871 6072
rect 5813 6063 5871 6069
rect 6086 6060 6092 6072
rect 6144 6060 6150 6112
rect 6641 6103 6699 6109
rect 6641 6069 6653 6103
rect 6687 6100 6699 6103
rect 6822 6100 6828 6112
rect 6687 6072 6828 6100
rect 6687 6069 6699 6072
rect 6641 6063 6699 6069
rect 6822 6060 6828 6072
rect 6880 6060 6886 6112
rect 7745 6103 7803 6109
rect 7745 6069 7757 6103
rect 7791 6100 7803 6103
rect 7834 6100 7840 6112
rect 7791 6072 7840 6100
rect 7791 6069 7803 6072
rect 7745 6063 7803 6069
rect 7834 6060 7840 6072
rect 7892 6060 7898 6112
rect 8297 6103 8355 6109
rect 8297 6069 8309 6103
rect 8343 6100 8355 6103
rect 8662 6100 8668 6112
rect 8343 6072 8668 6100
rect 8343 6069 8355 6072
rect 8297 6063 8355 6069
rect 8662 6060 8668 6072
rect 8720 6060 8726 6112
rect 9214 6060 9220 6112
rect 9272 6100 9278 6112
rect 9493 6103 9551 6109
rect 9493 6100 9505 6103
rect 9272 6072 9505 6100
rect 9272 6060 9278 6072
rect 9493 6069 9505 6072
rect 9539 6069 9551 6103
rect 9493 6063 9551 6069
rect 9674 6060 9680 6112
rect 9732 6100 9738 6112
rect 11606 6100 11612 6112
rect 9732 6072 11612 6100
rect 9732 6060 9738 6072
rect 11606 6060 11612 6072
rect 11664 6060 11670 6112
rect 11793 6103 11851 6109
rect 11793 6069 11805 6103
rect 11839 6100 11851 6103
rect 12066 6100 12072 6112
rect 11839 6072 12072 6100
rect 11839 6069 11851 6072
rect 11793 6063 11851 6069
rect 12066 6060 12072 6072
rect 12124 6060 12130 6112
rect 13630 6060 13636 6112
rect 13688 6100 13694 6112
rect 13832 6100 13860 6140
rect 15286 6128 15292 6140
rect 15344 6128 15350 6180
rect 15381 6171 15439 6177
rect 15381 6137 15393 6171
rect 15427 6168 15439 6171
rect 15427 6140 16528 6168
rect 15427 6137 15439 6140
rect 15381 6131 15439 6137
rect 13688 6072 13860 6100
rect 13688 6060 13694 6072
rect 14918 6060 14924 6112
rect 14976 6100 14982 6112
rect 15013 6103 15071 6109
rect 15013 6100 15025 6103
rect 14976 6072 15025 6100
rect 14976 6060 14982 6072
rect 15013 6069 15025 6072
rect 15059 6069 15071 6103
rect 15013 6063 15071 6069
rect 15562 6060 15568 6112
rect 15620 6100 15626 6112
rect 15933 6103 15991 6109
rect 15933 6100 15945 6103
rect 15620 6072 15945 6100
rect 15620 6060 15626 6072
rect 15933 6069 15945 6072
rect 15979 6069 15991 6103
rect 16500 6100 16528 6140
rect 16574 6128 16580 6180
rect 16632 6168 16638 6180
rect 17497 6171 17555 6177
rect 17497 6168 17509 6171
rect 16632 6140 17509 6168
rect 16632 6128 16638 6140
rect 17497 6137 17509 6140
rect 17543 6137 17555 6171
rect 17497 6131 17555 6137
rect 16850 6100 16856 6112
rect 16500 6072 16856 6100
rect 15933 6063 15991 6069
rect 16850 6060 16856 6072
rect 16908 6060 16914 6112
rect 17034 6100 17040 6112
rect 16995 6072 17040 6100
rect 17034 6060 17040 6072
rect 17092 6060 17098 6112
rect 19242 6060 19248 6112
rect 19300 6100 19306 6112
rect 19536 6100 19564 6199
rect 22922 6196 22928 6208
rect 22980 6236 22986 6248
rect 22980 6208 23244 6236
rect 22980 6196 22986 6208
rect 23216 6180 23244 6208
rect 20254 6128 20260 6180
rect 20312 6168 20318 6180
rect 21174 6168 21180 6180
rect 20312 6140 21180 6168
rect 20312 6128 20318 6140
rect 21174 6128 21180 6140
rect 21232 6128 21238 6180
rect 23198 6128 23204 6180
rect 23256 6128 23262 6180
rect 20438 6100 20444 6112
rect 19300 6072 19564 6100
rect 20399 6072 20444 6100
rect 19300 6060 19306 6072
rect 20438 6060 20444 6072
rect 20496 6060 20502 6112
rect 21266 6100 21272 6112
rect 21227 6072 21272 6100
rect 21266 6060 21272 6072
rect 21324 6060 21330 6112
rect 1104 6010 68816 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 65654 6010
rect 65706 5958 65718 6010
rect 65770 5958 65782 6010
rect 65834 5958 65846 6010
rect 65898 5958 65910 6010
rect 65962 5958 68816 6010
rect 1104 5936 68816 5958
rect 3970 5896 3976 5908
rect 3931 5868 3976 5896
rect 3970 5856 3976 5868
rect 4028 5856 4034 5908
rect 5445 5899 5503 5905
rect 5445 5865 5457 5899
rect 5491 5896 5503 5899
rect 5718 5896 5724 5908
rect 5491 5868 5724 5896
rect 5491 5865 5503 5868
rect 5445 5859 5503 5865
rect 5718 5856 5724 5868
rect 5776 5856 5782 5908
rect 7742 5896 7748 5908
rect 7703 5868 7748 5896
rect 7742 5856 7748 5868
rect 7800 5856 7806 5908
rect 8386 5856 8392 5908
rect 8444 5896 8450 5908
rect 8846 5896 8852 5908
rect 8444 5868 8852 5896
rect 8444 5856 8450 5868
rect 8846 5856 8852 5868
rect 8904 5896 8910 5908
rect 9030 5896 9036 5908
rect 8904 5868 9036 5896
rect 8904 5856 8910 5868
rect 9030 5856 9036 5868
rect 9088 5856 9094 5908
rect 9490 5896 9496 5908
rect 9451 5868 9496 5896
rect 9490 5856 9496 5868
rect 9548 5856 9554 5908
rect 11514 5856 11520 5908
rect 11572 5896 11578 5908
rect 13354 5896 13360 5908
rect 11572 5868 13360 5896
rect 11572 5856 11578 5868
rect 13354 5856 13360 5868
rect 13412 5856 13418 5908
rect 13814 5856 13820 5908
rect 13872 5896 13878 5908
rect 14826 5896 14832 5908
rect 13872 5868 14832 5896
rect 13872 5856 13878 5868
rect 14826 5856 14832 5868
rect 14884 5856 14890 5908
rect 14918 5856 14924 5908
rect 14976 5896 14982 5908
rect 15746 5896 15752 5908
rect 14976 5868 15021 5896
rect 15120 5868 15752 5896
rect 14976 5856 14982 5868
rect 4157 5831 4215 5837
rect 4157 5797 4169 5831
rect 4203 5828 4215 5831
rect 6454 5828 6460 5840
rect 4203 5800 6460 5828
rect 4203 5797 4215 5800
rect 4157 5791 4215 5797
rect 6454 5788 6460 5800
rect 6512 5788 6518 5840
rect 6546 5788 6552 5840
rect 6604 5828 6610 5840
rect 6604 5800 7696 5828
rect 6604 5788 6610 5800
rect 5442 5760 5448 5772
rect 5403 5732 5448 5760
rect 5442 5720 5448 5732
rect 5500 5720 5506 5772
rect 7558 5760 7564 5772
rect 5552 5732 7564 5760
rect 3786 5692 3792 5704
rect 3747 5664 3792 5692
rect 3786 5652 3792 5664
rect 3844 5652 3850 5704
rect 3973 5695 4031 5701
rect 3973 5661 3985 5695
rect 4019 5661 4031 5695
rect 3973 5655 4031 5661
rect 5261 5695 5319 5701
rect 5261 5661 5273 5695
rect 5307 5692 5319 5695
rect 5350 5692 5356 5704
rect 5307 5664 5356 5692
rect 5307 5661 5319 5664
rect 5261 5655 5319 5661
rect 3988 5624 4016 5655
rect 5350 5652 5356 5664
rect 5408 5652 5414 5704
rect 5552 5701 5580 5732
rect 7558 5720 7564 5732
rect 7616 5720 7622 5772
rect 7668 5760 7696 5800
rect 7834 5788 7840 5840
rect 7892 5828 7898 5840
rect 9674 5828 9680 5840
rect 7892 5800 9680 5828
rect 7892 5788 7898 5800
rect 9674 5788 9680 5800
rect 9732 5788 9738 5840
rect 12713 5831 12771 5837
rect 12713 5797 12725 5831
rect 12759 5828 12771 5831
rect 15120 5828 15148 5868
rect 15746 5856 15752 5868
rect 15804 5856 15810 5908
rect 16114 5856 16120 5908
rect 16172 5896 16178 5908
rect 16945 5899 17003 5905
rect 16945 5896 16957 5899
rect 16172 5868 16957 5896
rect 16172 5856 16178 5868
rect 16945 5865 16957 5868
rect 16991 5896 17003 5899
rect 18046 5896 18052 5908
rect 16991 5868 18052 5896
rect 16991 5865 17003 5868
rect 16945 5859 17003 5865
rect 18046 5856 18052 5868
rect 18104 5856 18110 5908
rect 20162 5856 20168 5908
rect 20220 5896 20226 5908
rect 20625 5899 20683 5905
rect 20625 5896 20637 5899
rect 20220 5868 20637 5896
rect 20220 5856 20226 5868
rect 20625 5865 20637 5868
rect 20671 5896 20683 5899
rect 23382 5896 23388 5908
rect 20671 5868 23388 5896
rect 20671 5865 20683 5868
rect 20625 5859 20683 5865
rect 23382 5856 23388 5868
rect 23440 5856 23446 5908
rect 23845 5899 23903 5905
rect 23845 5865 23857 5899
rect 23891 5896 23903 5899
rect 24302 5896 24308 5908
rect 23891 5868 24308 5896
rect 23891 5865 23903 5868
rect 23845 5859 23903 5865
rect 24302 5856 24308 5868
rect 24360 5856 24366 5908
rect 12759 5800 15148 5828
rect 12759 5797 12771 5800
rect 12713 5791 12771 5797
rect 15286 5788 15292 5840
rect 15344 5828 15350 5840
rect 17218 5828 17224 5840
rect 15344 5800 17224 5828
rect 15344 5788 15350 5800
rect 17218 5788 17224 5800
rect 17276 5788 17282 5840
rect 7668 5732 10180 5760
rect 10152 5704 10180 5732
rect 12066 5720 12072 5772
rect 12124 5760 12130 5772
rect 14090 5760 14096 5772
rect 12124 5732 14096 5760
rect 12124 5720 12130 5732
rect 14090 5720 14096 5732
rect 14148 5720 14154 5772
rect 14274 5720 14280 5772
rect 14332 5760 14338 5772
rect 14921 5763 14979 5769
rect 14921 5760 14933 5763
rect 14332 5732 14933 5760
rect 14332 5720 14338 5732
rect 14921 5729 14933 5732
rect 14967 5729 14979 5763
rect 14921 5723 14979 5729
rect 18046 5720 18052 5772
rect 18104 5760 18110 5772
rect 19242 5760 19248 5772
rect 18104 5732 19248 5760
rect 18104 5720 18110 5732
rect 19242 5720 19248 5732
rect 19300 5720 19306 5772
rect 21910 5760 21916 5772
rect 21871 5732 21916 5760
rect 21910 5720 21916 5732
rect 21968 5720 21974 5772
rect 22094 5720 22100 5772
rect 22152 5760 22158 5772
rect 22189 5763 22247 5769
rect 22189 5760 22201 5763
rect 22152 5732 22201 5760
rect 22152 5720 22158 5732
rect 22189 5729 22201 5732
rect 22235 5729 22247 5763
rect 22189 5723 22247 5729
rect 5537 5695 5595 5701
rect 5537 5661 5549 5695
rect 5583 5661 5595 5695
rect 5537 5655 5595 5661
rect 5626 5652 5632 5704
rect 5684 5692 5690 5704
rect 6178 5692 6184 5704
rect 5684 5664 6184 5692
rect 5684 5652 5690 5664
rect 6178 5652 6184 5664
rect 6236 5652 6242 5704
rect 6362 5692 6368 5704
rect 6323 5664 6368 5692
rect 6362 5652 6368 5664
rect 6420 5652 6426 5704
rect 6457 5695 6515 5701
rect 6457 5661 6469 5695
rect 6503 5661 6515 5695
rect 6457 5655 6515 5661
rect 6549 5695 6607 5701
rect 6549 5661 6561 5695
rect 6595 5692 6607 5695
rect 6730 5692 6736 5704
rect 6595 5664 6736 5692
rect 6595 5661 6607 5664
rect 6549 5655 6607 5661
rect 6270 5624 6276 5636
rect 3988 5596 6276 5624
rect 6270 5584 6276 5596
rect 6328 5584 6334 5636
rect 6472 5624 6500 5655
rect 6730 5652 6736 5664
rect 6788 5652 6794 5704
rect 7926 5692 7932 5704
rect 7887 5664 7932 5692
rect 7926 5652 7932 5664
rect 7984 5652 7990 5704
rect 9674 5692 9680 5704
rect 9635 5664 9680 5692
rect 9674 5652 9680 5664
rect 9732 5652 9738 5704
rect 10134 5692 10140 5704
rect 10095 5664 10140 5692
rect 10134 5652 10140 5664
rect 10192 5652 10198 5704
rect 10778 5692 10784 5704
rect 10691 5664 10784 5692
rect 10778 5652 10784 5664
rect 10836 5692 10842 5704
rect 12894 5692 12900 5704
rect 10836 5664 12900 5692
rect 10836 5652 10842 5664
rect 12894 5652 12900 5664
rect 12952 5652 12958 5704
rect 12986 5652 12992 5704
rect 13044 5692 13050 5704
rect 13173 5695 13231 5701
rect 13173 5692 13185 5695
rect 13044 5664 13185 5692
rect 13044 5652 13050 5664
rect 13173 5661 13185 5664
rect 13219 5661 13231 5695
rect 14182 5692 14188 5704
rect 14143 5664 14188 5692
rect 13173 5655 13231 5661
rect 14182 5652 14188 5664
rect 14240 5652 14246 5704
rect 14829 5695 14887 5701
rect 14829 5661 14841 5695
rect 14875 5661 14887 5695
rect 15654 5692 15660 5704
rect 15615 5664 15660 5692
rect 14829 5655 14887 5661
rect 6638 5624 6644 5636
rect 6472 5596 6644 5624
rect 6638 5584 6644 5596
rect 6696 5584 6702 5636
rect 11054 5633 11060 5636
rect 11048 5624 11060 5633
rect 11015 5596 11060 5624
rect 11048 5587 11060 5596
rect 11054 5584 11060 5587
rect 11112 5584 11118 5636
rect 12066 5624 12072 5636
rect 11532 5596 12072 5624
rect 5721 5559 5779 5565
rect 5721 5525 5733 5559
rect 5767 5556 5779 5559
rect 6546 5556 6552 5568
rect 5767 5528 6552 5556
rect 5767 5525 5779 5528
rect 5721 5519 5779 5525
rect 6546 5516 6552 5528
rect 6604 5516 6610 5568
rect 6825 5559 6883 5565
rect 6825 5525 6837 5559
rect 6871 5556 6883 5559
rect 7282 5556 7288 5568
rect 6871 5528 7288 5556
rect 6871 5525 6883 5528
rect 6825 5519 6883 5525
rect 7282 5516 7288 5528
rect 7340 5516 7346 5568
rect 10321 5559 10379 5565
rect 10321 5525 10333 5559
rect 10367 5556 10379 5559
rect 11532 5556 11560 5596
rect 12066 5584 12072 5596
rect 12124 5584 12130 5636
rect 10367 5528 11560 5556
rect 10367 5525 10379 5528
rect 10321 5519 10379 5525
rect 11606 5516 11612 5568
rect 11664 5556 11670 5568
rect 12161 5559 12219 5565
rect 12161 5556 12173 5559
rect 11664 5528 12173 5556
rect 11664 5516 11670 5528
rect 12161 5525 12173 5528
rect 12207 5525 12219 5559
rect 12161 5519 12219 5525
rect 13078 5516 13084 5568
rect 13136 5556 13142 5568
rect 13357 5559 13415 5565
rect 13357 5556 13369 5559
rect 13136 5528 13369 5556
rect 13136 5516 13142 5528
rect 13357 5525 13369 5528
rect 13403 5525 13415 5559
rect 13357 5519 13415 5525
rect 13722 5516 13728 5568
rect 13780 5556 13786 5568
rect 14369 5559 14427 5565
rect 14369 5556 14381 5559
rect 13780 5528 14381 5556
rect 13780 5516 13786 5528
rect 14369 5525 14381 5528
rect 14415 5556 14427 5559
rect 14844 5556 14872 5655
rect 15654 5652 15660 5664
rect 15712 5652 15718 5704
rect 17678 5652 17684 5704
rect 17736 5692 17742 5704
rect 17865 5695 17923 5701
rect 17865 5692 17877 5695
rect 17736 5664 17877 5692
rect 17736 5652 17742 5664
rect 17865 5661 17877 5664
rect 17911 5661 17923 5695
rect 17865 5655 17923 5661
rect 18509 5695 18567 5701
rect 18509 5661 18521 5695
rect 18555 5692 18567 5695
rect 19334 5692 19340 5704
rect 18555 5664 19340 5692
rect 18555 5661 18567 5664
rect 18509 5655 18567 5661
rect 19334 5652 19340 5664
rect 19392 5652 19398 5704
rect 20806 5692 20812 5704
rect 19444 5664 20812 5692
rect 19444 5624 19472 5664
rect 20806 5652 20812 5664
rect 20864 5652 20870 5704
rect 21174 5652 21180 5704
rect 21232 5692 21238 5704
rect 21269 5695 21327 5701
rect 21269 5692 21281 5695
rect 21232 5664 21281 5692
rect 21232 5652 21238 5664
rect 21269 5661 21281 5664
rect 21315 5661 21327 5695
rect 21269 5655 21327 5661
rect 18064 5596 19472 5624
rect 19512 5627 19570 5633
rect 14415 5528 14872 5556
rect 15197 5559 15255 5565
rect 14415 5525 14427 5528
rect 14369 5519 14427 5525
rect 15197 5525 15209 5559
rect 15243 5556 15255 5559
rect 15838 5556 15844 5568
rect 15243 5528 15844 5556
rect 15243 5525 15255 5528
rect 15197 5519 15255 5525
rect 15838 5516 15844 5528
rect 15896 5516 15902 5568
rect 18064 5565 18092 5596
rect 19512 5593 19524 5627
rect 19558 5624 19570 5627
rect 20254 5624 20260 5636
rect 19558 5596 20260 5624
rect 19558 5593 19570 5596
rect 19512 5587 19570 5593
rect 20254 5584 20260 5596
rect 20312 5584 20318 5636
rect 18049 5559 18107 5565
rect 18049 5525 18061 5559
rect 18095 5525 18107 5559
rect 18049 5519 18107 5525
rect 18693 5559 18751 5565
rect 18693 5525 18705 5559
rect 18739 5556 18751 5559
rect 20438 5556 20444 5568
rect 18739 5528 20444 5556
rect 18739 5525 18751 5528
rect 18693 5519 18751 5525
rect 20438 5516 20444 5528
rect 20496 5516 20502 5568
rect 23198 5556 23204 5568
rect 23159 5528 23204 5556
rect 23198 5516 23204 5528
rect 23256 5516 23262 5568
rect 1104 5466 68816 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 50294 5466
rect 50346 5414 50358 5466
rect 50410 5414 50422 5466
rect 50474 5414 50486 5466
rect 50538 5414 50550 5466
rect 50602 5414 68816 5466
rect 1104 5392 68816 5414
rect 4525 5355 4583 5361
rect 4525 5321 4537 5355
rect 4571 5352 4583 5355
rect 4798 5352 4804 5364
rect 4571 5324 4804 5352
rect 4571 5321 4583 5324
rect 4525 5315 4583 5321
rect 4798 5312 4804 5324
rect 4856 5352 4862 5364
rect 4856 5324 9720 5352
rect 4856 5312 4862 5324
rect 3513 5219 3571 5225
rect 3513 5185 3525 5219
rect 3559 5216 3571 5219
rect 3786 5216 3792 5228
rect 3559 5188 3792 5216
rect 3559 5185 3571 5188
rect 3513 5179 3571 5185
rect 3786 5176 3792 5188
rect 3844 5176 3850 5228
rect 5828 5225 5856 5324
rect 9582 5284 9588 5296
rect 9543 5256 9588 5284
rect 9582 5244 9588 5256
rect 9640 5244 9646 5296
rect 9692 5284 9720 5324
rect 10042 5312 10048 5364
rect 10100 5352 10106 5364
rect 10505 5355 10563 5361
rect 10505 5352 10517 5355
rect 10100 5324 10517 5352
rect 10100 5312 10106 5324
rect 10505 5321 10517 5324
rect 10551 5321 10563 5355
rect 11790 5352 11796 5364
rect 10505 5315 10563 5321
rect 10612 5324 11796 5352
rect 10612 5284 10640 5324
rect 11790 5312 11796 5324
rect 11848 5312 11854 5364
rect 12158 5312 12164 5364
rect 12216 5352 12222 5364
rect 14918 5352 14924 5364
rect 12216 5324 14924 5352
rect 12216 5312 12222 5324
rect 14918 5312 14924 5324
rect 14976 5312 14982 5364
rect 15749 5355 15807 5361
rect 15749 5321 15761 5355
rect 15795 5352 15807 5355
rect 16390 5352 16396 5364
rect 15795 5324 16396 5352
rect 15795 5321 15807 5324
rect 15749 5315 15807 5321
rect 16390 5312 16396 5324
rect 16448 5312 16454 5364
rect 16666 5352 16672 5364
rect 16627 5324 16672 5352
rect 16666 5312 16672 5324
rect 16724 5312 16730 5364
rect 19613 5355 19671 5361
rect 19613 5321 19625 5355
rect 19659 5352 19671 5355
rect 20622 5352 20628 5364
rect 19659 5324 20628 5352
rect 19659 5321 19671 5324
rect 19613 5315 19671 5321
rect 20622 5312 20628 5324
rect 20680 5312 20686 5364
rect 20993 5355 21051 5361
rect 20993 5321 21005 5355
rect 21039 5352 21051 5355
rect 21082 5352 21088 5364
rect 21039 5324 21088 5352
rect 21039 5321 21051 5324
rect 20993 5315 21051 5321
rect 21082 5312 21088 5324
rect 21140 5312 21146 5364
rect 23658 5312 23664 5364
rect 23716 5352 23722 5364
rect 23716 5324 23888 5352
rect 23716 5312 23722 5324
rect 9692 5256 10640 5284
rect 12066 5244 12072 5296
rect 12124 5284 12130 5296
rect 14550 5284 14556 5296
rect 12124 5256 14556 5284
rect 12124 5244 12130 5256
rect 14550 5244 14556 5256
rect 14608 5284 14614 5296
rect 15289 5287 15347 5293
rect 15289 5284 15301 5287
rect 14608 5256 15301 5284
rect 14608 5244 14614 5256
rect 15289 5253 15301 5256
rect 15335 5253 15347 5287
rect 15289 5247 15347 5253
rect 17804 5287 17862 5293
rect 17804 5253 17816 5287
rect 17850 5284 17862 5287
rect 20714 5284 20720 5296
rect 17850 5256 20720 5284
rect 17850 5253 17862 5256
rect 17804 5247 17862 5253
rect 20714 5244 20720 5256
rect 20772 5244 20778 5296
rect 23290 5244 23296 5296
rect 23348 5284 23354 5296
rect 23860 5284 23888 5324
rect 23348 5256 23704 5284
rect 23860 5256 23980 5284
rect 23348 5244 23354 5256
rect 5813 5219 5871 5225
rect 5813 5185 5825 5219
rect 5859 5185 5871 5219
rect 5813 5179 5871 5185
rect 6178 5176 6184 5228
rect 6236 5216 6242 5228
rect 6365 5219 6423 5225
rect 6365 5216 6377 5219
rect 6236 5188 6377 5216
rect 6236 5176 6242 5188
rect 6365 5185 6377 5188
rect 6411 5185 6423 5219
rect 6546 5216 6552 5228
rect 6507 5188 6552 5216
rect 6365 5179 6423 5185
rect 6546 5176 6552 5188
rect 6604 5176 6610 5228
rect 6641 5219 6699 5225
rect 6641 5185 6653 5219
rect 6687 5185 6699 5219
rect 6641 5179 6699 5185
rect 6733 5219 6791 5225
rect 6733 5185 6745 5219
rect 6779 5216 6791 5219
rect 6914 5216 6920 5228
rect 6779 5188 6920 5216
rect 6779 5185 6791 5188
rect 6733 5179 6791 5185
rect 3605 5151 3663 5157
rect 3605 5117 3617 5151
rect 3651 5148 3663 5151
rect 5166 5148 5172 5160
rect 3651 5120 5172 5148
rect 3651 5117 3663 5120
rect 3605 5111 3663 5117
rect 5166 5108 5172 5120
rect 5224 5108 5230 5160
rect 5537 5151 5595 5157
rect 5537 5117 5549 5151
rect 5583 5117 5595 5151
rect 5537 5111 5595 5117
rect 3881 5083 3939 5089
rect 3881 5049 3893 5083
rect 3927 5080 3939 5083
rect 4982 5080 4988 5092
rect 3927 5052 4988 5080
rect 3927 5049 3939 5052
rect 3881 5043 3939 5049
rect 4982 5040 4988 5052
rect 5040 5040 5046 5092
rect 3697 5015 3755 5021
rect 3697 4981 3709 5015
rect 3743 5012 3755 5015
rect 3970 5012 3976 5024
rect 3743 4984 3976 5012
rect 3743 4981 3755 4984
rect 3697 4975 3755 4981
rect 3970 4972 3976 4984
rect 4028 4972 4034 5024
rect 5166 4972 5172 5024
rect 5224 5012 5230 5024
rect 5552 5012 5580 5111
rect 6656 5092 6684 5179
rect 6914 5176 6920 5188
rect 6972 5176 6978 5228
rect 8386 5176 8392 5228
rect 8444 5216 8450 5228
rect 10045 5219 10103 5225
rect 10045 5216 10057 5219
rect 8444 5188 10057 5216
rect 8444 5176 8450 5188
rect 10045 5185 10057 5188
rect 10091 5185 10103 5219
rect 10045 5179 10103 5185
rect 10321 5219 10379 5225
rect 10321 5185 10333 5219
rect 10367 5216 10379 5219
rect 10410 5216 10416 5228
rect 10367 5188 10416 5216
rect 10367 5185 10379 5188
rect 10321 5179 10379 5185
rect 10410 5176 10416 5188
rect 10468 5176 10474 5228
rect 11698 5216 11704 5228
rect 11659 5188 11704 5216
rect 11698 5176 11704 5188
rect 11756 5176 11762 5228
rect 12802 5216 12808 5228
rect 12763 5188 12808 5216
rect 12802 5176 12808 5188
rect 12860 5176 12866 5228
rect 12897 5219 12955 5225
rect 12897 5185 12909 5219
rect 12943 5185 12955 5219
rect 12897 5179 12955 5185
rect 6932 5148 6960 5176
rect 10137 5151 10195 5157
rect 10137 5148 10149 5151
rect 6932 5120 10149 5148
rect 10137 5117 10149 5120
rect 10183 5117 10195 5151
rect 10428 5148 10456 5176
rect 11793 5151 11851 5157
rect 11793 5148 11805 5151
rect 10428 5120 11805 5148
rect 10137 5111 10195 5117
rect 11793 5117 11805 5120
rect 11839 5117 11851 5151
rect 11793 5111 11851 5117
rect 12434 5108 12440 5160
rect 12492 5148 12498 5160
rect 12912 5148 12940 5179
rect 12986 5176 12992 5228
rect 13044 5216 13050 5228
rect 13173 5219 13231 5225
rect 13044 5188 13089 5216
rect 13044 5176 13050 5188
rect 13173 5185 13185 5219
rect 13219 5185 13231 5219
rect 13630 5216 13636 5228
rect 13591 5188 13636 5216
rect 13173 5179 13231 5185
rect 12492 5120 12940 5148
rect 13188 5148 13216 5179
rect 13630 5176 13636 5188
rect 13688 5176 13694 5228
rect 15562 5216 15568 5228
rect 15523 5188 15568 5216
rect 15562 5176 15568 5188
rect 15620 5176 15626 5228
rect 18046 5216 18052 5228
rect 18007 5188 18052 5216
rect 18046 5176 18052 5188
rect 18104 5176 18110 5228
rect 19426 5176 19432 5228
rect 19484 5216 19490 5228
rect 19797 5219 19855 5225
rect 19797 5216 19809 5219
rect 19484 5188 19809 5216
rect 19484 5176 19490 5188
rect 19797 5185 19809 5188
rect 19843 5185 19855 5219
rect 20073 5219 20131 5225
rect 20073 5216 20085 5219
rect 19797 5179 19855 5185
rect 19904 5188 20085 5216
rect 13538 5148 13544 5160
rect 13188 5120 13544 5148
rect 12492 5108 12498 5120
rect 13538 5108 13544 5120
rect 13596 5148 13602 5160
rect 13909 5151 13967 5157
rect 13909 5148 13921 5151
rect 13596 5120 13921 5148
rect 13596 5108 13602 5120
rect 13909 5117 13921 5120
rect 13955 5117 13967 5151
rect 15470 5148 15476 5160
rect 15431 5120 15476 5148
rect 13909 5111 13967 5117
rect 15470 5108 15476 5120
rect 15528 5108 15534 5160
rect 6638 5040 6644 5092
rect 6696 5040 6702 5092
rect 9858 5040 9864 5092
rect 9916 5080 9922 5092
rect 12158 5080 12164 5092
rect 9916 5052 12164 5080
rect 9916 5040 9922 5052
rect 5224 4984 5580 5012
rect 5224 4972 5230 4984
rect 6822 4972 6828 5024
rect 6880 5012 6886 5024
rect 7009 5015 7067 5021
rect 7009 5012 7021 5015
rect 6880 4984 7021 5012
rect 6880 4972 6886 4984
rect 7009 4981 7021 4984
rect 7055 4981 7067 5015
rect 8294 5012 8300 5024
rect 8255 4984 8300 5012
rect 7009 4975 7067 4981
rect 8294 4972 8300 4984
rect 8352 4972 8358 5024
rect 10318 5012 10324 5024
rect 10279 4984 10324 5012
rect 10318 4972 10324 4984
rect 10376 5012 10382 5024
rect 11606 5012 11612 5024
rect 10376 4984 11612 5012
rect 10376 4972 10382 4984
rect 11606 4972 11612 4984
rect 11664 4972 11670 5024
rect 11716 5021 11744 5052
rect 12158 5040 12164 5052
rect 12216 5040 12222 5092
rect 19153 5083 19211 5089
rect 19153 5049 19165 5083
rect 19199 5080 19211 5083
rect 19702 5080 19708 5092
rect 19199 5052 19708 5080
rect 19199 5049 19211 5052
rect 19153 5043 19211 5049
rect 19702 5040 19708 5052
rect 19760 5040 19766 5092
rect 11701 5015 11759 5021
rect 11701 4981 11713 5015
rect 11747 4981 11759 5015
rect 11701 4975 11759 4981
rect 12069 5015 12127 5021
rect 12069 4981 12081 5015
rect 12115 5012 12127 5015
rect 12250 5012 12256 5024
rect 12115 4984 12256 5012
rect 12115 4981 12127 4984
rect 12069 4975 12127 4981
rect 12250 4972 12256 4984
rect 12308 4972 12314 5024
rect 12526 5012 12532 5024
rect 12487 4984 12532 5012
rect 12526 4972 12532 4984
rect 12584 4972 12590 5024
rect 15286 5012 15292 5024
rect 15247 4984 15292 5012
rect 15286 4972 15292 4984
rect 15344 4972 15350 5024
rect 19058 4972 19064 5024
rect 19116 5012 19122 5024
rect 19242 5012 19248 5024
rect 19116 4984 19248 5012
rect 19116 4972 19122 4984
rect 19242 4972 19248 4984
rect 19300 4972 19306 5024
rect 19794 4972 19800 5024
rect 19852 5012 19858 5024
rect 19904 5012 19932 5188
rect 20073 5185 20085 5188
rect 20119 5216 20131 5219
rect 20533 5219 20591 5225
rect 20533 5216 20545 5219
rect 20119 5188 20545 5216
rect 20119 5185 20131 5188
rect 20073 5179 20131 5185
rect 20533 5185 20545 5188
rect 20579 5216 20591 5219
rect 20579 5188 20760 5216
rect 20579 5185 20591 5188
rect 20533 5179 20591 5185
rect 19981 5151 20039 5157
rect 19981 5117 19993 5151
rect 20027 5148 20039 5151
rect 20438 5148 20444 5160
rect 20027 5120 20444 5148
rect 20027 5117 20039 5120
rect 19981 5111 20039 5117
rect 20438 5108 20444 5120
rect 20496 5148 20502 5160
rect 20625 5151 20683 5157
rect 20625 5148 20637 5151
rect 20496 5120 20637 5148
rect 20496 5108 20502 5120
rect 20625 5117 20637 5120
rect 20671 5117 20683 5151
rect 20732 5148 20760 5188
rect 20806 5176 20812 5228
rect 20864 5216 20870 5228
rect 21450 5216 21456 5228
rect 20864 5188 20909 5216
rect 21008 5188 21456 5216
rect 20864 5176 20870 5188
rect 21008 5148 21036 5188
rect 21450 5176 21456 5188
rect 21508 5176 21514 5228
rect 21542 5176 21548 5228
rect 21600 5216 21606 5228
rect 22005 5219 22063 5225
rect 22005 5216 22017 5219
rect 21600 5188 22017 5216
rect 21600 5176 21606 5188
rect 22005 5185 22017 5188
rect 22051 5216 22063 5219
rect 22051 5188 22692 5216
rect 22051 5185 22063 5188
rect 22005 5179 22063 5185
rect 20732 5120 21036 5148
rect 22664 5148 22692 5188
rect 22830 5176 22836 5228
rect 22888 5216 22894 5228
rect 23676 5225 23704 5256
rect 23569 5219 23627 5225
rect 23569 5216 23581 5219
rect 22888 5188 23581 5216
rect 22888 5176 22894 5188
rect 23569 5185 23581 5188
rect 23615 5185 23627 5219
rect 23569 5179 23627 5185
rect 23661 5219 23719 5225
rect 23661 5185 23673 5219
rect 23707 5185 23719 5219
rect 23661 5179 23719 5185
rect 23750 5176 23756 5228
rect 23808 5216 23814 5228
rect 23952 5225 23980 5256
rect 23937 5219 23995 5225
rect 23808 5188 23853 5216
rect 23808 5176 23814 5188
rect 23937 5185 23949 5219
rect 23983 5185 23995 5219
rect 23937 5179 23995 5185
rect 24397 5151 24455 5157
rect 24397 5148 24409 5151
rect 22664 5120 24409 5148
rect 20625 5111 20683 5117
rect 24397 5117 24409 5120
rect 24443 5117 24455 5151
rect 24397 5111 24455 5117
rect 20714 5040 20720 5092
rect 20772 5080 20778 5092
rect 23293 5083 23351 5089
rect 23293 5080 23305 5083
rect 20772 5052 23305 5080
rect 20772 5040 20778 5052
rect 23293 5049 23305 5052
rect 23339 5049 23351 5083
rect 23293 5043 23351 5049
rect 19852 4984 19932 5012
rect 20073 5015 20131 5021
rect 19852 4972 19858 4984
rect 20073 4981 20085 5015
rect 20119 5012 20131 5015
rect 20809 5015 20867 5021
rect 20809 5012 20821 5015
rect 20119 4984 20821 5012
rect 20119 4981 20131 4984
rect 20073 4975 20131 4981
rect 20809 4981 20821 4984
rect 20855 5012 20867 5015
rect 21266 5012 21272 5024
rect 20855 4984 21272 5012
rect 20855 4981 20867 4984
rect 20809 4975 20867 4981
rect 21266 4972 21272 4984
rect 21324 4972 21330 5024
rect 21818 5012 21824 5024
rect 21779 4984 21824 5012
rect 21818 4972 21824 4984
rect 21876 4972 21882 5024
rect 22278 4972 22284 5024
rect 22336 5012 22342 5024
rect 22465 5015 22523 5021
rect 22465 5012 22477 5015
rect 22336 4984 22477 5012
rect 22336 4972 22342 4984
rect 22465 4981 22477 4984
rect 22511 4981 22523 5015
rect 22465 4975 22523 4981
rect 1104 4922 68816 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 65654 4922
rect 65706 4870 65718 4922
rect 65770 4870 65782 4922
rect 65834 4870 65846 4922
rect 65898 4870 65910 4922
rect 65962 4870 68816 4922
rect 1104 4848 68816 4870
rect 3970 4808 3976 4820
rect 3931 4780 3976 4808
rect 3970 4768 3976 4780
rect 4028 4768 4034 4820
rect 4614 4768 4620 4820
rect 4672 4808 4678 4820
rect 4893 4811 4951 4817
rect 4893 4808 4905 4811
rect 4672 4780 4905 4808
rect 4672 4768 4678 4780
rect 4893 4777 4905 4780
rect 4939 4777 4951 4811
rect 5718 4808 5724 4820
rect 5679 4780 5724 4808
rect 4893 4771 4951 4777
rect 5718 4768 5724 4780
rect 5776 4768 5782 4820
rect 5905 4811 5963 4817
rect 5905 4777 5917 4811
rect 5951 4808 5963 4811
rect 6362 4808 6368 4820
rect 5951 4780 6368 4808
rect 5951 4777 5963 4780
rect 5905 4771 5963 4777
rect 6362 4768 6368 4780
rect 6420 4768 6426 4820
rect 8386 4808 8392 4820
rect 6748 4780 8392 4808
rect 6748 4752 6776 4780
rect 8386 4768 8392 4780
rect 8444 4768 8450 4820
rect 9677 4811 9735 4817
rect 9677 4777 9689 4811
rect 9723 4808 9735 4811
rect 12066 4808 12072 4820
rect 9723 4780 12072 4808
rect 9723 4777 9735 4780
rect 9677 4771 9735 4777
rect 12066 4768 12072 4780
rect 12124 4768 12130 4820
rect 12158 4768 12164 4820
rect 12216 4808 12222 4820
rect 12345 4811 12403 4817
rect 12345 4808 12357 4811
rect 12216 4780 12357 4808
rect 12216 4768 12222 4780
rect 12345 4777 12357 4780
rect 12391 4777 12403 4811
rect 12345 4771 12403 4777
rect 12713 4811 12771 4817
rect 12713 4777 12725 4811
rect 12759 4808 12771 4811
rect 12986 4808 12992 4820
rect 12759 4780 12992 4808
rect 12759 4777 12771 4780
rect 12713 4771 12771 4777
rect 12986 4768 12992 4780
rect 13044 4768 13050 4820
rect 14090 4768 14096 4820
rect 14148 4808 14154 4820
rect 14553 4811 14611 4817
rect 14553 4808 14565 4811
rect 14148 4780 14565 4808
rect 14148 4768 14154 4780
rect 14553 4777 14565 4780
rect 14599 4808 14611 4811
rect 15286 4808 15292 4820
rect 14599 4780 15292 4808
rect 14599 4777 14611 4780
rect 14553 4771 14611 4777
rect 15286 4768 15292 4780
rect 15344 4808 15350 4820
rect 15473 4811 15531 4817
rect 15473 4808 15485 4811
rect 15344 4780 15485 4808
rect 15344 4768 15350 4780
rect 15473 4777 15485 4780
rect 15519 4777 15531 4811
rect 15930 4808 15936 4820
rect 15891 4780 15936 4808
rect 15473 4771 15531 4777
rect 6730 4740 6736 4752
rect 3896 4712 6736 4740
rect 3896 4681 3924 4712
rect 6730 4700 6736 4712
rect 6788 4700 6794 4752
rect 15488 4740 15516 4771
rect 15930 4768 15936 4780
rect 15988 4768 15994 4820
rect 16393 4811 16451 4817
rect 16393 4777 16405 4811
rect 16439 4777 16451 4811
rect 16393 4771 16451 4777
rect 16853 4811 16911 4817
rect 16853 4777 16865 4811
rect 16899 4808 16911 4811
rect 17126 4808 17132 4820
rect 16899 4780 17132 4808
rect 16899 4777 16911 4780
rect 16853 4771 16911 4777
rect 16408 4740 16436 4771
rect 17126 4768 17132 4780
rect 17184 4768 17190 4820
rect 17313 4811 17371 4817
rect 17313 4777 17325 4811
rect 17359 4777 17371 4811
rect 17770 4808 17776 4820
rect 17731 4780 17776 4808
rect 17313 4771 17371 4777
rect 17328 4740 17356 4771
rect 17770 4768 17776 4780
rect 17828 4768 17834 4820
rect 18782 4768 18788 4820
rect 18840 4808 18846 4820
rect 19150 4808 19156 4820
rect 18840 4780 19156 4808
rect 18840 4768 18846 4780
rect 19150 4768 19156 4780
rect 19208 4768 19214 4820
rect 20257 4811 20315 4817
rect 20257 4808 20269 4811
rect 19306 4780 20269 4808
rect 15488 4712 17356 4740
rect 3881 4675 3939 4681
rect 3881 4641 3893 4675
rect 3927 4641 3939 4675
rect 5534 4672 5540 4684
rect 5495 4644 5540 4672
rect 3881 4635 3939 4641
rect 5534 4632 5540 4644
rect 5592 4632 5598 4684
rect 11606 4632 11612 4684
rect 11664 4672 11670 4684
rect 12437 4675 12495 4681
rect 12437 4672 12449 4675
rect 11664 4644 12449 4672
rect 11664 4632 11670 4644
rect 12437 4641 12449 4644
rect 12483 4641 12495 4675
rect 13722 4672 13728 4684
rect 12437 4635 12495 4641
rect 13096 4644 13728 4672
rect 3786 4604 3792 4616
rect 3747 4576 3792 4604
rect 3786 4564 3792 4576
rect 3844 4564 3850 4616
rect 4801 4607 4859 4613
rect 4801 4573 4813 4607
rect 4847 4604 4859 4607
rect 4890 4604 4896 4616
rect 4847 4576 4896 4604
rect 4847 4573 4859 4576
rect 4801 4567 4859 4573
rect 4890 4564 4896 4576
rect 4948 4564 4954 4616
rect 5350 4564 5356 4616
rect 5408 4604 5414 4616
rect 5445 4607 5503 4613
rect 5445 4604 5457 4607
rect 5408 4576 5457 4604
rect 5408 4564 5414 4576
rect 5445 4573 5457 4576
rect 5491 4573 5503 4607
rect 5718 4604 5724 4616
rect 5679 4576 5724 4604
rect 5445 4567 5503 4573
rect 5718 4564 5724 4576
rect 5776 4564 5782 4616
rect 6546 4604 6552 4616
rect 6507 4576 6552 4604
rect 6546 4564 6552 4576
rect 6604 4564 6610 4616
rect 7009 4607 7067 4613
rect 7009 4573 7021 4607
rect 7055 4604 7067 4607
rect 8294 4604 8300 4616
rect 7055 4576 8300 4604
rect 7055 4573 7067 4576
rect 7009 4567 7067 4573
rect 8294 4564 8300 4576
rect 8352 4564 8358 4616
rect 9490 4604 9496 4616
rect 9451 4576 9496 4604
rect 9490 4564 9496 4576
rect 9548 4564 9554 4616
rect 9582 4564 9588 4616
rect 9640 4604 9646 4616
rect 10137 4607 10195 4613
rect 10137 4604 10149 4607
rect 9640 4576 10149 4604
rect 9640 4564 9646 4576
rect 10137 4573 10149 4576
rect 10183 4604 10195 4607
rect 10778 4604 10784 4616
rect 10183 4576 10784 4604
rect 10183 4573 10195 4576
rect 10137 4567 10195 4573
rect 10778 4564 10784 4576
rect 10836 4564 10842 4616
rect 11698 4564 11704 4616
rect 11756 4604 11762 4616
rect 12345 4607 12403 4613
rect 12345 4604 12357 4607
rect 11756 4576 12357 4604
rect 11756 4564 11762 4576
rect 12345 4573 12357 4576
rect 12391 4604 12403 4607
rect 13096 4604 13124 4644
rect 13722 4632 13728 4644
rect 13780 4632 13786 4684
rect 14737 4675 14795 4681
rect 14737 4641 14749 4675
rect 14783 4672 14795 4675
rect 15470 4672 15476 4684
rect 14783 4644 15476 4672
rect 14783 4641 14795 4644
rect 14737 4635 14795 4641
rect 15470 4632 15476 4644
rect 15528 4672 15534 4684
rect 15657 4675 15715 4681
rect 15657 4672 15669 4675
rect 15528 4644 15669 4672
rect 15528 4632 15534 4644
rect 15657 4641 15669 4644
rect 15703 4672 15715 4675
rect 17497 4675 17555 4681
rect 17497 4672 17509 4675
rect 15703 4644 16620 4672
rect 15703 4641 15715 4644
rect 15657 4635 15715 4641
rect 13262 4604 13268 4616
rect 12391 4576 13124 4604
rect 13223 4576 13268 4604
rect 12391 4573 12403 4576
rect 12345 4567 12403 4573
rect 13262 4564 13268 4576
rect 13320 4564 13326 4616
rect 14550 4604 14556 4616
rect 14511 4576 14556 4604
rect 14550 4564 14556 4576
rect 14608 4564 14614 4616
rect 14829 4607 14887 4613
rect 14829 4573 14841 4607
rect 14875 4604 14887 4607
rect 15194 4604 15200 4616
rect 14875 4576 15200 4604
rect 14875 4573 14887 4576
rect 14829 4567 14887 4573
rect 15194 4564 15200 4576
rect 15252 4564 15258 4616
rect 15749 4607 15807 4613
rect 15749 4573 15761 4607
rect 15795 4604 15807 4607
rect 16482 4604 16488 4616
rect 15795 4576 16488 4604
rect 15795 4573 15807 4576
rect 15749 4567 15807 4573
rect 16482 4564 16488 4576
rect 16540 4564 16546 4616
rect 16592 4613 16620 4644
rect 16776 4644 17509 4672
rect 16577 4607 16635 4613
rect 16577 4573 16589 4607
rect 16623 4573 16635 4607
rect 16577 4567 16635 4573
rect 7282 4545 7288 4548
rect 7276 4536 7288 4545
rect 7243 4508 7288 4536
rect 7276 4499 7288 4508
rect 7282 4496 7288 4499
rect 7340 4496 7346 4548
rect 10404 4539 10462 4545
rect 10404 4505 10416 4539
rect 10450 4536 10462 4539
rect 12526 4536 12532 4548
rect 10450 4508 12532 4536
rect 10450 4505 10462 4508
rect 10404 4499 10462 4505
rect 12526 4496 12532 4508
rect 12584 4496 12590 4548
rect 14568 4536 14596 4564
rect 15473 4539 15531 4545
rect 15473 4536 15485 4539
rect 14568 4508 15485 4536
rect 15473 4505 15485 4508
rect 15519 4536 15531 4539
rect 16393 4539 16451 4545
rect 16393 4536 16405 4539
rect 15519 4508 16405 4536
rect 15519 4505 15531 4508
rect 15473 4499 15531 4505
rect 16393 4505 16405 4508
rect 16439 4505 16451 4539
rect 16592 4536 16620 4567
rect 16666 4564 16672 4616
rect 16724 4613 16730 4616
rect 16724 4607 16743 4613
rect 16731 4573 16743 4607
rect 16724 4567 16743 4573
rect 16724 4564 16730 4567
rect 16776 4536 16804 4644
rect 17497 4641 17509 4644
rect 17543 4672 17555 4675
rect 19306 4672 19334 4780
rect 20257 4777 20269 4780
rect 20303 4777 20315 4811
rect 20898 4808 20904 4820
rect 20859 4780 20904 4808
rect 20257 4771 20315 4777
rect 20898 4768 20904 4780
rect 20956 4768 20962 4820
rect 21266 4808 21272 4820
rect 21179 4780 21272 4808
rect 21266 4768 21272 4780
rect 21324 4808 21330 4820
rect 21910 4808 21916 4820
rect 21324 4780 21916 4808
rect 21324 4768 21330 4780
rect 21910 4768 21916 4780
rect 21968 4768 21974 4820
rect 19797 4743 19855 4749
rect 19797 4709 19809 4743
rect 19843 4740 19855 4743
rect 21358 4740 21364 4752
rect 19843 4712 21364 4740
rect 19843 4709 19855 4712
rect 19797 4703 19855 4709
rect 21358 4700 21364 4712
rect 21416 4700 21422 4752
rect 21634 4700 21640 4752
rect 21692 4740 21698 4752
rect 22281 4743 22339 4749
rect 22281 4740 22293 4743
rect 21692 4712 22293 4740
rect 21692 4700 21698 4712
rect 22281 4709 22293 4712
rect 22327 4709 22339 4743
rect 22281 4703 22339 4709
rect 23290 4700 23296 4752
rect 23348 4700 23354 4752
rect 17543 4644 19334 4672
rect 17543 4641 17555 4644
rect 17497 4635 17555 4641
rect 20530 4632 20536 4684
rect 20588 4672 20594 4684
rect 21177 4675 21235 4681
rect 21177 4672 21189 4675
rect 20588 4644 21189 4672
rect 20588 4632 20594 4644
rect 21177 4641 21189 4644
rect 21223 4672 21235 4675
rect 21913 4675 21971 4681
rect 21913 4672 21925 4675
rect 21223 4644 21925 4672
rect 21223 4641 21235 4644
rect 21177 4635 21235 4641
rect 21913 4641 21925 4644
rect 21959 4641 21971 4675
rect 23308 4672 23336 4700
rect 23308 4644 23428 4672
rect 21913 4635 21971 4641
rect 17586 4604 17592 4616
rect 17547 4576 17592 4604
rect 17586 4564 17592 4576
rect 17644 4564 17650 4616
rect 18414 4564 18420 4616
rect 18472 4604 18478 4616
rect 18509 4607 18567 4613
rect 18509 4604 18521 4607
rect 18472 4576 18521 4604
rect 18472 4564 18478 4576
rect 18509 4573 18521 4576
rect 18555 4573 18567 4607
rect 19610 4604 19616 4616
rect 19571 4576 19616 4604
rect 18509 4567 18567 4573
rect 19610 4564 19616 4576
rect 19668 4564 19674 4616
rect 20441 4607 20499 4613
rect 20441 4573 20453 4607
rect 20487 4604 20499 4607
rect 20622 4604 20628 4616
rect 20487 4576 20628 4604
rect 20487 4573 20499 4576
rect 20441 4567 20499 4573
rect 20622 4564 20628 4576
rect 20680 4564 20686 4616
rect 20990 4564 20996 4616
rect 21048 4604 21054 4616
rect 21085 4607 21143 4613
rect 21085 4604 21097 4607
rect 21048 4576 21097 4604
rect 21048 4564 21054 4576
rect 21085 4573 21097 4576
rect 21131 4573 21143 4607
rect 22094 4604 22100 4616
rect 21085 4567 21143 4573
rect 21192 4576 21956 4604
rect 22055 4576 22100 4604
rect 16592 4508 16804 4536
rect 17313 4539 17371 4545
rect 16393 4499 16451 4505
rect 17313 4505 17325 4539
rect 17359 4505 17371 4539
rect 17313 4499 17371 4505
rect 4062 4428 4068 4480
rect 4120 4468 4126 4480
rect 4157 4471 4215 4477
rect 4157 4468 4169 4471
rect 4120 4440 4169 4468
rect 4120 4428 4126 4440
rect 4157 4437 4169 4440
rect 4203 4437 4215 4471
rect 4157 4431 4215 4437
rect 9033 4471 9091 4477
rect 9033 4437 9045 4471
rect 9079 4468 9091 4471
rect 9398 4468 9404 4480
rect 9079 4440 9404 4468
rect 9079 4437 9091 4440
rect 9033 4431 9091 4437
rect 9398 4428 9404 4440
rect 9456 4468 9462 4480
rect 9674 4468 9680 4480
rect 9456 4440 9680 4468
rect 9456 4428 9462 4440
rect 9674 4428 9680 4440
rect 9732 4428 9738 4480
rect 11517 4471 11575 4477
rect 11517 4437 11529 4471
rect 11563 4468 11575 4471
rect 12802 4468 12808 4480
rect 11563 4440 12808 4468
rect 11563 4437 11575 4440
rect 11517 4431 11575 4437
rect 12802 4428 12808 4440
rect 12860 4428 12866 4480
rect 13449 4471 13507 4477
rect 13449 4437 13461 4471
rect 13495 4468 13507 4471
rect 13814 4468 13820 4480
rect 13495 4440 13820 4468
rect 13495 4437 13507 4440
rect 13449 4431 13507 4437
rect 13814 4428 13820 4440
rect 13872 4428 13878 4480
rect 15013 4471 15071 4477
rect 15013 4437 15025 4471
rect 15059 4468 15071 4471
rect 16298 4468 16304 4480
rect 15059 4440 16304 4468
rect 15059 4437 15071 4440
rect 15013 4431 15071 4437
rect 16298 4428 16304 4440
rect 16356 4428 16362 4480
rect 16408 4468 16436 4499
rect 17328 4468 17356 4499
rect 20898 4496 20904 4548
rect 20956 4536 20962 4548
rect 21192 4536 21220 4576
rect 20956 4508 21220 4536
rect 21361 4539 21419 4545
rect 20956 4496 20962 4508
rect 21361 4505 21373 4539
rect 21407 4536 21419 4539
rect 21450 4536 21456 4548
rect 21407 4508 21456 4536
rect 21407 4505 21419 4508
rect 21361 4499 21419 4505
rect 21450 4496 21456 4508
rect 21508 4536 21514 4548
rect 21821 4539 21879 4545
rect 21821 4536 21833 4539
rect 21508 4508 21833 4536
rect 21508 4496 21514 4508
rect 21821 4505 21833 4508
rect 21867 4505 21879 4539
rect 21928 4536 21956 4576
rect 22094 4564 22100 4576
rect 22152 4564 22158 4616
rect 23400 4613 23428 4644
rect 23293 4607 23351 4613
rect 23293 4573 23305 4607
rect 23339 4573 23351 4607
rect 23293 4567 23351 4573
rect 23382 4607 23440 4613
rect 23382 4573 23394 4607
rect 23428 4573 23440 4607
rect 23382 4567 23440 4573
rect 23477 4607 23535 4613
rect 23477 4573 23489 4607
rect 23523 4604 23535 4607
rect 23566 4604 23572 4616
rect 23523 4576 23572 4604
rect 23523 4573 23535 4576
rect 23477 4567 23535 4573
rect 23308 4536 23336 4567
rect 23566 4564 23572 4576
rect 23624 4564 23630 4616
rect 23658 4564 23664 4616
rect 23716 4604 23722 4616
rect 24394 4604 24400 4616
rect 23716 4576 23761 4604
rect 24355 4576 24400 4604
rect 23716 4564 23722 4576
rect 24394 4564 24400 4576
rect 24452 4564 24458 4616
rect 21928 4508 23336 4536
rect 21821 4499 21879 4505
rect 16408 4440 17356 4468
rect 17954 4428 17960 4480
rect 18012 4468 18018 4480
rect 18325 4471 18383 4477
rect 18325 4468 18337 4471
rect 18012 4440 18337 4468
rect 18012 4428 18018 4440
rect 18325 4437 18337 4440
rect 18371 4437 18383 4471
rect 18325 4431 18383 4437
rect 19702 4428 19708 4480
rect 19760 4468 19766 4480
rect 20346 4468 20352 4480
rect 19760 4440 20352 4468
rect 19760 4428 19766 4440
rect 20346 4428 20352 4440
rect 20404 4428 20410 4480
rect 20806 4428 20812 4480
rect 20864 4468 20870 4480
rect 23017 4471 23075 4477
rect 23017 4468 23029 4471
rect 20864 4440 23029 4468
rect 20864 4428 20870 4440
rect 23017 4437 23029 4440
rect 23063 4437 23075 4471
rect 23017 4431 23075 4437
rect 1104 4378 68816 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 50294 4378
rect 50346 4326 50358 4378
rect 50410 4326 50422 4378
rect 50474 4326 50486 4378
rect 50538 4326 50550 4378
rect 50602 4326 68816 4378
rect 1104 4304 68816 4326
rect 6914 4264 6920 4276
rect 5552 4236 6920 4264
rect 3252 4168 3924 4196
rect 2869 4131 2927 4137
rect 2869 4097 2881 4131
rect 2915 4128 2927 4131
rect 3252 4128 3280 4168
rect 2915 4100 3280 4128
rect 3329 4131 3387 4137
rect 2915 4097 2927 4100
rect 2869 4091 2927 4097
rect 3329 4097 3341 4131
rect 3375 4128 3387 4131
rect 3786 4128 3792 4140
rect 3375 4100 3792 4128
rect 3375 4097 3387 4100
rect 3329 4091 3387 4097
rect 3786 4088 3792 4100
rect 3844 4088 3850 4140
rect 3896 4128 3924 4168
rect 4154 4128 4160 4140
rect 3896 4100 4160 4128
rect 4154 4088 4160 4100
rect 4212 4088 4218 4140
rect 5552 4128 5580 4236
rect 6914 4224 6920 4236
rect 6972 4264 6978 4276
rect 7929 4267 7987 4273
rect 7929 4264 7941 4267
rect 6972 4236 7941 4264
rect 6972 4224 6978 4236
rect 7929 4233 7941 4236
rect 7975 4233 7987 4267
rect 7929 4227 7987 4233
rect 11609 4267 11667 4273
rect 11609 4233 11621 4267
rect 11655 4264 11667 4267
rect 11790 4264 11796 4276
rect 11655 4236 11796 4264
rect 11655 4233 11667 4236
rect 11609 4227 11667 4233
rect 11790 4224 11796 4236
rect 11848 4224 11854 4276
rect 12434 4264 12440 4276
rect 12360 4236 12440 4264
rect 8294 4196 8300 4208
rect 6748 4168 8300 4196
rect 4632 4100 5580 4128
rect 5629 4131 5687 4137
rect 3421 4063 3479 4069
rect 3421 4029 3433 4063
rect 3467 4060 3479 4063
rect 4632 4060 4660 4100
rect 5629 4097 5641 4131
rect 5675 4097 5687 4131
rect 5810 4128 5816 4140
rect 5771 4100 5816 4128
rect 5629 4091 5687 4097
rect 3467 4032 4660 4060
rect 4985 4063 5043 4069
rect 3467 4029 3479 4032
rect 3421 4023 3479 4029
rect 4985 4029 4997 4063
rect 5031 4060 5043 4063
rect 5074 4060 5080 4072
rect 5031 4032 5080 4060
rect 5031 4029 5043 4032
rect 4985 4023 5043 4029
rect 3970 3992 3976 4004
rect 3528 3964 3976 3992
rect 3528 3933 3556 3964
rect 3970 3952 3976 3964
rect 4028 3952 4034 4004
rect 4154 3952 4160 4004
rect 4212 3992 4218 4004
rect 5000 3992 5028 4023
rect 5074 4020 5080 4032
rect 5132 4020 5138 4072
rect 5644 4060 5672 4091
rect 5810 4088 5816 4100
rect 5868 4088 5874 4140
rect 6549 4131 6607 4137
rect 6549 4097 6561 4131
rect 6595 4128 6607 4131
rect 6748 4128 6776 4168
rect 8294 4156 8300 4168
rect 8352 4196 8358 4208
rect 9582 4196 9588 4208
rect 8352 4168 9588 4196
rect 8352 4156 8358 4168
rect 6822 4137 6828 4140
rect 6595 4100 6776 4128
rect 6595 4097 6607 4100
rect 6549 4091 6607 4097
rect 6816 4091 6828 4137
rect 6880 4128 6886 4140
rect 8404 4137 8432 4168
rect 9582 4156 9588 4168
rect 9640 4156 9646 4208
rect 10870 4196 10876 4208
rect 10831 4168 10876 4196
rect 10870 4156 10876 4168
rect 10928 4156 10934 4208
rect 8389 4131 8447 4137
rect 6880 4100 6916 4128
rect 6822 4088 6828 4091
rect 6880 4088 6886 4100
rect 8389 4097 8401 4131
rect 8435 4097 8447 4131
rect 8389 4091 8447 4097
rect 8478 4088 8484 4140
rect 8536 4128 8542 4140
rect 8645 4131 8703 4137
rect 8645 4128 8657 4131
rect 8536 4100 8657 4128
rect 8536 4088 8542 4100
rect 8645 4097 8657 4100
rect 8691 4097 8703 4131
rect 8645 4091 8703 4097
rect 9214 4088 9220 4140
rect 9272 4128 9278 4140
rect 12066 4128 12072 4140
rect 9272 4100 11928 4128
rect 12027 4100 12072 4128
rect 9272 4088 9278 4100
rect 6270 4060 6276 4072
rect 5644 4032 6276 4060
rect 6270 4020 6276 4032
rect 6328 4020 6334 4072
rect 10134 4020 10140 4072
rect 10192 4060 10198 4072
rect 10689 4063 10747 4069
rect 10689 4060 10701 4063
rect 10192 4032 10701 4060
rect 10192 4020 10198 4032
rect 10689 4029 10701 4032
rect 10735 4029 10747 4063
rect 11900 4060 11928 4100
rect 12066 4088 12072 4100
rect 12124 4088 12130 4140
rect 12250 4128 12256 4140
rect 12211 4100 12256 4128
rect 12250 4088 12256 4100
rect 12308 4088 12314 4140
rect 12360 4137 12388 4236
rect 12434 4224 12440 4236
rect 12492 4224 12498 4276
rect 20438 4264 20444 4276
rect 20399 4236 20444 4264
rect 20438 4224 20444 4236
rect 20496 4224 20502 4276
rect 20714 4196 20720 4208
rect 20548 4168 20720 4196
rect 12345 4131 12403 4137
rect 12345 4097 12357 4131
rect 12391 4097 12403 4131
rect 12345 4091 12403 4097
rect 12437 4131 12495 4137
rect 12437 4097 12449 4131
rect 12483 4097 12495 4131
rect 12437 4091 12495 4097
rect 12158 4060 12164 4072
rect 11900 4032 12164 4060
rect 10689 4023 10747 4029
rect 12158 4020 12164 4032
rect 12216 4020 12222 4072
rect 12360 4060 12388 4091
rect 12268 4032 12388 4060
rect 12268 4004 12296 4032
rect 4212 3964 5028 3992
rect 4212 3952 4218 3964
rect 9398 3952 9404 4004
rect 9456 3992 9462 4004
rect 11790 3992 11796 4004
rect 9456 3964 11796 3992
rect 9456 3952 9462 3964
rect 11790 3952 11796 3964
rect 11848 3952 11854 4004
rect 12250 3952 12256 4004
rect 12308 3952 12314 4004
rect 3513 3927 3571 3933
rect 3513 3893 3525 3927
rect 3559 3893 3571 3927
rect 3513 3887 3571 3893
rect 3697 3927 3755 3933
rect 3697 3893 3709 3927
rect 3743 3924 3755 3927
rect 4614 3924 4620 3936
rect 3743 3896 4620 3924
rect 3743 3893 3755 3896
rect 3697 3887 3755 3893
rect 4614 3884 4620 3896
rect 4672 3884 4678 3936
rect 4755 3927 4813 3933
rect 4755 3893 4767 3927
rect 4801 3924 4813 3927
rect 5442 3924 5448 3936
rect 4801 3896 5448 3924
rect 4801 3893 4813 3896
rect 4755 3887 4813 3893
rect 5442 3884 5448 3896
rect 5500 3884 5506 3936
rect 5721 3927 5779 3933
rect 5721 3893 5733 3927
rect 5767 3924 5779 3927
rect 6914 3924 6920 3936
rect 5767 3896 6920 3924
rect 5767 3893 5779 3896
rect 5721 3887 5779 3893
rect 6914 3884 6920 3896
rect 6972 3884 6978 3936
rect 9766 3924 9772 3936
rect 9727 3896 9772 3924
rect 9766 3884 9772 3896
rect 9824 3884 9830 3936
rect 12452 3924 12480 4091
rect 12894 4088 12900 4140
rect 12952 4128 12958 4140
rect 13173 4131 13231 4137
rect 13173 4128 13185 4131
rect 12952 4100 13185 4128
rect 12952 4088 12958 4100
rect 13173 4097 13185 4100
rect 13219 4097 13231 4131
rect 13429 4131 13487 4137
rect 13429 4128 13441 4131
rect 13173 4091 13231 4097
rect 13280 4100 13441 4128
rect 12713 4063 12771 4069
rect 12713 4029 12725 4063
rect 12759 4060 12771 4063
rect 13280 4060 13308 4100
rect 13429 4097 13441 4100
rect 13475 4097 13487 4131
rect 13429 4091 13487 4097
rect 13722 4088 13728 4140
rect 13780 4128 13786 4140
rect 15105 4131 15163 4137
rect 15105 4128 15117 4131
rect 13780 4100 15117 4128
rect 13780 4088 13786 4100
rect 15105 4097 15117 4100
rect 15151 4097 15163 4131
rect 15105 4091 15163 4097
rect 15841 4131 15899 4137
rect 15841 4097 15853 4131
rect 15887 4097 15899 4131
rect 17218 4128 17224 4140
rect 17179 4100 17224 4128
rect 15841 4091 15899 4097
rect 15856 4060 15884 4091
rect 17218 4088 17224 4100
rect 17276 4088 17282 4140
rect 17957 4131 18015 4137
rect 17957 4097 17969 4131
rect 18003 4128 18015 4131
rect 18046 4128 18052 4140
rect 18003 4100 18052 4128
rect 18003 4097 18015 4100
rect 17957 4091 18015 4097
rect 18046 4088 18052 4100
rect 18104 4088 18110 4140
rect 18224 4131 18282 4137
rect 18224 4097 18236 4131
rect 18270 4128 18282 4131
rect 20548 4128 20576 4168
rect 20714 4156 20720 4168
rect 20772 4156 20778 4208
rect 21450 4156 21456 4208
rect 21508 4196 21514 4208
rect 21821 4199 21879 4205
rect 21821 4196 21833 4199
rect 21508 4168 21833 4196
rect 21508 4156 21514 4168
rect 21821 4165 21833 4168
rect 21867 4165 21879 4199
rect 21821 4159 21879 4165
rect 18270 4100 20576 4128
rect 18270 4097 18282 4100
rect 18224 4091 18282 4097
rect 20622 4088 20628 4140
rect 20680 4128 20686 4140
rect 21085 4131 21143 4137
rect 20680 4100 20725 4128
rect 20680 4088 20686 4100
rect 21085 4097 21097 4131
rect 21131 4128 21143 4131
rect 21634 4128 21640 4140
rect 21131 4100 21640 4128
rect 21131 4097 21143 4100
rect 21085 4091 21143 4097
rect 21634 4088 21640 4100
rect 21692 4088 21698 4140
rect 22094 4128 22100 4140
rect 22055 4100 22100 4128
rect 22094 4088 22100 4100
rect 22152 4088 22158 4140
rect 12759 4032 13308 4060
rect 14568 4032 15884 4060
rect 12759 4029 12771 4032
rect 12713 4023 12771 4029
rect 14568 3933 14596 4032
rect 20438 4020 20444 4072
rect 20496 4060 20502 4072
rect 21913 4063 21971 4069
rect 21913 4060 21925 4063
rect 20496 4032 21925 4060
rect 20496 4020 20502 4032
rect 21913 4029 21925 4032
rect 21959 4029 21971 4063
rect 21913 4023 21971 4029
rect 22002 4020 22008 4072
rect 22060 4060 22066 4072
rect 23385 4063 23443 4069
rect 23385 4060 23397 4063
rect 22060 4032 23397 4060
rect 22060 4020 22066 4032
rect 23385 4029 23397 4032
rect 23431 4029 23443 4063
rect 23385 4023 23443 4029
rect 15746 3952 15752 4004
rect 15804 3992 15810 4004
rect 16666 3992 16672 4004
rect 15804 3964 16672 3992
rect 15804 3952 15810 3964
rect 16666 3952 16672 3964
rect 16724 3952 16730 4004
rect 16761 3995 16819 4001
rect 16761 3961 16773 3995
rect 16807 3992 16819 3995
rect 17678 3992 17684 4004
rect 16807 3964 17684 3992
rect 16807 3961 16819 3964
rect 16761 3955 16819 3961
rect 17678 3952 17684 3964
rect 17736 3992 17742 4004
rect 19981 3995 20039 4001
rect 17736 3964 18000 3992
rect 17736 3952 17742 3964
rect 14553 3927 14611 3933
rect 14553 3924 14565 3927
rect 12452 3896 14565 3924
rect 14553 3893 14565 3896
rect 14599 3893 14611 3927
rect 14553 3887 14611 3893
rect 15289 3927 15347 3933
rect 15289 3893 15301 3927
rect 15335 3924 15347 3927
rect 15930 3924 15936 3936
rect 15335 3896 15936 3924
rect 15335 3893 15347 3896
rect 15289 3887 15347 3893
rect 15930 3884 15936 3896
rect 15988 3884 15994 3936
rect 16025 3927 16083 3933
rect 16025 3893 16037 3927
rect 16071 3924 16083 3927
rect 16482 3924 16488 3936
rect 16071 3896 16488 3924
rect 16071 3893 16083 3896
rect 16025 3887 16083 3893
rect 16482 3884 16488 3896
rect 16540 3884 16546 3936
rect 17310 3884 17316 3936
rect 17368 3924 17374 3936
rect 17405 3927 17463 3933
rect 17405 3924 17417 3927
rect 17368 3896 17417 3924
rect 17368 3884 17374 3896
rect 17405 3893 17417 3896
rect 17451 3893 17463 3927
rect 17972 3924 18000 3964
rect 18892 3964 19472 3992
rect 18892 3924 18920 3964
rect 19334 3924 19340 3936
rect 17972 3896 18920 3924
rect 19295 3896 19340 3924
rect 17405 3887 17463 3893
rect 19334 3884 19340 3896
rect 19392 3884 19398 3936
rect 19444 3924 19472 3964
rect 19981 3961 19993 3995
rect 20027 3992 20039 3995
rect 21450 3992 21456 4004
rect 20027 3964 21456 3992
rect 20027 3961 20039 3964
rect 19981 3955 20039 3961
rect 21450 3952 21456 3964
rect 21508 3952 21514 4004
rect 22186 3952 22192 4004
rect 22244 3992 22250 4004
rect 22281 3995 22339 4001
rect 22281 3992 22293 3995
rect 22244 3964 22293 3992
rect 22244 3952 22250 3964
rect 22281 3961 22293 3964
rect 22327 3961 22339 3995
rect 22281 3955 22339 3961
rect 20530 3924 20536 3936
rect 19444 3896 20536 3924
rect 20530 3884 20536 3896
rect 20588 3884 20594 3936
rect 21269 3927 21327 3933
rect 21269 3893 21281 3927
rect 21315 3924 21327 3927
rect 21726 3924 21732 3936
rect 21315 3896 21732 3924
rect 21315 3893 21327 3896
rect 21269 3887 21327 3893
rect 21726 3884 21732 3896
rect 21784 3884 21790 3936
rect 21910 3924 21916 3936
rect 21871 3896 21916 3924
rect 21910 3884 21916 3896
rect 21968 3884 21974 3936
rect 22462 3884 22468 3936
rect 22520 3924 22526 3936
rect 22741 3927 22799 3933
rect 22741 3924 22753 3927
rect 22520 3896 22753 3924
rect 22520 3884 22526 3896
rect 22741 3893 22753 3896
rect 22787 3893 22799 3927
rect 24026 3924 24032 3936
rect 23987 3896 24032 3924
rect 22741 3887 22799 3893
rect 24026 3884 24032 3896
rect 24084 3884 24090 3936
rect 24670 3924 24676 3936
rect 24631 3896 24676 3924
rect 24670 3884 24676 3896
rect 24728 3884 24734 3936
rect 1104 3834 68816 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 65654 3834
rect 65706 3782 65718 3834
rect 65770 3782 65782 3834
rect 65834 3782 65846 3834
rect 65898 3782 65910 3834
rect 65962 3782 68816 3834
rect 1104 3760 68816 3782
rect 5905 3723 5963 3729
rect 5905 3689 5917 3723
rect 5951 3720 5963 3723
rect 8478 3720 8484 3732
rect 5951 3692 8484 3720
rect 5951 3689 5963 3692
rect 5905 3683 5963 3689
rect 8478 3680 8484 3692
rect 8536 3680 8542 3732
rect 8570 3680 8576 3732
rect 8628 3720 8634 3732
rect 8628 3692 11284 3720
rect 8628 3680 8634 3692
rect 4246 3652 4252 3664
rect 4207 3624 4252 3652
rect 4246 3612 4252 3624
rect 4304 3612 4310 3664
rect 5166 3612 5172 3664
rect 5224 3652 5230 3664
rect 6086 3652 6092 3664
rect 5224 3624 6092 3652
rect 5224 3612 5230 3624
rect 6086 3612 6092 3624
rect 6144 3612 6150 3664
rect 9766 3652 9772 3664
rect 6196 3624 9772 3652
rect 4982 3544 4988 3596
rect 5040 3584 5046 3596
rect 5040 3556 5375 3584
rect 5040 3544 5046 3556
rect 4154 3476 4160 3528
rect 4212 3516 4218 3528
rect 5166 3516 5172 3528
rect 4212 3488 5172 3516
rect 4212 3476 4218 3488
rect 5166 3476 5172 3488
rect 5224 3516 5230 3528
rect 5261 3519 5319 3525
rect 5261 3516 5273 3519
rect 5224 3488 5273 3516
rect 5224 3476 5230 3488
rect 5261 3485 5273 3488
rect 5307 3485 5319 3519
rect 5347 3516 5375 3556
rect 5424 3516 5482 3522
rect 5675 3519 5733 3525
rect 5347 3513 5396 3516
rect 5424 3513 5436 3516
rect 5347 3488 5436 3513
rect 5368 3485 5436 3488
rect 5261 3479 5319 3485
rect 5424 3482 5436 3485
rect 5470 3482 5482 3516
rect 5424 3476 5482 3482
rect 5524 3513 5582 3519
rect 5524 3479 5536 3513
rect 5570 3492 5582 3513
rect 5570 3479 5626 3492
rect 5675 3485 5687 3519
rect 5721 3516 5733 3519
rect 6196 3516 6224 3624
rect 9766 3612 9772 3624
rect 9824 3612 9830 3664
rect 11256 3652 11284 3692
rect 12066 3680 12072 3732
rect 12124 3720 12130 3732
rect 13538 3720 13544 3732
rect 12124 3692 13544 3720
rect 12124 3680 12130 3692
rect 13538 3680 13544 3692
rect 13596 3680 13602 3732
rect 15746 3720 15752 3732
rect 14108 3692 15752 3720
rect 14108 3652 14136 3692
rect 15746 3680 15752 3692
rect 15804 3680 15810 3732
rect 20254 3680 20260 3732
rect 20312 3720 20318 3732
rect 20438 3720 20444 3732
rect 20312 3692 20444 3720
rect 20312 3680 20318 3692
rect 20438 3680 20444 3692
rect 20496 3680 20502 3732
rect 21729 3723 21787 3729
rect 21729 3689 21741 3723
rect 21775 3720 21787 3723
rect 21818 3720 21824 3732
rect 21775 3692 21824 3720
rect 21775 3689 21787 3692
rect 21729 3683 21787 3689
rect 21818 3680 21824 3692
rect 21876 3680 21882 3732
rect 11256 3624 14136 3652
rect 14461 3655 14519 3661
rect 14461 3621 14473 3655
rect 14507 3652 14519 3655
rect 15562 3652 15568 3664
rect 14507 3624 15568 3652
rect 14507 3621 14519 3624
rect 14461 3615 14519 3621
rect 15562 3612 15568 3624
rect 15620 3612 15626 3664
rect 17221 3655 17279 3661
rect 17221 3621 17233 3655
rect 17267 3621 17279 3655
rect 17221 3615 17279 3621
rect 6914 3544 6920 3596
rect 6972 3584 6978 3596
rect 6972 3556 9536 3584
rect 6972 3544 6978 3556
rect 5721 3488 6224 3516
rect 6365 3519 6423 3525
rect 5721 3485 5733 3488
rect 5675 3479 5733 3485
rect 6365 3485 6377 3519
rect 6411 3485 6423 3519
rect 6365 3479 6423 3485
rect 5524 3473 5626 3479
rect 5552 3464 5626 3473
rect 4798 3380 4804 3392
rect 4759 3352 4804 3380
rect 4798 3340 4804 3352
rect 4856 3340 4862 3392
rect 5442 3340 5448 3392
rect 5500 3380 5506 3392
rect 5598 3380 5626 3464
rect 6086 3408 6092 3460
rect 6144 3448 6150 3460
rect 6380 3448 6408 3479
rect 6454 3476 6460 3528
rect 6512 3516 6518 3528
rect 6549 3519 6607 3525
rect 6549 3516 6561 3519
rect 6512 3488 6561 3516
rect 6512 3476 6518 3488
rect 6549 3485 6561 3488
rect 6595 3485 6607 3519
rect 6549 3479 6607 3485
rect 6641 3519 6699 3525
rect 6641 3485 6653 3519
rect 6687 3485 6699 3519
rect 6641 3479 6699 3485
rect 6733 3519 6791 3525
rect 6733 3485 6745 3519
rect 6779 3516 6791 3519
rect 7650 3516 7656 3528
rect 6779 3488 7656 3516
rect 6779 3485 6791 3488
rect 6733 3479 6791 3485
rect 6144 3420 6408 3448
rect 6144 3408 6150 3420
rect 6656 3380 6684 3479
rect 7650 3476 7656 3488
rect 7708 3476 7714 3528
rect 7745 3519 7803 3525
rect 7745 3485 7757 3519
rect 7791 3516 7803 3519
rect 8110 3516 8116 3528
rect 7791 3488 8116 3516
rect 7791 3485 7803 3488
rect 7745 3479 7803 3485
rect 8110 3476 8116 3488
rect 8168 3476 8174 3528
rect 8202 3476 8208 3528
rect 8260 3516 8266 3528
rect 8938 3516 8944 3528
rect 8260 3488 8305 3516
rect 8899 3488 8944 3516
rect 8260 3476 8266 3488
rect 8938 3476 8944 3488
rect 8996 3476 9002 3528
rect 9508 3525 9536 3556
rect 9582 3544 9588 3596
rect 9640 3584 9646 3596
rect 10321 3587 10379 3593
rect 10321 3584 10333 3587
rect 9640 3556 10333 3584
rect 9640 3544 9646 3556
rect 10321 3553 10333 3556
rect 10367 3553 10379 3587
rect 13262 3584 13268 3596
rect 13223 3556 13268 3584
rect 10321 3547 10379 3553
rect 13262 3544 13268 3556
rect 13320 3544 13326 3596
rect 14090 3584 14096 3596
rect 13372 3556 14096 3584
rect 9493 3519 9551 3525
rect 9493 3485 9505 3519
rect 9539 3516 9551 3519
rect 10870 3516 10876 3528
rect 9539 3488 10876 3516
rect 9539 3485 9551 3488
rect 9493 3479 9551 3485
rect 10870 3476 10876 3488
rect 10928 3476 10934 3528
rect 12250 3476 12256 3528
rect 12308 3516 12314 3528
rect 12989 3519 13047 3525
rect 12989 3516 13001 3519
rect 12308 3488 13001 3516
rect 12308 3476 12314 3488
rect 12989 3485 13001 3488
rect 13035 3516 13047 3519
rect 13372 3516 13400 3556
rect 14090 3544 14096 3556
rect 14148 3584 14154 3596
rect 14148 3556 16068 3584
rect 14148 3544 14154 3556
rect 13035 3488 13400 3516
rect 14277 3519 14335 3525
rect 13035 3485 13047 3488
rect 12989 3479 13047 3485
rect 14277 3485 14289 3519
rect 14323 3485 14335 3519
rect 15286 3516 15292 3528
rect 15247 3488 15292 3516
rect 14277 3479 14335 3485
rect 6822 3408 6828 3460
rect 6880 3448 6886 3460
rect 10566 3451 10624 3457
rect 10566 3448 10578 3451
rect 6880 3420 10578 3448
rect 6880 3408 6886 3420
rect 10566 3417 10578 3420
rect 10612 3417 10624 3451
rect 14292 3448 14320 3479
rect 15286 3476 15292 3488
rect 15344 3476 15350 3528
rect 15470 3476 15476 3528
rect 15528 3516 15534 3528
rect 15737 3519 15795 3525
rect 15737 3516 15749 3519
rect 15528 3488 15749 3516
rect 15528 3476 15534 3488
rect 15737 3485 15749 3488
rect 15783 3485 15795 3519
rect 15737 3479 15795 3485
rect 15838 3476 15844 3528
rect 15896 3516 15902 3528
rect 16040 3525 16068 3556
rect 16206 3525 16212 3528
rect 15933 3519 15991 3525
rect 15933 3516 15945 3519
rect 15896 3488 15945 3516
rect 15896 3476 15902 3488
rect 15933 3485 15945 3488
rect 15979 3485 15991 3519
rect 15933 3479 15991 3485
rect 16025 3519 16083 3525
rect 16025 3485 16037 3519
rect 16071 3485 16083 3519
rect 16025 3479 16083 3485
rect 16163 3519 16212 3525
rect 16163 3485 16175 3519
rect 16209 3485 16212 3519
rect 16163 3479 16212 3485
rect 15194 3448 15200 3460
rect 10566 3411 10624 3417
rect 11716 3420 14320 3448
rect 14384 3420 15200 3448
rect 11716 3392 11744 3420
rect 5500 3352 6684 3380
rect 7009 3383 7067 3389
rect 5500 3340 5506 3352
rect 7009 3349 7021 3383
rect 7055 3380 7067 3383
rect 7282 3380 7288 3392
rect 7055 3352 7288 3380
rect 7055 3349 7067 3352
rect 7009 3343 7067 3349
rect 7282 3340 7288 3352
rect 7340 3340 7346 3392
rect 7558 3380 7564 3392
rect 7519 3352 7564 3380
rect 7558 3340 7564 3352
rect 7616 3340 7622 3392
rect 8389 3383 8447 3389
rect 8389 3349 8401 3383
rect 8435 3380 8447 3383
rect 8754 3380 8760 3392
rect 8435 3352 8760 3380
rect 8435 3349 8447 3352
rect 8389 3343 8447 3349
rect 8754 3340 8760 3352
rect 8812 3340 8818 3392
rect 9674 3380 9680 3392
rect 9635 3352 9680 3380
rect 9674 3340 9680 3352
rect 9732 3340 9738 3392
rect 11698 3380 11704 3392
rect 11659 3352 11704 3380
rect 11698 3340 11704 3352
rect 11756 3340 11762 3392
rect 11790 3340 11796 3392
rect 11848 3380 11854 3392
rect 14384 3380 14412 3420
rect 15194 3408 15200 3420
rect 15252 3408 15258 3460
rect 16040 3448 16068 3479
rect 16206 3476 16212 3479
rect 16264 3516 16270 3528
rect 17236 3516 17264 3615
rect 18690 3612 18696 3664
rect 18748 3652 18754 3664
rect 20073 3655 20131 3661
rect 20073 3652 20085 3655
rect 18748 3624 20085 3652
rect 18748 3612 18754 3624
rect 20073 3621 20085 3624
rect 20119 3621 20131 3655
rect 20073 3615 20131 3621
rect 20622 3612 20628 3664
rect 20680 3652 20686 3664
rect 21913 3655 21971 3661
rect 21913 3652 21925 3655
rect 20680 3624 21925 3652
rect 20680 3612 20686 3624
rect 21913 3621 21925 3624
rect 21959 3621 21971 3655
rect 21913 3615 21971 3621
rect 51442 3612 51448 3664
rect 51500 3652 51506 3664
rect 52089 3655 52147 3661
rect 52089 3652 52101 3655
rect 51500 3624 52101 3652
rect 51500 3612 51506 3624
rect 52089 3621 52101 3624
rect 52135 3621 52147 3655
rect 52089 3615 52147 3621
rect 21818 3544 21824 3596
rect 21876 3584 21882 3596
rect 24397 3587 24455 3593
rect 24397 3584 24409 3587
rect 21876 3556 24409 3584
rect 21876 3544 21882 3556
rect 24397 3553 24409 3556
rect 24443 3553 24455 3587
rect 24397 3547 24455 3553
rect 16264 3488 17264 3516
rect 16264 3476 16270 3488
rect 18046 3476 18052 3528
rect 18104 3516 18110 3528
rect 18601 3519 18659 3525
rect 18601 3516 18613 3519
rect 18104 3488 18613 3516
rect 18104 3476 18110 3488
rect 18601 3485 18613 3488
rect 18647 3485 18659 3519
rect 18601 3479 18659 3485
rect 18966 3476 18972 3528
rect 19024 3516 19030 3528
rect 19521 3519 19579 3525
rect 19521 3516 19533 3519
rect 19024 3488 19533 3516
rect 19024 3476 19030 3488
rect 19521 3485 19533 3488
rect 19567 3485 19579 3519
rect 19521 3479 19579 3485
rect 20257 3519 20315 3525
rect 20257 3485 20269 3519
rect 20303 3516 20315 3519
rect 20898 3516 20904 3528
rect 20303 3488 20904 3516
rect 20303 3485 20315 3488
rect 20257 3479 20315 3485
rect 20898 3476 20904 3488
rect 20956 3476 20962 3528
rect 21266 3516 21272 3528
rect 21227 3488 21272 3516
rect 21266 3476 21272 3488
rect 21324 3476 21330 3528
rect 21358 3476 21364 3528
rect 21416 3516 21422 3528
rect 21726 3516 21732 3528
rect 21416 3488 21461 3516
rect 21687 3488 21732 3516
rect 21416 3476 21422 3488
rect 21726 3476 21732 3488
rect 21784 3476 21790 3528
rect 22738 3476 22744 3528
rect 22796 3516 22802 3528
rect 22833 3519 22891 3525
rect 22833 3516 22845 3519
rect 22796 3488 22845 3516
rect 22796 3476 22802 3488
rect 22833 3485 22845 3488
rect 22879 3485 22891 3519
rect 22833 3479 22891 3485
rect 23566 3476 23572 3528
rect 23624 3516 23630 3528
rect 23661 3519 23719 3525
rect 23661 3516 23673 3519
rect 23624 3488 23673 3516
rect 23624 3476 23630 3488
rect 23661 3485 23673 3488
rect 23707 3485 23719 3519
rect 23661 3479 23719 3485
rect 26050 3476 26056 3528
rect 26108 3516 26114 3528
rect 26145 3519 26203 3525
rect 26145 3516 26157 3519
rect 26108 3488 26157 3516
rect 26108 3476 26114 3488
rect 26145 3485 26157 3488
rect 26191 3485 26203 3519
rect 26145 3479 26203 3485
rect 27249 3519 27307 3525
rect 27249 3485 27261 3519
rect 27295 3516 27307 3519
rect 27430 3516 27436 3528
rect 27295 3488 27436 3516
rect 27295 3485 27307 3488
rect 27249 3479 27307 3485
rect 27430 3476 27436 3488
rect 27488 3476 27494 3528
rect 27706 3516 27712 3528
rect 27667 3488 27712 3516
rect 27706 3476 27712 3488
rect 27764 3476 27770 3528
rect 28258 3476 28264 3528
rect 28316 3516 28322 3528
rect 28353 3519 28411 3525
rect 28353 3516 28365 3519
rect 28316 3488 28365 3516
rect 28316 3476 28322 3488
rect 28353 3485 28365 3488
rect 28399 3485 28411 3519
rect 28353 3479 28411 3485
rect 29362 3476 29368 3528
rect 29420 3516 29426 3528
rect 29549 3519 29607 3525
rect 29549 3516 29561 3519
rect 29420 3488 29561 3516
rect 29420 3476 29426 3488
rect 29549 3485 29561 3488
rect 29595 3485 29607 3519
rect 29549 3479 29607 3485
rect 30190 3476 30196 3528
rect 30248 3516 30254 3528
rect 30285 3519 30343 3525
rect 30285 3516 30297 3519
rect 30248 3488 30297 3516
rect 30248 3476 30254 3488
rect 30285 3485 30297 3488
rect 30331 3485 30343 3519
rect 30285 3479 30343 3485
rect 31294 3476 31300 3528
rect 31352 3516 31358 3528
rect 31389 3519 31447 3525
rect 31389 3516 31401 3519
rect 31352 3488 31401 3516
rect 31352 3476 31358 3488
rect 31389 3485 31401 3488
rect 31435 3485 31447 3519
rect 31389 3479 31447 3485
rect 32122 3476 32128 3528
rect 32180 3516 32186 3528
rect 32217 3519 32275 3525
rect 32217 3516 32229 3519
rect 32180 3488 32229 3516
rect 32180 3476 32186 3488
rect 32217 3485 32229 3488
rect 32263 3485 32275 3519
rect 32217 3479 32275 3485
rect 32950 3476 32956 3528
rect 33008 3516 33014 3528
rect 33045 3519 33103 3525
rect 33045 3516 33057 3519
rect 33008 3488 33057 3516
rect 33008 3476 33014 3488
rect 33045 3485 33057 3488
rect 33091 3485 33103 3519
rect 33045 3479 33103 3485
rect 39850 3476 39856 3528
rect 39908 3516 39914 3528
rect 39945 3519 40003 3525
rect 39945 3516 39957 3519
rect 39908 3488 39957 3516
rect 39908 3476 39914 3488
rect 39945 3485 39957 3488
rect 39991 3485 40003 3519
rect 39945 3479 40003 3485
rect 40126 3476 40132 3528
rect 40184 3516 40190 3528
rect 40589 3519 40647 3525
rect 40589 3516 40601 3519
rect 40184 3488 40601 3516
rect 40184 3476 40190 3488
rect 40589 3485 40601 3488
rect 40635 3485 40647 3519
rect 40589 3479 40647 3485
rect 40954 3476 40960 3528
rect 41012 3516 41018 3528
rect 41233 3519 41291 3525
rect 41233 3516 41245 3519
rect 41012 3488 41245 3516
rect 41012 3476 41018 3488
rect 41233 3485 41245 3488
rect 41279 3485 41291 3519
rect 41233 3479 41291 3485
rect 41782 3476 41788 3528
rect 41840 3516 41846 3528
rect 41877 3519 41935 3525
rect 41877 3516 41889 3519
rect 41840 3488 41889 3516
rect 41840 3476 41846 3488
rect 41877 3485 41889 3488
rect 41923 3485 41935 3519
rect 41877 3479 41935 3485
rect 42610 3476 42616 3528
rect 42668 3516 42674 3528
rect 42705 3519 42763 3525
rect 42705 3516 42717 3519
rect 42668 3488 42717 3516
rect 42668 3476 42674 3488
rect 42705 3485 42717 3488
rect 42751 3485 42763 3519
rect 42705 3479 42763 3485
rect 43714 3476 43720 3528
rect 43772 3516 43778 3528
rect 43809 3519 43867 3525
rect 43809 3516 43821 3519
rect 43772 3488 43821 3516
rect 43772 3476 43778 3488
rect 43809 3485 43821 3488
rect 43855 3485 43867 3519
rect 43809 3479 43867 3485
rect 45094 3476 45100 3528
rect 45152 3516 45158 3528
rect 45189 3519 45247 3525
rect 45189 3516 45201 3519
rect 45152 3488 45201 3516
rect 45152 3476 45158 3488
rect 45189 3485 45201 3488
rect 45235 3485 45247 3519
rect 45189 3479 45247 3485
rect 45646 3476 45652 3528
rect 45704 3516 45710 3528
rect 45833 3519 45891 3525
rect 45833 3516 45845 3519
rect 45704 3488 45845 3516
rect 45704 3476 45710 3488
rect 45833 3485 45845 3488
rect 45879 3485 45891 3519
rect 45833 3479 45891 3485
rect 46198 3476 46204 3528
rect 46256 3516 46262 3528
rect 46477 3519 46535 3525
rect 46477 3516 46489 3519
rect 46256 3488 46489 3516
rect 46256 3476 46262 3488
rect 46477 3485 46489 3488
rect 46523 3485 46535 3519
rect 46477 3479 46535 3485
rect 47578 3476 47584 3528
rect 47636 3516 47642 3528
rect 47673 3519 47731 3525
rect 47673 3516 47685 3519
rect 47636 3488 47685 3516
rect 47636 3476 47642 3488
rect 47673 3485 47685 3488
rect 47719 3485 47731 3519
rect 47673 3479 47731 3485
rect 47854 3476 47860 3528
rect 47912 3516 47918 3528
rect 48317 3519 48375 3525
rect 48317 3516 48329 3519
rect 47912 3488 48329 3516
rect 47912 3476 47918 3488
rect 48317 3485 48329 3488
rect 48363 3485 48375 3519
rect 48317 3479 48375 3485
rect 49510 3476 49516 3528
rect 49568 3516 49574 3528
rect 50157 3519 50215 3525
rect 50157 3516 50169 3519
rect 49568 3488 50169 3516
rect 49568 3476 49574 3488
rect 50157 3485 50169 3488
rect 50203 3485 50215 3519
rect 50157 3479 50215 3485
rect 50614 3476 50620 3528
rect 50672 3516 50678 3528
rect 50801 3519 50859 3525
rect 50801 3516 50813 3519
rect 50672 3488 50813 3516
rect 50672 3476 50678 3488
rect 50801 3485 50813 3488
rect 50847 3485 50859 3519
rect 50801 3479 50859 3485
rect 51166 3476 51172 3528
rect 51224 3516 51230 3528
rect 51445 3519 51503 3525
rect 51445 3516 51457 3519
rect 51224 3488 51457 3516
rect 51224 3476 51230 3488
rect 51445 3485 51457 3488
rect 51491 3485 51503 3519
rect 51445 3479 51503 3485
rect 52822 3476 52828 3528
rect 52880 3516 52886 3528
rect 52917 3519 52975 3525
rect 52917 3516 52929 3519
rect 52880 3488 52929 3516
rect 52880 3476 52886 3488
rect 52917 3485 52929 3488
rect 52963 3485 52975 3519
rect 52917 3479 52975 3485
rect 53374 3476 53380 3528
rect 53432 3516 53438 3528
rect 53561 3519 53619 3525
rect 53561 3516 53573 3519
rect 53432 3488 53573 3516
rect 53432 3476 53438 3488
rect 53561 3485 53573 3488
rect 53607 3485 53619 3519
rect 53561 3479 53619 3485
rect 55306 3476 55312 3528
rect 55364 3516 55370 3528
rect 55401 3519 55459 3525
rect 55401 3516 55413 3519
rect 55364 3488 55413 3516
rect 55364 3476 55370 3488
rect 55401 3485 55413 3488
rect 55447 3485 55459 3519
rect 55401 3479 55459 3485
rect 55582 3476 55588 3528
rect 55640 3516 55646 3528
rect 56045 3519 56103 3525
rect 56045 3516 56057 3519
rect 55640 3488 56057 3516
rect 55640 3476 55646 3488
rect 56045 3485 56057 3488
rect 56091 3485 56103 3519
rect 56045 3479 56103 3485
rect 56410 3476 56416 3528
rect 56468 3516 56474 3528
rect 56689 3519 56747 3525
rect 56689 3516 56701 3519
rect 56468 3488 56701 3516
rect 56468 3476 56474 3488
rect 56689 3485 56701 3488
rect 56735 3485 56747 3519
rect 56689 3479 56747 3485
rect 57238 3476 57244 3528
rect 57296 3516 57302 3528
rect 57333 3519 57391 3525
rect 57333 3516 57345 3519
rect 57296 3488 57345 3516
rect 57296 3476 57302 3488
rect 57333 3485 57345 3488
rect 57379 3485 57391 3519
rect 57333 3479 57391 3485
rect 57514 3476 57520 3528
rect 57572 3516 57578 3528
rect 57977 3519 58035 3525
rect 57977 3516 57989 3519
rect 57572 3488 57989 3516
rect 57572 3476 57578 3488
rect 57977 3485 57989 3488
rect 58023 3485 58035 3519
rect 57977 3479 58035 3485
rect 16298 3448 16304 3460
rect 16040 3420 16304 3448
rect 16298 3408 16304 3420
rect 16356 3408 16362 3460
rect 16393 3451 16451 3457
rect 16393 3417 16405 3451
rect 16439 3448 16451 3451
rect 18334 3451 18392 3457
rect 18334 3448 18346 3451
rect 16439 3420 18346 3448
rect 16439 3417 16451 3420
rect 16393 3411 16451 3417
rect 18334 3417 18346 3420
rect 18380 3417 18392 3451
rect 18334 3411 18392 3417
rect 20622 3408 20628 3460
rect 20680 3448 20686 3460
rect 24026 3448 24032 3460
rect 20680 3420 24032 3448
rect 20680 3408 20686 3420
rect 24026 3408 24032 3420
rect 24084 3408 24090 3460
rect 11848 3352 14412 3380
rect 15105 3383 15163 3389
rect 11848 3340 11854 3352
rect 15105 3349 15117 3383
rect 15151 3380 15163 3383
rect 16758 3380 16764 3392
rect 15151 3352 16764 3380
rect 15151 3349 15163 3352
rect 15105 3343 15163 3349
rect 16758 3340 16764 3352
rect 16816 3340 16822 3392
rect 18966 3340 18972 3392
rect 19024 3380 19030 3392
rect 19337 3383 19395 3389
rect 19337 3380 19349 3383
rect 19024 3352 19349 3380
rect 19024 3340 19030 3352
rect 19337 3349 19349 3352
rect 19383 3349 19395 3383
rect 19337 3343 19395 3349
rect 21358 3340 21364 3392
rect 21416 3380 21422 3392
rect 24670 3380 24676 3392
rect 21416 3352 24676 3380
rect 21416 3340 21422 3352
rect 24670 3340 24676 3352
rect 24728 3340 24734 3392
rect 24946 3340 24952 3392
rect 25004 3380 25010 3392
rect 25041 3383 25099 3389
rect 25041 3380 25053 3383
rect 25004 3352 25053 3380
rect 25004 3340 25010 3352
rect 25041 3349 25053 3352
rect 25087 3349 25099 3383
rect 25041 3343 25099 3349
rect 1104 3290 68816 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 50294 3290
rect 50346 3238 50358 3290
rect 50410 3238 50422 3290
rect 50474 3238 50486 3290
rect 50538 3238 50550 3290
rect 50602 3238 68816 3290
rect 1104 3216 68816 3238
rect 3053 3179 3111 3185
rect 3053 3145 3065 3179
rect 3099 3176 3111 3179
rect 3878 3176 3884 3188
rect 3099 3148 3884 3176
rect 3099 3145 3111 3148
rect 3053 3139 3111 3145
rect 3878 3136 3884 3148
rect 3936 3136 3942 3188
rect 4062 3136 4068 3188
rect 4120 3176 4126 3188
rect 4709 3179 4767 3185
rect 4120 3148 4200 3176
rect 4120 3136 4126 3148
rect 4062 3040 4068 3052
rect 4023 3012 4068 3040
rect 4062 3000 4068 3012
rect 4120 3000 4126 3052
rect 4172 3040 4200 3148
rect 4709 3145 4721 3179
rect 4755 3176 4767 3179
rect 6822 3176 6828 3188
rect 4755 3148 6828 3176
rect 4755 3145 4767 3148
rect 4709 3139 4767 3145
rect 6822 3136 6828 3148
rect 6880 3136 6886 3188
rect 10689 3179 10747 3185
rect 10689 3176 10701 3179
rect 6932 3148 10701 3176
rect 4522 3108 4528 3120
rect 4448 3080 4528 3108
rect 4448 3049 4476 3080
rect 4522 3068 4528 3080
rect 4580 3068 4586 3120
rect 4614 3068 4620 3120
rect 4672 3108 4678 3120
rect 5902 3108 5908 3120
rect 4672 3080 5304 3108
rect 4672 3068 4678 3080
rect 4228 3043 4286 3049
rect 4228 3040 4240 3043
rect 4172 3012 4240 3040
rect 4228 3009 4240 3012
rect 4274 3009 4286 3043
rect 4228 3003 4286 3009
rect 4328 3043 4386 3049
rect 4328 3009 4340 3043
rect 4374 3009 4386 3043
rect 4328 3003 4386 3009
rect 4433 3043 4491 3049
rect 4433 3009 4445 3043
rect 4479 3009 4491 3043
rect 5166 3040 5172 3052
rect 5127 3012 5172 3040
rect 4433 3003 4491 3009
rect 4356 2972 4384 3003
rect 5166 3000 5172 3012
rect 5224 3000 5230 3052
rect 5276 3040 5304 3080
rect 5598 3080 5908 3108
rect 5332 3043 5390 3049
rect 5332 3040 5344 3043
rect 5276 3012 5344 3040
rect 5332 3009 5344 3012
rect 5378 3009 5390 3043
rect 5332 3003 5390 3009
rect 5442 3000 5448 3052
rect 5500 3040 5506 3052
rect 5598 3049 5626 3080
rect 5902 3068 5908 3080
rect 5960 3068 5966 3120
rect 5583 3043 5641 3049
rect 5500 3012 5545 3040
rect 5500 3000 5506 3012
rect 5583 3009 5595 3043
rect 5629 3009 5641 3043
rect 6730 3040 6736 3052
rect 5583 3003 5641 3009
rect 5736 3012 6736 3040
rect 5460 2972 5488 3000
rect 4356 2944 5488 2972
rect 3513 2839 3571 2845
rect 3513 2805 3525 2839
rect 3559 2836 3571 2839
rect 5736 2836 5764 3012
rect 6730 3000 6736 3012
rect 6788 3000 6794 3052
rect 5902 2932 5908 2984
rect 5960 2972 5966 2984
rect 6932 2972 6960 3148
rect 10689 3145 10701 3148
rect 10735 3176 10747 3179
rect 13722 3176 13728 3188
rect 10735 3148 13728 3176
rect 10735 3145 10747 3148
rect 10689 3139 10747 3145
rect 13722 3136 13728 3148
rect 13780 3136 13786 3188
rect 14090 3176 14096 3188
rect 13832 3148 14096 3176
rect 9398 3108 9404 3120
rect 7208 3080 9404 3108
rect 7208 3052 7236 3080
rect 7190 3040 7196 3052
rect 7103 3012 7196 3040
rect 7190 3000 7196 3012
rect 7248 3000 7254 3052
rect 7282 3000 7288 3052
rect 7340 3040 7346 3052
rect 7449 3043 7507 3049
rect 7449 3040 7461 3043
rect 7340 3012 7461 3040
rect 7340 3000 7346 3012
rect 7449 3009 7461 3012
rect 7495 3009 7507 3043
rect 7449 3003 7507 3009
rect 7742 3000 7748 3052
rect 7800 3040 7806 3052
rect 8570 3040 8576 3052
rect 7800 3012 8576 3040
rect 7800 3000 7806 3012
rect 8570 3000 8576 3012
rect 8628 3000 8634 3052
rect 9324 3049 9352 3080
rect 9398 3068 9404 3080
rect 9456 3068 9462 3120
rect 9766 3068 9772 3120
rect 9824 3068 9830 3120
rect 11882 3068 11888 3120
rect 11940 3108 11946 3120
rect 11940 3080 12940 3108
rect 11940 3068 11946 3080
rect 9309 3043 9367 3049
rect 9309 3009 9321 3043
rect 9355 3009 9367 3043
rect 9565 3043 9623 3049
rect 9565 3040 9577 3043
rect 9309 3003 9367 3009
rect 9416 3012 9577 3040
rect 9416 2972 9444 3012
rect 9565 3009 9577 3012
rect 9611 3009 9623 3043
rect 9784 3040 9812 3068
rect 11977 3043 12035 3049
rect 11977 3040 11989 3043
rect 9784 3012 11989 3040
rect 9565 3003 9623 3009
rect 11977 3009 11989 3012
rect 12023 3009 12035 3043
rect 11977 3003 12035 3009
rect 12158 3000 12164 3052
rect 12216 3040 12222 3052
rect 12912 3049 12940 3080
rect 13538 3049 13544 3052
rect 12713 3043 12771 3049
rect 12713 3040 12725 3043
rect 12216 3012 12725 3040
rect 12216 3000 12222 3012
rect 12713 3009 12725 3012
rect 12759 3009 12771 3043
rect 12713 3003 12771 3009
rect 12897 3043 12955 3049
rect 12897 3009 12909 3043
rect 12943 3009 12955 3043
rect 12897 3003 12955 3009
rect 13529 3043 13544 3049
rect 13529 3009 13541 3043
rect 13529 3003 13544 3009
rect 13538 3000 13544 3003
rect 13596 3000 13602 3052
rect 13630 3000 13636 3052
rect 13688 3043 13694 3052
rect 13832 3049 13860 3148
rect 14090 3136 14096 3148
rect 14148 3136 14154 3188
rect 15102 3136 15108 3188
rect 15160 3176 15166 3188
rect 16114 3176 16120 3188
rect 15160 3148 16120 3176
rect 15160 3136 15166 3148
rect 16114 3136 16120 3148
rect 16172 3136 16178 3188
rect 17957 3179 18015 3185
rect 17957 3145 17969 3179
rect 18003 3176 18015 3179
rect 21266 3176 21272 3188
rect 18003 3148 21272 3176
rect 18003 3145 18015 3148
rect 17957 3139 18015 3145
rect 21266 3136 21272 3148
rect 21324 3136 21330 3188
rect 14185 3111 14243 3117
rect 14185 3077 14197 3111
rect 14231 3108 14243 3111
rect 15758 3111 15816 3117
rect 15758 3108 15770 3111
rect 14231 3080 15770 3108
rect 14231 3077 14243 3080
rect 14185 3071 14243 3077
rect 15758 3077 15770 3080
rect 15804 3077 15816 3111
rect 15758 3071 15816 3077
rect 16298 3068 16304 3120
rect 16356 3108 16362 3120
rect 18684 3111 18742 3117
rect 16356 3080 16988 3108
rect 16356 3068 16362 3080
rect 13725 3043 13783 3049
rect 13688 3015 13737 3043
rect 13688 3000 13694 3015
rect 13725 3009 13737 3015
rect 13771 3009 13783 3043
rect 13725 3003 13783 3009
rect 13817 3043 13875 3049
rect 13817 3009 13829 3043
rect 13863 3009 13875 3043
rect 13817 3003 13875 3009
rect 13909 3043 13967 3049
rect 13909 3009 13921 3043
rect 13955 3024 13967 3043
rect 13955 3009 14044 3024
rect 13909 3003 14044 3009
rect 13924 2996 14044 3003
rect 15470 3000 15476 3052
rect 15528 3040 15534 3052
rect 16669 3043 16727 3049
rect 16669 3040 16681 3043
rect 15528 3012 16681 3040
rect 15528 3000 15534 3012
rect 16669 3009 16681 3012
rect 16715 3009 16727 3043
rect 16850 3040 16856 3052
rect 16811 3012 16856 3040
rect 16669 3003 16727 3009
rect 16850 3000 16856 3012
rect 16908 3000 16914 3052
rect 16960 3049 16988 3080
rect 18684 3077 18696 3111
rect 18730 3108 18742 3111
rect 20806 3108 20812 3120
rect 18730 3080 20812 3108
rect 18730 3077 18742 3080
rect 18684 3071 18742 3077
rect 20806 3068 20812 3080
rect 20864 3068 20870 3120
rect 16945 3043 17003 3049
rect 16945 3009 16957 3043
rect 16991 3009 17003 3043
rect 16945 3003 17003 3009
rect 17037 3043 17095 3049
rect 17037 3009 17049 3043
rect 17083 3040 17095 3043
rect 17218 3040 17224 3052
rect 17083 3012 17224 3040
rect 17083 3009 17095 3012
rect 17037 3003 17095 3009
rect 17218 3000 17224 3012
rect 17276 3000 17282 3052
rect 17773 3043 17831 3049
rect 17773 3009 17785 3043
rect 17819 3040 17831 3043
rect 20533 3043 20591 3049
rect 17819 3012 20484 3040
rect 17819 3009 17831 3012
rect 17773 3003 17831 3009
rect 5960 2944 6960 2972
rect 8404 2944 9444 2972
rect 14016 2972 14044 2996
rect 16025 2975 16083 2981
rect 14016 2944 14412 2972
rect 5960 2932 5966 2944
rect 5813 2907 5871 2913
rect 5813 2873 5825 2907
rect 5859 2904 5871 2907
rect 5859 2876 7236 2904
rect 5859 2873 5871 2876
rect 5813 2867 5871 2873
rect 3559 2808 5764 2836
rect 3559 2805 3571 2808
rect 3513 2799 3571 2805
rect 5994 2796 6000 2848
rect 6052 2836 6058 2848
rect 6549 2839 6607 2845
rect 6549 2836 6561 2839
rect 6052 2808 6561 2836
rect 6052 2796 6058 2808
rect 6549 2805 6561 2808
rect 6595 2805 6607 2839
rect 7208 2836 7236 2876
rect 8404 2836 8432 2944
rect 14384 2848 14412 2944
rect 16025 2941 16037 2975
rect 16071 2972 16083 2975
rect 18046 2972 18052 2984
rect 16071 2944 18052 2972
rect 16071 2941 16083 2944
rect 16025 2935 16083 2941
rect 18046 2932 18052 2944
rect 18104 2972 18110 2984
rect 18414 2972 18420 2984
rect 18104 2944 18420 2972
rect 18104 2932 18110 2944
rect 18414 2932 18420 2944
rect 18472 2932 18478 2984
rect 20456 2972 20484 3012
rect 20533 3009 20545 3043
rect 20579 3040 20591 3043
rect 20714 3040 20720 3052
rect 20579 3012 20720 3040
rect 20579 3009 20591 3012
rect 20533 3003 20591 3009
rect 20714 3000 20720 3012
rect 20772 3000 20778 3052
rect 21269 2975 21327 2981
rect 20456 2944 21220 2972
rect 16114 2864 16120 2916
rect 16172 2904 16178 2916
rect 18138 2904 18144 2916
rect 16172 2876 18144 2904
rect 16172 2864 16178 2876
rect 18138 2864 18144 2876
rect 18196 2864 18202 2916
rect 19426 2864 19432 2916
rect 19484 2904 19490 2916
rect 20349 2907 20407 2913
rect 20349 2904 20361 2907
rect 19484 2876 20361 2904
rect 19484 2864 19490 2876
rect 20349 2873 20361 2876
rect 20395 2873 20407 2907
rect 20349 2867 20407 2873
rect 20898 2864 20904 2916
rect 20956 2864 20962 2916
rect 7208 2808 8432 2836
rect 6549 2799 6607 2805
rect 8570 2796 8576 2848
rect 8628 2836 8634 2848
rect 10870 2836 10876 2848
rect 8628 2808 10876 2836
rect 8628 2796 8634 2808
rect 10870 2796 10876 2808
rect 10928 2796 10934 2848
rect 12158 2836 12164 2848
rect 12119 2808 12164 2836
rect 12158 2796 12164 2808
rect 12216 2796 12222 2848
rect 12805 2839 12863 2845
rect 12805 2805 12817 2839
rect 12851 2836 12863 2839
rect 12894 2836 12900 2848
rect 12851 2808 12900 2836
rect 12851 2805 12863 2808
rect 12805 2799 12863 2805
rect 12894 2796 12900 2808
rect 12952 2796 12958 2848
rect 14366 2796 14372 2848
rect 14424 2836 14430 2848
rect 14645 2839 14703 2845
rect 14645 2836 14657 2839
rect 14424 2808 14657 2836
rect 14424 2796 14430 2808
rect 14645 2805 14657 2808
rect 14691 2805 14703 2839
rect 14645 2799 14703 2805
rect 15286 2796 15292 2848
rect 15344 2836 15350 2848
rect 17034 2836 17040 2848
rect 15344 2808 17040 2836
rect 15344 2796 15350 2808
rect 17034 2796 17040 2808
rect 17092 2796 17098 2848
rect 17313 2839 17371 2845
rect 17313 2805 17325 2839
rect 17359 2836 17371 2839
rect 17678 2836 17684 2848
rect 17359 2808 17684 2836
rect 17359 2805 17371 2808
rect 17313 2799 17371 2805
rect 17678 2796 17684 2808
rect 17736 2796 17742 2848
rect 19797 2839 19855 2845
rect 19797 2805 19809 2839
rect 19843 2836 19855 2839
rect 20916 2836 20944 2864
rect 19843 2808 20944 2836
rect 21192 2836 21220 2944
rect 21269 2941 21281 2975
rect 21315 2972 21327 2975
rect 22186 2972 22192 2984
rect 21315 2944 22192 2972
rect 21315 2941 21327 2944
rect 21269 2935 21327 2941
rect 22186 2932 22192 2944
rect 22244 2932 22250 2984
rect 25133 2975 25191 2981
rect 25133 2941 25145 2975
rect 25179 2972 25191 2975
rect 25222 2972 25228 2984
rect 25179 2944 25228 2972
rect 25179 2941 25191 2944
rect 25133 2935 25191 2941
rect 25222 2932 25228 2944
rect 25280 2932 25286 2984
rect 37918 2932 37924 2984
rect 37976 2972 37982 2984
rect 38565 2975 38623 2981
rect 38565 2972 38577 2975
rect 37976 2944 38577 2972
rect 37976 2932 37982 2944
rect 38565 2941 38577 2944
rect 38611 2941 38623 2975
rect 38565 2935 38623 2941
rect 39574 2932 39580 2984
rect 39632 2972 39638 2984
rect 40497 2975 40555 2981
rect 40497 2972 40509 2975
rect 39632 2944 40509 2972
rect 39632 2932 39638 2944
rect 40497 2941 40509 2944
rect 40543 2941 40555 2975
rect 40497 2935 40555 2941
rect 43438 2932 43444 2984
rect 43496 2972 43502 2984
rect 44361 2975 44419 2981
rect 44361 2972 44373 2975
rect 43496 2944 44373 2972
rect 43496 2932 43502 2944
rect 44361 2941 44373 2944
rect 44407 2941 44419 2975
rect 44361 2935 44419 2941
rect 47302 2932 47308 2984
rect 47360 2972 47366 2984
rect 48225 2975 48283 2981
rect 48225 2972 48237 2975
rect 47360 2944 48237 2972
rect 47360 2932 47366 2944
rect 48225 2941 48237 2944
rect 48271 2941 48283 2975
rect 48225 2935 48283 2941
rect 49234 2932 49240 2984
rect 49292 2972 49298 2984
rect 50157 2975 50215 2981
rect 50157 2972 50169 2975
rect 49292 2944 50169 2972
rect 49292 2932 49298 2944
rect 50157 2941 50169 2944
rect 50203 2941 50215 2975
rect 50157 2935 50215 2941
rect 55030 2932 55036 2984
rect 55088 2972 55094 2984
rect 55953 2975 56011 2981
rect 55953 2972 55965 2975
rect 55088 2944 55965 2972
rect 55088 2932 55094 2944
rect 55953 2941 55965 2944
rect 55999 2941 56011 2975
rect 55953 2935 56011 2941
rect 38470 2864 38476 2916
rect 38528 2904 38534 2916
rect 39209 2907 39267 2913
rect 39209 2904 39221 2907
rect 38528 2876 39221 2904
rect 38528 2864 38534 2876
rect 39209 2873 39221 2876
rect 39255 2873 39267 2907
rect 39209 2867 39267 2873
rect 40402 2864 40408 2916
rect 40460 2904 40466 2916
rect 41141 2907 41199 2913
rect 41141 2904 41153 2907
rect 40460 2876 41153 2904
rect 40460 2864 40466 2876
rect 41141 2873 41153 2876
rect 41187 2873 41199 2907
rect 41141 2867 41199 2873
rect 42334 2864 42340 2916
rect 42392 2904 42398 2916
rect 43073 2907 43131 2913
rect 43073 2904 43085 2907
rect 42392 2876 43085 2904
rect 42392 2864 42398 2876
rect 43073 2873 43085 2876
rect 43119 2873 43131 2907
rect 43073 2867 43131 2873
rect 44266 2864 44272 2916
rect 44324 2904 44330 2916
rect 45005 2907 45063 2913
rect 45005 2904 45017 2907
rect 44324 2876 45017 2904
rect 44324 2864 44330 2876
rect 45005 2873 45017 2876
rect 45051 2873 45063 2907
rect 45005 2867 45063 2873
rect 45370 2864 45376 2916
rect 45428 2904 45434 2916
rect 46293 2907 46351 2913
rect 46293 2904 46305 2907
rect 45428 2876 46305 2904
rect 45428 2864 45434 2876
rect 46293 2873 46305 2876
rect 46339 2873 46351 2907
rect 46293 2867 46351 2873
rect 48130 2864 48136 2916
rect 48188 2904 48194 2916
rect 48869 2907 48927 2913
rect 48869 2904 48881 2907
rect 48188 2876 48881 2904
rect 48188 2864 48194 2876
rect 48869 2873 48881 2876
rect 48915 2873 48927 2907
rect 48869 2867 48927 2873
rect 50062 2864 50068 2916
rect 50120 2904 50126 2916
rect 50801 2907 50859 2913
rect 50801 2904 50813 2907
rect 50120 2876 50813 2904
rect 50120 2864 50126 2876
rect 50801 2873 50813 2876
rect 50847 2873 50859 2907
rect 50801 2867 50859 2873
rect 52546 2864 52552 2916
rect 52604 2904 52610 2916
rect 53377 2907 53435 2913
rect 53377 2904 53389 2907
rect 52604 2876 53389 2904
rect 52604 2864 52610 2876
rect 53377 2873 53389 2876
rect 53423 2873 53435 2907
rect 53377 2867 53435 2873
rect 53926 2864 53932 2916
rect 53984 2904 53990 2916
rect 54665 2907 54723 2913
rect 54665 2904 54677 2907
rect 53984 2876 54677 2904
rect 53984 2864 53990 2876
rect 54665 2873 54677 2876
rect 54711 2873 54723 2907
rect 54665 2867 54723 2873
rect 57606 2864 57612 2916
rect 57664 2904 57670 2916
rect 58529 2907 58587 2913
rect 58529 2904 58541 2907
rect 57664 2876 58541 2904
rect 57664 2864 57670 2876
rect 58529 2873 58541 2876
rect 58575 2873 58587 2907
rect 58529 2867 58587 2873
rect 21266 2836 21272 2848
rect 21192 2808 21272 2836
rect 19843 2805 19855 2808
rect 19797 2799 19855 2805
rect 21266 2796 21272 2808
rect 21324 2796 21330 2848
rect 21634 2796 21640 2848
rect 21692 2836 21698 2848
rect 21818 2836 21824 2848
rect 21692 2808 21824 2836
rect 21692 2796 21698 2808
rect 21818 2796 21824 2808
rect 21876 2796 21882 2848
rect 22557 2839 22615 2845
rect 22557 2805 22569 2839
rect 22603 2836 22615 2839
rect 23014 2836 23020 2848
rect 22603 2808 23020 2836
rect 22603 2805 22615 2808
rect 22557 2799 22615 2805
rect 23014 2796 23020 2808
rect 23072 2796 23078 2848
rect 23201 2839 23259 2845
rect 23201 2805 23213 2839
rect 23247 2836 23259 2839
rect 23290 2836 23296 2848
rect 23247 2808 23296 2836
rect 23247 2805 23259 2808
rect 23201 2799 23259 2805
rect 23290 2796 23296 2808
rect 23348 2796 23354 2848
rect 23845 2839 23903 2845
rect 23845 2805 23857 2839
rect 23891 2836 23903 2839
rect 24118 2836 24124 2848
rect 23891 2808 24124 2836
rect 23891 2805 23903 2808
rect 23845 2799 23903 2805
rect 24118 2796 24124 2808
rect 24176 2796 24182 2848
rect 24489 2839 24547 2845
rect 24489 2805 24501 2839
rect 24535 2836 24547 2839
rect 24670 2836 24676 2848
rect 24535 2808 24676 2836
rect 24535 2805 24547 2808
rect 24489 2799 24547 2805
rect 24670 2796 24676 2808
rect 24728 2796 24734 2848
rect 25774 2836 25780 2848
rect 25735 2808 25780 2836
rect 25774 2796 25780 2808
rect 25832 2796 25838 2848
rect 26237 2839 26295 2845
rect 26237 2805 26249 2839
rect 26283 2836 26295 2839
rect 26326 2836 26332 2848
rect 26283 2808 26332 2836
rect 26283 2805 26295 2808
rect 26237 2799 26295 2805
rect 26326 2796 26332 2808
rect 26384 2796 26390 2848
rect 26418 2796 26424 2848
rect 26476 2836 26482 2848
rect 26973 2839 27031 2845
rect 26973 2836 26985 2839
rect 26476 2808 26985 2836
rect 26476 2796 26482 2808
rect 26973 2805 26985 2808
rect 27019 2805 27031 2839
rect 26973 2799 27031 2805
rect 27709 2839 27767 2845
rect 27709 2805 27721 2839
rect 27755 2836 27767 2839
rect 27982 2836 27988 2848
rect 27755 2808 27988 2836
rect 27755 2805 27767 2808
rect 27709 2799 27767 2805
rect 27982 2796 27988 2808
rect 28040 2796 28046 2848
rect 28353 2839 28411 2845
rect 28353 2805 28365 2839
rect 28399 2836 28411 2839
rect 28534 2836 28540 2848
rect 28399 2808 28540 2836
rect 28399 2805 28411 2808
rect 28353 2799 28411 2805
rect 28534 2796 28540 2808
rect 28592 2796 28598 2848
rect 28997 2839 29055 2845
rect 28997 2805 29009 2839
rect 29043 2836 29055 2839
rect 29086 2836 29092 2848
rect 29043 2808 29092 2836
rect 29043 2805 29055 2808
rect 28997 2799 29055 2805
rect 29086 2796 29092 2808
rect 29144 2796 29150 2848
rect 29641 2839 29699 2845
rect 29641 2805 29653 2839
rect 29687 2836 29699 2839
rect 29914 2836 29920 2848
rect 29687 2808 29920 2836
rect 29687 2805 29699 2808
rect 29641 2799 29699 2805
rect 29914 2796 29920 2808
rect 29972 2796 29978 2848
rect 30285 2839 30343 2845
rect 30285 2805 30297 2839
rect 30331 2836 30343 2839
rect 30466 2836 30472 2848
rect 30331 2808 30472 2836
rect 30331 2805 30343 2808
rect 30285 2799 30343 2805
rect 30466 2796 30472 2808
rect 30524 2796 30530 2848
rect 30929 2839 30987 2845
rect 30929 2805 30941 2839
rect 30975 2836 30987 2839
rect 31018 2836 31024 2848
rect 30975 2808 31024 2836
rect 30975 2805 30987 2808
rect 30929 2799 30987 2805
rect 31018 2796 31024 2808
rect 31076 2796 31082 2848
rect 31573 2839 31631 2845
rect 31573 2805 31585 2839
rect 31619 2836 31631 2839
rect 31846 2836 31852 2848
rect 31619 2808 31852 2836
rect 31619 2805 31631 2808
rect 31573 2799 31631 2805
rect 31846 2796 31852 2808
rect 31904 2796 31910 2848
rect 32493 2839 32551 2845
rect 32493 2805 32505 2839
rect 32539 2836 32551 2839
rect 32674 2836 32680 2848
rect 32539 2808 32680 2836
rect 32539 2805 32551 2808
rect 32493 2799 32551 2805
rect 32674 2796 32680 2808
rect 32732 2796 32738 2848
rect 33137 2839 33195 2845
rect 33137 2805 33149 2839
rect 33183 2836 33195 2839
rect 33226 2836 33232 2848
rect 33183 2808 33232 2836
rect 33183 2805 33195 2808
rect 33137 2799 33195 2805
rect 33226 2796 33232 2808
rect 33284 2796 33290 2848
rect 33778 2836 33784 2848
rect 33739 2808 33784 2836
rect 33778 2796 33784 2808
rect 33836 2796 33842 2848
rect 34241 2839 34299 2845
rect 34241 2805 34253 2839
rect 34287 2836 34299 2839
rect 34330 2836 34336 2848
rect 34287 2808 34336 2836
rect 34287 2805 34299 2808
rect 34241 2799 34299 2805
rect 34330 2796 34336 2808
rect 34388 2796 34394 2848
rect 34790 2796 34796 2848
rect 34848 2836 34854 2848
rect 34885 2839 34943 2845
rect 34885 2836 34897 2839
rect 34848 2808 34897 2836
rect 34848 2796 34854 2808
rect 34885 2805 34897 2808
rect 34931 2805 34943 2839
rect 34885 2799 34943 2805
rect 35434 2796 35440 2848
rect 35492 2836 35498 2848
rect 35529 2839 35587 2845
rect 35529 2836 35541 2839
rect 35492 2808 35541 2836
rect 35492 2796 35498 2808
rect 35529 2805 35541 2808
rect 35575 2805 35587 2839
rect 35529 2799 35587 2805
rect 36262 2796 36268 2848
rect 36320 2836 36326 2848
rect 36357 2839 36415 2845
rect 36357 2836 36369 2839
rect 36320 2808 36369 2836
rect 36320 2796 36326 2808
rect 36357 2805 36369 2808
rect 36403 2805 36415 2839
rect 36357 2799 36415 2805
rect 36814 2796 36820 2848
rect 36872 2836 36878 2848
rect 37277 2839 37335 2845
rect 37277 2836 37289 2839
rect 36872 2808 37289 2836
rect 36872 2796 36878 2808
rect 37277 2805 37289 2808
rect 37323 2805 37335 2839
rect 37277 2799 37335 2805
rect 37366 2796 37372 2848
rect 37424 2836 37430 2848
rect 37921 2839 37979 2845
rect 37921 2836 37933 2839
rect 37424 2808 37933 2836
rect 37424 2796 37430 2808
rect 37921 2805 37933 2808
rect 37967 2805 37979 2839
rect 37921 2799 37979 2805
rect 39022 2796 39028 2848
rect 39080 2836 39086 2848
rect 39853 2839 39911 2845
rect 39853 2836 39865 2839
rect 39080 2808 39865 2836
rect 39080 2796 39086 2808
rect 39853 2805 39865 2808
rect 39899 2805 39911 2839
rect 39853 2799 39911 2805
rect 41506 2796 41512 2848
rect 41564 2836 41570 2848
rect 42429 2839 42487 2845
rect 42429 2836 42441 2839
rect 41564 2808 42441 2836
rect 41564 2796 41570 2808
rect 42429 2805 42441 2808
rect 42475 2805 42487 2839
rect 42429 2799 42487 2805
rect 42886 2796 42892 2848
rect 42944 2836 42950 2848
rect 43717 2839 43775 2845
rect 43717 2836 43729 2839
rect 42944 2808 43729 2836
rect 42944 2796 42950 2808
rect 43717 2805 43729 2808
rect 43763 2805 43775 2839
rect 43717 2799 43775 2805
rect 44818 2796 44824 2848
rect 44876 2836 44882 2848
rect 45649 2839 45707 2845
rect 45649 2836 45661 2839
rect 44876 2808 45661 2836
rect 44876 2796 44882 2808
rect 45649 2805 45661 2808
rect 45695 2805 45707 2839
rect 45649 2799 45707 2805
rect 46750 2796 46756 2848
rect 46808 2836 46814 2848
rect 47581 2839 47639 2845
rect 47581 2836 47593 2839
rect 46808 2808 47593 2836
rect 46808 2796 46814 2808
rect 47581 2805 47593 2808
rect 47627 2805 47639 2839
rect 47581 2799 47639 2805
rect 48682 2796 48688 2848
rect 48740 2836 48746 2848
rect 49513 2839 49571 2845
rect 49513 2836 49525 2839
rect 48740 2808 49525 2836
rect 48740 2796 48746 2808
rect 49513 2805 49525 2808
rect 49559 2805 49571 2839
rect 49513 2799 49571 2805
rect 50706 2796 50712 2848
rect 50764 2836 50770 2848
rect 51445 2839 51503 2845
rect 51445 2836 51457 2839
rect 50764 2808 51457 2836
rect 50764 2796 50770 2808
rect 51445 2805 51457 2808
rect 51491 2805 51503 2839
rect 51445 2799 51503 2805
rect 51994 2796 52000 2848
rect 52052 2836 52058 2848
rect 52733 2839 52791 2845
rect 52733 2836 52745 2839
rect 52052 2808 52745 2836
rect 52052 2796 52058 2808
rect 52733 2805 52745 2808
rect 52779 2805 52791 2839
rect 52733 2799 52791 2805
rect 53098 2796 53104 2848
rect 53156 2836 53162 2848
rect 54021 2839 54079 2845
rect 54021 2836 54033 2839
rect 53156 2808 54033 2836
rect 53156 2796 53162 2808
rect 54021 2805 54033 2808
rect 54067 2805 54079 2839
rect 54021 2799 54079 2805
rect 54478 2796 54484 2848
rect 54536 2836 54542 2848
rect 55309 2839 55367 2845
rect 55309 2836 55321 2839
rect 54536 2808 55321 2836
rect 54536 2796 54542 2808
rect 55309 2805 55321 2808
rect 55355 2805 55367 2839
rect 55309 2799 55367 2805
rect 55858 2796 55864 2848
rect 55916 2836 55922 2848
rect 56597 2839 56655 2845
rect 56597 2836 56609 2839
rect 55916 2808 56609 2836
rect 55916 2796 55922 2808
rect 56597 2805 56609 2808
rect 56643 2805 56655 2839
rect 56597 2799 56655 2805
rect 56962 2796 56968 2848
rect 57020 2836 57026 2848
rect 57885 2839 57943 2845
rect 57885 2836 57897 2839
rect 57020 2808 57897 2836
rect 57020 2796 57026 2808
rect 57885 2805 57897 2808
rect 57931 2805 57943 2839
rect 57885 2799 57943 2805
rect 1104 2746 68816 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 65654 2746
rect 65706 2694 65718 2746
rect 65770 2694 65782 2746
rect 65834 2694 65846 2746
rect 65898 2694 65910 2746
rect 65962 2694 68816 2746
rect 1104 2672 68816 2694
rect 4525 2635 4583 2641
rect 4525 2601 4537 2635
rect 4571 2632 4583 2635
rect 4706 2632 4712 2644
rect 4571 2604 4712 2632
rect 4571 2601 4583 2604
rect 4525 2595 4583 2601
rect 4706 2592 4712 2604
rect 4764 2592 4770 2644
rect 5810 2592 5816 2644
rect 5868 2632 5874 2644
rect 6365 2635 6423 2641
rect 6365 2632 6377 2635
rect 5868 2604 6377 2632
rect 5868 2592 5874 2604
rect 6365 2601 6377 2604
rect 6411 2601 6423 2635
rect 7190 2632 7196 2644
rect 6365 2595 6423 2601
rect 7024 2604 7196 2632
rect 4065 2567 4123 2573
rect 4065 2533 4077 2567
rect 4111 2564 4123 2567
rect 4890 2564 4896 2576
rect 4111 2536 4896 2564
rect 4111 2533 4123 2536
rect 4065 2527 4123 2533
rect 4890 2524 4896 2536
rect 4948 2524 4954 2576
rect 7024 2505 7052 2604
rect 7190 2592 7196 2604
rect 7248 2592 7254 2644
rect 9309 2635 9367 2641
rect 9309 2601 9321 2635
rect 9355 2632 9367 2635
rect 13446 2632 13452 2644
rect 9355 2604 13452 2632
rect 9355 2601 9367 2604
rect 9309 2595 9367 2601
rect 13446 2592 13452 2604
rect 13504 2592 13510 2644
rect 14553 2635 14611 2641
rect 14553 2601 14565 2635
rect 14599 2632 14611 2635
rect 15286 2632 15292 2644
rect 14599 2604 15292 2632
rect 14599 2601 14611 2604
rect 14553 2595 14611 2601
rect 15286 2592 15292 2604
rect 15344 2592 15350 2644
rect 17037 2635 17095 2641
rect 17037 2601 17049 2635
rect 17083 2632 17095 2635
rect 17218 2632 17224 2644
rect 17083 2604 17224 2632
rect 17083 2601 17095 2604
rect 17037 2595 17095 2601
rect 17218 2592 17224 2604
rect 17276 2592 17282 2644
rect 19058 2632 19064 2644
rect 17420 2604 19064 2632
rect 8389 2567 8447 2573
rect 8389 2533 8401 2567
rect 8435 2564 8447 2567
rect 11977 2567 12035 2573
rect 8435 2536 11836 2564
rect 8435 2533 8447 2536
rect 8389 2527 8447 2533
rect 7009 2499 7067 2505
rect 6472 2468 6776 2496
rect 3878 2428 3884 2440
rect 3839 2400 3884 2428
rect 3878 2388 3884 2400
rect 3936 2388 3942 2440
rect 4706 2428 4712 2440
rect 4667 2400 4712 2428
rect 4706 2388 4712 2400
rect 4764 2388 4770 2440
rect 5166 2428 5172 2440
rect 5127 2400 5172 2428
rect 5166 2388 5172 2400
rect 5224 2388 5230 2440
rect 5258 2388 5264 2440
rect 5316 2428 5322 2440
rect 5353 2431 5411 2437
rect 5353 2428 5365 2431
rect 5316 2400 5365 2428
rect 5316 2388 5322 2400
rect 5353 2397 5365 2400
rect 5399 2397 5411 2431
rect 5353 2391 5411 2397
rect 5442 2388 5448 2440
rect 5500 2428 5506 2440
rect 5583 2431 5641 2437
rect 5500 2400 5545 2428
rect 5500 2388 5506 2400
rect 5583 2397 5595 2431
rect 5629 2428 5641 2431
rect 6472 2428 6500 2468
rect 5629 2400 6500 2428
rect 5629 2397 5641 2400
rect 5583 2391 5641 2397
rect 6546 2388 6552 2440
rect 6604 2428 6610 2440
rect 6748 2428 6776 2468
rect 7009 2465 7021 2499
rect 7055 2465 7067 2499
rect 7009 2459 7067 2465
rect 8404 2428 8432 2527
rect 11330 2496 11336 2508
rect 10244 2468 11336 2496
rect 6604 2400 6649 2428
rect 6748 2400 8432 2428
rect 9493 2431 9551 2437
rect 6604 2388 6610 2400
rect 9493 2397 9505 2431
rect 9539 2428 9551 2431
rect 9950 2428 9956 2440
rect 9539 2400 9956 2428
rect 9539 2397 9551 2400
rect 9493 2391 9551 2397
rect 9950 2388 9956 2400
rect 10008 2388 10014 2440
rect 10244 2437 10272 2468
rect 11330 2456 11336 2468
rect 11388 2456 11394 2508
rect 10229 2431 10287 2437
rect 10229 2397 10241 2431
rect 10275 2397 10287 2431
rect 10229 2391 10287 2397
rect 10965 2431 11023 2437
rect 10965 2397 10977 2431
rect 11011 2428 11023 2431
rect 11698 2428 11704 2440
rect 11011 2400 11704 2428
rect 11011 2397 11023 2400
rect 10965 2391 11023 2397
rect 11698 2388 11704 2400
rect 11756 2388 11762 2440
rect 11808 2437 11836 2536
rect 11977 2533 11989 2567
rect 12023 2564 12035 2567
rect 12713 2567 12771 2573
rect 12023 2536 12434 2564
rect 12023 2533 12035 2536
rect 11977 2527 12035 2533
rect 12406 2496 12434 2536
rect 12713 2533 12725 2567
rect 12759 2564 12771 2567
rect 15378 2564 15384 2576
rect 12759 2536 15384 2564
rect 12759 2533 12771 2536
rect 12713 2527 12771 2533
rect 15378 2524 15384 2536
rect 15436 2524 15442 2576
rect 15102 2496 15108 2508
rect 12406 2468 15108 2496
rect 15102 2456 15108 2468
rect 15160 2456 15166 2508
rect 16574 2496 16580 2508
rect 15396 2468 16580 2496
rect 11793 2431 11851 2437
rect 11793 2397 11805 2431
rect 11839 2397 11851 2431
rect 12529 2431 12587 2437
rect 12529 2428 12541 2431
rect 11793 2391 11851 2397
rect 12406 2400 12541 2428
rect 2685 2363 2743 2369
rect 2685 2329 2697 2363
rect 2731 2360 2743 2363
rect 4724 2360 4752 2388
rect 2731 2332 4752 2360
rect 5813 2363 5871 2369
rect 2731 2329 2743 2332
rect 2685 2323 2743 2329
rect 5813 2329 5825 2363
rect 5859 2360 5871 2363
rect 7254 2363 7312 2369
rect 7254 2360 7266 2363
rect 5859 2332 7266 2360
rect 5859 2329 5871 2332
rect 5813 2323 5871 2329
rect 7254 2329 7266 2332
rect 7300 2329 7312 2363
rect 7254 2323 7312 2329
rect 10870 2320 10876 2372
rect 10928 2360 10934 2372
rect 12406 2360 12434 2400
rect 12529 2397 12541 2400
rect 12575 2397 12587 2431
rect 12529 2391 12587 2397
rect 12802 2388 12808 2440
rect 12860 2428 12866 2440
rect 13265 2431 13323 2437
rect 13265 2428 13277 2431
rect 12860 2400 13277 2428
rect 12860 2388 12866 2400
rect 13265 2397 13277 2400
rect 13311 2397 13323 2431
rect 14366 2428 14372 2440
rect 14327 2400 14372 2428
rect 13265 2391 13323 2397
rect 14366 2388 14372 2400
rect 14424 2388 14430 2440
rect 15286 2428 15292 2440
rect 15120 2400 15292 2428
rect 10928 2332 12434 2360
rect 10928 2320 10934 2332
rect 3237 2295 3295 2301
rect 3237 2261 3249 2295
rect 3283 2292 3295 2295
rect 6546 2292 6552 2304
rect 3283 2264 6552 2292
rect 3283 2261 3295 2264
rect 3237 2255 3295 2261
rect 6546 2252 6552 2264
rect 6604 2252 6610 2304
rect 10042 2292 10048 2304
rect 10003 2264 10048 2292
rect 10042 2252 10048 2264
rect 10100 2252 10106 2304
rect 10778 2292 10784 2304
rect 10739 2264 10784 2292
rect 10778 2252 10784 2264
rect 10836 2252 10842 2304
rect 13449 2295 13507 2301
rect 13449 2261 13461 2295
rect 13495 2292 13507 2295
rect 15120 2292 15148 2400
rect 15286 2388 15292 2400
rect 15344 2388 15350 2440
rect 15396 2437 15424 2468
rect 16574 2456 16580 2468
rect 16632 2456 16638 2508
rect 15381 2431 15439 2437
rect 15381 2397 15393 2431
rect 15427 2397 15439 2431
rect 15381 2391 15439 2397
rect 16117 2431 16175 2437
rect 16117 2397 16129 2431
rect 16163 2428 16175 2431
rect 17420 2428 17448 2604
rect 19058 2592 19064 2604
rect 19116 2592 19122 2644
rect 20898 2592 20904 2644
rect 20956 2632 20962 2644
rect 22278 2632 22284 2644
rect 20956 2604 22284 2632
rect 20956 2592 20962 2604
rect 22278 2592 22284 2604
rect 22336 2592 22342 2644
rect 19521 2567 19579 2573
rect 19521 2533 19533 2567
rect 19567 2564 19579 2567
rect 20254 2564 20260 2576
rect 19567 2536 20260 2564
rect 19567 2533 19579 2536
rect 19521 2527 19579 2533
rect 20254 2524 20260 2536
rect 20312 2524 20318 2576
rect 21913 2567 21971 2573
rect 21913 2564 21925 2567
rect 20364 2536 21925 2564
rect 18414 2496 18420 2508
rect 18375 2468 18420 2496
rect 18414 2456 18420 2468
rect 18472 2456 18478 2508
rect 20364 2496 20392 2536
rect 21913 2533 21925 2536
rect 21959 2533 21971 2567
rect 21913 2527 21971 2533
rect 23201 2567 23259 2573
rect 23201 2533 23213 2567
rect 23247 2564 23259 2567
rect 23842 2564 23848 2576
rect 23247 2536 23848 2564
rect 23247 2533 23259 2536
rect 23201 2527 23259 2533
rect 23842 2524 23848 2536
rect 23900 2524 23906 2576
rect 30929 2567 30987 2573
rect 30929 2533 30941 2567
rect 30975 2564 30987 2567
rect 31570 2564 31576 2576
rect 30975 2536 31576 2564
rect 30975 2533 30987 2536
rect 30929 2527 30987 2533
rect 31570 2524 31576 2536
rect 31628 2524 31634 2576
rect 32861 2567 32919 2573
rect 32861 2533 32873 2567
rect 32907 2564 32919 2567
rect 33502 2564 33508 2576
rect 32907 2536 33508 2564
rect 32907 2533 32919 2536
rect 32861 2527 32919 2533
rect 33502 2524 33508 2536
rect 33560 2524 33566 2576
rect 39298 2524 39304 2576
rect 39356 2564 39362 2576
rect 41141 2567 41199 2573
rect 41141 2564 41153 2567
rect 39356 2536 41153 2564
rect 39356 2524 39362 2536
rect 41141 2533 41153 2536
rect 41187 2533 41199 2567
rect 41141 2527 41199 2533
rect 43162 2524 43168 2576
rect 43220 2564 43226 2576
rect 45005 2567 45063 2573
rect 45005 2564 45017 2567
rect 43220 2536 45017 2564
rect 43220 2524 43226 2536
rect 45005 2533 45017 2536
rect 45051 2533 45063 2567
rect 45005 2527 45063 2533
rect 47026 2524 47032 2576
rect 47084 2564 47090 2576
rect 48869 2567 48927 2573
rect 48869 2564 48881 2567
rect 47084 2536 48881 2564
rect 47084 2524 47090 2536
rect 48869 2533 48881 2536
rect 48915 2533 48927 2567
rect 48869 2527 48927 2533
rect 50890 2524 50896 2576
rect 50948 2564 50954 2576
rect 52733 2567 52791 2573
rect 52733 2564 52745 2567
rect 50948 2536 52745 2564
rect 50948 2524 50954 2536
rect 52733 2533 52745 2536
rect 52779 2533 52791 2567
rect 52733 2527 52791 2533
rect 54754 2524 54760 2576
rect 54812 2564 54818 2576
rect 56597 2567 56655 2573
rect 56597 2564 56609 2567
rect 54812 2536 56609 2564
rect 54812 2524 54818 2536
rect 56597 2533 56609 2536
rect 56643 2533 56655 2567
rect 56597 2527 56655 2533
rect 56686 2524 56692 2576
rect 56744 2564 56750 2576
rect 58529 2567 58587 2573
rect 58529 2564 58541 2567
rect 56744 2536 58541 2564
rect 56744 2524 56750 2536
rect 58529 2533 58541 2536
rect 58575 2533 58587 2567
rect 58529 2527 58587 2533
rect 22646 2496 22652 2508
rect 19352 2468 20392 2496
rect 21192 2468 22652 2496
rect 16163 2400 17448 2428
rect 16163 2397 16175 2400
rect 16117 2391 16175 2397
rect 17678 2388 17684 2440
rect 17736 2428 17742 2440
rect 18150 2431 18208 2437
rect 18150 2428 18162 2431
rect 17736 2400 18162 2428
rect 17736 2388 17742 2400
rect 18150 2397 18162 2400
rect 18196 2397 18208 2431
rect 19352 2428 19380 2468
rect 18150 2391 18208 2397
rect 18248 2400 19380 2428
rect 19705 2431 19763 2437
rect 18248 2372 18276 2400
rect 19705 2397 19717 2431
rect 19751 2428 19763 2431
rect 20162 2428 20168 2440
rect 19751 2400 20168 2428
rect 19751 2397 19763 2400
rect 19705 2391 19763 2397
rect 20162 2388 20168 2400
rect 20220 2388 20226 2440
rect 20438 2428 20444 2440
rect 20399 2400 20444 2428
rect 20438 2388 20444 2400
rect 20496 2388 20502 2440
rect 21192 2437 21220 2468
rect 22646 2456 22652 2468
rect 22704 2456 22710 2508
rect 25685 2499 25743 2505
rect 25685 2465 25697 2499
rect 25731 2496 25743 2499
rect 27154 2496 27160 2508
rect 25731 2468 27160 2496
rect 25731 2465 25743 2468
rect 25685 2459 25743 2465
rect 27154 2456 27160 2468
rect 27212 2456 27218 2508
rect 37090 2456 37096 2508
rect 37148 2496 37154 2508
rect 37921 2499 37979 2505
rect 37921 2496 37933 2499
rect 37148 2468 37933 2496
rect 37148 2456 37154 2468
rect 37921 2465 37933 2468
rect 37967 2465 37979 2499
rect 37921 2459 37979 2465
rect 38194 2456 38200 2508
rect 38252 2496 38258 2508
rect 39853 2499 39911 2505
rect 39853 2496 39865 2499
rect 38252 2468 39865 2496
rect 38252 2456 38258 2468
rect 39853 2465 39865 2468
rect 39899 2465 39911 2499
rect 39853 2459 39911 2465
rect 40678 2456 40684 2508
rect 40736 2496 40742 2508
rect 42429 2499 42487 2505
rect 42429 2496 42441 2499
rect 40736 2468 42441 2496
rect 40736 2456 40742 2468
rect 42429 2465 42441 2468
rect 42475 2465 42487 2499
rect 42429 2459 42487 2465
rect 43990 2456 43996 2508
rect 44048 2496 44054 2508
rect 45649 2499 45707 2505
rect 45649 2496 45661 2499
rect 44048 2468 45661 2496
rect 44048 2456 44054 2468
rect 45649 2465 45661 2468
rect 45695 2465 45707 2499
rect 45649 2459 45707 2465
rect 45922 2456 45928 2508
rect 45980 2496 45986 2508
rect 47581 2499 47639 2505
rect 47581 2496 47593 2499
rect 45980 2468 47593 2496
rect 45980 2456 45986 2468
rect 47581 2465 47593 2468
rect 47627 2465 47639 2499
rect 47581 2459 47639 2465
rect 48406 2456 48412 2508
rect 48464 2496 48470 2508
rect 50157 2499 50215 2505
rect 50157 2496 50169 2499
rect 48464 2468 50169 2496
rect 48464 2456 48470 2468
rect 50157 2465 50169 2468
rect 50203 2465 50215 2499
rect 50157 2459 50215 2465
rect 51718 2456 51724 2508
rect 51776 2496 51782 2508
rect 53377 2499 53435 2505
rect 53377 2496 53389 2499
rect 51776 2468 53389 2496
rect 51776 2456 51782 2468
rect 53377 2465 53389 2468
rect 53423 2465 53435 2499
rect 53377 2459 53435 2465
rect 53650 2456 53656 2508
rect 53708 2496 53714 2508
rect 55309 2499 55367 2505
rect 55309 2496 55321 2499
rect 53708 2468 55321 2496
rect 53708 2456 53714 2468
rect 55309 2465 55321 2468
rect 55355 2465 55367 2499
rect 55309 2459 55367 2465
rect 57422 2456 57428 2508
rect 57480 2496 57486 2508
rect 59173 2499 59231 2505
rect 59173 2496 59185 2499
rect 57480 2468 59185 2496
rect 57480 2456 57486 2468
rect 59173 2465 59185 2468
rect 59219 2465 59231 2499
rect 59173 2459 59231 2465
rect 21177 2431 21235 2437
rect 21177 2397 21189 2431
rect 21223 2397 21235 2431
rect 21177 2391 21235 2397
rect 22097 2431 22155 2437
rect 22097 2397 22109 2431
rect 22143 2428 22155 2431
rect 22830 2428 22836 2440
rect 22143 2400 22836 2428
rect 22143 2397 22155 2400
rect 22097 2391 22155 2397
rect 22830 2388 22836 2400
rect 22888 2388 22894 2440
rect 23845 2431 23903 2437
rect 23845 2397 23857 2431
rect 23891 2428 23903 2431
rect 24394 2428 24400 2440
rect 23891 2400 24400 2428
rect 23891 2397 23903 2400
rect 23845 2391 23903 2397
rect 24394 2388 24400 2400
rect 24452 2388 24458 2440
rect 26145 2431 26203 2437
rect 26145 2397 26157 2431
rect 26191 2428 26203 2431
rect 26418 2428 26424 2440
rect 26191 2400 26424 2428
rect 26191 2397 26203 2400
rect 26145 2391 26203 2397
rect 26418 2388 26424 2400
rect 26476 2388 26482 2440
rect 26970 2428 26976 2440
rect 26931 2400 26976 2428
rect 26970 2388 26976 2400
rect 27028 2388 27034 2440
rect 28353 2431 28411 2437
rect 28353 2397 28365 2431
rect 28399 2428 28411 2431
rect 28810 2428 28816 2440
rect 28399 2400 28816 2428
rect 28399 2397 28411 2400
rect 28353 2391 28411 2397
rect 28810 2388 28816 2400
rect 28868 2388 28874 2440
rect 28997 2431 29055 2437
rect 28997 2397 29009 2431
rect 29043 2428 29055 2431
rect 29638 2428 29644 2440
rect 29043 2400 29644 2428
rect 29043 2397 29055 2400
rect 28997 2391 29055 2397
rect 29638 2388 29644 2400
rect 29696 2388 29702 2440
rect 30285 2431 30343 2437
rect 30285 2397 30297 2431
rect 30331 2428 30343 2431
rect 30742 2428 30748 2440
rect 30331 2400 30748 2428
rect 30331 2397 30343 2400
rect 30285 2391 30343 2397
rect 30742 2388 30748 2400
rect 30800 2388 30806 2440
rect 31573 2431 31631 2437
rect 31573 2397 31585 2431
rect 31619 2428 31631 2431
rect 32398 2428 32404 2440
rect 31619 2400 32404 2428
rect 31619 2397 31631 2400
rect 31573 2391 31631 2397
rect 32398 2388 32404 2400
rect 32456 2388 32462 2440
rect 33505 2431 33563 2437
rect 33505 2397 33517 2431
rect 33551 2428 33563 2431
rect 34054 2428 34060 2440
rect 33551 2400 34060 2428
rect 33551 2397 33563 2400
rect 33505 2391 33563 2397
rect 34054 2388 34060 2400
rect 34112 2388 34118 2440
rect 34149 2431 34207 2437
rect 34149 2397 34161 2431
rect 34195 2428 34207 2431
rect 34606 2428 34612 2440
rect 34195 2400 34612 2428
rect 34195 2397 34207 2400
rect 34149 2391 34207 2397
rect 34606 2388 34612 2400
rect 34664 2388 34670 2440
rect 34977 2431 35035 2437
rect 34977 2397 34989 2431
rect 35023 2428 35035 2431
rect 35158 2428 35164 2440
rect 35023 2400 35164 2428
rect 35023 2397 35035 2400
rect 34977 2391 35035 2397
rect 35158 2388 35164 2400
rect 35216 2388 35222 2440
rect 35621 2431 35679 2437
rect 35621 2397 35633 2431
rect 35667 2428 35679 2431
rect 35710 2428 35716 2440
rect 35667 2400 35716 2428
rect 35667 2397 35679 2400
rect 35621 2391 35679 2397
rect 35710 2388 35716 2400
rect 35768 2388 35774 2440
rect 35986 2388 35992 2440
rect 36044 2428 36050 2440
rect 36081 2431 36139 2437
rect 36081 2428 36093 2431
rect 36044 2400 36093 2428
rect 36044 2388 36050 2400
rect 36081 2397 36093 2400
rect 36127 2397 36139 2431
rect 36081 2391 36139 2397
rect 36538 2388 36544 2440
rect 36596 2428 36602 2440
rect 37277 2431 37335 2437
rect 37277 2428 37289 2431
rect 36596 2400 37289 2428
rect 36596 2388 36602 2400
rect 37277 2397 37289 2400
rect 37323 2397 37335 2431
rect 37277 2391 37335 2397
rect 37642 2388 37648 2440
rect 37700 2428 37706 2440
rect 38565 2431 38623 2437
rect 38565 2428 38577 2431
rect 37700 2400 38577 2428
rect 37700 2388 37706 2400
rect 38565 2397 38577 2400
rect 38611 2397 38623 2431
rect 38565 2391 38623 2397
rect 38746 2388 38752 2440
rect 38804 2428 38810 2440
rect 40497 2431 40555 2437
rect 40497 2428 40509 2431
rect 38804 2400 40509 2428
rect 38804 2388 38810 2400
rect 40497 2397 40509 2400
rect 40543 2397 40555 2431
rect 40497 2391 40555 2397
rect 41230 2388 41236 2440
rect 41288 2428 41294 2440
rect 43073 2431 43131 2437
rect 43073 2428 43085 2431
rect 41288 2400 43085 2428
rect 41288 2388 41294 2400
rect 43073 2397 43085 2400
rect 43119 2397 43131 2431
rect 43073 2391 43131 2397
rect 43717 2431 43775 2437
rect 43717 2397 43729 2431
rect 43763 2397 43775 2431
rect 46293 2431 46351 2437
rect 46293 2428 46305 2431
rect 43717 2391 43775 2397
rect 45526 2400 46305 2428
rect 17586 2360 17592 2372
rect 15212 2332 17592 2360
rect 15212 2301 15240 2332
rect 17586 2320 17592 2332
rect 17644 2320 17650 2372
rect 18230 2320 18236 2372
rect 18288 2320 18294 2372
rect 19242 2320 19248 2372
rect 19300 2360 19306 2372
rect 19300 2332 21036 2360
rect 19300 2320 19306 2332
rect 13495 2264 15148 2292
rect 15197 2295 15255 2301
rect 13495 2261 13507 2264
rect 13449 2255 13507 2261
rect 15197 2261 15209 2295
rect 15243 2261 15255 2295
rect 15197 2255 15255 2261
rect 15933 2295 15991 2301
rect 15933 2261 15945 2295
rect 15979 2292 15991 2295
rect 18414 2292 18420 2304
rect 15979 2264 18420 2292
rect 15979 2261 15991 2264
rect 15933 2255 15991 2261
rect 18414 2252 18420 2264
rect 18472 2252 18478 2304
rect 20070 2252 20076 2304
rect 20128 2292 20134 2304
rect 21008 2301 21036 2332
rect 42058 2320 42064 2372
rect 42116 2360 42122 2372
rect 43732 2360 43760 2391
rect 42116 2332 43760 2360
rect 42116 2320 42122 2332
rect 44542 2320 44548 2372
rect 44600 2360 44606 2372
rect 45526 2360 45554 2400
rect 46293 2397 46305 2400
rect 46339 2397 46351 2431
rect 46293 2391 46351 2397
rect 46474 2388 46480 2440
rect 46532 2428 46538 2440
rect 48225 2431 48283 2437
rect 48225 2428 48237 2431
rect 46532 2400 48237 2428
rect 46532 2388 46538 2400
rect 48225 2397 48237 2400
rect 48271 2397 48283 2431
rect 48225 2391 48283 2397
rect 48958 2388 48964 2440
rect 49016 2428 49022 2440
rect 50801 2431 50859 2437
rect 50801 2428 50813 2431
rect 49016 2400 50813 2428
rect 49016 2388 49022 2400
rect 50801 2397 50813 2400
rect 50847 2397 50859 2431
rect 50801 2391 50859 2397
rect 51445 2431 51503 2437
rect 51445 2397 51457 2431
rect 51491 2397 51503 2431
rect 51445 2391 51503 2397
rect 44600 2332 45554 2360
rect 44600 2320 44606 2332
rect 49786 2320 49792 2372
rect 49844 2360 49850 2372
rect 51460 2360 51488 2391
rect 52270 2388 52276 2440
rect 52328 2428 52334 2440
rect 54021 2431 54079 2437
rect 54021 2428 54033 2431
rect 52328 2400 54033 2428
rect 52328 2388 52334 2400
rect 54021 2397 54033 2400
rect 54067 2397 54079 2431
rect 54021 2391 54079 2397
rect 55953 2431 56011 2437
rect 55953 2397 55965 2431
rect 55999 2397 56011 2431
rect 55953 2391 56011 2397
rect 49844 2332 51488 2360
rect 49844 2320 49850 2332
rect 54202 2320 54208 2372
rect 54260 2360 54266 2372
rect 55968 2360 55996 2391
rect 56134 2388 56140 2440
rect 56192 2428 56198 2440
rect 57885 2431 57943 2437
rect 57885 2428 57897 2431
rect 56192 2400 57897 2428
rect 56192 2388 56198 2400
rect 57885 2397 57897 2400
rect 57931 2397 57943 2431
rect 57885 2391 57943 2397
rect 54260 2332 55996 2360
rect 54260 2320 54266 2332
rect 20257 2295 20315 2301
rect 20257 2292 20269 2295
rect 20128 2264 20269 2292
rect 20128 2252 20134 2264
rect 20257 2261 20269 2264
rect 20303 2261 20315 2295
rect 20257 2255 20315 2261
rect 20993 2295 21051 2301
rect 20993 2261 21005 2295
rect 21039 2261 21051 2295
rect 20993 2255 21051 2261
rect 25041 2295 25099 2301
rect 25041 2261 25053 2295
rect 25087 2292 25099 2295
rect 25498 2292 25504 2304
rect 25087 2264 25504 2292
rect 25087 2261 25099 2264
rect 25041 2255 25099 2261
rect 25498 2252 25504 2264
rect 25556 2252 25562 2304
rect 26329 2295 26387 2301
rect 26329 2261 26341 2295
rect 26375 2292 26387 2295
rect 26602 2292 26608 2304
rect 26375 2264 26608 2292
rect 26375 2261 26387 2264
rect 26329 2255 26387 2261
rect 26602 2252 26608 2264
rect 26660 2252 26666 2304
rect 26878 2252 26884 2304
rect 26936 2292 26942 2304
rect 27157 2295 27215 2301
rect 27157 2292 27169 2295
rect 26936 2264 27169 2292
rect 26936 2252 26942 2264
rect 27157 2261 27169 2264
rect 27203 2261 27215 2295
rect 27157 2255 27215 2261
rect 1104 2202 68816 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 50294 2202
rect 50346 2150 50358 2202
rect 50410 2150 50422 2202
rect 50474 2150 50486 2202
rect 50538 2150 50550 2202
rect 50602 2150 68816 2202
rect 1104 2128 68816 2150
rect 10778 2048 10784 2100
rect 10836 2088 10842 2100
rect 14550 2088 14556 2100
rect 10836 2060 14556 2088
rect 10836 2048 10842 2060
rect 14550 2048 14556 2060
rect 14608 2048 14614 2100
rect 4706 1980 4712 2032
rect 4764 2020 4770 2032
rect 14090 2020 14096 2032
rect 4764 1992 14096 2020
rect 4764 1980 4770 1992
rect 14090 1980 14096 1992
rect 14148 1980 14154 2032
rect 6546 1912 6552 1964
rect 6604 1952 6610 1964
rect 12802 1952 12808 1964
rect 6604 1924 12808 1952
rect 6604 1912 6610 1924
rect 12802 1912 12808 1924
rect 12860 1912 12866 1964
rect 8202 1844 8208 1896
rect 8260 1884 8266 1896
rect 16390 1884 16396 1896
rect 8260 1856 16396 1884
rect 8260 1844 8266 1856
rect 16390 1844 16396 1856
rect 16448 1844 16454 1896
rect 10042 1776 10048 1828
rect 10100 1816 10106 1828
rect 14182 1816 14188 1828
rect 10100 1788 14188 1816
rect 10100 1776 10106 1788
rect 14182 1776 14188 1788
rect 14240 1776 14246 1828
rect 15286 1504 15292 1556
rect 15344 1544 15350 1556
rect 16206 1544 16212 1556
rect 15344 1516 16212 1544
rect 15344 1504 15350 1516
rect 16206 1504 16212 1516
rect 16264 1504 16270 1556
rect 12158 1436 12164 1488
rect 12216 1476 12222 1488
rect 14826 1476 14832 1488
rect 12216 1448 14832 1476
rect 12216 1436 12222 1448
rect 14826 1436 14832 1448
rect 14884 1436 14890 1488
rect 20254 1408 20260 1420
rect 19812 1380 20260 1408
rect 19812 1352 19840 1380
rect 20254 1368 20260 1380
rect 20312 1368 20318 1420
rect 19794 1300 19800 1352
rect 19852 1300 19858 1352
rect 19978 1300 19984 1352
rect 20036 1340 20042 1352
rect 20530 1340 20536 1352
rect 20036 1312 20536 1340
rect 20036 1300 20042 1312
rect 20530 1300 20536 1312
rect 20588 1300 20594 1352
<< via1 >>
rect 19574 57638 19626 57690
rect 19638 57638 19690 57690
rect 19702 57638 19754 57690
rect 19766 57638 19818 57690
rect 19830 57638 19882 57690
rect 50294 57638 50346 57690
rect 50358 57638 50410 57690
rect 50422 57638 50474 57690
rect 50486 57638 50538 57690
rect 50550 57638 50602 57690
rect 3516 57400 3568 57452
rect 4160 57443 4212 57452
rect 4160 57409 4169 57443
rect 4169 57409 4203 57443
rect 4203 57409 4212 57443
rect 4160 57400 4212 57409
rect 5172 57443 5224 57452
rect 5172 57409 5181 57443
rect 5181 57409 5215 57443
rect 5215 57409 5224 57443
rect 5172 57400 5224 57409
rect 5724 57400 5776 57452
rect 6828 57443 6880 57452
rect 6828 57409 6837 57443
rect 6837 57409 6871 57443
rect 6871 57409 6880 57443
rect 6828 57400 6880 57409
rect 7380 57400 7432 57452
rect 8484 57400 8536 57452
rect 9036 57400 9088 57452
rect 10140 57443 10192 57452
rect 10140 57409 10149 57443
rect 10149 57409 10183 57443
rect 10183 57409 10192 57443
rect 10140 57400 10192 57409
rect 10692 57400 10744 57452
rect 11796 57443 11848 57452
rect 11796 57409 11805 57443
rect 11805 57409 11839 57443
rect 11839 57409 11848 57443
rect 11796 57400 11848 57409
rect 12440 57443 12492 57452
rect 12440 57409 12449 57443
rect 12449 57409 12483 57443
rect 12483 57409 12492 57443
rect 12440 57400 12492 57409
rect 13452 57400 13504 57452
rect 14004 57400 14056 57452
rect 15108 57443 15160 57452
rect 15108 57409 15117 57443
rect 15117 57409 15151 57443
rect 15151 57409 15160 57443
rect 15108 57400 15160 57409
rect 15660 57400 15712 57452
rect 16764 57443 16816 57452
rect 16764 57409 16773 57443
rect 16773 57409 16807 57443
rect 16807 57409 16816 57443
rect 16764 57400 16816 57409
rect 17316 57400 17368 57452
rect 18420 57400 18472 57452
rect 18972 57400 19024 57452
rect 20076 57443 20128 57452
rect 20076 57409 20085 57443
rect 20085 57409 20119 57443
rect 20119 57409 20128 57443
rect 20076 57400 20128 57409
rect 20720 57443 20772 57452
rect 20720 57409 20729 57443
rect 20729 57409 20763 57443
rect 20763 57409 20772 57443
rect 20720 57400 20772 57409
rect 22284 57400 22336 57452
rect 23480 57443 23532 57452
rect 23480 57409 23489 57443
rect 23489 57409 23523 57443
rect 23523 57409 23532 57443
rect 23480 57400 23532 57409
rect 23940 57400 23992 57452
rect 25044 57443 25096 57452
rect 25044 57409 25053 57443
rect 25053 57409 25087 57443
rect 25087 57409 25096 57443
rect 25044 57400 25096 57409
rect 25596 57400 25648 57452
rect 27252 57400 27304 57452
rect 28356 57443 28408 57452
rect 28356 57409 28365 57443
rect 28365 57409 28399 57443
rect 28399 57409 28408 57443
rect 28356 57400 28408 57409
rect 28908 57400 28960 57452
rect 30012 57443 30064 57452
rect 30012 57409 30021 57443
rect 30021 57409 30055 57443
rect 30055 57409 30064 57443
rect 30012 57400 30064 57409
rect 30564 57400 30616 57452
rect 31668 57400 31720 57452
rect 32220 57400 32272 57452
rect 33324 57443 33376 57452
rect 33324 57409 33333 57443
rect 33333 57409 33367 57443
rect 33367 57409 33376 57443
rect 33324 57400 33376 57409
rect 33876 57400 33928 57452
rect 34980 57443 35032 57452
rect 34980 57409 34989 57443
rect 34989 57409 35023 57443
rect 35023 57409 35032 57443
rect 34980 57400 35032 57409
rect 35532 57400 35584 57452
rect 36636 57400 36688 57452
rect 38292 57400 38344 57452
rect 40040 57443 40092 57452
rect 40040 57409 40049 57443
rect 40049 57409 40083 57443
rect 40083 57409 40092 57443
rect 40040 57400 40092 57409
rect 40500 57400 40552 57452
rect 41604 57400 41656 57452
rect 42156 57400 42208 57452
rect 43260 57400 43312 57452
rect 43812 57400 43864 57452
rect 44916 57400 44968 57452
rect 46572 57400 46624 57452
rect 47124 57400 47176 57452
rect 48320 57443 48372 57452
rect 48320 57409 48329 57443
rect 48329 57409 48363 57443
rect 48363 57409 48372 57443
rect 48320 57400 48372 57409
rect 48780 57400 48832 57452
rect 49884 57400 49936 57452
rect 50620 57400 50672 57452
rect 51540 57400 51592 57452
rect 52460 57400 52512 57452
rect 53196 57400 53248 57452
rect 53840 57400 53892 57452
rect 54852 57400 54904 57452
rect 55404 57400 55456 57452
rect 56600 57443 56652 57452
rect 56600 57409 56609 57443
rect 56609 57409 56643 57443
rect 56643 57409 56652 57443
rect 56600 57400 56652 57409
rect 57060 57400 57112 57452
rect 58164 57400 58216 57452
rect 58716 57400 58768 57452
rect 59820 57400 59872 57452
rect 60740 57400 60792 57452
rect 61476 57400 61528 57452
rect 63132 57400 63184 57452
rect 63684 57400 63736 57452
rect 65340 57400 65392 57452
rect 66996 57400 67048 57452
rect 45468 57332 45520 57384
rect 64788 57332 64840 57384
rect 37280 57264 37332 57316
rect 4214 57094 4266 57146
rect 4278 57094 4330 57146
rect 4342 57094 4394 57146
rect 4406 57094 4458 57146
rect 4470 57094 4522 57146
rect 34934 57094 34986 57146
rect 34998 57094 35050 57146
rect 35062 57094 35114 57146
rect 35126 57094 35178 57146
rect 35190 57094 35242 57146
rect 65654 57094 65706 57146
rect 65718 57094 65770 57146
rect 65782 57094 65834 57146
rect 65846 57094 65898 57146
rect 65910 57094 65962 57146
rect 21732 56992 21784 57044
rect 26700 56992 26752 57044
rect 38844 56992 38896 57044
rect 62120 57035 62172 57044
rect 62120 57001 62129 57035
rect 62129 57001 62163 57035
rect 62163 57001 62172 57035
rect 62120 56992 62172 57001
rect 19574 56550 19626 56602
rect 19638 56550 19690 56602
rect 19702 56550 19754 56602
rect 19766 56550 19818 56602
rect 19830 56550 19882 56602
rect 50294 56550 50346 56602
rect 50358 56550 50410 56602
rect 50422 56550 50474 56602
rect 50486 56550 50538 56602
rect 50550 56550 50602 56602
rect 4214 56006 4266 56058
rect 4278 56006 4330 56058
rect 4342 56006 4394 56058
rect 4406 56006 4458 56058
rect 4470 56006 4522 56058
rect 34934 56006 34986 56058
rect 34998 56006 35050 56058
rect 35062 56006 35114 56058
rect 35126 56006 35178 56058
rect 35190 56006 35242 56058
rect 65654 56006 65706 56058
rect 65718 56006 65770 56058
rect 65782 56006 65834 56058
rect 65846 56006 65898 56058
rect 65910 56006 65962 56058
rect 19574 55462 19626 55514
rect 19638 55462 19690 55514
rect 19702 55462 19754 55514
rect 19766 55462 19818 55514
rect 19830 55462 19882 55514
rect 50294 55462 50346 55514
rect 50358 55462 50410 55514
rect 50422 55462 50474 55514
rect 50486 55462 50538 55514
rect 50550 55462 50602 55514
rect 4214 54918 4266 54970
rect 4278 54918 4330 54970
rect 4342 54918 4394 54970
rect 4406 54918 4458 54970
rect 4470 54918 4522 54970
rect 34934 54918 34986 54970
rect 34998 54918 35050 54970
rect 35062 54918 35114 54970
rect 35126 54918 35178 54970
rect 35190 54918 35242 54970
rect 65654 54918 65706 54970
rect 65718 54918 65770 54970
rect 65782 54918 65834 54970
rect 65846 54918 65898 54970
rect 65910 54918 65962 54970
rect 19574 54374 19626 54426
rect 19638 54374 19690 54426
rect 19702 54374 19754 54426
rect 19766 54374 19818 54426
rect 19830 54374 19882 54426
rect 50294 54374 50346 54426
rect 50358 54374 50410 54426
rect 50422 54374 50474 54426
rect 50486 54374 50538 54426
rect 50550 54374 50602 54426
rect 4214 53830 4266 53882
rect 4278 53830 4330 53882
rect 4342 53830 4394 53882
rect 4406 53830 4458 53882
rect 4470 53830 4522 53882
rect 34934 53830 34986 53882
rect 34998 53830 35050 53882
rect 35062 53830 35114 53882
rect 35126 53830 35178 53882
rect 35190 53830 35242 53882
rect 65654 53830 65706 53882
rect 65718 53830 65770 53882
rect 65782 53830 65834 53882
rect 65846 53830 65898 53882
rect 65910 53830 65962 53882
rect 19574 53286 19626 53338
rect 19638 53286 19690 53338
rect 19702 53286 19754 53338
rect 19766 53286 19818 53338
rect 19830 53286 19882 53338
rect 50294 53286 50346 53338
rect 50358 53286 50410 53338
rect 50422 53286 50474 53338
rect 50486 53286 50538 53338
rect 50550 53286 50602 53338
rect 4214 52742 4266 52794
rect 4278 52742 4330 52794
rect 4342 52742 4394 52794
rect 4406 52742 4458 52794
rect 4470 52742 4522 52794
rect 34934 52742 34986 52794
rect 34998 52742 35050 52794
rect 35062 52742 35114 52794
rect 35126 52742 35178 52794
rect 35190 52742 35242 52794
rect 65654 52742 65706 52794
rect 65718 52742 65770 52794
rect 65782 52742 65834 52794
rect 65846 52742 65898 52794
rect 65910 52742 65962 52794
rect 19574 52198 19626 52250
rect 19638 52198 19690 52250
rect 19702 52198 19754 52250
rect 19766 52198 19818 52250
rect 19830 52198 19882 52250
rect 50294 52198 50346 52250
rect 50358 52198 50410 52250
rect 50422 52198 50474 52250
rect 50486 52198 50538 52250
rect 50550 52198 50602 52250
rect 4214 51654 4266 51706
rect 4278 51654 4330 51706
rect 4342 51654 4394 51706
rect 4406 51654 4458 51706
rect 4470 51654 4522 51706
rect 34934 51654 34986 51706
rect 34998 51654 35050 51706
rect 35062 51654 35114 51706
rect 35126 51654 35178 51706
rect 35190 51654 35242 51706
rect 65654 51654 65706 51706
rect 65718 51654 65770 51706
rect 65782 51654 65834 51706
rect 65846 51654 65898 51706
rect 65910 51654 65962 51706
rect 19574 51110 19626 51162
rect 19638 51110 19690 51162
rect 19702 51110 19754 51162
rect 19766 51110 19818 51162
rect 19830 51110 19882 51162
rect 50294 51110 50346 51162
rect 50358 51110 50410 51162
rect 50422 51110 50474 51162
rect 50486 51110 50538 51162
rect 50550 51110 50602 51162
rect 4214 50566 4266 50618
rect 4278 50566 4330 50618
rect 4342 50566 4394 50618
rect 4406 50566 4458 50618
rect 4470 50566 4522 50618
rect 34934 50566 34986 50618
rect 34998 50566 35050 50618
rect 35062 50566 35114 50618
rect 35126 50566 35178 50618
rect 35190 50566 35242 50618
rect 65654 50566 65706 50618
rect 65718 50566 65770 50618
rect 65782 50566 65834 50618
rect 65846 50566 65898 50618
rect 65910 50566 65962 50618
rect 19574 50022 19626 50074
rect 19638 50022 19690 50074
rect 19702 50022 19754 50074
rect 19766 50022 19818 50074
rect 19830 50022 19882 50074
rect 50294 50022 50346 50074
rect 50358 50022 50410 50074
rect 50422 50022 50474 50074
rect 50486 50022 50538 50074
rect 50550 50022 50602 50074
rect 4214 49478 4266 49530
rect 4278 49478 4330 49530
rect 4342 49478 4394 49530
rect 4406 49478 4458 49530
rect 4470 49478 4522 49530
rect 34934 49478 34986 49530
rect 34998 49478 35050 49530
rect 35062 49478 35114 49530
rect 35126 49478 35178 49530
rect 35190 49478 35242 49530
rect 65654 49478 65706 49530
rect 65718 49478 65770 49530
rect 65782 49478 65834 49530
rect 65846 49478 65898 49530
rect 65910 49478 65962 49530
rect 19574 48934 19626 48986
rect 19638 48934 19690 48986
rect 19702 48934 19754 48986
rect 19766 48934 19818 48986
rect 19830 48934 19882 48986
rect 50294 48934 50346 48986
rect 50358 48934 50410 48986
rect 50422 48934 50474 48986
rect 50486 48934 50538 48986
rect 50550 48934 50602 48986
rect 4214 48390 4266 48442
rect 4278 48390 4330 48442
rect 4342 48390 4394 48442
rect 4406 48390 4458 48442
rect 4470 48390 4522 48442
rect 34934 48390 34986 48442
rect 34998 48390 35050 48442
rect 35062 48390 35114 48442
rect 35126 48390 35178 48442
rect 35190 48390 35242 48442
rect 65654 48390 65706 48442
rect 65718 48390 65770 48442
rect 65782 48390 65834 48442
rect 65846 48390 65898 48442
rect 65910 48390 65962 48442
rect 19574 47846 19626 47898
rect 19638 47846 19690 47898
rect 19702 47846 19754 47898
rect 19766 47846 19818 47898
rect 19830 47846 19882 47898
rect 50294 47846 50346 47898
rect 50358 47846 50410 47898
rect 50422 47846 50474 47898
rect 50486 47846 50538 47898
rect 50550 47846 50602 47898
rect 4214 47302 4266 47354
rect 4278 47302 4330 47354
rect 4342 47302 4394 47354
rect 4406 47302 4458 47354
rect 4470 47302 4522 47354
rect 34934 47302 34986 47354
rect 34998 47302 35050 47354
rect 35062 47302 35114 47354
rect 35126 47302 35178 47354
rect 35190 47302 35242 47354
rect 65654 47302 65706 47354
rect 65718 47302 65770 47354
rect 65782 47302 65834 47354
rect 65846 47302 65898 47354
rect 65910 47302 65962 47354
rect 19574 46758 19626 46810
rect 19638 46758 19690 46810
rect 19702 46758 19754 46810
rect 19766 46758 19818 46810
rect 19830 46758 19882 46810
rect 50294 46758 50346 46810
rect 50358 46758 50410 46810
rect 50422 46758 50474 46810
rect 50486 46758 50538 46810
rect 50550 46758 50602 46810
rect 4214 46214 4266 46266
rect 4278 46214 4330 46266
rect 4342 46214 4394 46266
rect 4406 46214 4458 46266
rect 4470 46214 4522 46266
rect 34934 46214 34986 46266
rect 34998 46214 35050 46266
rect 35062 46214 35114 46266
rect 35126 46214 35178 46266
rect 35190 46214 35242 46266
rect 65654 46214 65706 46266
rect 65718 46214 65770 46266
rect 65782 46214 65834 46266
rect 65846 46214 65898 46266
rect 65910 46214 65962 46266
rect 19574 45670 19626 45722
rect 19638 45670 19690 45722
rect 19702 45670 19754 45722
rect 19766 45670 19818 45722
rect 19830 45670 19882 45722
rect 50294 45670 50346 45722
rect 50358 45670 50410 45722
rect 50422 45670 50474 45722
rect 50486 45670 50538 45722
rect 50550 45670 50602 45722
rect 4214 45126 4266 45178
rect 4278 45126 4330 45178
rect 4342 45126 4394 45178
rect 4406 45126 4458 45178
rect 4470 45126 4522 45178
rect 34934 45126 34986 45178
rect 34998 45126 35050 45178
rect 35062 45126 35114 45178
rect 35126 45126 35178 45178
rect 35190 45126 35242 45178
rect 65654 45126 65706 45178
rect 65718 45126 65770 45178
rect 65782 45126 65834 45178
rect 65846 45126 65898 45178
rect 65910 45126 65962 45178
rect 19574 44582 19626 44634
rect 19638 44582 19690 44634
rect 19702 44582 19754 44634
rect 19766 44582 19818 44634
rect 19830 44582 19882 44634
rect 50294 44582 50346 44634
rect 50358 44582 50410 44634
rect 50422 44582 50474 44634
rect 50486 44582 50538 44634
rect 50550 44582 50602 44634
rect 4214 44038 4266 44090
rect 4278 44038 4330 44090
rect 4342 44038 4394 44090
rect 4406 44038 4458 44090
rect 4470 44038 4522 44090
rect 34934 44038 34986 44090
rect 34998 44038 35050 44090
rect 35062 44038 35114 44090
rect 35126 44038 35178 44090
rect 35190 44038 35242 44090
rect 65654 44038 65706 44090
rect 65718 44038 65770 44090
rect 65782 44038 65834 44090
rect 65846 44038 65898 44090
rect 65910 44038 65962 44090
rect 19574 43494 19626 43546
rect 19638 43494 19690 43546
rect 19702 43494 19754 43546
rect 19766 43494 19818 43546
rect 19830 43494 19882 43546
rect 50294 43494 50346 43546
rect 50358 43494 50410 43546
rect 50422 43494 50474 43546
rect 50486 43494 50538 43546
rect 50550 43494 50602 43546
rect 4214 42950 4266 43002
rect 4278 42950 4330 43002
rect 4342 42950 4394 43002
rect 4406 42950 4458 43002
rect 4470 42950 4522 43002
rect 34934 42950 34986 43002
rect 34998 42950 35050 43002
rect 35062 42950 35114 43002
rect 35126 42950 35178 43002
rect 35190 42950 35242 43002
rect 65654 42950 65706 43002
rect 65718 42950 65770 43002
rect 65782 42950 65834 43002
rect 65846 42950 65898 43002
rect 65910 42950 65962 43002
rect 19574 42406 19626 42458
rect 19638 42406 19690 42458
rect 19702 42406 19754 42458
rect 19766 42406 19818 42458
rect 19830 42406 19882 42458
rect 50294 42406 50346 42458
rect 50358 42406 50410 42458
rect 50422 42406 50474 42458
rect 50486 42406 50538 42458
rect 50550 42406 50602 42458
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 34934 41862 34986 41914
rect 34998 41862 35050 41914
rect 35062 41862 35114 41914
rect 35126 41862 35178 41914
rect 35190 41862 35242 41914
rect 65654 41862 65706 41914
rect 65718 41862 65770 41914
rect 65782 41862 65834 41914
rect 65846 41862 65898 41914
rect 65910 41862 65962 41914
rect 19574 41318 19626 41370
rect 19638 41318 19690 41370
rect 19702 41318 19754 41370
rect 19766 41318 19818 41370
rect 19830 41318 19882 41370
rect 50294 41318 50346 41370
rect 50358 41318 50410 41370
rect 50422 41318 50474 41370
rect 50486 41318 50538 41370
rect 50550 41318 50602 41370
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 34934 40774 34986 40826
rect 34998 40774 35050 40826
rect 35062 40774 35114 40826
rect 35126 40774 35178 40826
rect 35190 40774 35242 40826
rect 65654 40774 65706 40826
rect 65718 40774 65770 40826
rect 65782 40774 65834 40826
rect 65846 40774 65898 40826
rect 65910 40774 65962 40826
rect 19574 40230 19626 40282
rect 19638 40230 19690 40282
rect 19702 40230 19754 40282
rect 19766 40230 19818 40282
rect 19830 40230 19882 40282
rect 50294 40230 50346 40282
rect 50358 40230 50410 40282
rect 50422 40230 50474 40282
rect 50486 40230 50538 40282
rect 50550 40230 50602 40282
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 65654 39686 65706 39738
rect 65718 39686 65770 39738
rect 65782 39686 65834 39738
rect 65846 39686 65898 39738
rect 65910 39686 65962 39738
rect 19574 39142 19626 39194
rect 19638 39142 19690 39194
rect 19702 39142 19754 39194
rect 19766 39142 19818 39194
rect 19830 39142 19882 39194
rect 50294 39142 50346 39194
rect 50358 39142 50410 39194
rect 50422 39142 50474 39194
rect 50486 39142 50538 39194
rect 50550 39142 50602 39194
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 65654 38598 65706 38650
rect 65718 38598 65770 38650
rect 65782 38598 65834 38650
rect 65846 38598 65898 38650
rect 65910 38598 65962 38650
rect 19574 38054 19626 38106
rect 19638 38054 19690 38106
rect 19702 38054 19754 38106
rect 19766 38054 19818 38106
rect 19830 38054 19882 38106
rect 50294 38054 50346 38106
rect 50358 38054 50410 38106
rect 50422 38054 50474 38106
rect 50486 38054 50538 38106
rect 50550 38054 50602 38106
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 65654 37510 65706 37562
rect 65718 37510 65770 37562
rect 65782 37510 65834 37562
rect 65846 37510 65898 37562
rect 65910 37510 65962 37562
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 50294 36966 50346 37018
rect 50358 36966 50410 37018
rect 50422 36966 50474 37018
rect 50486 36966 50538 37018
rect 50550 36966 50602 37018
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 65654 36422 65706 36474
rect 65718 36422 65770 36474
rect 65782 36422 65834 36474
rect 65846 36422 65898 36474
rect 65910 36422 65962 36474
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 50294 35878 50346 35930
rect 50358 35878 50410 35930
rect 50422 35878 50474 35930
rect 50486 35878 50538 35930
rect 50550 35878 50602 35930
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 65654 35334 65706 35386
rect 65718 35334 65770 35386
rect 65782 35334 65834 35386
rect 65846 35334 65898 35386
rect 65910 35334 65962 35386
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 50294 34790 50346 34842
rect 50358 34790 50410 34842
rect 50422 34790 50474 34842
rect 50486 34790 50538 34842
rect 50550 34790 50602 34842
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 65654 34246 65706 34298
rect 65718 34246 65770 34298
rect 65782 34246 65834 34298
rect 65846 34246 65898 34298
rect 65910 34246 65962 34298
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 50294 33702 50346 33754
rect 50358 33702 50410 33754
rect 50422 33702 50474 33754
rect 50486 33702 50538 33754
rect 50550 33702 50602 33754
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 65654 33158 65706 33210
rect 65718 33158 65770 33210
rect 65782 33158 65834 33210
rect 65846 33158 65898 33210
rect 65910 33158 65962 33210
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 50294 32614 50346 32666
rect 50358 32614 50410 32666
rect 50422 32614 50474 32666
rect 50486 32614 50538 32666
rect 50550 32614 50602 32666
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 65654 32070 65706 32122
rect 65718 32070 65770 32122
rect 65782 32070 65834 32122
rect 65846 32070 65898 32122
rect 65910 32070 65962 32122
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 50294 31526 50346 31578
rect 50358 31526 50410 31578
rect 50422 31526 50474 31578
rect 50486 31526 50538 31578
rect 50550 31526 50602 31578
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 65654 30982 65706 31034
rect 65718 30982 65770 31034
rect 65782 30982 65834 31034
rect 65846 30982 65898 31034
rect 65910 30982 65962 31034
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 50294 30438 50346 30490
rect 50358 30438 50410 30490
rect 50422 30438 50474 30490
rect 50486 30438 50538 30490
rect 50550 30438 50602 30490
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 65654 29894 65706 29946
rect 65718 29894 65770 29946
rect 65782 29894 65834 29946
rect 65846 29894 65898 29946
rect 65910 29894 65962 29946
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 50294 29350 50346 29402
rect 50358 29350 50410 29402
rect 50422 29350 50474 29402
rect 50486 29350 50538 29402
rect 50550 29350 50602 29402
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 65654 28806 65706 28858
rect 65718 28806 65770 28858
rect 65782 28806 65834 28858
rect 65846 28806 65898 28858
rect 65910 28806 65962 28858
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 50294 28262 50346 28314
rect 50358 28262 50410 28314
rect 50422 28262 50474 28314
rect 50486 28262 50538 28314
rect 50550 28262 50602 28314
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 65654 27718 65706 27770
rect 65718 27718 65770 27770
rect 65782 27718 65834 27770
rect 65846 27718 65898 27770
rect 65910 27718 65962 27770
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 50294 27174 50346 27226
rect 50358 27174 50410 27226
rect 50422 27174 50474 27226
rect 50486 27174 50538 27226
rect 50550 27174 50602 27226
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 65654 26630 65706 26682
rect 65718 26630 65770 26682
rect 65782 26630 65834 26682
rect 65846 26630 65898 26682
rect 65910 26630 65962 26682
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 50294 26086 50346 26138
rect 50358 26086 50410 26138
rect 50422 26086 50474 26138
rect 50486 26086 50538 26138
rect 50550 26086 50602 26138
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 65654 25542 65706 25594
rect 65718 25542 65770 25594
rect 65782 25542 65834 25594
rect 65846 25542 65898 25594
rect 65910 25542 65962 25594
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 50294 24998 50346 25050
rect 50358 24998 50410 25050
rect 50422 24998 50474 25050
rect 50486 24998 50538 25050
rect 50550 24998 50602 25050
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 65654 24454 65706 24506
rect 65718 24454 65770 24506
rect 65782 24454 65834 24506
rect 65846 24454 65898 24506
rect 65910 24454 65962 24506
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 50294 23910 50346 23962
rect 50358 23910 50410 23962
rect 50422 23910 50474 23962
rect 50486 23910 50538 23962
rect 50550 23910 50602 23962
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 65654 23366 65706 23418
rect 65718 23366 65770 23418
rect 65782 23366 65834 23418
rect 65846 23366 65898 23418
rect 65910 23366 65962 23418
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 50294 22822 50346 22874
rect 50358 22822 50410 22874
rect 50422 22822 50474 22874
rect 50486 22822 50538 22874
rect 50550 22822 50602 22874
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 65654 22278 65706 22330
rect 65718 22278 65770 22330
rect 65782 22278 65834 22330
rect 65846 22278 65898 22330
rect 65910 22278 65962 22330
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 50294 21734 50346 21786
rect 50358 21734 50410 21786
rect 50422 21734 50474 21786
rect 50486 21734 50538 21786
rect 50550 21734 50602 21786
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 65654 21190 65706 21242
rect 65718 21190 65770 21242
rect 65782 21190 65834 21242
rect 65846 21190 65898 21242
rect 65910 21190 65962 21242
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 50294 20646 50346 20698
rect 50358 20646 50410 20698
rect 50422 20646 50474 20698
rect 50486 20646 50538 20698
rect 50550 20646 50602 20698
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 65654 20102 65706 20154
rect 65718 20102 65770 20154
rect 65782 20102 65834 20154
rect 65846 20102 65898 20154
rect 65910 20102 65962 20154
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 50294 19558 50346 19610
rect 50358 19558 50410 19610
rect 50422 19558 50474 19610
rect 50486 19558 50538 19610
rect 50550 19558 50602 19610
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 65654 19014 65706 19066
rect 65718 19014 65770 19066
rect 65782 19014 65834 19066
rect 65846 19014 65898 19066
rect 65910 19014 65962 19066
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 50294 18470 50346 18522
rect 50358 18470 50410 18522
rect 50422 18470 50474 18522
rect 50486 18470 50538 18522
rect 50550 18470 50602 18522
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 65654 17926 65706 17978
rect 65718 17926 65770 17978
rect 65782 17926 65834 17978
rect 65846 17926 65898 17978
rect 65910 17926 65962 17978
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 50294 17382 50346 17434
rect 50358 17382 50410 17434
rect 50422 17382 50474 17434
rect 50486 17382 50538 17434
rect 50550 17382 50602 17434
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 65654 16838 65706 16890
rect 65718 16838 65770 16890
rect 65782 16838 65834 16890
rect 65846 16838 65898 16890
rect 65910 16838 65962 16890
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 50294 16294 50346 16346
rect 50358 16294 50410 16346
rect 50422 16294 50474 16346
rect 50486 16294 50538 16346
rect 50550 16294 50602 16346
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 65654 15750 65706 15802
rect 65718 15750 65770 15802
rect 65782 15750 65834 15802
rect 65846 15750 65898 15802
rect 65910 15750 65962 15802
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 50294 15206 50346 15258
rect 50358 15206 50410 15258
rect 50422 15206 50474 15258
rect 50486 15206 50538 15258
rect 50550 15206 50602 15258
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 65654 14662 65706 14714
rect 65718 14662 65770 14714
rect 65782 14662 65834 14714
rect 65846 14662 65898 14714
rect 65910 14662 65962 14714
rect 11704 14424 11756 14476
rect 10508 14356 10560 14408
rect 10416 14288 10468 14340
rect 4344 14220 4396 14272
rect 5080 14220 5132 14272
rect 11428 14220 11480 14272
rect 11612 14263 11664 14272
rect 11612 14229 11621 14263
rect 11621 14229 11655 14263
rect 11655 14229 11664 14263
rect 11612 14220 11664 14229
rect 12440 14356 12492 14408
rect 15200 14356 15252 14408
rect 15016 14263 15068 14272
rect 15016 14229 15025 14263
rect 15025 14229 15059 14263
rect 15059 14229 15068 14263
rect 15016 14220 15068 14229
rect 16856 14356 16908 14408
rect 16304 14288 16356 14340
rect 15660 14220 15712 14272
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 50294 14118 50346 14170
rect 50358 14118 50410 14170
rect 50422 14118 50474 14170
rect 50486 14118 50538 14170
rect 50550 14118 50602 14170
rect 4344 14059 4396 14068
rect 4344 14025 4353 14059
rect 4353 14025 4387 14059
rect 4387 14025 4396 14059
rect 4344 14016 4396 14025
rect 11428 14016 11480 14068
rect 14740 14016 14792 14068
rect 12900 13948 12952 14000
rect 5816 13880 5868 13932
rect 8852 13923 8904 13932
rect 8852 13889 8861 13923
rect 8861 13889 8895 13923
rect 8895 13889 8904 13923
rect 8852 13880 8904 13889
rect 10600 13923 10652 13932
rect 10600 13889 10609 13923
rect 10609 13889 10643 13923
rect 10643 13889 10652 13923
rect 10600 13880 10652 13889
rect 8116 13855 8168 13864
rect 8116 13821 8125 13855
rect 8125 13821 8159 13855
rect 8159 13821 8168 13855
rect 8116 13812 8168 13821
rect 8760 13812 8812 13864
rect 9864 13812 9916 13864
rect 11152 13880 11204 13932
rect 12440 13880 12492 13932
rect 13084 13923 13136 13932
rect 13084 13889 13093 13923
rect 13093 13889 13127 13923
rect 13127 13889 13136 13923
rect 13084 13880 13136 13889
rect 10876 13812 10928 13864
rect 11520 13812 11572 13864
rect 12716 13812 12768 13864
rect 7288 13744 7340 13796
rect 10784 13744 10836 13796
rect 11704 13744 11756 13796
rect 12164 13744 12216 13796
rect 13728 13855 13780 13864
rect 13728 13821 13737 13855
rect 13737 13821 13771 13855
rect 13771 13821 13780 13855
rect 13728 13812 13780 13821
rect 14740 13855 14792 13864
rect 14740 13821 14749 13855
rect 14749 13821 14783 13855
rect 14783 13821 14792 13855
rect 14740 13812 14792 13821
rect 21548 13812 21600 13864
rect 9036 13719 9088 13728
rect 9036 13685 9045 13719
rect 9045 13685 9079 13719
rect 9079 13685 9088 13719
rect 9036 13676 9088 13685
rect 13084 13676 13136 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 65654 13574 65706 13626
rect 65718 13574 65770 13626
rect 65782 13574 65834 13626
rect 65846 13574 65898 13626
rect 65910 13574 65962 13626
rect 9036 13515 9088 13524
rect 9036 13481 9045 13515
rect 9045 13481 9079 13515
rect 9079 13481 9088 13515
rect 9036 13472 9088 13481
rect 10416 13472 10468 13524
rect 7288 13311 7340 13320
rect 7288 13277 7297 13311
rect 7297 13277 7331 13311
rect 7331 13277 7340 13311
rect 7288 13268 7340 13277
rect 8576 13268 8628 13320
rect 8944 13311 8996 13320
rect 8944 13277 8953 13311
rect 8953 13277 8987 13311
rect 8987 13277 8996 13311
rect 8944 13268 8996 13277
rect 9220 13268 9272 13320
rect 10784 13404 10836 13456
rect 11520 13515 11572 13524
rect 11520 13481 11529 13515
rect 11529 13481 11563 13515
rect 11563 13481 11572 13515
rect 11520 13472 11572 13481
rect 12716 13472 12768 13524
rect 12900 13404 12952 13456
rect 10805 13305 10857 13314
rect 10805 13271 10814 13305
rect 10814 13271 10848 13305
rect 10848 13271 10857 13305
rect 10805 13262 10857 13271
rect 11152 13268 11204 13320
rect 13084 13336 13136 13388
rect 10324 13175 10376 13184
rect 10324 13141 10333 13175
rect 10333 13141 10367 13175
rect 10367 13141 10376 13175
rect 10324 13132 10376 13141
rect 11428 13132 11480 13184
rect 12532 13175 12584 13184
rect 12532 13141 12541 13175
rect 12541 13141 12575 13175
rect 12575 13141 12584 13175
rect 12532 13132 12584 13141
rect 13176 13311 13228 13320
rect 13176 13277 13197 13311
rect 13197 13277 13228 13311
rect 13176 13268 13228 13277
rect 15292 13268 15344 13320
rect 15660 13336 15712 13388
rect 16856 13404 16908 13456
rect 16396 13268 16448 13320
rect 16672 13311 16724 13320
rect 16672 13277 16686 13311
rect 16686 13277 16720 13311
rect 16720 13277 16724 13311
rect 16672 13268 16724 13277
rect 16856 13311 16908 13320
rect 16856 13277 16865 13311
rect 16865 13277 16899 13311
rect 16899 13277 16908 13311
rect 16856 13268 16908 13277
rect 17316 13268 17368 13320
rect 13268 13132 13320 13184
rect 14924 13132 14976 13184
rect 16212 13175 16264 13184
rect 16212 13141 16221 13175
rect 16221 13141 16255 13175
rect 16255 13141 16264 13175
rect 16212 13132 16264 13141
rect 16396 13132 16448 13184
rect 16580 13132 16632 13184
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 50294 13030 50346 13082
rect 50358 13030 50410 13082
rect 50422 13030 50474 13082
rect 50486 13030 50538 13082
rect 50550 13030 50602 13082
rect 10784 12928 10836 12980
rect 15660 12928 15712 12980
rect 16580 12928 16632 12980
rect 15016 12860 15068 12912
rect 4712 12835 4764 12844
rect 4712 12801 4721 12835
rect 4721 12801 4755 12835
rect 4755 12801 4764 12835
rect 4712 12792 4764 12801
rect 4620 12724 4672 12776
rect 8760 12792 8812 12844
rect 8944 12792 8996 12844
rect 13544 12792 13596 12844
rect 21732 12792 21784 12844
rect 6184 12724 6236 12776
rect 8392 12724 8444 12776
rect 16120 12767 16172 12776
rect 16120 12733 16129 12767
rect 16129 12733 16163 12767
rect 16163 12733 16172 12767
rect 16120 12724 16172 12733
rect 10140 12656 10192 12708
rect 7288 12588 7340 12640
rect 8852 12588 8904 12640
rect 9036 12631 9088 12640
rect 9036 12597 9045 12631
rect 9045 12597 9079 12631
rect 9079 12597 9088 12631
rect 9036 12588 9088 12597
rect 15200 12588 15252 12640
rect 20076 12588 20128 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 65654 12486 65706 12538
rect 65718 12486 65770 12538
rect 65782 12486 65834 12538
rect 65846 12486 65898 12538
rect 65910 12486 65962 12538
rect 4712 12248 4764 12300
rect 5540 12223 5592 12232
rect 5540 12189 5549 12223
rect 5549 12189 5583 12223
rect 5583 12189 5592 12223
rect 5540 12180 5592 12189
rect 7104 12180 7156 12232
rect 11704 12180 11756 12232
rect 12532 12180 12584 12232
rect 14648 12180 14700 12232
rect 16948 12180 17000 12232
rect 5356 12112 5408 12164
rect 10416 12155 10468 12164
rect 10416 12121 10450 12155
rect 10450 12121 10468 12155
rect 10416 12112 10468 12121
rect 20904 12316 20956 12368
rect 20812 12248 20864 12300
rect 8392 12087 8444 12096
rect 8392 12053 8401 12087
rect 8401 12053 8435 12087
rect 8435 12053 8444 12087
rect 8392 12044 8444 12053
rect 11428 12044 11480 12096
rect 13268 12044 13320 12096
rect 16856 12087 16908 12096
rect 16856 12053 16865 12087
rect 16865 12053 16899 12087
rect 16899 12053 16908 12087
rect 16856 12044 16908 12053
rect 16948 12044 17000 12096
rect 17868 12180 17920 12232
rect 18420 12180 18472 12232
rect 20536 12112 20588 12164
rect 21272 12180 21324 12232
rect 21732 12223 21784 12232
rect 21732 12189 21741 12223
rect 21741 12189 21775 12223
rect 21775 12189 21784 12223
rect 21732 12180 21784 12189
rect 22376 12223 22428 12232
rect 22376 12189 22380 12223
rect 22380 12189 22414 12223
rect 22414 12189 22428 12223
rect 22376 12180 22428 12189
rect 18696 12087 18748 12096
rect 18696 12053 18705 12087
rect 18705 12053 18739 12087
rect 18739 12053 18748 12087
rect 18696 12044 18748 12053
rect 21640 12044 21692 12096
rect 22560 12044 22612 12096
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 50294 11942 50346 11994
rect 50358 11942 50410 11994
rect 50422 11942 50474 11994
rect 50486 11942 50538 11994
rect 50550 11942 50602 11994
rect 5356 11883 5408 11892
rect 5356 11849 5365 11883
rect 5365 11849 5399 11883
rect 5399 11849 5408 11883
rect 5356 11840 5408 11849
rect 5540 11840 5592 11892
rect 4712 11747 4764 11756
rect 4712 11713 4721 11747
rect 4721 11713 4755 11747
rect 4755 11713 4764 11747
rect 4712 11704 4764 11713
rect 8392 11772 8444 11824
rect 8760 11840 8812 11892
rect 12716 11840 12768 11892
rect 16120 11840 16172 11892
rect 20536 11840 20588 11892
rect 10140 11815 10192 11824
rect 10140 11781 10158 11815
rect 10158 11781 10192 11815
rect 14924 11815 14976 11824
rect 10140 11772 10192 11781
rect 14924 11781 14958 11815
rect 14958 11781 14976 11815
rect 14924 11772 14976 11781
rect 16856 11772 16908 11824
rect 22560 11772 22612 11824
rect 6368 11704 6420 11756
rect 13544 11704 13596 11756
rect 14648 11747 14700 11756
rect 14648 11713 14657 11747
rect 14657 11713 14691 11747
rect 14691 11713 14700 11747
rect 14648 11704 14700 11713
rect 18420 11747 18472 11756
rect 18420 11713 18429 11747
rect 18429 11713 18463 11747
rect 18463 11713 18472 11747
rect 18420 11704 18472 11713
rect 20444 11704 20496 11756
rect 20904 11747 20956 11756
rect 20904 11713 20913 11747
rect 20913 11713 20947 11747
rect 20947 11713 20956 11747
rect 20904 11704 20956 11713
rect 6184 11636 6236 11688
rect 7196 11679 7248 11688
rect 7196 11645 7205 11679
rect 7205 11645 7239 11679
rect 7239 11645 7248 11679
rect 7196 11636 7248 11645
rect 4804 11568 4856 11620
rect 8576 11543 8628 11552
rect 8576 11509 8585 11543
rect 8585 11509 8619 11543
rect 8619 11509 8628 11543
rect 8576 11500 8628 11509
rect 9496 11500 9548 11552
rect 11704 11636 11756 11688
rect 20812 11636 20864 11688
rect 21088 11747 21140 11756
rect 21088 11713 21097 11747
rect 21097 11713 21131 11747
rect 21131 11713 21140 11747
rect 21088 11704 21140 11713
rect 21272 11747 21324 11756
rect 21272 11713 21281 11747
rect 21281 11713 21315 11747
rect 21315 11713 21324 11747
rect 21272 11704 21324 11713
rect 21732 11704 21784 11756
rect 15292 11500 15344 11552
rect 16028 11543 16080 11552
rect 16028 11509 16037 11543
rect 16037 11509 16071 11543
rect 16071 11509 16080 11543
rect 16028 11500 16080 11509
rect 19800 11543 19852 11552
rect 19800 11509 19809 11543
rect 19809 11509 19843 11543
rect 19843 11509 19852 11543
rect 19800 11500 19852 11509
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 65654 11398 65706 11450
rect 65718 11398 65770 11450
rect 65782 11398 65834 11450
rect 65846 11398 65898 11450
rect 65910 11398 65962 11450
rect 4436 11339 4488 11348
rect 4436 11305 4445 11339
rect 4445 11305 4479 11339
rect 4479 11305 4488 11339
rect 4436 11296 4488 11305
rect 4620 11339 4672 11348
rect 4620 11305 4629 11339
rect 4629 11305 4663 11339
rect 4663 11305 4672 11339
rect 4620 11296 4672 11305
rect 6368 11339 6420 11348
rect 6368 11305 6377 11339
rect 6377 11305 6411 11339
rect 6411 11305 6420 11339
rect 6368 11296 6420 11305
rect 9956 11296 10008 11348
rect 10508 11296 10560 11348
rect 12164 11339 12216 11348
rect 12164 11305 12173 11339
rect 12173 11305 12207 11339
rect 12207 11305 12216 11339
rect 12164 11296 12216 11305
rect 22100 11296 22152 11348
rect 23204 11339 23256 11348
rect 4344 11135 4396 11144
rect 4344 11101 4353 11135
rect 4353 11101 4387 11135
rect 4387 11101 4396 11135
rect 4344 11092 4396 11101
rect 5448 11160 5500 11212
rect 4712 11092 4764 11144
rect 5724 11135 5776 11144
rect 5724 11101 5733 11135
rect 5733 11101 5767 11135
rect 5767 11101 5776 11135
rect 5724 11092 5776 11101
rect 6184 11160 6236 11212
rect 8576 11092 8628 11144
rect 4160 11067 4212 11076
rect 4160 11033 4169 11067
rect 4169 11033 4203 11067
rect 4203 11033 4212 11067
rect 4160 11024 4212 11033
rect 19800 11228 19852 11280
rect 20628 11228 20680 11280
rect 23204 11305 23213 11339
rect 23213 11305 23247 11339
rect 23247 11305 23256 11339
rect 23204 11296 23256 11305
rect 23112 11228 23164 11280
rect 11704 11203 11756 11212
rect 11704 11169 11713 11203
rect 11713 11169 11747 11203
rect 11747 11169 11756 11203
rect 11704 11160 11756 11169
rect 13544 11203 13596 11212
rect 13544 11169 13553 11203
rect 13553 11169 13587 11203
rect 13587 11169 13596 11203
rect 13544 11160 13596 11169
rect 18696 11160 18748 11212
rect 21364 11160 21416 11212
rect 23848 11228 23900 11280
rect 11612 11092 11664 11144
rect 13728 11092 13780 11144
rect 22376 11135 22428 11144
rect 22376 11101 22385 11135
rect 22385 11101 22419 11135
rect 22419 11101 22428 11135
rect 22376 11092 22428 11101
rect 23020 11092 23072 11144
rect 23572 11092 23624 11144
rect 10692 11024 10744 11076
rect 16028 11024 16080 11076
rect 24492 11024 24544 11076
rect 23664 10999 23716 11008
rect 23664 10965 23673 10999
rect 23673 10965 23707 10999
rect 23707 10965 23716 10999
rect 23664 10956 23716 10965
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 50294 10854 50346 10906
rect 50358 10854 50410 10906
rect 50422 10854 50474 10906
rect 50486 10854 50538 10906
rect 50550 10854 50602 10906
rect 4804 10752 4856 10804
rect 4160 10727 4212 10736
rect 4160 10693 4169 10727
rect 4169 10693 4203 10727
rect 4203 10693 4212 10727
rect 4160 10684 4212 10693
rect 4712 10616 4764 10668
rect 4988 10616 5040 10668
rect 6000 10684 6052 10736
rect 10600 10752 10652 10804
rect 7196 10684 7248 10736
rect 9864 10727 9916 10736
rect 5724 10616 5776 10668
rect 9864 10693 9898 10727
rect 9898 10693 9916 10727
rect 9864 10684 9916 10693
rect 4344 10591 4396 10600
rect 4344 10557 4353 10591
rect 4353 10557 4387 10591
rect 4387 10557 4396 10591
rect 4344 10548 4396 10557
rect 5172 10548 5224 10600
rect 6184 10548 6236 10600
rect 4436 10455 4488 10464
rect 4436 10421 4445 10455
rect 4445 10421 4479 10455
rect 4479 10421 4488 10455
rect 4436 10412 4488 10421
rect 5264 10412 5316 10464
rect 6368 10412 6420 10464
rect 9496 10616 9548 10668
rect 9220 10412 9272 10464
rect 20444 10795 20496 10804
rect 13544 10684 13596 10736
rect 20444 10761 20453 10795
rect 20453 10761 20487 10795
rect 20487 10761 20496 10795
rect 20444 10752 20496 10761
rect 19156 10684 19208 10736
rect 20812 10752 20864 10804
rect 20904 10752 20956 10804
rect 17316 10659 17368 10668
rect 15660 10480 15712 10532
rect 16948 10480 17000 10532
rect 17316 10625 17325 10659
rect 17325 10625 17359 10659
rect 17359 10625 17368 10659
rect 17316 10616 17368 10625
rect 17868 10616 17920 10668
rect 20168 10616 20220 10668
rect 20628 10616 20680 10668
rect 20904 10662 20956 10671
rect 20904 10628 20913 10662
rect 20913 10628 20947 10662
rect 20947 10628 20956 10662
rect 20904 10619 20956 10628
rect 17776 10548 17828 10600
rect 20996 10548 21048 10600
rect 21272 10616 21324 10668
rect 23664 10684 23716 10736
rect 22376 10616 22428 10668
rect 22652 10616 22704 10668
rect 23848 10659 23900 10668
rect 23848 10625 23857 10659
rect 23857 10625 23891 10659
rect 23891 10625 23900 10659
rect 23848 10616 23900 10625
rect 22560 10548 22612 10600
rect 20536 10480 20588 10532
rect 12992 10412 13044 10464
rect 20444 10412 20496 10464
rect 20720 10412 20772 10464
rect 22100 10455 22152 10464
rect 22100 10421 22109 10455
rect 22109 10421 22143 10455
rect 22143 10421 22152 10455
rect 22100 10412 22152 10421
rect 23388 10455 23440 10464
rect 23388 10421 23397 10455
rect 23397 10421 23431 10455
rect 23431 10421 23440 10455
rect 23388 10412 23440 10421
rect 26976 10412 27028 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 65654 10310 65706 10362
rect 65718 10310 65770 10362
rect 65782 10310 65834 10362
rect 65846 10310 65898 10362
rect 65910 10310 65962 10362
rect 5264 10251 5316 10260
rect 5264 10217 5273 10251
rect 5273 10217 5307 10251
rect 5307 10217 5316 10251
rect 5264 10208 5316 10217
rect 5448 10251 5500 10260
rect 5448 10217 5457 10251
rect 5457 10217 5491 10251
rect 5491 10217 5500 10251
rect 5448 10208 5500 10217
rect 5448 10072 5500 10124
rect 5172 10047 5224 10056
rect 5172 10013 5181 10047
rect 5181 10013 5215 10047
rect 5215 10013 5224 10047
rect 5172 10004 5224 10013
rect 5264 10047 5316 10056
rect 5264 10013 5273 10047
rect 5273 10013 5307 10047
rect 5307 10013 5316 10047
rect 5264 10004 5316 10013
rect 5724 10004 5776 10056
rect 4988 9979 5040 9988
rect 4988 9945 4997 9979
rect 4997 9945 5031 9979
rect 5031 9945 5040 9979
rect 4988 9936 5040 9945
rect 8116 10208 8168 10260
rect 16488 10208 16540 10260
rect 20168 10251 20220 10260
rect 20168 10217 20177 10251
rect 20177 10217 20211 10251
rect 20211 10217 20220 10251
rect 20168 10208 20220 10217
rect 22100 10208 22152 10260
rect 22560 10140 22612 10192
rect 23572 10140 23624 10192
rect 23204 10072 23256 10124
rect 7104 10004 7156 10056
rect 16580 10004 16632 10056
rect 17868 10004 17920 10056
rect 20444 10047 20496 10056
rect 20444 10013 20453 10047
rect 20453 10013 20487 10047
rect 20487 10013 20496 10047
rect 20444 10004 20496 10013
rect 16212 9936 16264 9988
rect 19248 9936 19300 9988
rect 6092 9868 6144 9920
rect 6184 9868 6236 9920
rect 11244 9868 11296 9920
rect 12440 9868 12492 9920
rect 13084 9911 13136 9920
rect 13084 9877 13093 9911
rect 13093 9877 13127 9911
rect 13127 9877 13136 9911
rect 13084 9868 13136 9877
rect 14188 9911 14240 9920
rect 14188 9877 14197 9911
rect 14197 9877 14231 9911
rect 14231 9877 14240 9911
rect 14188 9868 14240 9877
rect 14740 9911 14792 9920
rect 14740 9877 14749 9911
rect 14749 9877 14783 9911
rect 14783 9877 14792 9911
rect 14740 9868 14792 9877
rect 15568 9868 15620 9920
rect 20628 10047 20680 10056
rect 20628 10013 20637 10047
rect 20637 10013 20671 10047
rect 20671 10013 20680 10047
rect 20628 10004 20680 10013
rect 20996 10004 21048 10056
rect 22652 10047 22704 10056
rect 22652 10013 22661 10047
rect 22661 10013 22695 10047
rect 22695 10013 22704 10047
rect 22652 10004 22704 10013
rect 20812 9868 20864 9920
rect 21732 9911 21784 9920
rect 21732 9877 21741 9911
rect 21741 9877 21775 9911
rect 21775 9877 21784 9911
rect 21732 9868 21784 9877
rect 23204 9868 23256 9920
rect 23296 9868 23348 9920
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 50294 9766 50346 9818
rect 50358 9766 50410 9818
rect 50422 9766 50474 9818
rect 50486 9766 50538 9818
rect 50550 9766 50602 9818
rect 6092 9664 6144 9716
rect 16488 9664 16540 9716
rect 23020 9664 23072 9716
rect 4988 9596 5040 9648
rect 12900 9596 12952 9648
rect 3332 9571 3384 9580
rect 3332 9537 3341 9571
rect 3341 9537 3375 9571
rect 3375 9537 3384 9571
rect 3332 9528 3384 9537
rect 6092 9528 6144 9580
rect 4620 9460 4672 9512
rect 5172 9460 5224 9512
rect 7748 9528 7800 9580
rect 12808 9571 12860 9580
rect 12808 9537 12817 9571
rect 12817 9537 12851 9571
rect 12851 9537 12860 9571
rect 19248 9596 19300 9648
rect 12808 9528 12860 9537
rect 12624 9460 12676 9512
rect 15568 9503 15620 9512
rect 15568 9469 15577 9503
rect 15577 9469 15611 9503
rect 15611 9469 15620 9503
rect 15568 9460 15620 9469
rect 20812 9528 20864 9580
rect 16948 9503 17000 9512
rect 16948 9469 16957 9503
rect 16957 9469 16991 9503
rect 16991 9469 17000 9503
rect 16948 9460 17000 9469
rect 20444 9460 20496 9512
rect 21732 9460 21784 9512
rect 22560 9528 22612 9580
rect 22928 9460 22980 9512
rect 23204 9571 23256 9580
rect 23204 9537 23213 9571
rect 23213 9537 23247 9571
rect 23247 9537 23256 9571
rect 23204 9528 23256 9537
rect 9036 9392 9088 9444
rect 19984 9392 20036 9444
rect 22100 9392 22152 9444
rect 23204 9392 23256 9444
rect 5632 9324 5684 9376
rect 6368 9367 6420 9376
rect 6368 9333 6377 9367
rect 6377 9333 6411 9367
rect 6411 9333 6420 9367
rect 6368 9324 6420 9333
rect 7840 9367 7892 9376
rect 7840 9333 7849 9367
rect 7849 9333 7883 9367
rect 7883 9333 7892 9367
rect 7840 9324 7892 9333
rect 9312 9367 9364 9376
rect 9312 9333 9321 9367
rect 9321 9333 9355 9367
rect 9355 9333 9364 9367
rect 9312 9324 9364 9333
rect 11520 9324 11572 9376
rect 13452 9367 13504 9376
rect 13452 9333 13461 9367
rect 13461 9333 13495 9367
rect 13495 9333 13504 9367
rect 13452 9324 13504 9333
rect 15200 9324 15252 9376
rect 18236 9324 18288 9376
rect 22652 9324 22704 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 65654 9222 65706 9274
rect 65718 9222 65770 9274
rect 65782 9222 65834 9274
rect 65846 9222 65898 9274
rect 65910 9222 65962 9274
rect 12808 9120 12860 9172
rect 20444 9120 20496 9172
rect 9496 8984 9548 9036
rect 2688 8959 2740 8968
rect 2688 8925 2697 8959
rect 2697 8925 2731 8959
rect 2731 8925 2740 8959
rect 2688 8916 2740 8925
rect 3332 8916 3384 8968
rect 3884 8916 3936 8968
rect 6184 8916 6236 8968
rect 6644 8916 6696 8968
rect 7104 8916 7156 8968
rect 9312 8916 9364 8968
rect 12532 8984 12584 9036
rect 12716 8959 12768 8968
rect 12716 8925 12725 8959
rect 12725 8925 12759 8959
rect 12759 8925 12768 8959
rect 12716 8916 12768 8925
rect 16580 8916 16632 8968
rect 20168 8916 20220 8968
rect 22100 9120 22152 9172
rect 23204 9052 23256 9104
rect 20720 8959 20772 8968
rect 20720 8925 20729 8959
rect 20729 8925 20763 8959
rect 20763 8925 20772 8959
rect 20720 8916 20772 8925
rect 21272 8916 21324 8968
rect 7288 8891 7340 8900
rect 7288 8857 7322 8891
rect 7322 8857 7340 8891
rect 7288 8848 7340 8857
rect 10140 8848 10192 8900
rect 3700 8780 3752 8832
rect 6276 8780 6328 8832
rect 6920 8780 6972 8832
rect 9588 8823 9640 8832
rect 9588 8789 9597 8823
rect 9597 8789 9631 8823
rect 9631 8789 9640 8823
rect 9588 8780 9640 8789
rect 10416 8780 10468 8832
rect 12348 8780 12400 8832
rect 13176 8848 13228 8900
rect 15476 8823 15528 8832
rect 15476 8789 15485 8823
rect 15485 8789 15519 8823
rect 15519 8789 15528 8823
rect 15476 8780 15528 8789
rect 20352 8848 20404 8900
rect 22100 8848 22152 8900
rect 22928 8848 22980 8900
rect 23296 8916 23348 8968
rect 16672 8780 16724 8832
rect 17868 8823 17920 8832
rect 17868 8789 17877 8823
rect 17877 8789 17911 8823
rect 17911 8789 17920 8823
rect 17868 8780 17920 8789
rect 18512 8780 18564 8832
rect 19432 8780 19484 8832
rect 22744 8823 22796 8832
rect 22744 8789 22753 8823
rect 22753 8789 22787 8823
rect 22787 8789 22796 8823
rect 22744 8780 22796 8789
rect 23296 8780 23348 8832
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 50294 8678 50346 8730
rect 50358 8678 50410 8730
rect 50422 8678 50474 8730
rect 50486 8678 50538 8730
rect 50550 8678 50602 8730
rect 2688 8304 2740 8356
rect 5908 8576 5960 8628
rect 5632 8508 5684 8560
rect 7288 8576 7340 8628
rect 5448 8440 5500 8492
rect 6184 8372 6236 8424
rect 6647 8483 6699 8492
rect 6647 8449 6656 8483
rect 6656 8449 6690 8483
rect 6690 8449 6699 8483
rect 6647 8440 6699 8449
rect 6920 8440 6972 8492
rect 7840 8440 7892 8492
rect 5540 8304 5592 8356
rect 9312 8576 9364 8628
rect 10140 8619 10192 8628
rect 10140 8585 10149 8619
rect 10149 8585 10183 8619
rect 10183 8585 10192 8619
rect 10140 8576 10192 8585
rect 9036 8483 9088 8492
rect 9036 8449 9045 8483
rect 9045 8449 9079 8483
rect 9079 8449 9088 8483
rect 9036 8440 9088 8449
rect 12900 8576 12952 8628
rect 13176 8619 13228 8628
rect 13176 8585 13185 8619
rect 13185 8585 13219 8619
rect 13219 8585 13228 8619
rect 13176 8576 13228 8585
rect 15108 8576 15160 8628
rect 15476 8576 15528 8628
rect 10416 8483 10468 8492
rect 10416 8449 10425 8483
rect 10425 8449 10459 8483
rect 10459 8449 10468 8483
rect 10416 8440 10468 8449
rect 10324 8372 10376 8424
rect 10784 8483 10836 8492
rect 10784 8449 10793 8483
rect 10793 8449 10827 8483
rect 10827 8449 10836 8483
rect 11612 8483 11664 8492
rect 10784 8440 10836 8449
rect 11612 8449 11621 8483
rect 11621 8449 11655 8483
rect 11655 8449 11664 8483
rect 11612 8440 11664 8449
rect 12256 8440 12308 8492
rect 12532 8483 12584 8492
rect 12532 8449 12541 8483
rect 12541 8449 12575 8483
rect 12575 8449 12584 8483
rect 12532 8440 12584 8449
rect 13544 8508 13596 8560
rect 10876 8372 10928 8424
rect 11796 8415 11848 8424
rect 11796 8381 11805 8415
rect 11805 8381 11839 8415
rect 11839 8381 11848 8415
rect 11796 8372 11848 8381
rect 5448 8236 5500 8288
rect 5724 8279 5776 8288
rect 5724 8245 5733 8279
rect 5733 8245 5767 8279
rect 5767 8245 5776 8279
rect 9680 8279 9732 8288
rect 5724 8236 5776 8245
rect 9680 8245 9689 8279
rect 9689 8245 9723 8279
rect 9723 8245 9732 8279
rect 9680 8236 9732 8245
rect 10048 8236 10100 8288
rect 10784 8236 10836 8288
rect 11612 8279 11664 8288
rect 11612 8245 11621 8279
rect 11621 8245 11655 8279
rect 11655 8245 11664 8279
rect 11612 8236 11664 8245
rect 13176 8440 13228 8492
rect 13452 8440 13504 8492
rect 18144 8483 18196 8492
rect 18144 8449 18153 8483
rect 18153 8449 18187 8483
rect 18187 8449 18196 8483
rect 18144 8440 18196 8449
rect 18972 8576 19024 8628
rect 20352 8576 20404 8628
rect 20536 8576 20588 8628
rect 22744 8508 22796 8560
rect 23296 8508 23348 8560
rect 20260 8483 20312 8492
rect 20260 8449 20269 8483
rect 20269 8449 20303 8483
rect 20303 8449 20312 8483
rect 20260 8440 20312 8449
rect 20444 8440 20496 8492
rect 16120 8372 16172 8424
rect 16672 8415 16724 8424
rect 16672 8381 16681 8415
rect 16681 8381 16715 8415
rect 16715 8381 16724 8415
rect 16672 8372 16724 8381
rect 17316 8372 17368 8424
rect 19156 8372 19208 8424
rect 21272 8415 21324 8424
rect 21272 8381 21281 8415
rect 21281 8381 21315 8415
rect 21315 8381 21324 8415
rect 21272 8372 21324 8381
rect 21548 8440 21600 8492
rect 21916 8440 21968 8492
rect 22100 8483 22152 8492
rect 22100 8449 22109 8483
rect 22109 8449 22143 8483
rect 22143 8449 22152 8483
rect 22100 8440 22152 8449
rect 23204 8483 23256 8492
rect 23204 8449 23213 8483
rect 23213 8449 23247 8483
rect 23247 8449 23256 8483
rect 23204 8440 23256 8449
rect 23388 8483 23440 8492
rect 23388 8449 23397 8483
rect 23397 8449 23431 8483
rect 23431 8449 23440 8483
rect 23388 8440 23440 8449
rect 24308 8483 24360 8492
rect 24308 8449 24317 8483
rect 24317 8449 24351 8483
rect 24351 8449 24360 8483
rect 24308 8440 24360 8449
rect 13636 8347 13688 8356
rect 13636 8313 13645 8347
rect 13645 8313 13679 8347
rect 13679 8313 13688 8347
rect 13636 8304 13688 8313
rect 14280 8347 14332 8356
rect 14280 8313 14289 8347
rect 14289 8313 14323 8347
rect 14323 8313 14332 8347
rect 14280 8304 14332 8313
rect 19340 8304 19392 8356
rect 12624 8236 12676 8288
rect 12808 8236 12860 8288
rect 20076 8279 20128 8288
rect 20076 8245 20085 8279
rect 20085 8245 20119 8279
rect 20119 8245 20128 8279
rect 20076 8236 20128 8245
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 65654 8134 65706 8186
rect 65718 8134 65770 8186
rect 65782 8134 65834 8186
rect 65846 8134 65898 8186
rect 65910 8134 65962 8186
rect 5448 8032 5500 8084
rect 8392 8075 8444 8084
rect 4068 7964 4120 8016
rect 8392 8041 8401 8075
rect 8401 8041 8435 8075
rect 8435 8041 8444 8075
rect 8392 8032 8444 8041
rect 9588 8075 9640 8084
rect 9588 8041 9597 8075
rect 9597 8041 9631 8075
rect 9631 8041 9640 8075
rect 9588 8032 9640 8041
rect 10876 8032 10928 8084
rect 11612 8032 11664 8084
rect 5540 7896 5592 7948
rect 5632 7871 5684 7880
rect 5632 7837 5641 7871
rect 5641 7837 5675 7871
rect 5675 7837 5684 7871
rect 5632 7828 5684 7837
rect 9680 7896 9732 7948
rect 11796 7896 11848 7948
rect 4620 7760 4672 7812
rect 4804 7692 4856 7744
rect 7104 7828 7156 7880
rect 9404 7871 9456 7880
rect 9404 7837 9413 7871
rect 9413 7837 9447 7871
rect 9447 7837 9456 7871
rect 9404 7828 9456 7837
rect 8760 7760 8812 7812
rect 13360 8032 13412 8084
rect 13544 8075 13596 8084
rect 13544 8041 13553 8075
rect 13553 8041 13587 8075
rect 13587 8041 13596 8075
rect 13544 8032 13596 8041
rect 16580 8032 16632 8084
rect 21548 8075 21600 8084
rect 21548 8041 21557 8075
rect 21557 8041 21591 8075
rect 21591 8041 21600 8075
rect 21548 8032 21600 8041
rect 21732 8032 21784 8084
rect 15476 7964 15528 8016
rect 20352 7964 20404 8016
rect 12808 7896 12860 7948
rect 12532 7828 12584 7880
rect 10508 7760 10560 7812
rect 11704 7760 11756 7812
rect 14280 7828 14332 7880
rect 15200 7871 15252 7880
rect 15200 7837 15209 7871
rect 15209 7837 15243 7871
rect 15243 7837 15252 7871
rect 15200 7828 15252 7837
rect 16028 7828 16080 7880
rect 17868 7828 17920 7880
rect 18144 7828 18196 7880
rect 20076 7828 20128 7880
rect 21456 7871 21508 7880
rect 21456 7837 21465 7871
rect 21465 7837 21499 7871
rect 21499 7837 21508 7871
rect 21456 7828 21508 7837
rect 23296 7964 23348 8016
rect 23204 7896 23256 7948
rect 23112 7871 23164 7880
rect 23112 7837 23121 7871
rect 23121 7837 23155 7871
rect 23155 7837 23164 7871
rect 23112 7828 23164 7837
rect 6644 7692 6696 7744
rect 10232 7692 10284 7744
rect 11888 7692 11940 7744
rect 14740 7760 14792 7812
rect 15384 7760 15436 7812
rect 15660 7803 15712 7812
rect 15660 7769 15669 7803
rect 15669 7769 15703 7803
rect 15703 7769 15712 7803
rect 15660 7760 15712 7769
rect 14372 7735 14424 7744
rect 14372 7701 14381 7735
rect 14381 7701 14415 7735
rect 14415 7701 14424 7735
rect 14372 7692 14424 7701
rect 15016 7735 15068 7744
rect 15016 7701 15025 7735
rect 15025 7701 15059 7735
rect 15059 7701 15068 7735
rect 15016 7692 15068 7701
rect 15200 7692 15252 7744
rect 18880 7692 18932 7744
rect 20352 7692 20404 7744
rect 22284 7692 22336 7744
rect 24400 7735 24452 7744
rect 24400 7701 24409 7735
rect 24409 7701 24443 7735
rect 24443 7701 24452 7735
rect 24400 7692 24452 7701
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 50294 7590 50346 7642
rect 50358 7590 50410 7642
rect 50422 7590 50474 7642
rect 50486 7590 50538 7642
rect 50550 7590 50602 7642
rect 5632 7488 5684 7540
rect 6184 7488 6236 7540
rect 10324 7488 10376 7540
rect 11704 7488 11756 7540
rect 12440 7488 12492 7540
rect 16948 7488 17000 7540
rect 5356 7420 5408 7472
rect 7104 7420 7156 7472
rect 10784 7420 10836 7472
rect 3884 7352 3936 7404
rect 4988 7395 5040 7404
rect 4988 7361 4997 7395
rect 4997 7361 5031 7395
rect 5031 7361 5040 7395
rect 4988 7352 5040 7361
rect 6092 7352 6144 7404
rect 9496 7352 9548 7404
rect 9588 7395 9640 7404
rect 9588 7361 9597 7395
rect 9597 7361 9631 7395
rect 9631 7361 9640 7395
rect 10048 7395 10100 7404
rect 9588 7352 9640 7361
rect 10048 7361 10057 7395
rect 10057 7361 10091 7395
rect 10091 7361 10100 7395
rect 10048 7352 10100 7361
rect 10232 7395 10284 7404
rect 10232 7361 10236 7395
rect 10236 7361 10270 7395
rect 10270 7361 10284 7395
rect 10232 7352 10284 7361
rect 11888 7420 11940 7472
rect 12808 7420 12860 7472
rect 20444 7488 20496 7540
rect 19340 7420 19392 7472
rect 5540 7284 5592 7336
rect 10324 7216 10376 7268
rect 12716 7352 12768 7404
rect 15936 7395 15988 7404
rect 11704 7216 11756 7268
rect 12164 7216 12216 7268
rect 12716 7216 12768 7268
rect 15936 7361 15945 7395
rect 15945 7361 15979 7395
rect 15979 7361 15988 7395
rect 15936 7352 15988 7361
rect 16856 7352 16908 7404
rect 17132 7395 17184 7404
rect 17132 7361 17141 7395
rect 17141 7361 17175 7395
rect 17175 7361 17184 7395
rect 17132 7352 17184 7361
rect 17316 7395 17368 7404
rect 17316 7361 17325 7395
rect 17325 7361 17359 7395
rect 17359 7361 17368 7395
rect 18144 7395 18196 7404
rect 17316 7352 17368 7361
rect 18144 7361 18153 7395
rect 18153 7361 18187 7395
rect 18187 7361 18196 7395
rect 18144 7352 18196 7361
rect 19156 7352 19208 7404
rect 21456 7488 21508 7540
rect 22008 7395 22060 7404
rect 22008 7361 22017 7395
rect 22017 7361 22051 7395
rect 22051 7361 22060 7395
rect 22008 7352 22060 7361
rect 23756 7488 23808 7540
rect 23296 7395 23348 7404
rect 23296 7361 23305 7395
rect 23305 7361 23339 7395
rect 23339 7361 23348 7395
rect 23296 7352 23348 7361
rect 17500 7284 17552 7336
rect 22560 7327 22612 7336
rect 22560 7293 22569 7327
rect 22569 7293 22603 7327
rect 22603 7293 22612 7327
rect 22560 7284 22612 7293
rect 23020 7284 23072 7336
rect 5724 7148 5776 7200
rect 7932 7148 7984 7200
rect 11060 7148 11112 7200
rect 11888 7148 11940 7200
rect 12348 7148 12400 7200
rect 17592 7216 17644 7268
rect 21456 7216 21508 7268
rect 12900 7191 12952 7200
rect 12900 7157 12909 7191
rect 12909 7157 12943 7191
rect 12943 7157 12952 7191
rect 14648 7191 14700 7200
rect 12900 7148 12952 7157
rect 14648 7157 14657 7191
rect 14657 7157 14691 7191
rect 14691 7157 14700 7191
rect 14648 7148 14700 7157
rect 15660 7148 15712 7200
rect 16672 7191 16724 7200
rect 16672 7157 16681 7191
rect 16681 7157 16715 7191
rect 16715 7157 16724 7191
rect 16672 7148 16724 7157
rect 20720 7148 20772 7200
rect 21548 7148 21600 7200
rect 24400 7284 24452 7336
rect 23572 7148 23624 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 65654 7046 65706 7098
rect 65718 7046 65770 7098
rect 65782 7046 65834 7098
rect 65846 7046 65898 7098
rect 65910 7046 65962 7098
rect 6092 6944 6144 6996
rect 8392 6944 8444 6996
rect 10508 6944 10560 6996
rect 13360 6987 13412 6996
rect 13360 6953 13369 6987
rect 13369 6953 13403 6987
rect 13403 6953 13412 6987
rect 13360 6944 13412 6953
rect 14924 6987 14976 6996
rect 14924 6953 14933 6987
rect 14933 6953 14967 6987
rect 14967 6953 14976 6987
rect 14924 6944 14976 6953
rect 15476 6987 15528 6996
rect 15476 6953 15485 6987
rect 15485 6953 15519 6987
rect 15519 6953 15528 6987
rect 15476 6944 15528 6953
rect 16856 6944 16908 6996
rect 20260 6944 20312 6996
rect 20812 6944 20864 6996
rect 24400 6987 24452 6996
rect 24400 6953 24409 6987
rect 24409 6953 24443 6987
rect 24443 6953 24452 6987
rect 24400 6944 24452 6953
rect 12532 6876 12584 6928
rect 2688 6808 2740 6860
rect 5172 6808 5224 6860
rect 5448 6740 5500 6792
rect 5632 6740 5684 6792
rect 6092 6783 6144 6792
rect 6092 6749 6101 6783
rect 6101 6749 6135 6783
rect 6135 6749 6144 6783
rect 6092 6740 6144 6749
rect 6644 6672 6696 6724
rect 10784 6808 10836 6860
rect 14280 6808 14332 6860
rect 15936 6808 15988 6860
rect 16120 6851 16172 6860
rect 16120 6817 16129 6851
rect 16129 6817 16163 6851
rect 16163 6817 16172 6851
rect 16120 6808 16172 6817
rect 22008 6876 22060 6928
rect 20996 6808 21048 6860
rect 23296 6808 23348 6860
rect 24492 6851 24544 6860
rect 8300 6740 8352 6792
rect 9220 6783 9272 6792
rect 9220 6749 9229 6783
rect 9229 6749 9263 6783
rect 9263 6749 9272 6783
rect 9220 6740 9272 6749
rect 10140 6783 10192 6792
rect 9220 6604 9272 6656
rect 10140 6749 10149 6783
rect 10149 6749 10183 6783
rect 10183 6749 10192 6783
rect 10140 6740 10192 6749
rect 11244 6740 11296 6792
rect 11520 6740 11572 6792
rect 10048 6672 10100 6724
rect 10600 6604 10652 6656
rect 10692 6604 10744 6656
rect 11336 6604 11388 6656
rect 12072 6647 12124 6656
rect 12072 6613 12081 6647
rect 12081 6613 12115 6647
rect 12115 6613 12124 6647
rect 12072 6604 12124 6613
rect 13544 6783 13596 6792
rect 13544 6749 13553 6783
rect 13553 6749 13587 6783
rect 13587 6749 13596 6783
rect 13544 6740 13596 6749
rect 14096 6740 14148 6792
rect 15016 6783 15068 6792
rect 15016 6749 15025 6783
rect 15025 6749 15059 6783
rect 15059 6749 15068 6783
rect 15016 6740 15068 6749
rect 15752 6740 15804 6792
rect 16672 6740 16724 6792
rect 18880 6740 18932 6792
rect 13084 6672 13136 6724
rect 14740 6672 14792 6724
rect 18788 6672 18840 6724
rect 13820 6604 13872 6656
rect 13912 6604 13964 6656
rect 16672 6604 16724 6656
rect 20536 6672 20588 6724
rect 21456 6783 21508 6792
rect 21456 6749 21465 6783
rect 21465 6749 21499 6783
rect 21499 6749 21508 6783
rect 21456 6740 21508 6749
rect 22468 6740 22520 6792
rect 23388 6783 23440 6792
rect 23388 6749 23397 6783
rect 23397 6749 23431 6783
rect 23431 6749 23440 6783
rect 23388 6740 23440 6749
rect 22100 6672 22152 6724
rect 23296 6672 23348 6724
rect 19432 6647 19484 6656
rect 19432 6613 19441 6647
rect 19441 6613 19475 6647
rect 19475 6613 19484 6647
rect 19432 6604 19484 6613
rect 20720 6604 20772 6656
rect 21180 6604 21232 6656
rect 23664 6740 23716 6792
rect 24492 6817 24501 6851
rect 24501 6817 24535 6851
rect 24535 6817 24544 6851
rect 24492 6808 24544 6817
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 50294 6502 50346 6554
rect 50358 6502 50410 6554
rect 50422 6502 50474 6554
rect 50486 6502 50538 6554
rect 50550 6502 50602 6554
rect 2688 6307 2740 6316
rect 2688 6273 2697 6307
rect 2697 6273 2731 6307
rect 2731 6273 2740 6307
rect 2688 6264 2740 6273
rect 3700 6332 3752 6384
rect 8392 6400 8444 6452
rect 10048 6400 10100 6452
rect 10232 6443 10284 6452
rect 10232 6409 10241 6443
rect 10241 6409 10275 6443
rect 10275 6409 10284 6443
rect 10232 6400 10284 6409
rect 5356 6375 5408 6384
rect 5356 6341 5365 6375
rect 5365 6341 5399 6375
rect 5399 6341 5408 6375
rect 5356 6332 5408 6341
rect 12532 6400 12584 6452
rect 12808 6400 12860 6452
rect 14096 6400 14148 6452
rect 3792 6264 3844 6316
rect 4068 6307 4120 6316
rect 4068 6273 4077 6307
rect 4077 6273 4111 6307
rect 4111 6273 4120 6307
rect 5540 6307 5592 6316
rect 4068 6264 4120 6273
rect 5540 6273 5549 6307
rect 5549 6273 5583 6307
rect 5583 6273 5592 6307
rect 5540 6264 5592 6273
rect 6276 6264 6328 6316
rect 9220 6264 9272 6316
rect 3884 6196 3936 6248
rect 5264 6128 5316 6180
rect 5448 6196 5500 6248
rect 9864 6196 9916 6248
rect 6552 6128 6604 6180
rect 10048 6307 10100 6316
rect 10048 6273 10057 6307
rect 10057 6273 10091 6307
rect 10091 6273 10100 6307
rect 10048 6264 10100 6273
rect 10600 6332 10652 6384
rect 10692 6264 10744 6316
rect 12164 6332 12216 6384
rect 11612 6307 11664 6316
rect 11612 6273 11621 6307
rect 11621 6273 11655 6307
rect 11655 6273 11664 6307
rect 11612 6264 11664 6273
rect 11704 6264 11756 6316
rect 12716 6332 12768 6384
rect 12900 6332 12952 6384
rect 13544 6332 13596 6384
rect 14188 6332 14240 6384
rect 16948 6400 17000 6452
rect 18420 6400 18472 6452
rect 12808 6264 12860 6316
rect 13728 6264 13780 6316
rect 15016 6307 15068 6316
rect 15016 6273 15025 6307
rect 15025 6273 15059 6307
rect 15059 6273 15068 6307
rect 15016 6264 15068 6273
rect 15108 6307 15160 6316
rect 15108 6273 15117 6307
rect 15117 6273 15151 6307
rect 15151 6273 15160 6307
rect 15108 6264 15160 6273
rect 12900 6239 12952 6248
rect 12900 6205 12909 6239
rect 12909 6205 12943 6239
rect 12943 6205 12952 6239
rect 12900 6196 12952 6205
rect 18512 6264 18564 6316
rect 19064 6332 19116 6384
rect 19984 6264 20036 6316
rect 20536 6264 20588 6316
rect 20812 6264 20864 6316
rect 22100 6400 22152 6452
rect 22284 6307 22336 6316
rect 22284 6273 22293 6307
rect 22293 6273 22327 6307
rect 22327 6273 22336 6307
rect 22284 6264 22336 6273
rect 22468 6307 22520 6316
rect 22468 6273 22477 6307
rect 22477 6273 22511 6307
rect 22511 6273 22520 6307
rect 22468 6264 22520 6273
rect 23664 6264 23716 6316
rect 18236 6196 18288 6248
rect 22928 6239 22980 6248
rect 12256 6171 12308 6180
rect 12256 6137 12265 6171
rect 12265 6137 12299 6171
rect 12299 6137 12308 6171
rect 12256 6128 12308 6137
rect 12624 6128 12676 6180
rect 3792 6060 3844 6112
rect 3976 6103 4028 6112
rect 3976 6069 3985 6103
rect 3985 6069 4019 6103
rect 4019 6069 4028 6103
rect 3976 6060 4028 6069
rect 5724 6060 5776 6112
rect 6092 6060 6144 6112
rect 6828 6060 6880 6112
rect 7840 6060 7892 6112
rect 8668 6060 8720 6112
rect 9220 6060 9272 6112
rect 9680 6060 9732 6112
rect 11612 6060 11664 6112
rect 12072 6060 12124 6112
rect 13636 6060 13688 6112
rect 15292 6128 15344 6180
rect 14924 6060 14976 6112
rect 15568 6060 15620 6112
rect 16580 6128 16632 6180
rect 16856 6060 16908 6112
rect 17040 6103 17092 6112
rect 17040 6069 17049 6103
rect 17049 6069 17083 6103
rect 17083 6069 17092 6103
rect 17040 6060 17092 6069
rect 19248 6060 19300 6112
rect 22928 6205 22937 6239
rect 22937 6205 22971 6239
rect 22971 6205 22980 6239
rect 22928 6196 22980 6205
rect 20260 6128 20312 6180
rect 21180 6128 21232 6180
rect 23204 6128 23256 6180
rect 20444 6103 20496 6112
rect 20444 6069 20453 6103
rect 20453 6069 20487 6103
rect 20487 6069 20496 6103
rect 20444 6060 20496 6069
rect 21272 6103 21324 6112
rect 21272 6069 21281 6103
rect 21281 6069 21315 6103
rect 21315 6069 21324 6103
rect 21272 6060 21324 6069
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 65654 5958 65706 6010
rect 65718 5958 65770 6010
rect 65782 5958 65834 6010
rect 65846 5958 65898 6010
rect 65910 5958 65962 6010
rect 3976 5899 4028 5908
rect 3976 5865 3985 5899
rect 3985 5865 4019 5899
rect 4019 5865 4028 5899
rect 3976 5856 4028 5865
rect 5724 5856 5776 5908
rect 7748 5899 7800 5908
rect 7748 5865 7757 5899
rect 7757 5865 7791 5899
rect 7791 5865 7800 5899
rect 7748 5856 7800 5865
rect 8392 5856 8444 5908
rect 8852 5856 8904 5908
rect 9036 5899 9088 5908
rect 9036 5865 9045 5899
rect 9045 5865 9079 5899
rect 9079 5865 9088 5899
rect 9036 5856 9088 5865
rect 9496 5899 9548 5908
rect 9496 5865 9505 5899
rect 9505 5865 9539 5899
rect 9539 5865 9548 5899
rect 9496 5856 9548 5865
rect 11520 5856 11572 5908
rect 13360 5856 13412 5908
rect 13820 5856 13872 5908
rect 14832 5856 14884 5908
rect 14924 5899 14976 5908
rect 14924 5865 14933 5899
rect 14933 5865 14967 5899
rect 14967 5865 14976 5899
rect 14924 5856 14976 5865
rect 6460 5788 6512 5840
rect 6552 5788 6604 5840
rect 5448 5763 5500 5772
rect 5448 5729 5457 5763
rect 5457 5729 5491 5763
rect 5491 5729 5500 5763
rect 5448 5720 5500 5729
rect 3792 5695 3844 5704
rect 3792 5661 3801 5695
rect 3801 5661 3835 5695
rect 3835 5661 3844 5695
rect 3792 5652 3844 5661
rect 5356 5652 5408 5704
rect 7564 5720 7616 5772
rect 7840 5788 7892 5840
rect 9680 5788 9732 5840
rect 15752 5856 15804 5908
rect 16120 5856 16172 5908
rect 18052 5856 18104 5908
rect 20168 5856 20220 5908
rect 23388 5856 23440 5908
rect 24308 5856 24360 5908
rect 15292 5788 15344 5840
rect 17224 5788 17276 5840
rect 12072 5720 12124 5772
rect 14096 5720 14148 5772
rect 14280 5720 14332 5772
rect 18052 5720 18104 5772
rect 19248 5763 19300 5772
rect 19248 5729 19257 5763
rect 19257 5729 19291 5763
rect 19291 5729 19300 5763
rect 19248 5720 19300 5729
rect 21916 5763 21968 5772
rect 21916 5729 21925 5763
rect 21925 5729 21959 5763
rect 21959 5729 21968 5763
rect 21916 5720 21968 5729
rect 22100 5720 22152 5772
rect 5632 5652 5684 5704
rect 6184 5695 6236 5704
rect 6184 5661 6193 5695
rect 6193 5661 6227 5695
rect 6227 5661 6236 5695
rect 6184 5652 6236 5661
rect 6368 5695 6420 5704
rect 6368 5661 6377 5695
rect 6377 5661 6411 5695
rect 6411 5661 6420 5695
rect 6368 5652 6420 5661
rect 6276 5584 6328 5636
rect 6736 5652 6788 5704
rect 7932 5695 7984 5704
rect 7932 5661 7941 5695
rect 7941 5661 7975 5695
rect 7975 5661 7984 5695
rect 7932 5652 7984 5661
rect 9680 5695 9732 5704
rect 9680 5661 9689 5695
rect 9689 5661 9723 5695
rect 9723 5661 9732 5695
rect 9680 5652 9732 5661
rect 10140 5695 10192 5704
rect 10140 5661 10149 5695
rect 10149 5661 10183 5695
rect 10183 5661 10192 5695
rect 10140 5652 10192 5661
rect 10784 5695 10836 5704
rect 10784 5661 10793 5695
rect 10793 5661 10827 5695
rect 10827 5661 10836 5695
rect 10784 5652 10836 5661
rect 12900 5652 12952 5704
rect 12992 5652 13044 5704
rect 14188 5695 14240 5704
rect 14188 5661 14197 5695
rect 14197 5661 14231 5695
rect 14231 5661 14240 5695
rect 14188 5652 14240 5661
rect 15660 5695 15712 5704
rect 6644 5584 6696 5636
rect 11060 5627 11112 5636
rect 11060 5593 11094 5627
rect 11094 5593 11112 5627
rect 11060 5584 11112 5593
rect 6552 5516 6604 5568
rect 7288 5516 7340 5568
rect 12072 5584 12124 5636
rect 11612 5516 11664 5568
rect 13084 5516 13136 5568
rect 13728 5516 13780 5568
rect 15660 5661 15669 5695
rect 15669 5661 15703 5695
rect 15703 5661 15712 5695
rect 15660 5652 15712 5661
rect 17684 5652 17736 5704
rect 19340 5652 19392 5704
rect 20812 5652 20864 5704
rect 21180 5652 21232 5704
rect 15844 5516 15896 5568
rect 20260 5584 20312 5636
rect 20444 5516 20496 5568
rect 23204 5559 23256 5568
rect 23204 5525 23213 5559
rect 23213 5525 23247 5559
rect 23247 5525 23256 5559
rect 23204 5516 23256 5525
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 50294 5414 50346 5466
rect 50358 5414 50410 5466
rect 50422 5414 50474 5466
rect 50486 5414 50538 5466
rect 50550 5414 50602 5466
rect 4804 5312 4856 5364
rect 3792 5176 3844 5228
rect 9588 5287 9640 5296
rect 9588 5253 9597 5287
rect 9597 5253 9631 5287
rect 9631 5253 9640 5287
rect 9588 5244 9640 5253
rect 10048 5312 10100 5364
rect 11796 5312 11848 5364
rect 12164 5312 12216 5364
rect 14924 5312 14976 5364
rect 16396 5312 16448 5364
rect 16672 5355 16724 5364
rect 16672 5321 16681 5355
rect 16681 5321 16715 5355
rect 16715 5321 16724 5355
rect 16672 5312 16724 5321
rect 20628 5312 20680 5364
rect 21088 5312 21140 5364
rect 23664 5312 23716 5364
rect 12072 5244 12124 5296
rect 14556 5244 14608 5296
rect 20720 5244 20772 5296
rect 23296 5244 23348 5296
rect 6184 5176 6236 5228
rect 6552 5219 6604 5228
rect 6552 5185 6561 5219
rect 6561 5185 6595 5219
rect 6595 5185 6604 5219
rect 6552 5176 6604 5185
rect 5172 5108 5224 5160
rect 4988 5040 5040 5092
rect 3976 4972 4028 5024
rect 5172 4972 5224 5024
rect 6920 5176 6972 5228
rect 8392 5176 8444 5228
rect 10416 5176 10468 5228
rect 11704 5219 11756 5228
rect 11704 5185 11713 5219
rect 11713 5185 11747 5219
rect 11747 5185 11756 5219
rect 11704 5176 11756 5185
rect 12808 5219 12860 5228
rect 12808 5185 12817 5219
rect 12817 5185 12851 5219
rect 12851 5185 12860 5219
rect 12808 5176 12860 5185
rect 12440 5108 12492 5160
rect 12992 5219 13044 5228
rect 12992 5185 13001 5219
rect 13001 5185 13035 5219
rect 13035 5185 13044 5219
rect 12992 5176 13044 5185
rect 13636 5219 13688 5228
rect 13636 5185 13645 5219
rect 13645 5185 13679 5219
rect 13679 5185 13688 5219
rect 13636 5176 13688 5185
rect 15568 5219 15620 5228
rect 15568 5185 15577 5219
rect 15577 5185 15611 5219
rect 15611 5185 15620 5219
rect 15568 5176 15620 5185
rect 18052 5219 18104 5228
rect 18052 5185 18061 5219
rect 18061 5185 18095 5219
rect 18095 5185 18104 5219
rect 18052 5176 18104 5185
rect 19432 5176 19484 5228
rect 13544 5108 13596 5160
rect 15476 5151 15528 5160
rect 15476 5117 15485 5151
rect 15485 5117 15519 5151
rect 15519 5117 15528 5151
rect 15476 5108 15528 5117
rect 6644 5040 6696 5092
rect 9864 5040 9916 5092
rect 6828 4972 6880 5024
rect 8300 5015 8352 5024
rect 8300 4981 8309 5015
rect 8309 4981 8343 5015
rect 8343 4981 8352 5015
rect 8300 4972 8352 4981
rect 10324 5015 10376 5024
rect 10324 4981 10333 5015
rect 10333 4981 10367 5015
rect 10367 4981 10376 5015
rect 10324 4972 10376 4981
rect 11612 4972 11664 5024
rect 12164 5040 12216 5092
rect 19708 5040 19760 5092
rect 12256 4972 12308 5024
rect 12532 5015 12584 5024
rect 12532 4981 12541 5015
rect 12541 4981 12575 5015
rect 12575 4981 12584 5015
rect 12532 4972 12584 4981
rect 15292 5015 15344 5024
rect 15292 4981 15301 5015
rect 15301 4981 15335 5015
rect 15335 4981 15344 5015
rect 15292 4972 15344 4981
rect 19064 4972 19116 5024
rect 19248 4972 19300 5024
rect 19800 4972 19852 5024
rect 20444 5108 20496 5160
rect 20812 5219 20864 5228
rect 20812 5185 20821 5219
rect 20821 5185 20855 5219
rect 20855 5185 20864 5219
rect 20812 5176 20864 5185
rect 21456 5176 21508 5228
rect 21548 5176 21600 5228
rect 22836 5176 22888 5228
rect 23756 5219 23808 5228
rect 23756 5185 23765 5219
rect 23765 5185 23799 5219
rect 23799 5185 23808 5219
rect 23756 5176 23808 5185
rect 20720 5040 20772 5092
rect 21272 4972 21324 5024
rect 21824 5015 21876 5024
rect 21824 4981 21833 5015
rect 21833 4981 21867 5015
rect 21867 4981 21876 5015
rect 21824 4972 21876 4981
rect 22284 4972 22336 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 65654 4870 65706 4922
rect 65718 4870 65770 4922
rect 65782 4870 65834 4922
rect 65846 4870 65898 4922
rect 65910 4870 65962 4922
rect 3976 4811 4028 4820
rect 3976 4777 3985 4811
rect 3985 4777 4019 4811
rect 4019 4777 4028 4811
rect 3976 4768 4028 4777
rect 4620 4768 4672 4820
rect 5724 4811 5776 4820
rect 5724 4777 5733 4811
rect 5733 4777 5767 4811
rect 5767 4777 5776 4811
rect 5724 4768 5776 4777
rect 6368 4768 6420 4820
rect 8392 4811 8444 4820
rect 8392 4777 8401 4811
rect 8401 4777 8435 4811
rect 8435 4777 8444 4811
rect 8392 4768 8444 4777
rect 12072 4768 12124 4820
rect 12164 4768 12216 4820
rect 12992 4768 13044 4820
rect 14096 4768 14148 4820
rect 15292 4768 15344 4820
rect 15936 4811 15988 4820
rect 6736 4700 6788 4752
rect 15936 4777 15945 4811
rect 15945 4777 15979 4811
rect 15979 4777 15988 4811
rect 15936 4768 15988 4777
rect 17132 4768 17184 4820
rect 17776 4811 17828 4820
rect 17776 4777 17785 4811
rect 17785 4777 17819 4811
rect 17819 4777 17828 4811
rect 17776 4768 17828 4777
rect 18788 4768 18840 4820
rect 19156 4768 19208 4820
rect 5540 4675 5592 4684
rect 5540 4641 5549 4675
rect 5549 4641 5583 4675
rect 5583 4641 5592 4675
rect 5540 4632 5592 4641
rect 11612 4632 11664 4684
rect 3792 4607 3844 4616
rect 3792 4573 3801 4607
rect 3801 4573 3835 4607
rect 3835 4573 3844 4607
rect 3792 4564 3844 4573
rect 4896 4564 4948 4616
rect 5356 4564 5408 4616
rect 5724 4607 5776 4616
rect 5724 4573 5733 4607
rect 5733 4573 5767 4607
rect 5767 4573 5776 4607
rect 5724 4564 5776 4573
rect 6552 4607 6604 4616
rect 6552 4573 6561 4607
rect 6561 4573 6595 4607
rect 6595 4573 6604 4607
rect 6552 4564 6604 4573
rect 8300 4564 8352 4616
rect 9496 4607 9548 4616
rect 9496 4573 9505 4607
rect 9505 4573 9539 4607
rect 9539 4573 9548 4607
rect 9496 4564 9548 4573
rect 9588 4564 9640 4616
rect 10784 4564 10836 4616
rect 11704 4564 11756 4616
rect 13728 4632 13780 4684
rect 15476 4632 15528 4684
rect 13268 4607 13320 4616
rect 13268 4573 13277 4607
rect 13277 4573 13311 4607
rect 13311 4573 13320 4607
rect 13268 4564 13320 4573
rect 14556 4607 14608 4616
rect 14556 4573 14565 4607
rect 14565 4573 14599 4607
rect 14599 4573 14608 4607
rect 14556 4564 14608 4573
rect 15200 4564 15252 4616
rect 16488 4564 16540 4616
rect 7288 4539 7340 4548
rect 7288 4505 7322 4539
rect 7322 4505 7340 4539
rect 7288 4496 7340 4505
rect 12532 4496 12584 4548
rect 16672 4607 16724 4616
rect 16672 4573 16697 4607
rect 16697 4573 16724 4607
rect 16672 4564 16724 4573
rect 20904 4811 20956 4820
rect 20904 4777 20913 4811
rect 20913 4777 20947 4811
rect 20947 4777 20956 4811
rect 20904 4768 20956 4777
rect 21272 4811 21324 4820
rect 21272 4777 21281 4811
rect 21281 4777 21315 4811
rect 21315 4777 21324 4811
rect 21916 4811 21968 4820
rect 21272 4768 21324 4777
rect 21916 4777 21925 4811
rect 21925 4777 21959 4811
rect 21959 4777 21968 4811
rect 21916 4768 21968 4777
rect 21364 4700 21416 4752
rect 21640 4700 21692 4752
rect 23296 4700 23348 4752
rect 20536 4632 20588 4684
rect 17592 4607 17644 4616
rect 17592 4573 17601 4607
rect 17601 4573 17635 4607
rect 17635 4573 17644 4607
rect 17592 4564 17644 4573
rect 18420 4564 18472 4616
rect 19616 4607 19668 4616
rect 19616 4573 19625 4607
rect 19625 4573 19659 4607
rect 19659 4573 19668 4607
rect 19616 4564 19668 4573
rect 20628 4564 20680 4616
rect 20996 4564 21048 4616
rect 22100 4607 22152 4616
rect 4068 4428 4120 4480
rect 9404 4428 9456 4480
rect 9680 4428 9732 4480
rect 12808 4428 12860 4480
rect 13820 4428 13872 4480
rect 16304 4428 16356 4480
rect 20904 4496 20956 4548
rect 21456 4496 21508 4548
rect 22100 4573 22109 4607
rect 22109 4573 22143 4607
rect 22143 4573 22152 4607
rect 22100 4564 22152 4573
rect 23572 4564 23624 4616
rect 23664 4607 23716 4616
rect 23664 4573 23673 4607
rect 23673 4573 23707 4607
rect 23707 4573 23716 4607
rect 24400 4607 24452 4616
rect 23664 4564 23716 4573
rect 24400 4573 24409 4607
rect 24409 4573 24443 4607
rect 24443 4573 24452 4607
rect 24400 4564 24452 4573
rect 17960 4428 18012 4480
rect 19708 4428 19760 4480
rect 20352 4428 20404 4480
rect 20812 4428 20864 4480
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 50294 4326 50346 4378
rect 50358 4326 50410 4378
rect 50422 4326 50474 4378
rect 50486 4326 50538 4378
rect 50550 4326 50602 4378
rect 3792 4088 3844 4140
rect 4160 4088 4212 4140
rect 6920 4224 6972 4276
rect 11796 4224 11848 4276
rect 5816 4131 5868 4140
rect 3976 3952 4028 4004
rect 4160 3952 4212 4004
rect 5080 4020 5132 4072
rect 5816 4097 5825 4131
rect 5825 4097 5859 4131
rect 5859 4097 5868 4131
rect 5816 4088 5868 4097
rect 8300 4156 8352 4208
rect 6828 4131 6880 4140
rect 6828 4097 6862 4131
rect 6862 4097 6880 4131
rect 9588 4156 9640 4208
rect 10876 4199 10928 4208
rect 10876 4165 10885 4199
rect 10885 4165 10919 4199
rect 10919 4165 10928 4199
rect 10876 4156 10928 4165
rect 6828 4088 6880 4097
rect 8484 4088 8536 4140
rect 9220 4088 9272 4140
rect 12072 4131 12124 4140
rect 6276 4020 6328 4072
rect 10140 4020 10192 4072
rect 12072 4097 12081 4131
rect 12081 4097 12115 4131
rect 12115 4097 12124 4131
rect 12072 4088 12124 4097
rect 12256 4131 12308 4140
rect 12256 4097 12265 4131
rect 12265 4097 12299 4131
rect 12299 4097 12308 4131
rect 12256 4088 12308 4097
rect 12440 4224 12492 4276
rect 20444 4267 20496 4276
rect 20444 4233 20453 4267
rect 20453 4233 20487 4267
rect 20487 4233 20496 4267
rect 20444 4224 20496 4233
rect 12164 4020 12216 4072
rect 9404 3952 9456 4004
rect 11796 3952 11848 4004
rect 12256 3952 12308 4004
rect 4620 3884 4672 3936
rect 5448 3884 5500 3936
rect 6920 3884 6972 3936
rect 9772 3927 9824 3936
rect 9772 3893 9781 3927
rect 9781 3893 9815 3927
rect 9815 3893 9824 3927
rect 9772 3884 9824 3893
rect 12900 4088 12952 4140
rect 13728 4088 13780 4140
rect 17224 4131 17276 4140
rect 17224 4097 17233 4131
rect 17233 4097 17267 4131
rect 17267 4097 17276 4131
rect 17224 4088 17276 4097
rect 18052 4088 18104 4140
rect 20720 4156 20772 4208
rect 21456 4156 21508 4208
rect 20628 4131 20680 4140
rect 20628 4097 20637 4131
rect 20637 4097 20671 4131
rect 20671 4097 20680 4131
rect 20628 4088 20680 4097
rect 21640 4088 21692 4140
rect 22100 4131 22152 4140
rect 22100 4097 22109 4131
rect 22109 4097 22143 4131
rect 22143 4097 22152 4131
rect 22100 4088 22152 4097
rect 20444 4020 20496 4072
rect 22008 4020 22060 4072
rect 15752 3952 15804 4004
rect 16672 3952 16724 4004
rect 17684 3952 17736 4004
rect 15936 3884 15988 3936
rect 16488 3884 16540 3936
rect 17316 3884 17368 3936
rect 19340 3927 19392 3936
rect 19340 3893 19349 3927
rect 19349 3893 19383 3927
rect 19383 3893 19392 3927
rect 19340 3884 19392 3893
rect 21456 3952 21508 4004
rect 22192 3952 22244 4004
rect 20536 3884 20588 3936
rect 21732 3884 21784 3936
rect 21916 3927 21968 3936
rect 21916 3893 21925 3927
rect 21925 3893 21959 3927
rect 21959 3893 21968 3927
rect 21916 3884 21968 3893
rect 22468 3884 22520 3936
rect 24032 3927 24084 3936
rect 24032 3893 24041 3927
rect 24041 3893 24075 3927
rect 24075 3893 24084 3927
rect 24032 3884 24084 3893
rect 24676 3927 24728 3936
rect 24676 3893 24685 3927
rect 24685 3893 24719 3927
rect 24719 3893 24728 3927
rect 24676 3884 24728 3893
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 65654 3782 65706 3834
rect 65718 3782 65770 3834
rect 65782 3782 65834 3834
rect 65846 3782 65898 3834
rect 65910 3782 65962 3834
rect 8484 3680 8536 3732
rect 8576 3680 8628 3732
rect 4252 3655 4304 3664
rect 4252 3621 4261 3655
rect 4261 3621 4295 3655
rect 4295 3621 4304 3655
rect 4252 3612 4304 3621
rect 5172 3612 5224 3664
rect 6092 3612 6144 3664
rect 4988 3544 5040 3596
rect 4160 3476 4212 3528
rect 5172 3476 5224 3528
rect 9772 3612 9824 3664
rect 12072 3680 12124 3732
rect 13544 3680 13596 3732
rect 15752 3680 15804 3732
rect 20260 3680 20312 3732
rect 20444 3680 20496 3732
rect 21824 3680 21876 3732
rect 15568 3612 15620 3664
rect 6920 3544 6972 3596
rect 4804 3383 4856 3392
rect 4804 3349 4813 3383
rect 4813 3349 4847 3383
rect 4847 3349 4856 3383
rect 4804 3340 4856 3349
rect 5448 3340 5500 3392
rect 6092 3408 6144 3460
rect 6460 3476 6512 3528
rect 7656 3476 7708 3528
rect 8116 3476 8168 3528
rect 8208 3519 8260 3528
rect 8208 3485 8217 3519
rect 8217 3485 8251 3519
rect 8251 3485 8260 3519
rect 8944 3519 8996 3528
rect 8208 3476 8260 3485
rect 8944 3485 8953 3519
rect 8953 3485 8987 3519
rect 8987 3485 8996 3519
rect 8944 3476 8996 3485
rect 9588 3544 9640 3596
rect 13268 3587 13320 3596
rect 13268 3553 13277 3587
rect 13277 3553 13311 3587
rect 13311 3553 13320 3587
rect 13268 3544 13320 3553
rect 10876 3476 10928 3528
rect 12256 3476 12308 3528
rect 14096 3544 14148 3596
rect 15292 3519 15344 3528
rect 6828 3408 6880 3460
rect 15292 3485 15301 3519
rect 15301 3485 15335 3519
rect 15335 3485 15344 3519
rect 15292 3476 15344 3485
rect 15476 3476 15528 3528
rect 15844 3476 15896 3528
rect 7288 3340 7340 3392
rect 7564 3383 7616 3392
rect 7564 3349 7573 3383
rect 7573 3349 7607 3383
rect 7607 3349 7616 3383
rect 7564 3340 7616 3349
rect 8760 3340 8812 3392
rect 9680 3383 9732 3392
rect 9680 3349 9689 3383
rect 9689 3349 9723 3383
rect 9723 3349 9732 3383
rect 9680 3340 9732 3349
rect 11704 3383 11756 3392
rect 11704 3349 11713 3383
rect 11713 3349 11747 3383
rect 11747 3349 11756 3383
rect 11704 3340 11756 3349
rect 11796 3340 11848 3392
rect 15200 3408 15252 3460
rect 16212 3476 16264 3528
rect 18696 3612 18748 3664
rect 20628 3612 20680 3664
rect 51448 3612 51500 3664
rect 21824 3544 21876 3596
rect 18052 3476 18104 3528
rect 18972 3476 19024 3528
rect 20904 3476 20956 3528
rect 21272 3519 21324 3528
rect 21272 3485 21281 3519
rect 21281 3485 21315 3519
rect 21315 3485 21324 3519
rect 21272 3476 21324 3485
rect 21364 3519 21416 3528
rect 21364 3485 21373 3519
rect 21373 3485 21407 3519
rect 21407 3485 21416 3519
rect 21732 3519 21784 3528
rect 21364 3476 21416 3485
rect 21732 3485 21741 3519
rect 21741 3485 21775 3519
rect 21775 3485 21784 3519
rect 21732 3476 21784 3485
rect 22744 3476 22796 3528
rect 23572 3476 23624 3528
rect 26056 3476 26108 3528
rect 27436 3476 27488 3528
rect 27712 3519 27764 3528
rect 27712 3485 27721 3519
rect 27721 3485 27755 3519
rect 27755 3485 27764 3519
rect 27712 3476 27764 3485
rect 28264 3476 28316 3528
rect 29368 3476 29420 3528
rect 30196 3476 30248 3528
rect 31300 3476 31352 3528
rect 32128 3476 32180 3528
rect 32956 3476 33008 3528
rect 39856 3476 39908 3528
rect 40132 3476 40184 3528
rect 40960 3476 41012 3528
rect 41788 3476 41840 3528
rect 42616 3476 42668 3528
rect 43720 3476 43772 3528
rect 45100 3476 45152 3528
rect 45652 3476 45704 3528
rect 46204 3476 46256 3528
rect 47584 3476 47636 3528
rect 47860 3476 47912 3528
rect 49516 3476 49568 3528
rect 50620 3476 50672 3528
rect 51172 3476 51224 3528
rect 52828 3476 52880 3528
rect 53380 3476 53432 3528
rect 55312 3476 55364 3528
rect 55588 3476 55640 3528
rect 56416 3476 56468 3528
rect 57244 3476 57296 3528
rect 57520 3476 57572 3528
rect 16304 3408 16356 3460
rect 20628 3408 20680 3460
rect 24032 3408 24084 3460
rect 16764 3340 16816 3392
rect 18972 3340 19024 3392
rect 21364 3340 21416 3392
rect 24676 3340 24728 3392
rect 24952 3340 25004 3392
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 50294 3238 50346 3290
rect 50358 3238 50410 3290
rect 50422 3238 50474 3290
rect 50486 3238 50538 3290
rect 50550 3238 50602 3290
rect 3884 3136 3936 3188
rect 4068 3136 4120 3188
rect 4068 3043 4120 3052
rect 4068 3009 4077 3043
rect 4077 3009 4111 3043
rect 4111 3009 4120 3043
rect 4068 3000 4120 3009
rect 6828 3136 6880 3188
rect 4528 3068 4580 3120
rect 4620 3068 4672 3120
rect 5172 3043 5224 3052
rect 5172 3009 5181 3043
rect 5181 3009 5215 3043
rect 5215 3009 5224 3043
rect 5172 3000 5224 3009
rect 5448 3043 5500 3052
rect 5448 3009 5457 3043
rect 5457 3009 5491 3043
rect 5491 3009 5500 3043
rect 5908 3068 5960 3120
rect 5448 3000 5500 3009
rect 6736 3043 6788 3052
rect 6736 3009 6745 3043
rect 6745 3009 6779 3043
rect 6779 3009 6788 3043
rect 6736 3000 6788 3009
rect 5908 2932 5960 2984
rect 13728 3136 13780 3188
rect 7196 3043 7248 3052
rect 7196 3009 7205 3043
rect 7205 3009 7239 3043
rect 7239 3009 7248 3043
rect 7196 3000 7248 3009
rect 7288 3000 7340 3052
rect 7748 3000 7800 3052
rect 8576 3000 8628 3052
rect 9404 3068 9456 3120
rect 9772 3068 9824 3120
rect 11888 3068 11940 3120
rect 12164 3000 12216 3052
rect 13544 3043 13596 3052
rect 13544 3009 13575 3043
rect 13575 3009 13596 3043
rect 13544 3000 13596 3009
rect 13636 3000 13688 3052
rect 14096 3136 14148 3188
rect 15108 3136 15160 3188
rect 16120 3136 16172 3188
rect 21272 3136 21324 3188
rect 16304 3068 16356 3120
rect 15476 3000 15528 3052
rect 16856 3043 16908 3052
rect 16856 3009 16865 3043
rect 16865 3009 16899 3043
rect 16899 3009 16908 3043
rect 16856 3000 16908 3009
rect 20812 3068 20864 3120
rect 17224 3000 17276 3052
rect 6000 2796 6052 2848
rect 18052 2932 18104 2984
rect 18420 2975 18472 2984
rect 18420 2941 18429 2975
rect 18429 2941 18463 2975
rect 18463 2941 18472 2975
rect 18420 2932 18472 2941
rect 20720 3000 20772 3052
rect 16120 2864 16172 2916
rect 18144 2864 18196 2916
rect 19432 2864 19484 2916
rect 20904 2864 20956 2916
rect 8576 2839 8628 2848
rect 8576 2805 8585 2839
rect 8585 2805 8619 2839
rect 8619 2805 8628 2839
rect 8576 2796 8628 2805
rect 10876 2796 10928 2848
rect 12164 2839 12216 2848
rect 12164 2805 12173 2839
rect 12173 2805 12207 2839
rect 12207 2805 12216 2839
rect 12164 2796 12216 2805
rect 12900 2796 12952 2848
rect 14372 2796 14424 2848
rect 15292 2796 15344 2848
rect 17040 2796 17092 2848
rect 17684 2796 17736 2848
rect 22192 2932 22244 2984
rect 25228 2932 25280 2984
rect 37924 2932 37976 2984
rect 39580 2932 39632 2984
rect 43444 2932 43496 2984
rect 47308 2932 47360 2984
rect 49240 2932 49292 2984
rect 55036 2932 55088 2984
rect 38476 2864 38528 2916
rect 40408 2864 40460 2916
rect 42340 2864 42392 2916
rect 44272 2864 44324 2916
rect 45376 2864 45428 2916
rect 48136 2864 48188 2916
rect 50068 2864 50120 2916
rect 52552 2864 52604 2916
rect 53932 2864 53984 2916
rect 57612 2864 57664 2916
rect 21272 2796 21324 2848
rect 21640 2796 21692 2848
rect 21824 2839 21876 2848
rect 21824 2805 21833 2839
rect 21833 2805 21867 2839
rect 21867 2805 21876 2839
rect 21824 2796 21876 2805
rect 23020 2796 23072 2848
rect 23296 2796 23348 2848
rect 24124 2796 24176 2848
rect 24676 2796 24728 2848
rect 25780 2839 25832 2848
rect 25780 2805 25789 2839
rect 25789 2805 25823 2839
rect 25823 2805 25832 2839
rect 25780 2796 25832 2805
rect 26332 2796 26384 2848
rect 26424 2796 26476 2848
rect 27988 2796 28040 2848
rect 28540 2796 28592 2848
rect 29092 2796 29144 2848
rect 29920 2796 29972 2848
rect 30472 2796 30524 2848
rect 31024 2796 31076 2848
rect 31852 2796 31904 2848
rect 32680 2796 32732 2848
rect 33232 2796 33284 2848
rect 33784 2839 33836 2848
rect 33784 2805 33793 2839
rect 33793 2805 33827 2839
rect 33827 2805 33836 2839
rect 33784 2796 33836 2805
rect 34336 2796 34388 2848
rect 34796 2796 34848 2848
rect 35440 2796 35492 2848
rect 36268 2796 36320 2848
rect 36820 2796 36872 2848
rect 37372 2796 37424 2848
rect 39028 2796 39080 2848
rect 41512 2796 41564 2848
rect 42892 2796 42944 2848
rect 44824 2796 44876 2848
rect 46756 2796 46808 2848
rect 48688 2796 48740 2848
rect 50712 2796 50764 2848
rect 52000 2796 52052 2848
rect 53104 2796 53156 2848
rect 54484 2796 54536 2848
rect 55864 2796 55916 2848
rect 56968 2796 57020 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 65654 2694 65706 2746
rect 65718 2694 65770 2746
rect 65782 2694 65834 2746
rect 65846 2694 65898 2746
rect 65910 2694 65962 2746
rect 4712 2592 4764 2644
rect 5816 2592 5868 2644
rect 4896 2524 4948 2576
rect 7196 2592 7248 2644
rect 13452 2592 13504 2644
rect 15292 2592 15344 2644
rect 17224 2592 17276 2644
rect 3884 2431 3936 2440
rect 3884 2397 3893 2431
rect 3893 2397 3927 2431
rect 3927 2397 3936 2431
rect 3884 2388 3936 2397
rect 4712 2431 4764 2440
rect 4712 2397 4721 2431
rect 4721 2397 4755 2431
rect 4755 2397 4764 2431
rect 4712 2388 4764 2397
rect 5172 2431 5224 2440
rect 5172 2397 5181 2431
rect 5181 2397 5215 2431
rect 5215 2397 5224 2431
rect 5172 2388 5224 2397
rect 5264 2388 5316 2440
rect 5448 2431 5500 2440
rect 5448 2397 5457 2431
rect 5457 2397 5491 2431
rect 5491 2397 5500 2431
rect 5448 2388 5500 2397
rect 6552 2431 6604 2440
rect 6552 2397 6561 2431
rect 6561 2397 6595 2431
rect 6595 2397 6604 2431
rect 6552 2388 6604 2397
rect 9956 2388 10008 2440
rect 11336 2456 11388 2508
rect 11704 2388 11756 2440
rect 15384 2524 15436 2576
rect 15108 2456 15160 2508
rect 10876 2320 10928 2372
rect 12808 2388 12860 2440
rect 14372 2431 14424 2440
rect 14372 2397 14381 2431
rect 14381 2397 14415 2431
rect 14415 2397 14424 2431
rect 14372 2388 14424 2397
rect 6552 2252 6604 2304
rect 10048 2295 10100 2304
rect 10048 2261 10057 2295
rect 10057 2261 10091 2295
rect 10091 2261 10100 2295
rect 10048 2252 10100 2261
rect 10784 2295 10836 2304
rect 10784 2261 10793 2295
rect 10793 2261 10827 2295
rect 10827 2261 10836 2295
rect 10784 2252 10836 2261
rect 15292 2388 15344 2440
rect 16580 2456 16632 2508
rect 19064 2592 19116 2644
rect 20904 2592 20956 2644
rect 22284 2592 22336 2644
rect 20260 2524 20312 2576
rect 18420 2499 18472 2508
rect 18420 2465 18429 2499
rect 18429 2465 18463 2499
rect 18463 2465 18472 2499
rect 18420 2456 18472 2465
rect 23848 2524 23900 2576
rect 31576 2524 31628 2576
rect 33508 2524 33560 2576
rect 39304 2524 39356 2576
rect 43168 2524 43220 2576
rect 47032 2524 47084 2576
rect 50896 2524 50948 2576
rect 54760 2524 54812 2576
rect 56692 2524 56744 2576
rect 17684 2388 17736 2440
rect 20168 2388 20220 2440
rect 20444 2431 20496 2440
rect 20444 2397 20453 2431
rect 20453 2397 20487 2431
rect 20487 2397 20496 2431
rect 20444 2388 20496 2397
rect 22652 2456 22704 2508
rect 27160 2456 27212 2508
rect 37096 2456 37148 2508
rect 38200 2456 38252 2508
rect 40684 2456 40736 2508
rect 43996 2456 44048 2508
rect 45928 2456 45980 2508
rect 48412 2456 48464 2508
rect 51724 2456 51776 2508
rect 53656 2456 53708 2508
rect 57428 2456 57480 2508
rect 22836 2388 22888 2440
rect 24400 2388 24452 2440
rect 26424 2388 26476 2440
rect 26976 2431 27028 2440
rect 26976 2397 26985 2431
rect 26985 2397 27019 2431
rect 27019 2397 27028 2431
rect 26976 2388 27028 2397
rect 28816 2388 28868 2440
rect 29644 2388 29696 2440
rect 30748 2388 30800 2440
rect 32404 2388 32456 2440
rect 34060 2388 34112 2440
rect 34612 2388 34664 2440
rect 35164 2388 35216 2440
rect 35716 2388 35768 2440
rect 35992 2388 36044 2440
rect 36544 2388 36596 2440
rect 37648 2388 37700 2440
rect 38752 2388 38804 2440
rect 41236 2388 41288 2440
rect 17592 2320 17644 2372
rect 18236 2320 18288 2372
rect 19248 2320 19300 2372
rect 18420 2252 18472 2304
rect 20076 2252 20128 2304
rect 42064 2320 42116 2372
rect 44548 2320 44600 2372
rect 46480 2388 46532 2440
rect 48964 2388 49016 2440
rect 49792 2320 49844 2372
rect 52276 2388 52328 2440
rect 54208 2320 54260 2372
rect 56140 2388 56192 2440
rect 25504 2252 25556 2304
rect 26608 2252 26660 2304
rect 26884 2252 26936 2304
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 50294 2150 50346 2202
rect 50358 2150 50410 2202
rect 50422 2150 50474 2202
rect 50486 2150 50538 2202
rect 50550 2150 50602 2202
rect 10784 2048 10836 2100
rect 14556 2048 14608 2100
rect 4712 1980 4764 2032
rect 14096 1980 14148 2032
rect 6552 1912 6604 1964
rect 12808 1912 12860 1964
rect 8208 1844 8260 1896
rect 16396 1844 16448 1896
rect 10048 1776 10100 1828
rect 14188 1776 14240 1828
rect 15292 1504 15344 1556
rect 16212 1504 16264 1556
rect 12164 1436 12216 1488
rect 14832 1436 14884 1488
rect 20260 1368 20312 1420
rect 19800 1300 19852 1352
rect 19984 1300 20036 1352
rect 20536 1300 20588 1352
<< metal2 >>
rect 2962 59200 3018 60000
rect 3514 59200 3570 60000
rect 4066 59200 4122 60000
rect 4618 59200 4674 60000
rect 5170 59200 5226 60000
rect 5722 59200 5778 60000
rect 6274 59200 6330 60000
rect 6826 59200 6882 60000
rect 7378 59200 7434 60000
rect 7930 59200 7986 60000
rect 8482 59200 8538 60000
rect 9034 59200 9090 60000
rect 9586 59200 9642 60000
rect 10138 59200 10194 60000
rect 10690 59200 10746 60000
rect 11242 59200 11298 60000
rect 11794 59200 11850 60000
rect 12346 59200 12402 60000
rect 12898 59200 12954 60000
rect 13450 59200 13506 60000
rect 14002 59200 14058 60000
rect 14554 59200 14610 60000
rect 15106 59200 15162 60000
rect 15658 59200 15714 60000
rect 16210 59200 16266 60000
rect 16762 59200 16818 60000
rect 17314 59200 17370 60000
rect 17866 59200 17922 60000
rect 18418 59200 18474 60000
rect 18970 59200 19026 60000
rect 19522 59200 19578 60000
rect 20074 59200 20130 60000
rect 20626 59200 20682 60000
rect 21178 59200 21234 60000
rect 21730 59200 21786 60000
rect 22282 59200 22338 60000
rect 22834 59200 22890 60000
rect 23386 59200 23442 60000
rect 23938 59200 23994 60000
rect 24490 59200 24546 60000
rect 25042 59200 25098 60000
rect 25594 59200 25650 60000
rect 26146 59200 26202 60000
rect 26698 59200 26754 60000
rect 27250 59200 27306 60000
rect 27802 59200 27858 60000
rect 28354 59200 28410 60000
rect 28906 59200 28962 60000
rect 29458 59200 29514 60000
rect 30010 59200 30066 60000
rect 30562 59200 30618 60000
rect 31114 59200 31170 60000
rect 31666 59200 31722 60000
rect 32218 59200 32274 60000
rect 32770 59200 32826 60000
rect 33322 59200 33378 60000
rect 33874 59200 33930 60000
rect 34426 59200 34482 60000
rect 34978 59200 35034 60000
rect 35530 59200 35586 60000
rect 36082 59200 36138 60000
rect 36634 59200 36690 60000
rect 37186 59200 37242 60000
rect 37738 59200 37794 60000
rect 38290 59200 38346 60000
rect 38842 59200 38898 60000
rect 39394 59200 39450 60000
rect 39946 59200 40002 60000
rect 40498 59200 40554 60000
rect 41050 59200 41106 60000
rect 41602 59200 41658 60000
rect 42154 59200 42210 60000
rect 42706 59200 42762 60000
rect 43258 59200 43314 60000
rect 43810 59200 43866 60000
rect 44362 59200 44418 60000
rect 44914 59200 44970 60000
rect 45466 59200 45522 60000
rect 46018 59200 46074 60000
rect 46570 59200 46626 60000
rect 47122 59200 47178 60000
rect 47674 59200 47730 60000
rect 48226 59200 48282 60000
rect 48778 59200 48834 60000
rect 49330 59200 49386 60000
rect 49882 59200 49938 60000
rect 50434 59200 50490 60000
rect 50986 59200 51042 60000
rect 51538 59200 51594 60000
rect 52090 59200 52146 60000
rect 52196 59214 52408 59242
rect 3528 57458 3556 59200
rect 4080 57882 4108 59200
rect 4080 57854 4200 57882
rect 4172 57458 4200 57854
rect 5184 57458 5212 59200
rect 5736 57458 5764 59200
rect 6840 57458 6868 59200
rect 7392 57458 7420 59200
rect 8496 57458 8524 59200
rect 9048 57458 9076 59200
rect 10152 57458 10180 59200
rect 10704 57458 10732 59200
rect 11808 57458 11836 59200
rect 3516 57452 3568 57458
rect 3516 57394 3568 57400
rect 4160 57452 4212 57458
rect 4160 57394 4212 57400
rect 5172 57452 5224 57458
rect 5172 57394 5224 57400
rect 5724 57452 5776 57458
rect 5724 57394 5776 57400
rect 6828 57452 6880 57458
rect 6828 57394 6880 57400
rect 7380 57452 7432 57458
rect 7380 57394 7432 57400
rect 8484 57452 8536 57458
rect 8484 57394 8536 57400
rect 9036 57452 9088 57458
rect 9036 57394 9088 57400
rect 10140 57452 10192 57458
rect 10140 57394 10192 57400
rect 10692 57452 10744 57458
rect 10692 57394 10744 57400
rect 11796 57452 11848 57458
rect 12360 57440 12388 59200
rect 13464 57458 13492 59200
rect 14016 57458 14044 59200
rect 15120 57458 15148 59200
rect 15672 57458 15700 59200
rect 16776 57458 16804 59200
rect 17328 57458 17356 59200
rect 18432 57458 18460 59200
rect 18984 57458 19012 59200
rect 19574 57692 19882 57701
rect 19574 57690 19580 57692
rect 19636 57690 19660 57692
rect 19716 57690 19740 57692
rect 19796 57690 19820 57692
rect 19876 57690 19882 57692
rect 19636 57638 19638 57690
rect 19818 57638 19820 57690
rect 19574 57636 19580 57638
rect 19636 57636 19660 57638
rect 19716 57636 19740 57638
rect 19796 57636 19820 57638
rect 19876 57636 19882 57638
rect 19574 57627 19882 57636
rect 20088 57458 20116 59200
rect 20640 57882 20668 59200
rect 20640 57854 20760 57882
rect 20732 57458 20760 57854
rect 12440 57452 12492 57458
rect 12360 57412 12440 57440
rect 11796 57394 11848 57400
rect 12440 57394 12492 57400
rect 13452 57452 13504 57458
rect 13452 57394 13504 57400
rect 14004 57452 14056 57458
rect 14004 57394 14056 57400
rect 15108 57452 15160 57458
rect 15108 57394 15160 57400
rect 15660 57452 15712 57458
rect 15660 57394 15712 57400
rect 16764 57452 16816 57458
rect 16764 57394 16816 57400
rect 17316 57452 17368 57458
rect 17316 57394 17368 57400
rect 18420 57452 18472 57458
rect 18420 57394 18472 57400
rect 18972 57452 19024 57458
rect 18972 57394 19024 57400
rect 20076 57452 20128 57458
rect 20076 57394 20128 57400
rect 20720 57452 20772 57458
rect 20720 57394 20772 57400
rect 4214 57148 4522 57157
rect 4214 57146 4220 57148
rect 4276 57146 4300 57148
rect 4356 57146 4380 57148
rect 4436 57146 4460 57148
rect 4516 57146 4522 57148
rect 4276 57094 4278 57146
rect 4458 57094 4460 57146
rect 4214 57092 4220 57094
rect 4276 57092 4300 57094
rect 4356 57092 4380 57094
rect 4436 57092 4460 57094
rect 4516 57092 4522 57094
rect 4214 57083 4522 57092
rect 21744 57050 21772 59200
rect 22296 57458 22324 59200
rect 23400 57882 23428 59200
rect 23400 57854 23520 57882
rect 23492 57458 23520 57854
rect 23952 57458 23980 59200
rect 25056 57458 25084 59200
rect 25608 57458 25636 59200
rect 22284 57452 22336 57458
rect 22284 57394 22336 57400
rect 23480 57452 23532 57458
rect 23480 57394 23532 57400
rect 23940 57452 23992 57458
rect 23940 57394 23992 57400
rect 25044 57452 25096 57458
rect 25044 57394 25096 57400
rect 25596 57452 25648 57458
rect 25596 57394 25648 57400
rect 26712 57050 26740 59200
rect 27264 57458 27292 59200
rect 28368 57458 28396 59200
rect 28920 57458 28948 59200
rect 30024 57458 30052 59200
rect 30576 57458 30604 59200
rect 31680 57458 31708 59200
rect 32232 57458 32260 59200
rect 33336 57458 33364 59200
rect 33888 57458 33916 59200
rect 34992 57458 35020 59200
rect 35544 57458 35572 59200
rect 36648 57458 36676 59200
rect 27252 57452 27304 57458
rect 27252 57394 27304 57400
rect 28356 57452 28408 57458
rect 28356 57394 28408 57400
rect 28908 57452 28960 57458
rect 28908 57394 28960 57400
rect 30012 57452 30064 57458
rect 30012 57394 30064 57400
rect 30564 57452 30616 57458
rect 30564 57394 30616 57400
rect 31668 57452 31720 57458
rect 31668 57394 31720 57400
rect 32220 57452 32272 57458
rect 32220 57394 32272 57400
rect 33324 57452 33376 57458
rect 33324 57394 33376 57400
rect 33876 57452 33928 57458
rect 33876 57394 33928 57400
rect 34980 57452 35032 57458
rect 34980 57394 35032 57400
rect 35532 57452 35584 57458
rect 35532 57394 35584 57400
rect 36636 57452 36688 57458
rect 36636 57394 36688 57400
rect 37200 57338 37228 59200
rect 38304 57458 38332 59200
rect 38292 57452 38344 57458
rect 38292 57394 38344 57400
rect 37200 57322 37320 57338
rect 37200 57316 37332 57322
rect 37200 57310 37280 57316
rect 37280 57258 37332 57264
rect 34934 57148 35242 57157
rect 34934 57146 34940 57148
rect 34996 57146 35020 57148
rect 35076 57146 35100 57148
rect 35156 57146 35180 57148
rect 35236 57146 35242 57148
rect 34996 57094 34998 57146
rect 35178 57094 35180 57146
rect 34934 57092 34940 57094
rect 34996 57092 35020 57094
rect 35076 57092 35100 57094
rect 35156 57092 35180 57094
rect 35236 57092 35242 57094
rect 34934 57083 35242 57092
rect 38856 57050 38884 59200
rect 39960 57440 39988 59200
rect 40512 57458 40540 59200
rect 41616 57458 41644 59200
rect 42168 57458 42196 59200
rect 43272 57458 43300 59200
rect 43824 57458 43852 59200
rect 44928 57458 44956 59200
rect 40040 57452 40092 57458
rect 39960 57412 40040 57440
rect 40040 57394 40092 57400
rect 40500 57452 40552 57458
rect 40500 57394 40552 57400
rect 41604 57452 41656 57458
rect 41604 57394 41656 57400
rect 42156 57452 42208 57458
rect 42156 57394 42208 57400
rect 43260 57452 43312 57458
rect 43260 57394 43312 57400
rect 43812 57452 43864 57458
rect 43812 57394 43864 57400
rect 44916 57452 44968 57458
rect 44916 57394 44968 57400
rect 45480 57390 45508 59200
rect 46584 57458 46612 59200
rect 47136 57458 47164 59200
rect 46572 57452 46624 57458
rect 46572 57394 46624 57400
rect 47124 57452 47176 57458
rect 48240 57440 48268 59200
rect 48792 57458 48820 59200
rect 49896 57458 49924 59200
rect 50448 57882 50476 59200
rect 50448 57854 50660 57882
rect 50294 57692 50602 57701
rect 50294 57690 50300 57692
rect 50356 57690 50380 57692
rect 50436 57690 50460 57692
rect 50516 57690 50540 57692
rect 50596 57690 50602 57692
rect 50356 57638 50358 57690
rect 50538 57638 50540 57690
rect 50294 57636 50300 57638
rect 50356 57636 50380 57638
rect 50436 57636 50460 57638
rect 50516 57636 50540 57638
rect 50596 57636 50602 57638
rect 50294 57627 50602 57636
rect 50632 57458 50660 57854
rect 51552 57458 51580 59200
rect 52104 59106 52132 59200
rect 52196 59106 52224 59214
rect 52104 59078 52224 59106
rect 48320 57452 48372 57458
rect 48240 57412 48320 57440
rect 47124 57394 47176 57400
rect 48320 57394 48372 57400
rect 48780 57452 48832 57458
rect 48780 57394 48832 57400
rect 49884 57452 49936 57458
rect 49884 57394 49936 57400
rect 50620 57452 50672 57458
rect 50620 57394 50672 57400
rect 51540 57452 51592 57458
rect 52380 57440 52408 59214
rect 52642 59200 52698 60000
rect 53194 59200 53250 60000
rect 53746 59200 53802 60000
rect 54298 59200 54354 60000
rect 54850 59200 54906 60000
rect 55402 59200 55458 60000
rect 55954 59200 56010 60000
rect 56506 59200 56562 60000
rect 57058 59200 57114 60000
rect 57610 59200 57666 60000
rect 58162 59200 58218 60000
rect 58714 59200 58770 60000
rect 59266 59200 59322 60000
rect 59818 59200 59874 60000
rect 60370 59200 60426 60000
rect 60476 59214 60688 59242
rect 53208 57458 53236 59200
rect 52460 57452 52512 57458
rect 52380 57412 52460 57440
rect 51540 57394 51592 57400
rect 52460 57394 52512 57400
rect 53196 57452 53248 57458
rect 53760 57440 53788 59200
rect 54864 57458 54892 59200
rect 55416 57458 55444 59200
rect 56520 57882 56548 59200
rect 56520 57854 56640 57882
rect 56612 57458 56640 57854
rect 57072 57458 57100 59200
rect 58176 57458 58204 59200
rect 58728 57458 58756 59200
rect 59832 57458 59860 59200
rect 60384 59106 60412 59200
rect 60476 59106 60504 59214
rect 60384 59078 60504 59106
rect 60660 57474 60688 59214
rect 60922 59200 60978 60000
rect 61474 59200 61530 60000
rect 62026 59200 62082 60000
rect 62578 59200 62634 60000
rect 63130 59200 63186 60000
rect 63682 59200 63738 60000
rect 64234 59200 64290 60000
rect 64786 59200 64842 60000
rect 65338 59200 65394 60000
rect 65890 59200 65946 60000
rect 66442 59200 66498 60000
rect 66994 59200 67050 60000
rect 60660 57458 60780 57474
rect 61488 57458 61516 59200
rect 62040 57882 62068 59200
rect 62040 57854 62160 57882
rect 53840 57452 53892 57458
rect 53760 57412 53840 57440
rect 53196 57394 53248 57400
rect 53840 57394 53892 57400
rect 54852 57452 54904 57458
rect 54852 57394 54904 57400
rect 55404 57452 55456 57458
rect 55404 57394 55456 57400
rect 56600 57452 56652 57458
rect 56600 57394 56652 57400
rect 57060 57452 57112 57458
rect 57060 57394 57112 57400
rect 58164 57452 58216 57458
rect 58164 57394 58216 57400
rect 58716 57452 58768 57458
rect 58716 57394 58768 57400
rect 59820 57452 59872 57458
rect 60660 57452 60792 57458
rect 60660 57446 60740 57452
rect 59820 57394 59872 57400
rect 60740 57394 60792 57400
rect 61476 57452 61528 57458
rect 61476 57394 61528 57400
rect 45468 57384 45520 57390
rect 45468 57326 45520 57332
rect 62132 57050 62160 57854
rect 63144 57458 63172 59200
rect 63696 57458 63724 59200
rect 63132 57452 63184 57458
rect 63132 57394 63184 57400
rect 63684 57452 63736 57458
rect 63684 57394 63736 57400
rect 64800 57390 64828 59200
rect 65352 57458 65380 59200
rect 67008 57458 67036 59200
rect 65340 57452 65392 57458
rect 65340 57394 65392 57400
rect 66996 57452 67048 57458
rect 66996 57394 67048 57400
rect 64788 57384 64840 57390
rect 64788 57326 64840 57332
rect 65654 57148 65962 57157
rect 65654 57146 65660 57148
rect 65716 57146 65740 57148
rect 65796 57146 65820 57148
rect 65876 57146 65900 57148
rect 65956 57146 65962 57148
rect 65716 57094 65718 57146
rect 65898 57094 65900 57146
rect 65654 57092 65660 57094
rect 65716 57092 65740 57094
rect 65796 57092 65820 57094
rect 65876 57092 65900 57094
rect 65956 57092 65962 57094
rect 65654 57083 65962 57092
rect 21732 57044 21784 57050
rect 21732 56986 21784 56992
rect 26700 57044 26752 57050
rect 26700 56986 26752 56992
rect 38844 57044 38896 57050
rect 38844 56986 38896 56992
rect 62120 57044 62172 57050
rect 62120 56986 62172 56992
rect 19574 56604 19882 56613
rect 19574 56602 19580 56604
rect 19636 56602 19660 56604
rect 19716 56602 19740 56604
rect 19796 56602 19820 56604
rect 19876 56602 19882 56604
rect 19636 56550 19638 56602
rect 19818 56550 19820 56602
rect 19574 56548 19580 56550
rect 19636 56548 19660 56550
rect 19716 56548 19740 56550
rect 19796 56548 19820 56550
rect 19876 56548 19882 56550
rect 19574 56539 19882 56548
rect 50294 56604 50602 56613
rect 50294 56602 50300 56604
rect 50356 56602 50380 56604
rect 50436 56602 50460 56604
rect 50516 56602 50540 56604
rect 50596 56602 50602 56604
rect 50356 56550 50358 56602
rect 50538 56550 50540 56602
rect 50294 56548 50300 56550
rect 50356 56548 50380 56550
rect 50436 56548 50460 56550
rect 50516 56548 50540 56550
rect 50596 56548 50602 56550
rect 50294 56539 50602 56548
rect 4214 56060 4522 56069
rect 4214 56058 4220 56060
rect 4276 56058 4300 56060
rect 4356 56058 4380 56060
rect 4436 56058 4460 56060
rect 4516 56058 4522 56060
rect 4276 56006 4278 56058
rect 4458 56006 4460 56058
rect 4214 56004 4220 56006
rect 4276 56004 4300 56006
rect 4356 56004 4380 56006
rect 4436 56004 4460 56006
rect 4516 56004 4522 56006
rect 4214 55995 4522 56004
rect 34934 56060 35242 56069
rect 34934 56058 34940 56060
rect 34996 56058 35020 56060
rect 35076 56058 35100 56060
rect 35156 56058 35180 56060
rect 35236 56058 35242 56060
rect 34996 56006 34998 56058
rect 35178 56006 35180 56058
rect 34934 56004 34940 56006
rect 34996 56004 35020 56006
rect 35076 56004 35100 56006
rect 35156 56004 35180 56006
rect 35236 56004 35242 56006
rect 34934 55995 35242 56004
rect 65654 56060 65962 56069
rect 65654 56058 65660 56060
rect 65716 56058 65740 56060
rect 65796 56058 65820 56060
rect 65876 56058 65900 56060
rect 65956 56058 65962 56060
rect 65716 56006 65718 56058
rect 65898 56006 65900 56058
rect 65654 56004 65660 56006
rect 65716 56004 65740 56006
rect 65796 56004 65820 56006
rect 65876 56004 65900 56006
rect 65956 56004 65962 56006
rect 65654 55995 65962 56004
rect 19574 55516 19882 55525
rect 19574 55514 19580 55516
rect 19636 55514 19660 55516
rect 19716 55514 19740 55516
rect 19796 55514 19820 55516
rect 19876 55514 19882 55516
rect 19636 55462 19638 55514
rect 19818 55462 19820 55514
rect 19574 55460 19580 55462
rect 19636 55460 19660 55462
rect 19716 55460 19740 55462
rect 19796 55460 19820 55462
rect 19876 55460 19882 55462
rect 19574 55451 19882 55460
rect 50294 55516 50602 55525
rect 50294 55514 50300 55516
rect 50356 55514 50380 55516
rect 50436 55514 50460 55516
rect 50516 55514 50540 55516
rect 50596 55514 50602 55516
rect 50356 55462 50358 55514
rect 50538 55462 50540 55514
rect 50294 55460 50300 55462
rect 50356 55460 50380 55462
rect 50436 55460 50460 55462
rect 50516 55460 50540 55462
rect 50596 55460 50602 55462
rect 50294 55451 50602 55460
rect 4214 54972 4522 54981
rect 4214 54970 4220 54972
rect 4276 54970 4300 54972
rect 4356 54970 4380 54972
rect 4436 54970 4460 54972
rect 4516 54970 4522 54972
rect 4276 54918 4278 54970
rect 4458 54918 4460 54970
rect 4214 54916 4220 54918
rect 4276 54916 4300 54918
rect 4356 54916 4380 54918
rect 4436 54916 4460 54918
rect 4516 54916 4522 54918
rect 4214 54907 4522 54916
rect 34934 54972 35242 54981
rect 34934 54970 34940 54972
rect 34996 54970 35020 54972
rect 35076 54970 35100 54972
rect 35156 54970 35180 54972
rect 35236 54970 35242 54972
rect 34996 54918 34998 54970
rect 35178 54918 35180 54970
rect 34934 54916 34940 54918
rect 34996 54916 35020 54918
rect 35076 54916 35100 54918
rect 35156 54916 35180 54918
rect 35236 54916 35242 54918
rect 34934 54907 35242 54916
rect 65654 54972 65962 54981
rect 65654 54970 65660 54972
rect 65716 54970 65740 54972
rect 65796 54970 65820 54972
rect 65876 54970 65900 54972
rect 65956 54970 65962 54972
rect 65716 54918 65718 54970
rect 65898 54918 65900 54970
rect 65654 54916 65660 54918
rect 65716 54916 65740 54918
rect 65796 54916 65820 54918
rect 65876 54916 65900 54918
rect 65956 54916 65962 54918
rect 65654 54907 65962 54916
rect 19574 54428 19882 54437
rect 19574 54426 19580 54428
rect 19636 54426 19660 54428
rect 19716 54426 19740 54428
rect 19796 54426 19820 54428
rect 19876 54426 19882 54428
rect 19636 54374 19638 54426
rect 19818 54374 19820 54426
rect 19574 54372 19580 54374
rect 19636 54372 19660 54374
rect 19716 54372 19740 54374
rect 19796 54372 19820 54374
rect 19876 54372 19882 54374
rect 19574 54363 19882 54372
rect 50294 54428 50602 54437
rect 50294 54426 50300 54428
rect 50356 54426 50380 54428
rect 50436 54426 50460 54428
rect 50516 54426 50540 54428
rect 50596 54426 50602 54428
rect 50356 54374 50358 54426
rect 50538 54374 50540 54426
rect 50294 54372 50300 54374
rect 50356 54372 50380 54374
rect 50436 54372 50460 54374
rect 50516 54372 50540 54374
rect 50596 54372 50602 54374
rect 50294 54363 50602 54372
rect 4214 53884 4522 53893
rect 4214 53882 4220 53884
rect 4276 53882 4300 53884
rect 4356 53882 4380 53884
rect 4436 53882 4460 53884
rect 4516 53882 4522 53884
rect 4276 53830 4278 53882
rect 4458 53830 4460 53882
rect 4214 53828 4220 53830
rect 4276 53828 4300 53830
rect 4356 53828 4380 53830
rect 4436 53828 4460 53830
rect 4516 53828 4522 53830
rect 4214 53819 4522 53828
rect 34934 53884 35242 53893
rect 34934 53882 34940 53884
rect 34996 53882 35020 53884
rect 35076 53882 35100 53884
rect 35156 53882 35180 53884
rect 35236 53882 35242 53884
rect 34996 53830 34998 53882
rect 35178 53830 35180 53882
rect 34934 53828 34940 53830
rect 34996 53828 35020 53830
rect 35076 53828 35100 53830
rect 35156 53828 35180 53830
rect 35236 53828 35242 53830
rect 34934 53819 35242 53828
rect 65654 53884 65962 53893
rect 65654 53882 65660 53884
rect 65716 53882 65740 53884
rect 65796 53882 65820 53884
rect 65876 53882 65900 53884
rect 65956 53882 65962 53884
rect 65716 53830 65718 53882
rect 65898 53830 65900 53882
rect 65654 53828 65660 53830
rect 65716 53828 65740 53830
rect 65796 53828 65820 53830
rect 65876 53828 65900 53830
rect 65956 53828 65962 53830
rect 65654 53819 65962 53828
rect 19574 53340 19882 53349
rect 19574 53338 19580 53340
rect 19636 53338 19660 53340
rect 19716 53338 19740 53340
rect 19796 53338 19820 53340
rect 19876 53338 19882 53340
rect 19636 53286 19638 53338
rect 19818 53286 19820 53338
rect 19574 53284 19580 53286
rect 19636 53284 19660 53286
rect 19716 53284 19740 53286
rect 19796 53284 19820 53286
rect 19876 53284 19882 53286
rect 19574 53275 19882 53284
rect 50294 53340 50602 53349
rect 50294 53338 50300 53340
rect 50356 53338 50380 53340
rect 50436 53338 50460 53340
rect 50516 53338 50540 53340
rect 50596 53338 50602 53340
rect 50356 53286 50358 53338
rect 50538 53286 50540 53338
rect 50294 53284 50300 53286
rect 50356 53284 50380 53286
rect 50436 53284 50460 53286
rect 50516 53284 50540 53286
rect 50596 53284 50602 53286
rect 50294 53275 50602 53284
rect 4214 52796 4522 52805
rect 4214 52794 4220 52796
rect 4276 52794 4300 52796
rect 4356 52794 4380 52796
rect 4436 52794 4460 52796
rect 4516 52794 4522 52796
rect 4276 52742 4278 52794
rect 4458 52742 4460 52794
rect 4214 52740 4220 52742
rect 4276 52740 4300 52742
rect 4356 52740 4380 52742
rect 4436 52740 4460 52742
rect 4516 52740 4522 52742
rect 4214 52731 4522 52740
rect 34934 52796 35242 52805
rect 34934 52794 34940 52796
rect 34996 52794 35020 52796
rect 35076 52794 35100 52796
rect 35156 52794 35180 52796
rect 35236 52794 35242 52796
rect 34996 52742 34998 52794
rect 35178 52742 35180 52794
rect 34934 52740 34940 52742
rect 34996 52740 35020 52742
rect 35076 52740 35100 52742
rect 35156 52740 35180 52742
rect 35236 52740 35242 52742
rect 34934 52731 35242 52740
rect 65654 52796 65962 52805
rect 65654 52794 65660 52796
rect 65716 52794 65740 52796
rect 65796 52794 65820 52796
rect 65876 52794 65900 52796
rect 65956 52794 65962 52796
rect 65716 52742 65718 52794
rect 65898 52742 65900 52794
rect 65654 52740 65660 52742
rect 65716 52740 65740 52742
rect 65796 52740 65820 52742
rect 65876 52740 65900 52742
rect 65956 52740 65962 52742
rect 65654 52731 65962 52740
rect 19574 52252 19882 52261
rect 19574 52250 19580 52252
rect 19636 52250 19660 52252
rect 19716 52250 19740 52252
rect 19796 52250 19820 52252
rect 19876 52250 19882 52252
rect 19636 52198 19638 52250
rect 19818 52198 19820 52250
rect 19574 52196 19580 52198
rect 19636 52196 19660 52198
rect 19716 52196 19740 52198
rect 19796 52196 19820 52198
rect 19876 52196 19882 52198
rect 19574 52187 19882 52196
rect 50294 52252 50602 52261
rect 50294 52250 50300 52252
rect 50356 52250 50380 52252
rect 50436 52250 50460 52252
rect 50516 52250 50540 52252
rect 50596 52250 50602 52252
rect 50356 52198 50358 52250
rect 50538 52198 50540 52250
rect 50294 52196 50300 52198
rect 50356 52196 50380 52198
rect 50436 52196 50460 52198
rect 50516 52196 50540 52198
rect 50596 52196 50602 52198
rect 50294 52187 50602 52196
rect 4214 51708 4522 51717
rect 4214 51706 4220 51708
rect 4276 51706 4300 51708
rect 4356 51706 4380 51708
rect 4436 51706 4460 51708
rect 4516 51706 4522 51708
rect 4276 51654 4278 51706
rect 4458 51654 4460 51706
rect 4214 51652 4220 51654
rect 4276 51652 4300 51654
rect 4356 51652 4380 51654
rect 4436 51652 4460 51654
rect 4516 51652 4522 51654
rect 4214 51643 4522 51652
rect 34934 51708 35242 51717
rect 34934 51706 34940 51708
rect 34996 51706 35020 51708
rect 35076 51706 35100 51708
rect 35156 51706 35180 51708
rect 35236 51706 35242 51708
rect 34996 51654 34998 51706
rect 35178 51654 35180 51706
rect 34934 51652 34940 51654
rect 34996 51652 35020 51654
rect 35076 51652 35100 51654
rect 35156 51652 35180 51654
rect 35236 51652 35242 51654
rect 34934 51643 35242 51652
rect 65654 51708 65962 51717
rect 65654 51706 65660 51708
rect 65716 51706 65740 51708
rect 65796 51706 65820 51708
rect 65876 51706 65900 51708
rect 65956 51706 65962 51708
rect 65716 51654 65718 51706
rect 65898 51654 65900 51706
rect 65654 51652 65660 51654
rect 65716 51652 65740 51654
rect 65796 51652 65820 51654
rect 65876 51652 65900 51654
rect 65956 51652 65962 51654
rect 65654 51643 65962 51652
rect 19574 51164 19882 51173
rect 19574 51162 19580 51164
rect 19636 51162 19660 51164
rect 19716 51162 19740 51164
rect 19796 51162 19820 51164
rect 19876 51162 19882 51164
rect 19636 51110 19638 51162
rect 19818 51110 19820 51162
rect 19574 51108 19580 51110
rect 19636 51108 19660 51110
rect 19716 51108 19740 51110
rect 19796 51108 19820 51110
rect 19876 51108 19882 51110
rect 19574 51099 19882 51108
rect 50294 51164 50602 51173
rect 50294 51162 50300 51164
rect 50356 51162 50380 51164
rect 50436 51162 50460 51164
rect 50516 51162 50540 51164
rect 50596 51162 50602 51164
rect 50356 51110 50358 51162
rect 50538 51110 50540 51162
rect 50294 51108 50300 51110
rect 50356 51108 50380 51110
rect 50436 51108 50460 51110
rect 50516 51108 50540 51110
rect 50596 51108 50602 51110
rect 50294 51099 50602 51108
rect 4214 50620 4522 50629
rect 4214 50618 4220 50620
rect 4276 50618 4300 50620
rect 4356 50618 4380 50620
rect 4436 50618 4460 50620
rect 4516 50618 4522 50620
rect 4276 50566 4278 50618
rect 4458 50566 4460 50618
rect 4214 50564 4220 50566
rect 4276 50564 4300 50566
rect 4356 50564 4380 50566
rect 4436 50564 4460 50566
rect 4516 50564 4522 50566
rect 4214 50555 4522 50564
rect 34934 50620 35242 50629
rect 34934 50618 34940 50620
rect 34996 50618 35020 50620
rect 35076 50618 35100 50620
rect 35156 50618 35180 50620
rect 35236 50618 35242 50620
rect 34996 50566 34998 50618
rect 35178 50566 35180 50618
rect 34934 50564 34940 50566
rect 34996 50564 35020 50566
rect 35076 50564 35100 50566
rect 35156 50564 35180 50566
rect 35236 50564 35242 50566
rect 34934 50555 35242 50564
rect 65654 50620 65962 50629
rect 65654 50618 65660 50620
rect 65716 50618 65740 50620
rect 65796 50618 65820 50620
rect 65876 50618 65900 50620
rect 65956 50618 65962 50620
rect 65716 50566 65718 50618
rect 65898 50566 65900 50618
rect 65654 50564 65660 50566
rect 65716 50564 65740 50566
rect 65796 50564 65820 50566
rect 65876 50564 65900 50566
rect 65956 50564 65962 50566
rect 65654 50555 65962 50564
rect 19574 50076 19882 50085
rect 19574 50074 19580 50076
rect 19636 50074 19660 50076
rect 19716 50074 19740 50076
rect 19796 50074 19820 50076
rect 19876 50074 19882 50076
rect 19636 50022 19638 50074
rect 19818 50022 19820 50074
rect 19574 50020 19580 50022
rect 19636 50020 19660 50022
rect 19716 50020 19740 50022
rect 19796 50020 19820 50022
rect 19876 50020 19882 50022
rect 19574 50011 19882 50020
rect 50294 50076 50602 50085
rect 50294 50074 50300 50076
rect 50356 50074 50380 50076
rect 50436 50074 50460 50076
rect 50516 50074 50540 50076
rect 50596 50074 50602 50076
rect 50356 50022 50358 50074
rect 50538 50022 50540 50074
rect 50294 50020 50300 50022
rect 50356 50020 50380 50022
rect 50436 50020 50460 50022
rect 50516 50020 50540 50022
rect 50596 50020 50602 50022
rect 50294 50011 50602 50020
rect 4214 49532 4522 49541
rect 4214 49530 4220 49532
rect 4276 49530 4300 49532
rect 4356 49530 4380 49532
rect 4436 49530 4460 49532
rect 4516 49530 4522 49532
rect 4276 49478 4278 49530
rect 4458 49478 4460 49530
rect 4214 49476 4220 49478
rect 4276 49476 4300 49478
rect 4356 49476 4380 49478
rect 4436 49476 4460 49478
rect 4516 49476 4522 49478
rect 4214 49467 4522 49476
rect 34934 49532 35242 49541
rect 34934 49530 34940 49532
rect 34996 49530 35020 49532
rect 35076 49530 35100 49532
rect 35156 49530 35180 49532
rect 35236 49530 35242 49532
rect 34996 49478 34998 49530
rect 35178 49478 35180 49530
rect 34934 49476 34940 49478
rect 34996 49476 35020 49478
rect 35076 49476 35100 49478
rect 35156 49476 35180 49478
rect 35236 49476 35242 49478
rect 34934 49467 35242 49476
rect 65654 49532 65962 49541
rect 65654 49530 65660 49532
rect 65716 49530 65740 49532
rect 65796 49530 65820 49532
rect 65876 49530 65900 49532
rect 65956 49530 65962 49532
rect 65716 49478 65718 49530
rect 65898 49478 65900 49530
rect 65654 49476 65660 49478
rect 65716 49476 65740 49478
rect 65796 49476 65820 49478
rect 65876 49476 65900 49478
rect 65956 49476 65962 49478
rect 65654 49467 65962 49476
rect 19574 48988 19882 48997
rect 19574 48986 19580 48988
rect 19636 48986 19660 48988
rect 19716 48986 19740 48988
rect 19796 48986 19820 48988
rect 19876 48986 19882 48988
rect 19636 48934 19638 48986
rect 19818 48934 19820 48986
rect 19574 48932 19580 48934
rect 19636 48932 19660 48934
rect 19716 48932 19740 48934
rect 19796 48932 19820 48934
rect 19876 48932 19882 48934
rect 19574 48923 19882 48932
rect 50294 48988 50602 48997
rect 50294 48986 50300 48988
rect 50356 48986 50380 48988
rect 50436 48986 50460 48988
rect 50516 48986 50540 48988
rect 50596 48986 50602 48988
rect 50356 48934 50358 48986
rect 50538 48934 50540 48986
rect 50294 48932 50300 48934
rect 50356 48932 50380 48934
rect 50436 48932 50460 48934
rect 50516 48932 50540 48934
rect 50596 48932 50602 48934
rect 50294 48923 50602 48932
rect 4214 48444 4522 48453
rect 4214 48442 4220 48444
rect 4276 48442 4300 48444
rect 4356 48442 4380 48444
rect 4436 48442 4460 48444
rect 4516 48442 4522 48444
rect 4276 48390 4278 48442
rect 4458 48390 4460 48442
rect 4214 48388 4220 48390
rect 4276 48388 4300 48390
rect 4356 48388 4380 48390
rect 4436 48388 4460 48390
rect 4516 48388 4522 48390
rect 4214 48379 4522 48388
rect 34934 48444 35242 48453
rect 34934 48442 34940 48444
rect 34996 48442 35020 48444
rect 35076 48442 35100 48444
rect 35156 48442 35180 48444
rect 35236 48442 35242 48444
rect 34996 48390 34998 48442
rect 35178 48390 35180 48442
rect 34934 48388 34940 48390
rect 34996 48388 35020 48390
rect 35076 48388 35100 48390
rect 35156 48388 35180 48390
rect 35236 48388 35242 48390
rect 34934 48379 35242 48388
rect 65654 48444 65962 48453
rect 65654 48442 65660 48444
rect 65716 48442 65740 48444
rect 65796 48442 65820 48444
rect 65876 48442 65900 48444
rect 65956 48442 65962 48444
rect 65716 48390 65718 48442
rect 65898 48390 65900 48442
rect 65654 48388 65660 48390
rect 65716 48388 65740 48390
rect 65796 48388 65820 48390
rect 65876 48388 65900 48390
rect 65956 48388 65962 48390
rect 65654 48379 65962 48388
rect 19574 47900 19882 47909
rect 19574 47898 19580 47900
rect 19636 47898 19660 47900
rect 19716 47898 19740 47900
rect 19796 47898 19820 47900
rect 19876 47898 19882 47900
rect 19636 47846 19638 47898
rect 19818 47846 19820 47898
rect 19574 47844 19580 47846
rect 19636 47844 19660 47846
rect 19716 47844 19740 47846
rect 19796 47844 19820 47846
rect 19876 47844 19882 47846
rect 19574 47835 19882 47844
rect 50294 47900 50602 47909
rect 50294 47898 50300 47900
rect 50356 47898 50380 47900
rect 50436 47898 50460 47900
rect 50516 47898 50540 47900
rect 50596 47898 50602 47900
rect 50356 47846 50358 47898
rect 50538 47846 50540 47898
rect 50294 47844 50300 47846
rect 50356 47844 50380 47846
rect 50436 47844 50460 47846
rect 50516 47844 50540 47846
rect 50596 47844 50602 47846
rect 50294 47835 50602 47844
rect 4214 47356 4522 47365
rect 4214 47354 4220 47356
rect 4276 47354 4300 47356
rect 4356 47354 4380 47356
rect 4436 47354 4460 47356
rect 4516 47354 4522 47356
rect 4276 47302 4278 47354
rect 4458 47302 4460 47354
rect 4214 47300 4220 47302
rect 4276 47300 4300 47302
rect 4356 47300 4380 47302
rect 4436 47300 4460 47302
rect 4516 47300 4522 47302
rect 4214 47291 4522 47300
rect 34934 47356 35242 47365
rect 34934 47354 34940 47356
rect 34996 47354 35020 47356
rect 35076 47354 35100 47356
rect 35156 47354 35180 47356
rect 35236 47354 35242 47356
rect 34996 47302 34998 47354
rect 35178 47302 35180 47354
rect 34934 47300 34940 47302
rect 34996 47300 35020 47302
rect 35076 47300 35100 47302
rect 35156 47300 35180 47302
rect 35236 47300 35242 47302
rect 34934 47291 35242 47300
rect 65654 47356 65962 47365
rect 65654 47354 65660 47356
rect 65716 47354 65740 47356
rect 65796 47354 65820 47356
rect 65876 47354 65900 47356
rect 65956 47354 65962 47356
rect 65716 47302 65718 47354
rect 65898 47302 65900 47354
rect 65654 47300 65660 47302
rect 65716 47300 65740 47302
rect 65796 47300 65820 47302
rect 65876 47300 65900 47302
rect 65956 47300 65962 47302
rect 65654 47291 65962 47300
rect 19574 46812 19882 46821
rect 19574 46810 19580 46812
rect 19636 46810 19660 46812
rect 19716 46810 19740 46812
rect 19796 46810 19820 46812
rect 19876 46810 19882 46812
rect 19636 46758 19638 46810
rect 19818 46758 19820 46810
rect 19574 46756 19580 46758
rect 19636 46756 19660 46758
rect 19716 46756 19740 46758
rect 19796 46756 19820 46758
rect 19876 46756 19882 46758
rect 19574 46747 19882 46756
rect 50294 46812 50602 46821
rect 50294 46810 50300 46812
rect 50356 46810 50380 46812
rect 50436 46810 50460 46812
rect 50516 46810 50540 46812
rect 50596 46810 50602 46812
rect 50356 46758 50358 46810
rect 50538 46758 50540 46810
rect 50294 46756 50300 46758
rect 50356 46756 50380 46758
rect 50436 46756 50460 46758
rect 50516 46756 50540 46758
rect 50596 46756 50602 46758
rect 50294 46747 50602 46756
rect 4214 46268 4522 46277
rect 4214 46266 4220 46268
rect 4276 46266 4300 46268
rect 4356 46266 4380 46268
rect 4436 46266 4460 46268
rect 4516 46266 4522 46268
rect 4276 46214 4278 46266
rect 4458 46214 4460 46266
rect 4214 46212 4220 46214
rect 4276 46212 4300 46214
rect 4356 46212 4380 46214
rect 4436 46212 4460 46214
rect 4516 46212 4522 46214
rect 4214 46203 4522 46212
rect 34934 46268 35242 46277
rect 34934 46266 34940 46268
rect 34996 46266 35020 46268
rect 35076 46266 35100 46268
rect 35156 46266 35180 46268
rect 35236 46266 35242 46268
rect 34996 46214 34998 46266
rect 35178 46214 35180 46266
rect 34934 46212 34940 46214
rect 34996 46212 35020 46214
rect 35076 46212 35100 46214
rect 35156 46212 35180 46214
rect 35236 46212 35242 46214
rect 34934 46203 35242 46212
rect 65654 46268 65962 46277
rect 65654 46266 65660 46268
rect 65716 46266 65740 46268
rect 65796 46266 65820 46268
rect 65876 46266 65900 46268
rect 65956 46266 65962 46268
rect 65716 46214 65718 46266
rect 65898 46214 65900 46266
rect 65654 46212 65660 46214
rect 65716 46212 65740 46214
rect 65796 46212 65820 46214
rect 65876 46212 65900 46214
rect 65956 46212 65962 46214
rect 65654 46203 65962 46212
rect 19574 45724 19882 45733
rect 19574 45722 19580 45724
rect 19636 45722 19660 45724
rect 19716 45722 19740 45724
rect 19796 45722 19820 45724
rect 19876 45722 19882 45724
rect 19636 45670 19638 45722
rect 19818 45670 19820 45722
rect 19574 45668 19580 45670
rect 19636 45668 19660 45670
rect 19716 45668 19740 45670
rect 19796 45668 19820 45670
rect 19876 45668 19882 45670
rect 19574 45659 19882 45668
rect 50294 45724 50602 45733
rect 50294 45722 50300 45724
rect 50356 45722 50380 45724
rect 50436 45722 50460 45724
rect 50516 45722 50540 45724
rect 50596 45722 50602 45724
rect 50356 45670 50358 45722
rect 50538 45670 50540 45722
rect 50294 45668 50300 45670
rect 50356 45668 50380 45670
rect 50436 45668 50460 45670
rect 50516 45668 50540 45670
rect 50596 45668 50602 45670
rect 50294 45659 50602 45668
rect 4214 45180 4522 45189
rect 4214 45178 4220 45180
rect 4276 45178 4300 45180
rect 4356 45178 4380 45180
rect 4436 45178 4460 45180
rect 4516 45178 4522 45180
rect 4276 45126 4278 45178
rect 4458 45126 4460 45178
rect 4214 45124 4220 45126
rect 4276 45124 4300 45126
rect 4356 45124 4380 45126
rect 4436 45124 4460 45126
rect 4516 45124 4522 45126
rect 4214 45115 4522 45124
rect 34934 45180 35242 45189
rect 34934 45178 34940 45180
rect 34996 45178 35020 45180
rect 35076 45178 35100 45180
rect 35156 45178 35180 45180
rect 35236 45178 35242 45180
rect 34996 45126 34998 45178
rect 35178 45126 35180 45178
rect 34934 45124 34940 45126
rect 34996 45124 35020 45126
rect 35076 45124 35100 45126
rect 35156 45124 35180 45126
rect 35236 45124 35242 45126
rect 34934 45115 35242 45124
rect 65654 45180 65962 45189
rect 65654 45178 65660 45180
rect 65716 45178 65740 45180
rect 65796 45178 65820 45180
rect 65876 45178 65900 45180
rect 65956 45178 65962 45180
rect 65716 45126 65718 45178
rect 65898 45126 65900 45178
rect 65654 45124 65660 45126
rect 65716 45124 65740 45126
rect 65796 45124 65820 45126
rect 65876 45124 65900 45126
rect 65956 45124 65962 45126
rect 65654 45115 65962 45124
rect 19574 44636 19882 44645
rect 19574 44634 19580 44636
rect 19636 44634 19660 44636
rect 19716 44634 19740 44636
rect 19796 44634 19820 44636
rect 19876 44634 19882 44636
rect 19636 44582 19638 44634
rect 19818 44582 19820 44634
rect 19574 44580 19580 44582
rect 19636 44580 19660 44582
rect 19716 44580 19740 44582
rect 19796 44580 19820 44582
rect 19876 44580 19882 44582
rect 19574 44571 19882 44580
rect 50294 44636 50602 44645
rect 50294 44634 50300 44636
rect 50356 44634 50380 44636
rect 50436 44634 50460 44636
rect 50516 44634 50540 44636
rect 50596 44634 50602 44636
rect 50356 44582 50358 44634
rect 50538 44582 50540 44634
rect 50294 44580 50300 44582
rect 50356 44580 50380 44582
rect 50436 44580 50460 44582
rect 50516 44580 50540 44582
rect 50596 44580 50602 44582
rect 50294 44571 50602 44580
rect 4214 44092 4522 44101
rect 4214 44090 4220 44092
rect 4276 44090 4300 44092
rect 4356 44090 4380 44092
rect 4436 44090 4460 44092
rect 4516 44090 4522 44092
rect 4276 44038 4278 44090
rect 4458 44038 4460 44090
rect 4214 44036 4220 44038
rect 4276 44036 4300 44038
rect 4356 44036 4380 44038
rect 4436 44036 4460 44038
rect 4516 44036 4522 44038
rect 4214 44027 4522 44036
rect 34934 44092 35242 44101
rect 34934 44090 34940 44092
rect 34996 44090 35020 44092
rect 35076 44090 35100 44092
rect 35156 44090 35180 44092
rect 35236 44090 35242 44092
rect 34996 44038 34998 44090
rect 35178 44038 35180 44090
rect 34934 44036 34940 44038
rect 34996 44036 35020 44038
rect 35076 44036 35100 44038
rect 35156 44036 35180 44038
rect 35236 44036 35242 44038
rect 34934 44027 35242 44036
rect 65654 44092 65962 44101
rect 65654 44090 65660 44092
rect 65716 44090 65740 44092
rect 65796 44090 65820 44092
rect 65876 44090 65900 44092
rect 65956 44090 65962 44092
rect 65716 44038 65718 44090
rect 65898 44038 65900 44090
rect 65654 44036 65660 44038
rect 65716 44036 65740 44038
rect 65796 44036 65820 44038
rect 65876 44036 65900 44038
rect 65956 44036 65962 44038
rect 65654 44027 65962 44036
rect 19574 43548 19882 43557
rect 19574 43546 19580 43548
rect 19636 43546 19660 43548
rect 19716 43546 19740 43548
rect 19796 43546 19820 43548
rect 19876 43546 19882 43548
rect 19636 43494 19638 43546
rect 19818 43494 19820 43546
rect 19574 43492 19580 43494
rect 19636 43492 19660 43494
rect 19716 43492 19740 43494
rect 19796 43492 19820 43494
rect 19876 43492 19882 43494
rect 19574 43483 19882 43492
rect 50294 43548 50602 43557
rect 50294 43546 50300 43548
rect 50356 43546 50380 43548
rect 50436 43546 50460 43548
rect 50516 43546 50540 43548
rect 50596 43546 50602 43548
rect 50356 43494 50358 43546
rect 50538 43494 50540 43546
rect 50294 43492 50300 43494
rect 50356 43492 50380 43494
rect 50436 43492 50460 43494
rect 50516 43492 50540 43494
rect 50596 43492 50602 43494
rect 50294 43483 50602 43492
rect 4214 43004 4522 43013
rect 4214 43002 4220 43004
rect 4276 43002 4300 43004
rect 4356 43002 4380 43004
rect 4436 43002 4460 43004
rect 4516 43002 4522 43004
rect 4276 42950 4278 43002
rect 4458 42950 4460 43002
rect 4214 42948 4220 42950
rect 4276 42948 4300 42950
rect 4356 42948 4380 42950
rect 4436 42948 4460 42950
rect 4516 42948 4522 42950
rect 4214 42939 4522 42948
rect 34934 43004 35242 43013
rect 34934 43002 34940 43004
rect 34996 43002 35020 43004
rect 35076 43002 35100 43004
rect 35156 43002 35180 43004
rect 35236 43002 35242 43004
rect 34996 42950 34998 43002
rect 35178 42950 35180 43002
rect 34934 42948 34940 42950
rect 34996 42948 35020 42950
rect 35076 42948 35100 42950
rect 35156 42948 35180 42950
rect 35236 42948 35242 42950
rect 34934 42939 35242 42948
rect 65654 43004 65962 43013
rect 65654 43002 65660 43004
rect 65716 43002 65740 43004
rect 65796 43002 65820 43004
rect 65876 43002 65900 43004
rect 65956 43002 65962 43004
rect 65716 42950 65718 43002
rect 65898 42950 65900 43002
rect 65654 42948 65660 42950
rect 65716 42948 65740 42950
rect 65796 42948 65820 42950
rect 65876 42948 65900 42950
rect 65956 42948 65962 42950
rect 65654 42939 65962 42948
rect 19574 42460 19882 42469
rect 19574 42458 19580 42460
rect 19636 42458 19660 42460
rect 19716 42458 19740 42460
rect 19796 42458 19820 42460
rect 19876 42458 19882 42460
rect 19636 42406 19638 42458
rect 19818 42406 19820 42458
rect 19574 42404 19580 42406
rect 19636 42404 19660 42406
rect 19716 42404 19740 42406
rect 19796 42404 19820 42406
rect 19876 42404 19882 42406
rect 19574 42395 19882 42404
rect 50294 42460 50602 42469
rect 50294 42458 50300 42460
rect 50356 42458 50380 42460
rect 50436 42458 50460 42460
rect 50516 42458 50540 42460
rect 50596 42458 50602 42460
rect 50356 42406 50358 42458
rect 50538 42406 50540 42458
rect 50294 42404 50300 42406
rect 50356 42404 50380 42406
rect 50436 42404 50460 42406
rect 50516 42404 50540 42406
rect 50596 42404 50602 42406
rect 50294 42395 50602 42404
rect 4214 41916 4522 41925
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41851 4522 41860
rect 34934 41916 35242 41925
rect 34934 41914 34940 41916
rect 34996 41914 35020 41916
rect 35076 41914 35100 41916
rect 35156 41914 35180 41916
rect 35236 41914 35242 41916
rect 34996 41862 34998 41914
rect 35178 41862 35180 41914
rect 34934 41860 34940 41862
rect 34996 41860 35020 41862
rect 35076 41860 35100 41862
rect 35156 41860 35180 41862
rect 35236 41860 35242 41862
rect 34934 41851 35242 41860
rect 65654 41916 65962 41925
rect 65654 41914 65660 41916
rect 65716 41914 65740 41916
rect 65796 41914 65820 41916
rect 65876 41914 65900 41916
rect 65956 41914 65962 41916
rect 65716 41862 65718 41914
rect 65898 41862 65900 41914
rect 65654 41860 65660 41862
rect 65716 41860 65740 41862
rect 65796 41860 65820 41862
rect 65876 41860 65900 41862
rect 65956 41860 65962 41862
rect 65654 41851 65962 41860
rect 19574 41372 19882 41381
rect 19574 41370 19580 41372
rect 19636 41370 19660 41372
rect 19716 41370 19740 41372
rect 19796 41370 19820 41372
rect 19876 41370 19882 41372
rect 19636 41318 19638 41370
rect 19818 41318 19820 41370
rect 19574 41316 19580 41318
rect 19636 41316 19660 41318
rect 19716 41316 19740 41318
rect 19796 41316 19820 41318
rect 19876 41316 19882 41318
rect 19574 41307 19882 41316
rect 50294 41372 50602 41381
rect 50294 41370 50300 41372
rect 50356 41370 50380 41372
rect 50436 41370 50460 41372
rect 50516 41370 50540 41372
rect 50596 41370 50602 41372
rect 50356 41318 50358 41370
rect 50538 41318 50540 41370
rect 50294 41316 50300 41318
rect 50356 41316 50380 41318
rect 50436 41316 50460 41318
rect 50516 41316 50540 41318
rect 50596 41316 50602 41318
rect 50294 41307 50602 41316
rect 4214 40828 4522 40837
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40763 4522 40772
rect 34934 40828 35242 40837
rect 34934 40826 34940 40828
rect 34996 40826 35020 40828
rect 35076 40826 35100 40828
rect 35156 40826 35180 40828
rect 35236 40826 35242 40828
rect 34996 40774 34998 40826
rect 35178 40774 35180 40826
rect 34934 40772 34940 40774
rect 34996 40772 35020 40774
rect 35076 40772 35100 40774
rect 35156 40772 35180 40774
rect 35236 40772 35242 40774
rect 34934 40763 35242 40772
rect 65654 40828 65962 40837
rect 65654 40826 65660 40828
rect 65716 40826 65740 40828
rect 65796 40826 65820 40828
rect 65876 40826 65900 40828
rect 65956 40826 65962 40828
rect 65716 40774 65718 40826
rect 65898 40774 65900 40826
rect 65654 40772 65660 40774
rect 65716 40772 65740 40774
rect 65796 40772 65820 40774
rect 65876 40772 65900 40774
rect 65956 40772 65962 40774
rect 65654 40763 65962 40772
rect 19574 40284 19882 40293
rect 19574 40282 19580 40284
rect 19636 40282 19660 40284
rect 19716 40282 19740 40284
rect 19796 40282 19820 40284
rect 19876 40282 19882 40284
rect 19636 40230 19638 40282
rect 19818 40230 19820 40282
rect 19574 40228 19580 40230
rect 19636 40228 19660 40230
rect 19716 40228 19740 40230
rect 19796 40228 19820 40230
rect 19876 40228 19882 40230
rect 19574 40219 19882 40228
rect 50294 40284 50602 40293
rect 50294 40282 50300 40284
rect 50356 40282 50380 40284
rect 50436 40282 50460 40284
rect 50516 40282 50540 40284
rect 50596 40282 50602 40284
rect 50356 40230 50358 40282
rect 50538 40230 50540 40282
rect 50294 40228 50300 40230
rect 50356 40228 50380 40230
rect 50436 40228 50460 40230
rect 50516 40228 50540 40230
rect 50596 40228 50602 40230
rect 50294 40219 50602 40228
rect 4214 39740 4522 39749
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39675 4522 39684
rect 34934 39740 35242 39749
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39675 35242 39684
rect 65654 39740 65962 39749
rect 65654 39738 65660 39740
rect 65716 39738 65740 39740
rect 65796 39738 65820 39740
rect 65876 39738 65900 39740
rect 65956 39738 65962 39740
rect 65716 39686 65718 39738
rect 65898 39686 65900 39738
rect 65654 39684 65660 39686
rect 65716 39684 65740 39686
rect 65796 39684 65820 39686
rect 65876 39684 65900 39686
rect 65956 39684 65962 39686
rect 65654 39675 65962 39684
rect 19574 39196 19882 39205
rect 19574 39194 19580 39196
rect 19636 39194 19660 39196
rect 19716 39194 19740 39196
rect 19796 39194 19820 39196
rect 19876 39194 19882 39196
rect 19636 39142 19638 39194
rect 19818 39142 19820 39194
rect 19574 39140 19580 39142
rect 19636 39140 19660 39142
rect 19716 39140 19740 39142
rect 19796 39140 19820 39142
rect 19876 39140 19882 39142
rect 19574 39131 19882 39140
rect 50294 39196 50602 39205
rect 50294 39194 50300 39196
rect 50356 39194 50380 39196
rect 50436 39194 50460 39196
rect 50516 39194 50540 39196
rect 50596 39194 50602 39196
rect 50356 39142 50358 39194
rect 50538 39142 50540 39194
rect 50294 39140 50300 39142
rect 50356 39140 50380 39142
rect 50436 39140 50460 39142
rect 50516 39140 50540 39142
rect 50596 39140 50602 39142
rect 50294 39131 50602 39140
rect 4214 38652 4522 38661
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38587 4522 38596
rect 34934 38652 35242 38661
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38587 35242 38596
rect 65654 38652 65962 38661
rect 65654 38650 65660 38652
rect 65716 38650 65740 38652
rect 65796 38650 65820 38652
rect 65876 38650 65900 38652
rect 65956 38650 65962 38652
rect 65716 38598 65718 38650
rect 65898 38598 65900 38650
rect 65654 38596 65660 38598
rect 65716 38596 65740 38598
rect 65796 38596 65820 38598
rect 65876 38596 65900 38598
rect 65956 38596 65962 38598
rect 65654 38587 65962 38596
rect 19574 38108 19882 38117
rect 19574 38106 19580 38108
rect 19636 38106 19660 38108
rect 19716 38106 19740 38108
rect 19796 38106 19820 38108
rect 19876 38106 19882 38108
rect 19636 38054 19638 38106
rect 19818 38054 19820 38106
rect 19574 38052 19580 38054
rect 19636 38052 19660 38054
rect 19716 38052 19740 38054
rect 19796 38052 19820 38054
rect 19876 38052 19882 38054
rect 19574 38043 19882 38052
rect 50294 38108 50602 38117
rect 50294 38106 50300 38108
rect 50356 38106 50380 38108
rect 50436 38106 50460 38108
rect 50516 38106 50540 38108
rect 50596 38106 50602 38108
rect 50356 38054 50358 38106
rect 50538 38054 50540 38106
rect 50294 38052 50300 38054
rect 50356 38052 50380 38054
rect 50436 38052 50460 38054
rect 50516 38052 50540 38054
rect 50596 38052 50602 38054
rect 50294 38043 50602 38052
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 65654 37564 65962 37573
rect 65654 37562 65660 37564
rect 65716 37562 65740 37564
rect 65796 37562 65820 37564
rect 65876 37562 65900 37564
rect 65956 37562 65962 37564
rect 65716 37510 65718 37562
rect 65898 37510 65900 37562
rect 65654 37508 65660 37510
rect 65716 37508 65740 37510
rect 65796 37508 65820 37510
rect 65876 37508 65900 37510
rect 65956 37508 65962 37510
rect 65654 37499 65962 37508
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 50294 37020 50602 37029
rect 50294 37018 50300 37020
rect 50356 37018 50380 37020
rect 50436 37018 50460 37020
rect 50516 37018 50540 37020
rect 50596 37018 50602 37020
rect 50356 36966 50358 37018
rect 50538 36966 50540 37018
rect 50294 36964 50300 36966
rect 50356 36964 50380 36966
rect 50436 36964 50460 36966
rect 50516 36964 50540 36966
rect 50596 36964 50602 36966
rect 50294 36955 50602 36964
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 65654 36476 65962 36485
rect 65654 36474 65660 36476
rect 65716 36474 65740 36476
rect 65796 36474 65820 36476
rect 65876 36474 65900 36476
rect 65956 36474 65962 36476
rect 65716 36422 65718 36474
rect 65898 36422 65900 36474
rect 65654 36420 65660 36422
rect 65716 36420 65740 36422
rect 65796 36420 65820 36422
rect 65876 36420 65900 36422
rect 65956 36420 65962 36422
rect 65654 36411 65962 36420
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 50294 35932 50602 35941
rect 50294 35930 50300 35932
rect 50356 35930 50380 35932
rect 50436 35930 50460 35932
rect 50516 35930 50540 35932
rect 50596 35930 50602 35932
rect 50356 35878 50358 35930
rect 50538 35878 50540 35930
rect 50294 35876 50300 35878
rect 50356 35876 50380 35878
rect 50436 35876 50460 35878
rect 50516 35876 50540 35878
rect 50596 35876 50602 35878
rect 50294 35867 50602 35876
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 65654 35388 65962 35397
rect 65654 35386 65660 35388
rect 65716 35386 65740 35388
rect 65796 35386 65820 35388
rect 65876 35386 65900 35388
rect 65956 35386 65962 35388
rect 65716 35334 65718 35386
rect 65898 35334 65900 35386
rect 65654 35332 65660 35334
rect 65716 35332 65740 35334
rect 65796 35332 65820 35334
rect 65876 35332 65900 35334
rect 65956 35332 65962 35334
rect 65654 35323 65962 35332
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 50294 34844 50602 34853
rect 50294 34842 50300 34844
rect 50356 34842 50380 34844
rect 50436 34842 50460 34844
rect 50516 34842 50540 34844
rect 50596 34842 50602 34844
rect 50356 34790 50358 34842
rect 50538 34790 50540 34842
rect 50294 34788 50300 34790
rect 50356 34788 50380 34790
rect 50436 34788 50460 34790
rect 50516 34788 50540 34790
rect 50596 34788 50602 34790
rect 50294 34779 50602 34788
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 65654 34300 65962 34309
rect 65654 34298 65660 34300
rect 65716 34298 65740 34300
rect 65796 34298 65820 34300
rect 65876 34298 65900 34300
rect 65956 34298 65962 34300
rect 65716 34246 65718 34298
rect 65898 34246 65900 34298
rect 65654 34244 65660 34246
rect 65716 34244 65740 34246
rect 65796 34244 65820 34246
rect 65876 34244 65900 34246
rect 65956 34244 65962 34246
rect 65654 34235 65962 34244
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 50294 33756 50602 33765
rect 50294 33754 50300 33756
rect 50356 33754 50380 33756
rect 50436 33754 50460 33756
rect 50516 33754 50540 33756
rect 50596 33754 50602 33756
rect 50356 33702 50358 33754
rect 50538 33702 50540 33754
rect 50294 33700 50300 33702
rect 50356 33700 50380 33702
rect 50436 33700 50460 33702
rect 50516 33700 50540 33702
rect 50596 33700 50602 33702
rect 50294 33691 50602 33700
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 65654 33212 65962 33221
rect 65654 33210 65660 33212
rect 65716 33210 65740 33212
rect 65796 33210 65820 33212
rect 65876 33210 65900 33212
rect 65956 33210 65962 33212
rect 65716 33158 65718 33210
rect 65898 33158 65900 33210
rect 65654 33156 65660 33158
rect 65716 33156 65740 33158
rect 65796 33156 65820 33158
rect 65876 33156 65900 33158
rect 65956 33156 65962 33158
rect 65654 33147 65962 33156
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 50294 32668 50602 32677
rect 50294 32666 50300 32668
rect 50356 32666 50380 32668
rect 50436 32666 50460 32668
rect 50516 32666 50540 32668
rect 50596 32666 50602 32668
rect 50356 32614 50358 32666
rect 50538 32614 50540 32666
rect 50294 32612 50300 32614
rect 50356 32612 50380 32614
rect 50436 32612 50460 32614
rect 50516 32612 50540 32614
rect 50596 32612 50602 32614
rect 50294 32603 50602 32612
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 65654 32124 65962 32133
rect 65654 32122 65660 32124
rect 65716 32122 65740 32124
rect 65796 32122 65820 32124
rect 65876 32122 65900 32124
rect 65956 32122 65962 32124
rect 65716 32070 65718 32122
rect 65898 32070 65900 32122
rect 65654 32068 65660 32070
rect 65716 32068 65740 32070
rect 65796 32068 65820 32070
rect 65876 32068 65900 32070
rect 65956 32068 65962 32070
rect 65654 32059 65962 32068
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 50294 31580 50602 31589
rect 50294 31578 50300 31580
rect 50356 31578 50380 31580
rect 50436 31578 50460 31580
rect 50516 31578 50540 31580
rect 50596 31578 50602 31580
rect 50356 31526 50358 31578
rect 50538 31526 50540 31578
rect 50294 31524 50300 31526
rect 50356 31524 50380 31526
rect 50436 31524 50460 31526
rect 50516 31524 50540 31526
rect 50596 31524 50602 31526
rect 50294 31515 50602 31524
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 65654 31036 65962 31045
rect 65654 31034 65660 31036
rect 65716 31034 65740 31036
rect 65796 31034 65820 31036
rect 65876 31034 65900 31036
rect 65956 31034 65962 31036
rect 65716 30982 65718 31034
rect 65898 30982 65900 31034
rect 65654 30980 65660 30982
rect 65716 30980 65740 30982
rect 65796 30980 65820 30982
rect 65876 30980 65900 30982
rect 65956 30980 65962 30982
rect 65654 30971 65962 30980
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 50294 30492 50602 30501
rect 50294 30490 50300 30492
rect 50356 30490 50380 30492
rect 50436 30490 50460 30492
rect 50516 30490 50540 30492
rect 50596 30490 50602 30492
rect 50356 30438 50358 30490
rect 50538 30438 50540 30490
rect 50294 30436 50300 30438
rect 50356 30436 50380 30438
rect 50436 30436 50460 30438
rect 50516 30436 50540 30438
rect 50596 30436 50602 30438
rect 50294 30427 50602 30436
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 65654 29948 65962 29957
rect 65654 29946 65660 29948
rect 65716 29946 65740 29948
rect 65796 29946 65820 29948
rect 65876 29946 65900 29948
rect 65956 29946 65962 29948
rect 65716 29894 65718 29946
rect 65898 29894 65900 29946
rect 65654 29892 65660 29894
rect 65716 29892 65740 29894
rect 65796 29892 65820 29894
rect 65876 29892 65900 29894
rect 65956 29892 65962 29894
rect 65654 29883 65962 29892
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 50294 29404 50602 29413
rect 50294 29402 50300 29404
rect 50356 29402 50380 29404
rect 50436 29402 50460 29404
rect 50516 29402 50540 29404
rect 50596 29402 50602 29404
rect 50356 29350 50358 29402
rect 50538 29350 50540 29402
rect 50294 29348 50300 29350
rect 50356 29348 50380 29350
rect 50436 29348 50460 29350
rect 50516 29348 50540 29350
rect 50596 29348 50602 29350
rect 50294 29339 50602 29348
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 65654 28860 65962 28869
rect 65654 28858 65660 28860
rect 65716 28858 65740 28860
rect 65796 28858 65820 28860
rect 65876 28858 65900 28860
rect 65956 28858 65962 28860
rect 65716 28806 65718 28858
rect 65898 28806 65900 28858
rect 65654 28804 65660 28806
rect 65716 28804 65740 28806
rect 65796 28804 65820 28806
rect 65876 28804 65900 28806
rect 65956 28804 65962 28806
rect 65654 28795 65962 28804
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 50294 28316 50602 28325
rect 50294 28314 50300 28316
rect 50356 28314 50380 28316
rect 50436 28314 50460 28316
rect 50516 28314 50540 28316
rect 50596 28314 50602 28316
rect 50356 28262 50358 28314
rect 50538 28262 50540 28314
rect 50294 28260 50300 28262
rect 50356 28260 50380 28262
rect 50436 28260 50460 28262
rect 50516 28260 50540 28262
rect 50596 28260 50602 28262
rect 50294 28251 50602 28260
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 65654 27772 65962 27781
rect 65654 27770 65660 27772
rect 65716 27770 65740 27772
rect 65796 27770 65820 27772
rect 65876 27770 65900 27772
rect 65956 27770 65962 27772
rect 65716 27718 65718 27770
rect 65898 27718 65900 27770
rect 65654 27716 65660 27718
rect 65716 27716 65740 27718
rect 65796 27716 65820 27718
rect 65876 27716 65900 27718
rect 65956 27716 65962 27718
rect 65654 27707 65962 27716
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 50294 27228 50602 27237
rect 50294 27226 50300 27228
rect 50356 27226 50380 27228
rect 50436 27226 50460 27228
rect 50516 27226 50540 27228
rect 50596 27226 50602 27228
rect 50356 27174 50358 27226
rect 50538 27174 50540 27226
rect 50294 27172 50300 27174
rect 50356 27172 50380 27174
rect 50436 27172 50460 27174
rect 50516 27172 50540 27174
rect 50596 27172 50602 27174
rect 50294 27163 50602 27172
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 65654 26684 65962 26693
rect 65654 26682 65660 26684
rect 65716 26682 65740 26684
rect 65796 26682 65820 26684
rect 65876 26682 65900 26684
rect 65956 26682 65962 26684
rect 65716 26630 65718 26682
rect 65898 26630 65900 26682
rect 65654 26628 65660 26630
rect 65716 26628 65740 26630
rect 65796 26628 65820 26630
rect 65876 26628 65900 26630
rect 65956 26628 65962 26630
rect 65654 26619 65962 26628
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 50294 26140 50602 26149
rect 50294 26138 50300 26140
rect 50356 26138 50380 26140
rect 50436 26138 50460 26140
rect 50516 26138 50540 26140
rect 50596 26138 50602 26140
rect 50356 26086 50358 26138
rect 50538 26086 50540 26138
rect 50294 26084 50300 26086
rect 50356 26084 50380 26086
rect 50436 26084 50460 26086
rect 50516 26084 50540 26086
rect 50596 26084 50602 26086
rect 50294 26075 50602 26084
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 65654 25596 65962 25605
rect 65654 25594 65660 25596
rect 65716 25594 65740 25596
rect 65796 25594 65820 25596
rect 65876 25594 65900 25596
rect 65956 25594 65962 25596
rect 65716 25542 65718 25594
rect 65898 25542 65900 25594
rect 65654 25540 65660 25542
rect 65716 25540 65740 25542
rect 65796 25540 65820 25542
rect 65876 25540 65900 25542
rect 65956 25540 65962 25542
rect 65654 25531 65962 25540
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 50294 25052 50602 25061
rect 50294 25050 50300 25052
rect 50356 25050 50380 25052
rect 50436 25050 50460 25052
rect 50516 25050 50540 25052
rect 50596 25050 50602 25052
rect 50356 24998 50358 25050
rect 50538 24998 50540 25050
rect 50294 24996 50300 24998
rect 50356 24996 50380 24998
rect 50436 24996 50460 24998
rect 50516 24996 50540 24998
rect 50596 24996 50602 24998
rect 50294 24987 50602 24996
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 65654 24508 65962 24517
rect 65654 24506 65660 24508
rect 65716 24506 65740 24508
rect 65796 24506 65820 24508
rect 65876 24506 65900 24508
rect 65956 24506 65962 24508
rect 65716 24454 65718 24506
rect 65898 24454 65900 24506
rect 65654 24452 65660 24454
rect 65716 24452 65740 24454
rect 65796 24452 65820 24454
rect 65876 24452 65900 24454
rect 65956 24452 65962 24454
rect 65654 24443 65962 24452
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 50294 23964 50602 23973
rect 50294 23962 50300 23964
rect 50356 23962 50380 23964
rect 50436 23962 50460 23964
rect 50516 23962 50540 23964
rect 50596 23962 50602 23964
rect 50356 23910 50358 23962
rect 50538 23910 50540 23962
rect 50294 23908 50300 23910
rect 50356 23908 50380 23910
rect 50436 23908 50460 23910
rect 50516 23908 50540 23910
rect 50596 23908 50602 23910
rect 50294 23899 50602 23908
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 65654 23420 65962 23429
rect 65654 23418 65660 23420
rect 65716 23418 65740 23420
rect 65796 23418 65820 23420
rect 65876 23418 65900 23420
rect 65956 23418 65962 23420
rect 65716 23366 65718 23418
rect 65898 23366 65900 23418
rect 65654 23364 65660 23366
rect 65716 23364 65740 23366
rect 65796 23364 65820 23366
rect 65876 23364 65900 23366
rect 65956 23364 65962 23366
rect 65654 23355 65962 23364
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 50294 22876 50602 22885
rect 50294 22874 50300 22876
rect 50356 22874 50380 22876
rect 50436 22874 50460 22876
rect 50516 22874 50540 22876
rect 50596 22874 50602 22876
rect 50356 22822 50358 22874
rect 50538 22822 50540 22874
rect 50294 22820 50300 22822
rect 50356 22820 50380 22822
rect 50436 22820 50460 22822
rect 50516 22820 50540 22822
rect 50596 22820 50602 22822
rect 50294 22811 50602 22820
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 65654 22332 65962 22341
rect 65654 22330 65660 22332
rect 65716 22330 65740 22332
rect 65796 22330 65820 22332
rect 65876 22330 65900 22332
rect 65956 22330 65962 22332
rect 65716 22278 65718 22330
rect 65898 22278 65900 22330
rect 65654 22276 65660 22278
rect 65716 22276 65740 22278
rect 65796 22276 65820 22278
rect 65876 22276 65900 22278
rect 65956 22276 65962 22278
rect 65654 22267 65962 22276
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 50294 21788 50602 21797
rect 50294 21786 50300 21788
rect 50356 21786 50380 21788
rect 50436 21786 50460 21788
rect 50516 21786 50540 21788
rect 50596 21786 50602 21788
rect 50356 21734 50358 21786
rect 50538 21734 50540 21786
rect 50294 21732 50300 21734
rect 50356 21732 50380 21734
rect 50436 21732 50460 21734
rect 50516 21732 50540 21734
rect 50596 21732 50602 21734
rect 50294 21723 50602 21732
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 65654 21244 65962 21253
rect 65654 21242 65660 21244
rect 65716 21242 65740 21244
rect 65796 21242 65820 21244
rect 65876 21242 65900 21244
rect 65956 21242 65962 21244
rect 65716 21190 65718 21242
rect 65898 21190 65900 21242
rect 65654 21188 65660 21190
rect 65716 21188 65740 21190
rect 65796 21188 65820 21190
rect 65876 21188 65900 21190
rect 65956 21188 65962 21190
rect 65654 21179 65962 21188
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 50294 20700 50602 20709
rect 50294 20698 50300 20700
rect 50356 20698 50380 20700
rect 50436 20698 50460 20700
rect 50516 20698 50540 20700
rect 50596 20698 50602 20700
rect 50356 20646 50358 20698
rect 50538 20646 50540 20698
rect 50294 20644 50300 20646
rect 50356 20644 50380 20646
rect 50436 20644 50460 20646
rect 50516 20644 50540 20646
rect 50596 20644 50602 20646
rect 50294 20635 50602 20644
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 65654 20156 65962 20165
rect 65654 20154 65660 20156
rect 65716 20154 65740 20156
rect 65796 20154 65820 20156
rect 65876 20154 65900 20156
rect 65956 20154 65962 20156
rect 65716 20102 65718 20154
rect 65898 20102 65900 20154
rect 65654 20100 65660 20102
rect 65716 20100 65740 20102
rect 65796 20100 65820 20102
rect 65876 20100 65900 20102
rect 65956 20100 65962 20102
rect 65654 20091 65962 20100
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 50294 19612 50602 19621
rect 50294 19610 50300 19612
rect 50356 19610 50380 19612
rect 50436 19610 50460 19612
rect 50516 19610 50540 19612
rect 50596 19610 50602 19612
rect 50356 19558 50358 19610
rect 50538 19558 50540 19610
rect 50294 19556 50300 19558
rect 50356 19556 50380 19558
rect 50436 19556 50460 19558
rect 50516 19556 50540 19558
rect 50596 19556 50602 19558
rect 50294 19547 50602 19556
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 65654 19068 65962 19077
rect 65654 19066 65660 19068
rect 65716 19066 65740 19068
rect 65796 19066 65820 19068
rect 65876 19066 65900 19068
rect 65956 19066 65962 19068
rect 65716 19014 65718 19066
rect 65898 19014 65900 19066
rect 65654 19012 65660 19014
rect 65716 19012 65740 19014
rect 65796 19012 65820 19014
rect 65876 19012 65900 19014
rect 65956 19012 65962 19014
rect 65654 19003 65962 19012
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 50294 18524 50602 18533
rect 50294 18522 50300 18524
rect 50356 18522 50380 18524
rect 50436 18522 50460 18524
rect 50516 18522 50540 18524
rect 50596 18522 50602 18524
rect 50356 18470 50358 18522
rect 50538 18470 50540 18522
rect 50294 18468 50300 18470
rect 50356 18468 50380 18470
rect 50436 18468 50460 18470
rect 50516 18468 50540 18470
rect 50596 18468 50602 18470
rect 50294 18459 50602 18468
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 65654 17980 65962 17989
rect 65654 17978 65660 17980
rect 65716 17978 65740 17980
rect 65796 17978 65820 17980
rect 65876 17978 65900 17980
rect 65956 17978 65962 17980
rect 65716 17926 65718 17978
rect 65898 17926 65900 17978
rect 65654 17924 65660 17926
rect 65716 17924 65740 17926
rect 65796 17924 65820 17926
rect 65876 17924 65900 17926
rect 65956 17924 65962 17926
rect 65654 17915 65962 17924
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 50294 17436 50602 17445
rect 50294 17434 50300 17436
rect 50356 17434 50380 17436
rect 50436 17434 50460 17436
rect 50516 17434 50540 17436
rect 50596 17434 50602 17436
rect 50356 17382 50358 17434
rect 50538 17382 50540 17434
rect 50294 17380 50300 17382
rect 50356 17380 50380 17382
rect 50436 17380 50460 17382
rect 50516 17380 50540 17382
rect 50596 17380 50602 17382
rect 50294 17371 50602 17380
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 65654 16892 65962 16901
rect 65654 16890 65660 16892
rect 65716 16890 65740 16892
rect 65796 16890 65820 16892
rect 65876 16890 65900 16892
rect 65956 16890 65962 16892
rect 65716 16838 65718 16890
rect 65898 16838 65900 16890
rect 65654 16836 65660 16838
rect 65716 16836 65740 16838
rect 65796 16836 65820 16838
rect 65876 16836 65900 16838
rect 65956 16836 65962 16838
rect 65654 16827 65962 16836
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 50294 16348 50602 16357
rect 50294 16346 50300 16348
rect 50356 16346 50380 16348
rect 50436 16346 50460 16348
rect 50516 16346 50540 16348
rect 50596 16346 50602 16348
rect 50356 16294 50358 16346
rect 50538 16294 50540 16346
rect 50294 16292 50300 16294
rect 50356 16292 50380 16294
rect 50436 16292 50460 16294
rect 50516 16292 50540 16294
rect 50596 16292 50602 16294
rect 50294 16283 50602 16292
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 65654 15804 65962 15813
rect 65654 15802 65660 15804
rect 65716 15802 65740 15804
rect 65796 15802 65820 15804
rect 65876 15802 65900 15804
rect 65956 15802 65962 15804
rect 65716 15750 65718 15802
rect 65898 15750 65900 15802
rect 65654 15748 65660 15750
rect 65716 15748 65740 15750
rect 65796 15748 65820 15750
rect 65876 15748 65900 15750
rect 65956 15748 65962 15750
rect 65654 15739 65962 15748
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 50294 15260 50602 15269
rect 50294 15258 50300 15260
rect 50356 15258 50380 15260
rect 50436 15258 50460 15260
rect 50516 15258 50540 15260
rect 50596 15258 50602 15260
rect 50356 15206 50358 15258
rect 50538 15206 50540 15258
rect 50294 15204 50300 15206
rect 50356 15204 50380 15206
rect 50436 15204 50460 15206
rect 50516 15204 50540 15206
rect 50596 15204 50602 15206
rect 50294 15195 50602 15204
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 65654 14716 65962 14725
rect 65654 14714 65660 14716
rect 65716 14714 65740 14716
rect 65796 14714 65820 14716
rect 65876 14714 65900 14716
rect 65956 14714 65962 14716
rect 65716 14662 65718 14714
rect 65898 14662 65900 14714
rect 65654 14660 65660 14662
rect 65716 14660 65740 14662
rect 65796 14660 65820 14662
rect 65876 14660 65900 14662
rect 65956 14660 65962 14662
rect 65654 14651 65962 14660
rect 11704 14476 11756 14482
rect 11704 14418 11756 14424
rect 10508 14408 10560 14414
rect 10508 14350 10560 14356
rect 10416 14340 10468 14346
rect 10416 14282 10468 14288
rect 4344 14272 4396 14278
rect 4344 14214 4396 14220
rect 5080 14272 5132 14278
rect 5080 14214 5132 14220
rect 4356 14074 4384 14214
rect 4344 14068 4396 14074
rect 4344 14010 4396 14016
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4712 12844 4764 12850
rect 4712 12786 4764 12792
rect 4620 12776 4672 12782
rect 4620 12718 4672 12724
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4632 11354 4660 12718
rect 4724 12306 4752 12786
rect 4712 12300 4764 12306
rect 4712 12242 4764 12248
rect 4724 11762 4752 12242
rect 4712 11756 4764 11762
rect 4712 11698 4764 11704
rect 4436 11348 4488 11354
rect 4436 11290 4488 11296
rect 4620 11348 4672 11354
rect 4620 11290 4672 11296
rect 4344 11144 4396 11150
rect 4344 11086 4396 11092
rect 4160 11076 4212 11082
rect 4160 11018 4212 11024
rect 4172 10742 4200 11018
rect 4160 10736 4212 10742
rect 4160 10678 4212 10684
rect 4356 10606 4384 11086
rect 4344 10600 4396 10606
rect 4344 10542 4396 10548
rect 4448 10470 4476 11290
rect 4724 11150 4752 11698
rect 4804 11620 4856 11626
rect 4804 11562 4856 11568
rect 4712 11144 4764 11150
rect 4712 11086 4764 11092
rect 4816 10810 4844 11562
rect 4804 10804 4856 10810
rect 4804 10746 4856 10752
rect 4712 10668 4764 10674
rect 4712 10610 4764 10616
rect 4988 10668 5040 10674
rect 4988 10610 5040 10616
rect 4436 10464 4488 10470
rect 4436 10406 4488 10412
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 3332 9580 3384 9586
rect 3332 9522 3384 9528
rect 3344 8974 3372 9522
rect 4620 9512 4672 9518
rect 4620 9454 4672 9460
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 2688 8968 2740 8974
rect 2688 8910 2740 8916
rect 3332 8968 3384 8974
rect 3332 8910 3384 8916
rect 3884 8968 3936 8974
rect 3884 8910 3936 8916
rect 2700 8362 2728 8910
rect 3700 8832 3752 8838
rect 3700 8774 3752 8780
rect 2688 8356 2740 8362
rect 2688 8298 2740 8304
rect 2700 6866 2728 8298
rect 2688 6860 2740 6866
rect 2688 6802 2740 6808
rect 2700 6322 2728 6802
rect 3712 6390 3740 8774
rect 3896 7410 3924 8910
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4068 8016 4120 8022
rect 4068 7958 4120 7964
rect 3884 7404 3936 7410
rect 3884 7346 3936 7352
rect 3700 6384 3752 6390
rect 3700 6326 3752 6332
rect 2688 6316 2740 6322
rect 2688 6258 2740 6264
rect 3792 6316 3844 6322
rect 3792 6258 3844 6264
rect 3804 6118 3832 6258
rect 3896 6254 3924 7346
rect 4080 6322 4108 7958
rect 4632 7818 4660 9454
rect 4620 7812 4672 7818
rect 4620 7754 4672 7760
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4068 6316 4120 6322
rect 4068 6258 4120 6264
rect 3884 6248 3936 6254
rect 3884 6190 3936 6196
rect 3792 6112 3844 6118
rect 3792 6054 3844 6060
rect 3976 6112 4028 6118
rect 3976 6054 4028 6060
rect 3804 5710 3832 6054
rect 3988 5914 4016 6054
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 3976 5908 4028 5914
rect 3976 5850 4028 5856
rect 3792 5704 3844 5710
rect 3792 5646 3844 5652
rect 3804 5234 3832 5646
rect 3792 5228 3844 5234
rect 3792 5170 3844 5176
rect 3804 4622 3832 5170
rect 3988 5030 4016 5850
rect 3976 5024 4028 5030
rect 3976 4966 4028 4972
rect 3988 4826 4016 4966
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4632 4826 4660 7754
rect 3976 4820 4028 4826
rect 3976 4762 4028 4768
rect 4620 4820 4672 4826
rect 4620 4762 4672 4768
rect 3792 4616 3844 4622
rect 3792 4558 3844 4564
rect 3804 4146 3832 4558
rect 3882 4176 3938 4185
rect 3792 4140 3844 4146
rect 3882 4111 3938 4120
rect 3792 4082 3844 4088
rect 3896 3194 3924 4111
rect 3988 4010 4016 4762
rect 4068 4480 4120 4486
rect 4068 4422 4120 4428
rect 3976 4004 4028 4010
rect 3976 3946 4028 3952
rect 4080 3194 4108 4422
rect 4160 4140 4212 4146
rect 4160 4082 4212 4088
rect 4172 4010 4200 4082
rect 4160 4004 4212 4010
rect 4160 3946 4212 3952
rect 4620 3936 4672 3942
rect 4620 3878 4672 3884
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4252 3664 4304 3670
rect 4250 3632 4252 3641
rect 4304 3632 4306 3641
rect 4250 3567 4306 3576
rect 4160 3528 4212 3534
rect 4160 3470 4212 3476
rect 3884 3188 3936 3194
rect 3884 3130 3936 3136
rect 4068 3188 4120 3194
rect 4068 3130 4120 3136
rect 3896 2446 3924 3130
rect 4068 3052 4120 3058
rect 4172 3040 4200 3470
rect 4526 3360 4582 3369
rect 4526 3295 4582 3304
rect 4540 3126 4568 3295
rect 4632 3126 4660 3878
rect 4528 3120 4580 3126
rect 4528 3062 4580 3068
rect 4620 3120 4672 3126
rect 4620 3062 4672 3068
rect 4120 3012 4200 3040
rect 4068 2994 4120 3000
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 4724 2650 4752 10610
rect 5000 9994 5028 10610
rect 4988 9988 5040 9994
rect 4988 9930 5040 9936
rect 5000 9654 5028 9930
rect 4988 9648 5040 9654
rect 4988 9590 5040 9596
rect 4804 7744 4856 7750
rect 4804 7686 4856 7692
rect 4816 5370 4844 7686
rect 4988 7404 5040 7410
rect 4988 7346 5040 7352
rect 5000 6769 5028 7346
rect 4986 6760 5042 6769
rect 4986 6695 5042 6704
rect 4804 5364 4856 5370
rect 4804 5306 4856 5312
rect 4988 5092 5040 5098
rect 4988 5034 5040 5040
rect 4896 4616 4948 4622
rect 4896 4558 4948 4564
rect 4802 3496 4858 3505
rect 4802 3431 4858 3440
rect 4816 3398 4844 3431
rect 4804 3392 4856 3398
rect 4804 3334 4856 3340
rect 4712 2644 4764 2650
rect 4712 2586 4764 2592
rect 4908 2582 4936 4558
rect 5000 3602 5028 5034
rect 5092 4078 5120 14214
rect 5816 13932 5868 13938
rect 5816 13874 5868 13880
rect 8852 13932 8904 13938
rect 8852 13874 8904 13880
rect 5540 12232 5592 12238
rect 5540 12174 5592 12180
rect 5356 12164 5408 12170
rect 5356 12106 5408 12112
rect 5368 11898 5396 12106
rect 5552 11898 5580 12174
rect 5356 11892 5408 11898
rect 5356 11834 5408 11840
rect 5540 11892 5592 11898
rect 5592 11852 5672 11880
rect 5540 11834 5592 11840
rect 5448 11212 5500 11218
rect 5448 11154 5500 11160
rect 5172 10600 5224 10606
rect 5172 10542 5224 10548
rect 5184 10062 5212 10542
rect 5264 10464 5316 10470
rect 5264 10406 5316 10412
rect 5276 10266 5304 10406
rect 5460 10266 5488 11154
rect 5264 10260 5316 10266
rect 5264 10202 5316 10208
rect 5448 10260 5500 10266
rect 5448 10202 5500 10208
rect 5448 10124 5500 10130
rect 5448 10066 5500 10072
rect 5172 10056 5224 10062
rect 5172 9998 5224 10004
rect 5264 10056 5316 10062
rect 5264 9998 5316 10004
rect 5184 9518 5212 9998
rect 5172 9512 5224 9518
rect 5172 9454 5224 9460
rect 5276 6905 5304 9998
rect 5460 8498 5488 10066
rect 5644 9382 5672 11852
rect 5724 11144 5776 11150
rect 5724 11086 5776 11092
rect 5736 10674 5764 11086
rect 5724 10668 5776 10674
rect 5724 10610 5776 10616
rect 5736 10062 5764 10610
rect 5724 10056 5776 10062
rect 5724 9998 5776 10004
rect 5828 9738 5856 13874
rect 8116 13864 8168 13870
rect 8116 13806 8168 13812
rect 8760 13864 8812 13870
rect 8760 13806 8812 13812
rect 7288 13796 7340 13802
rect 7288 13738 7340 13744
rect 7300 13326 7328 13738
rect 7288 13320 7340 13326
rect 7288 13262 7340 13268
rect 6184 12776 6236 12782
rect 6184 12718 6236 12724
rect 6196 11694 6224 12718
rect 7300 12646 7328 13262
rect 7288 12640 7340 12646
rect 7288 12582 7340 12588
rect 7104 12232 7156 12238
rect 7156 12192 7236 12220
rect 7104 12174 7156 12180
rect 6368 11756 6420 11762
rect 6368 11698 6420 11704
rect 6184 11688 6236 11694
rect 6184 11630 6236 11636
rect 6196 11218 6224 11630
rect 6380 11354 6408 11698
rect 7208 11694 7236 12192
rect 7196 11688 7248 11694
rect 7196 11630 7248 11636
rect 6368 11348 6420 11354
rect 6368 11290 6420 11296
rect 6184 11212 6236 11218
rect 6184 11154 6236 11160
rect 6000 10736 6052 10742
rect 6000 10678 6052 10684
rect 5828 9710 5948 9738
rect 5632 9376 5684 9382
rect 5632 9318 5684 9324
rect 5644 8566 5672 9318
rect 5920 8634 5948 9710
rect 5908 8628 5960 8634
rect 5908 8570 5960 8576
rect 5632 8560 5684 8566
rect 5632 8502 5684 8508
rect 5448 8492 5500 8498
rect 5448 8434 5500 8440
rect 5460 8294 5488 8434
rect 5540 8356 5592 8362
rect 5540 8298 5592 8304
rect 5448 8288 5500 8294
rect 5448 8230 5500 8236
rect 5460 8090 5488 8230
rect 5448 8084 5500 8090
rect 5448 8026 5500 8032
rect 5552 7954 5580 8298
rect 5724 8288 5776 8294
rect 5724 8230 5776 8236
rect 5540 7948 5592 7954
rect 5540 7890 5592 7896
rect 5356 7472 5408 7478
rect 5356 7414 5408 7420
rect 5552 7426 5580 7890
rect 5632 7880 5684 7886
rect 5632 7822 5684 7828
rect 5644 7546 5672 7822
rect 5632 7540 5684 7546
rect 5632 7482 5684 7488
rect 5262 6896 5318 6905
rect 5172 6860 5224 6866
rect 5262 6831 5318 6840
rect 5172 6802 5224 6808
rect 5184 5166 5212 6802
rect 5368 6390 5396 7414
rect 5552 7398 5672 7426
rect 5540 7336 5592 7342
rect 5540 7278 5592 7284
rect 5448 6792 5500 6798
rect 5448 6734 5500 6740
rect 5356 6384 5408 6390
rect 5356 6326 5408 6332
rect 5264 6180 5316 6186
rect 5264 6122 5316 6128
rect 5172 5160 5224 5166
rect 5172 5102 5224 5108
rect 5172 5024 5224 5030
rect 5172 4966 5224 4972
rect 5080 4072 5132 4078
rect 5080 4014 5132 4020
rect 5092 3777 5120 4014
rect 5078 3768 5134 3777
rect 5078 3703 5134 3712
rect 5184 3670 5212 4966
rect 5172 3664 5224 3670
rect 5172 3606 5224 3612
rect 4988 3596 5040 3602
rect 4988 3538 5040 3544
rect 5184 3534 5212 3606
rect 5172 3528 5224 3534
rect 5172 3470 5224 3476
rect 5184 3058 5212 3470
rect 5172 3052 5224 3058
rect 5172 2994 5224 3000
rect 4896 2576 4948 2582
rect 4896 2518 4948 2524
rect 5184 2446 5212 2994
rect 5276 2446 5304 6122
rect 5368 5710 5396 6326
rect 5460 6254 5488 6734
rect 5552 6322 5580 7278
rect 5644 6798 5672 7398
rect 5736 7206 5764 8230
rect 5724 7200 5776 7206
rect 5724 7142 5776 7148
rect 5632 6792 5684 6798
rect 5632 6734 5684 6740
rect 5540 6316 5592 6322
rect 5540 6258 5592 6264
rect 5448 6248 5500 6254
rect 5448 6190 5500 6196
rect 5552 5794 5580 6258
rect 5460 5778 5580 5794
rect 5448 5772 5580 5778
rect 5500 5766 5580 5772
rect 5448 5714 5500 5720
rect 5356 5704 5408 5710
rect 5356 5646 5408 5652
rect 5368 4622 5396 5646
rect 5552 4690 5580 5766
rect 5644 5710 5672 6734
rect 5736 6118 5764 7142
rect 5724 6112 5776 6118
rect 5724 6054 5776 6060
rect 5736 5914 5764 6054
rect 5724 5908 5776 5914
rect 5724 5850 5776 5856
rect 5632 5704 5684 5710
rect 5632 5646 5684 5652
rect 5736 4826 5764 5850
rect 5724 4820 5776 4826
rect 5724 4762 5776 4768
rect 5722 4720 5778 4729
rect 5540 4684 5592 4690
rect 5722 4655 5778 4664
rect 5540 4626 5592 4632
rect 5736 4622 5764 4655
rect 5356 4616 5408 4622
rect 5356 4558 5408 4564
rect 5724 4616 5776 4622
rect 5724 4558 5776 4564
rect 5816 4140 5868 4146
rect 5816 4082 5868 4088
rect 5448 3936 5500 3942
rect 5448 3878 5500 3884
rect 5460 3398 5488 3878
rect 5448 3392 5500 3398
rect 5448 3334 5500 3340
rect 5460 3058 5488 3334
rect 5448 3052 5500 3058
rect 5448 2994 5500 3000
rect 5460 2446 5488 2994
rect 5828 2650 5856 4082
rect 5908 3120 5960 3126
rect 5908 3062 5960 3068
rect 5920 2990 5948 3062
rect 5908 2984 5960 2990
rect 5908 2926 5960 2932
rect 6012 2854 6040 10678
rect 6196 10606 6224 11154
rect 7208 10742 7236 11630
rect 7196 10736 7248 10742
rect 7196 10678 7248 10684
rect 6184 10600 6236 10606
rect 6184 10542 6236 10548
rect 6196 9926 6224 10542
rect 6368 10464 6420 10470
rect 6368 10406 6420 10412
rect 6092 9920 6144 9926
rect 6092 9862 6144 9868
rect 6184 9920 6236 9926
rect 6184 9862 6236 9868
rect 6104 9722 6132 9862
rect 6092 9716 6144 9722
rect 6092 9658 6144 9664
rect 6092 9580 6144 9586
rect 6092 9522 6144 9528
rect 6104 7410 6132 9522
rect 6196 8974 6224 9862
rect 6380 9382 6408 10406
rect 7208 10146 7236 10678
rect 8128 10266 8156 13806
rect 8576 13320 8628 13326
rect 8576 13262 8628 13268
rect 8392 12776 8444 12782
rect 8392 12718 8444 12724
rect 8404 12102 8432 12718
rect 8392 12096 8444 12102
rect 8392 12038 8444 12044
rect 8404 11830 8432 12038
rect 8392 11824 8444 11830
rect 8392 11766 8444 11772
rect 8588 11558 8616 13262
rect 8772 12850 8800 13806
rect 8864 13308 8892 13874
rect 9864 13864 9916 13870
rect 9864 13806 9916 13812
rect 9036 13728 9088 13734
rect 9036 13670 9088 13676
rect 9048 13530 9076 13670
rect 9036 13524 9088 13530
rect 9036 13466 9088 13472
rect 8944 13320 8996 13326
rect 8864 13280 8944 13308
rect 8944 13262 8996 13268
rect 8956 12850 8984 13262
rect 8760 12844 8812 12850
rect 8760 12786 8812 12792
rect 8944 12844 8996 12850
rect 8944 12786 8996 12792
rect 8772 11898 8800 12786
rect 9048 12646 9076 13466
rect 9220 13320 9272 13326
rect 9220 13262 9272 13268
rect 8852 12640 8904 12646
rect 8852 12582 8904 12588
rect 9036 12640 9088 12646
rect 9036 12582 9088 12588
rect 8760 11892 8812 11898
rect 8760 11834 8812 11840
rect 8576 11552 8628 11558
rect 8576 11494 8628 11500
rect 8588 11150 8616 11494
rect 8576 11144 8628 11150
rect 8576 11086 8628 11092
rect 8116 10260 8168 10266
rect 8116 10202 8168 10208
rect 7116 10118 7236 10146
rect 7116 10062 7144 10118
rect 7104 10056 7156 10062
rect 7104 9998 7156 10004
rect 6368 9376 6420 9382
rect 6368 9318 6420 9324
rect 7116 8974 7144 9998
rect 7748 9580 7800 9586
rect 7748 9522 7800 9528
rect 6184 8968 6236 8974
rect 6184 8910 6236 8916
rect 6644 8968 6696 8974
rect 6644 8910 6696 8916
rect 7104 8968 7156 8974
rect 7104 8910 7156 8916
rect 6276 8832 6328 8838
rect 6276 8774 6328 8780
rect 6184 8424 6236 8430
rect 6184 8366 6236 8372
rect 6196 7546 6224 8366
rect 6184 7540 6236 7546
rect 6184 7482 6236 7488
rect 6092 7404 6144 7410
rect 6092 7346 6144 7352
rect 6104 7002 6132 7346
rect 6092 6996 6144 7002
rect 6092 6938 6144 6944
rect 6092 6792 6144 6798
rect 6092 6734 6144 6740
rect 6104 6118 6132 6734
rect 6288 6322 6316 8774
rect 6656 8560 6684 8910
rect 6920 8832 6972 8838
rect 6920 8774 6972 8780
rect 6656 8498 6687 8560
rect 6932 8498 6960 8774
rect 6647 8492 6699 8498
rect 6647 8434 6699 8440
rect 6920 8492 6972 8498
rect 6920 8434 6972 8440
rect 6656 7750 6684 8434
rect 7116 7886 7144 8910
rect 7288 8900 7340 8906
rect 7288 8842 7340 8848
rect 7300 8634 7328 8842
rect 7288 8628 7340 8634
rect 7288 8570 7340 8576
rect 7104 7880 7156 7886
rect 7104 7822 7156 7828
rect 6644 7744 6696 7750
rect 6644 7686 6696 7692
rect 6656 6730 6684 7686
rect 7116 7478 7144 7822
rect 7104 7472 7156 7478
rect 7104 7414 7156 7420
rect 6644 6724 6696 6730
rect 6644 6666 6696 6672
rect 6276 6316 6328 6322
rect 6276 6258 6328 6264
rect 6092 6112 6144 6118
rect 6092 6054 6144 6060
rect 6184 5704 6236 5710
rect 6184 5646 6236 5652
rect 6196 5234 6224 5646
rect 6288 5642 6316 6258
rect 6552 6180 6604 6186
rect 6552 6122 6604 6128
rect 6564 5846 6592 6122
rect 6460 5840 6512 5846
rect 6460 5782 6512 5788
rect 6552 5840 6604 5846
rect 6552 5782 6604 5788
rect 6368 5704 6420 5710
rect 6368 5646 6420 5652
rect 6276 5636 6328 5642
rect 6276 5578 6328 5584
rect 6184 5228 6236 5234
rect 6184 5170 6236 5176
rect 6380 4826 6408 5646
rect 6368 4820 6420 4826
rect 6368 4762 6420 4768
rect 6276 4072 6328 4078
rect 6274 4040 6276 4049
rect 6328 4040 6330 4049
rect 6274 3975 6330 3984
rect 6092 3664 6144 3670
rect 6092 3606 6144 3612
rect 6104 3466 6132 3606
rect 6472 3534 6500 5782
rect 6656 5642 6684 6666
rect 6828 6112 6880 6118
rect 6828 6054 6880 6060
rect 6736 5704 6788 5710
rect 6840 5681 6868 6054
rect 7760 5914 7788 9522
rect 7840 9376 7892 9382
rect 7840 9318 7892 9324
rect 7852 8498 7880 9318
rect 7840 8492 7892 8498
rect 7840 8434 7892 8440
rect 7852 6118 7880 8434
rect 8392 8084 8444 8090
rect 8392 8026 8444 8032
rect 7932 7200 7984 7206
rect 7932 7142 7984 7148
rect 7840 6112 7892 6118
rect 7840 6054 7892 6060
rect 7748 5908 7800 5914
rect 7748 5850 7800 5856
rect 7852 5846 7880 6054
rect 7840 5840 7892 5846
rect 7840 5782 7892 5788
rect 7564 5772 7616 5778
rect 7564 5714 7616 5720
rect 6736 5646 6788 5652
rect 6826 5672 6882 5681
rect 6644 5636 6696 5642
rect 6644 5578 6696 5584
rect 6552 5568 6604 5574
rect 6552 5510 6604 5516
rect 6564 5234 6592 5510
rect 6552 5228 6604 5234
rect 6552 5170 6604 5176
rect 6656 5098 6684 5578
rect 6644 5092 6696 5098
rect 6644 5034 6696 5040
rect 6748 4758 6776 5646
rect 6826 5607 6882 5616
rect 7288 5568 7340 5574
rect 7288 5510 7340 5516
rect 6920 5228 6972 5234
rect 6920 5170 6972 5176
rect 6828 5024 6880 5030
rect 6828 4966 6880 4972
rect 6736 4752 6788 4758
rect 6736 4694 6788 4700
rect 6552 4616 6604 4622
rect 6552 4558 6604 4564
rect 6564 4457 6592 4558
rect 6550 4448 6606 4457
rect 6550 4383 6606 4392
rect 6840 4146 6868 4966
rect 6932 4282 6960 5170
rect 7300 4554 7328 5510
rect 7288 4548 7340 4554
rect 7288 4490 7340 4496
rect 6920 4276 6972 4282
rect 6920 4218 6972 4224
rect 6828 4140 6880 4146
rect 6828 4082 6880 4088
rect 6920 3936 6972 3942
rect 6920 3878 6972 3884
rect 6932 3602 6960 3878
rect 6920 3596 6972 3602
rect 6920 3538 6972 3544
rect 6460 3528 6512 3534
rect 6460 3470 6512 3476
rect 6092 3460 6144 3466
rect 6092 3402 6144 3408
rect 6828 3460 6880 3466
rect 6828 3402 6880 3408
rect 6840 3194 6868 3402
rect 7576 3398 7604 5714
rect 7944 5710 7972 7142
rect 8404 7002 8432 8026
rect 8760 7812 8812 7818
rect 8760 7754 8812 7760
rect 8392 6996 8444 7002
rect 8392 6938 8444 6944
rect 8300 6792 8352 6798
rect 8300 6734 8352 6740
rect 7932 5704 7984 5710
rect 7932 5646 7984 5652
rect 7944 4321 7972 5646
rect 8312 5030 8340 6734
rect 8392 6452 8444 6458
rect 8392 6394 8444 6400
rect 8404 5914 8432 6394
rect 8668 6112 8720 6118
rect 8666 6080 8668 6089
rect 8720 6080 8722 6089
rect 8666 6015 8722 6024
rect 8392 5908 8444 5914
rect 8392 5850 8444 5856
rect 8392 5228 8444 5234
rect 8392 5170 8444 5176
rect 8300 5024 8352 5030
rect 8300 4966 8352 4972
rect 8312 4622 8340 4966
rect 8404 4826 8432 5170
rect 8392 4820 8444 4826
rect 8392 4762 8444 4768
rect 8300 4616 8352 4622
rect 8300 4558 8352 4564
rect 7930 4312 7986 4321
rect 7930 4247 7986 4256
rect 8312 4214 8340 4558
rect 8300 4208 8352 4214
rect 8300 4150 8352 4156
rect 8484 4140 8536 4146
rect 8484 4082 8536 4088
rect 8496 3738 8524 4082
rect 8484 3732 8536 3738
rect 8484 3674 8536 3680
rect 8576 3732 8628 3738
rect 8576 3674 8628 3680
rect 8114 3632 8170 3641
rect 8588 3618 8616 3674
rect 8170 3590 8616 3618
rect 8114 3567 8170 3576
rect 8128 3534 8156 3567
rect 7656 3528 7708 3534
rect 8116 3528 8168 3534
rect 7708 3476 7788 3482
rect 7656 3470 7788 3476
rect 8208 3528 8260 3534
rect 8116 3470 8168 3476
rect 8206 3496 8208 3505
rect 8260 3496 8262 3505
rect 7668 3454 7788 3470
rect 7288 3392 7340 3398
rect 7288 3334 7340 3340
rect 7564 3392 7616 3398
rect 7564 3334 7616 3340
rect 6828 3188 6880 3194
rect 6828 3130 6880 3136
rect 7300 3058 7328 3334
rect 7760 3058 7788 3454
rect 8206 3431 8262 3440
rect 6736 3052 6788 3058
rect 6736 2994 6788 3000
rect 7196 3052 7248 3058
rect 7196 2994 7248 3000
rect 7288 3052 7340 3058
rect 7288 2994 7340 3000
rect 7748 3052 7800 3058
rect 7748 2994 7800 3000
rect 6000 2848 6052 2854
rect 6748 2825 6776 2994
rect 6000 2790 6052 2796
rect 6734 2816 6790 2825
rect 6734 2751 6790 2760
rect 7208 2650 7236 2994
rect 5816 2644 5868 2650
rect 5816 2586 5868 2592
rect 7196 2644 7248 2650
rect 7196 2586 7248 2592
rect 3884 2440 3936 2446
rect 3884 2382 3936 2388
rect 4712 2440 4764 2446
rect 4712 2382 4764 2388
rect 5172 2440 5224 2446
rect 5172 2382 5224 2388
rect 5264 2440 5316 2446
rect 5264 2382 5316 2388
rect 5448 2440 5500 2446
rect 5448 2382 5500 2388
rect 6552 2440 6604 2446
rect 6552 2382 6604 2388
rect 4724 2038 4752 2382
rect 6564 2310 6592 2382
rect 6552 2304 6604 2310
rect 6552 2246 6604 2252
rect 4712 2032 4764 2038
rect 4712 1974 4764 1980
rect 6564 1970 6592 2246
rect 6552 1964 6604 1970
rect 6552 1906 6604 1912
rect 8220 1902 8248 3431
rect 8772 3398 8800 7754
rect 8864 5914 8892 12582
rect 9232 10470 9260 13262
rect 9496 11552 9548 11558
rect 9496 11494 9548 11500
rect 9508 10674 9536 11494
rect 9876 10742 9904 13806
rect 10428 13530 10456 14282
rect 10416 13524 10468 13530
rect 10416 13466 10468 13472
rect 10324 13184 10376 13190
rect 10324 13126 10376 13132
rect 10140 12708 10192 12714
rect 10140 12650 10192 12656
rect 10152 11830 10180 12650
rect 10336 12434 10364 13126
rect 10336 12406 10456 12434
rect 10428 12170 10456 12406
rect 10416 12164 10468 12170
rect 10416 12106 10468 12112
rect 10140 11824 10192 11830
rect 10140 11766 10192 11772
rect 10520 11354 10548 14350
rect 11428 14272 11480 14278
rect 11428 14214 11480 14220
rect 11612 14272 11664 14278
rect 11612 14214 11664 14220
rect 11440 14074 11468 14214
rect 11428 14068 11480 14074
rect 11428 14010 11480 14016
rect 10600 13932 10652 13938
rect 10600 13874 10652 13880
rect 11152 13932 11204 13938
rect 11152 13874 11204 13880
rect 9956 11348 10008 11354
rect 9956 11290 10008 11296
rect 10508 11348 10560 11354
rect 10508 11290 10560 11296
rect 9864 10736 9916 10742
rect 9864 10678 9916 10684
rect 9496 10668 9548 10674
rect 9496 10610 9548 10616
rect 9220 10464 9272 10470
rect 9220 10406 9272 10412
rect 9036 9444 9088 9450
rect 9036 9386 9088 9392
rect 9048 8498 9076 9386
rect 9036 8492 9088 8498
rect 9036 8434 9088 8440
rect 9232 6798 9260 10406
rect 9312 9376 9364 9382
rect 9312 9318 9364 9324
rect 9324 8974 9352 9318
rect 9508 9042 9536 10610
rect 9496 9036 9548 9042
rect 9496 8978 9548 8984
rect 9312 8968 9364 8974
rect 9312 8910 9364 8916
rect 9324 8634 9352 8910
rect 9588 8832 9640 8838
rect 9588 8774 9640 8780
rect 9312 8628 9364 8634
rect 9312 8570 9364 8576
rect 9600 8090 9628 8774
rect 9680 8288 9732 8294
rect 9680 8230 9732 8236
rect 9588 8084 9640 8090
rect 9588 8026 9640 8032
rect 9692 7954 9720 8230
rect 9680 7948 9732 7954
rect 9680 7890 9732 7896
rect 9404 7880 9456 7886
rect 9402 7848 9404 7857
rect 9456 7848 9458 7857
rect 9402 7783 9458 7792
rect 9496 7404 9548 7410
rect 9496 7346 9548 7352
rect 9588 7404 9640 7410
rect 9588 7346 9640 7352
rect 9220 6792 9272 6798
rect 9220 6734 9272 6740
rect 9220 6656 9272 6662
rect 9220 6598 9272 6604
rect 9232 6322 9260 6598
rect 9220 6316 9272 6322
rect 9220 6258 9272 6264
rect 9220 6112 9272 6118
rect 9220 6054 9272 6060
rect 8852 5908 8904 5914
rect 8852 5850 8904 5856
rect 9036 5908 9088 5914
rect 9036 5850 9088 5856
rect 9048 5817 9076 5850
rect 9034 5808 9090 5817
rect 9034 5743 9090 5752
rect 9232 4146 9260 6054
rect 9508 5914 9536 7346
rect 9600 7177 9628 7346
rect 9586 7168 9642 7177
rect 9586 7103 9642 7112
rect 9496 5908 9548 5914
rect 9496 5850 9548 5856
rect 9494 5672 9550 5681
rect 9494 5607 9550 5616
rect 9508 4622 9536 5607
rect 9600 5302 9628 7103
rect 9864 6248 9916 6254
rect 9864 6190 9916 6196
rect 9680 6112 9732 6118
rect 9680 6054 9732 6060
rect 9692 5846 9720 6054
rect 9680 5840 9732 5846
rect 9680 5782 9732 5788
rect 9680 5704 9732 5710
rect 9680 5646 9732 5652
rect 9588 5296 9640 5302
rect 9588 5238 9640 5244
rect 9496 4616 9548 4622
rect 9494 4584 9496 4593
rect 9588 4616 9640 4622
rect 9548 4584 9550 4593
rect 9588 4558 9640 4564
rect 9494 4519 9550 4528
rect 9404 4480 9456 4486
rect 9404 4422 9456 4428
rect 9220 4140 9272 4146
rect 9220 4082 9272 4088
rect 9416 4010 9444 4422
rect 9600 4214 9628 4558
rect 9692 4486 9720 5646
rect 9876 5098 9904 6190
rect 9864 5092 9916 5098
rect 9864 5034 9916 5040
rect 9680 4480 9732 4486
rect 9680 4422 9732 4428
rect 9588 4208 9640 4214
rect 9588 4150 9640 4156
rect 9404 4004 9456 4010
rect 9404 3946 9456 3952
rect 8942 3768 8998 3777
rect 8942 3703 8998 3712
rect 8956 3534 8984 3703
rect 9600 3602 9628 4150
rect 9772 3936 9824 3942
rect 9772 3878 9824 3884
rect 9784 3670 9812 3878
rect 9772 3664 9824 3670
rect 9772 3606 9824 3612
rect 9588 3596 9640 3602
rect 9588 3538 9640 3544
rect 8944 3528 8996 3534
rect 8944 3470 8996 3476
rect 8760 3392 8812 3398
rect 8760 3334 8812 3340
rect 9600 3210 9628 3538
rect 9678 3496 9734 3505
rect 9678 3431 9734 3440
rect 9692 3398 9720 3431
rect 9680 3392 9732 3398
rect 9680 3334 9732 3340
rect 9416 3182 9628 3210
rect 9416 3126 9444 3182
rect 9784 3126 9812 3606
rect 9404 3120 9456 3126
rect 9404 3062 9456 3068
rect 9772 3120 9824 3126
rect 9772 3062 9824 3068
rect 8576 3052 8628 3058
rect 8576 2994 8628 3000
rect 8588 2854 8616 2994
rect 8576 2848 8628 2854
rect 8576 2790 8628 2796
rect 9968 2446 9996 11290
rect 10612 10810 10640 13874
rect 10876 13864 10928 13870
rect 10796 13812 10876 13814
rect 10796 13806 10928 13812
rect 10796 13802 10916 13806
rect 10784 13796 10916 13802
rect 10836 13786 10916 13796
rect 10784 13738 10836 13744
rect 10796 13462 10824 13738
rect 10784 13456 10836 13462
rect 10784 13398 10836 13404
rect 11164 13326 11192 13874
rect 11520 13864 11572 13870
rect 11520 13806 11572 13812
rect 11532 13530 11560 13806
rect 11520 13524 11572 13530
rect 11520 13466 11572 13472
rect 11152 13320 11204 13326
rect 10805 13314 10857 13320
rect 10796 13262 10805 13308
rect 11152 13262 11204 13268
rect 10796 13256 10857 13262
rect 10796 12986 10824 13256
rect 11428 13184 11480 13190
rect 11428 13126 11480 13132
rect 10784 12980 10836 12986
rect 10784 12922 10836 12928
rect 11440 12102 11468 13126
rect 11428 12096 11480 12102
rect 11428 12038 11480 12044
rect 10692 11076 10744 11082
rect 10692 11018 10744 11024
rect 10600 10804 10652 10810
rect 10600 10746 10652 10752
rect 10140 8900 10192 8906
rect 10140 8842 10192 8848
rect 10152 8634 10180 8842
rect 10416 8832 10468 8838
rect 10416 8774 10468 8780
rect 10140 8628 10192 8634
rect 10140 8570 10192 8576
rect 10428 8498 10456 8774
rect 10416 8492 10468 8498
rect 10416 8434 10468 8440
rect 10324 8424 10376 8430
rect 10324 8366 10376 8372
rect 10048 8288 10100 8294
rect 10048 8230 10100 8236
rect 10060 7410 10088 8230
rect 10232 7744 10284 7750
rect 10232 7686 10284 7692
rect 10244 7410 10272 7686
rect 10336 7546 10364 8366
rect 10324 7540 10376 7546
rect 10324 7482 10376 7488
rect 10048 7404 10100 7410
rect 10048 7346 10100 7352
rect 10232 7404 10284 7410
rect 10232 7346 10284 7352
rect 10324 7268 10376 7274
rect 10324 7210 10376 7216
rect 10140 6792 10192 6798
rect 10140 6734 10192 6740
rect 10048 6724 10100 6730
rect 10048 6666 10100 6672
rect 10060 6458 10088 6666
rect 10048 6452 10100 6458
rect 10048 6394 10100 6400
rect 10048 6316 10100 6322
rect 10048 6258 10100 6264
rect 10060 5370 10088 6258
rect 10152 5710 10180 6734
rect 10232 6452 10284 6458
rect 10232 6394 10284 6400
rect 10140 5704 10192 5710
rect 10140 5646 10192 5652
rect 10048 5364 10100 5370
rect 10048 5306 10100 5312
rect 10152 4078 10180 5646
rect 10140 4072 10192 4078
rect 10140 4014 10192 4020
rect 10244 2961 10272 6394
rect 10336 5030 10364 7210
rect 10428 5234 10456 8434
rect 10508 7812 10560 7818
rect 10508 7754 10560 7760
rect 10520 7002 10548 7754
rect 10508 6996 10560 7002
rect 10508 6938 10560 6944
rect 10704 6662 10732 11018
rect 11244 9920 11296 9926
rect 11244 9862 11296 9868
rect 10784 8492 10836 8498
rect 10784 8434 10836 8440
rect 10796 8294 10824 8434
rect 10876 8424 10928 8430
rect 10876 8366 10928 8372
rect 10784 8288 10836 8294
rect 10784 8230 10836 8236
rect 10796 7478 10824 8230
rect 10888 8090 10916 8366
rect 10876 8084 10928 8090
rect 10876 8026 10928 8032
rect 10784 7472 10836 7478
rect 10784 7414 10836 7420
rect 11060 7200 11112 7206
rect 11060 7142 11112 7148
rect 10784 6860 10836 6866
rect 10784 6802 10836 6808
rect 10600 6656 10652 6662
rect 10600 6598 10652 6604
rect 10692 6656 10744 6662
rect 10692 6598 10744 6604
rect 10612 6390 10640 6598
rect 10796 6474 10824 6802
rect 10704 6446 10824 6474
rect 10600 6384 10652 6390
rect 10600 6326 10652 6332
rect 10704 6322 10732 6446
rect 10692 6316 10744 6322
rect 10692 6258 10744 6264
rect 10784 5704 10836 5710
rect 10784 5646 10836 5652
rect 10416 5228 10468 5234
rect 10416 5170 10468 5176
rect 10324 5024 10376 5030
rect 10324 4966 10376 4972
rect 10796 4622 10824 5646
rect 11072 5642 11100 7142
rect 11256 6798 11284 9862
rect 11334 6896 11390 6905
rect 11334 6831 11390 6840
rect 11244 6792 11296 6798
rect 11244 6734 11296 6740
rect 11256 5681 11284 6734
rect 11348 6662 11376 6831
rect 11336 6656 11388 6662
rect 11336 6598 11388 6604
rect 11242 5672 11298 5681
rect 11060 5636 11112 5642
rect 11242 5607 11298 5616
rect 11060 5578 11112 5584
rect 10784 4616 10836 4622
rect 10784 4558 10836 4564
rect 10876 4208 10928 4214
rect 10876 4150 10928 4156
rect 10888 3534 10916 4150
rect 10876 3528 10928 3534
rect 10876 3470 10928 3476
rect 10230 2952 10286 2961
rect 10230 2887 10286 2896
rect 10876 2848 10928 2854
rect 10876 2790 10928 2796
rect 9956 2440 10008 2446
rect 9956 2382 10008 2388
rect 10888 2378 10916 2790
rect 11440 2774 11468 12038
rect 11532 9466 11560 13466
rect 11624 11150 11652 14214
rect 11716 13802 11744 14418
rect 12440 14408 12492 14414
rect 12440 14350 12492 14356
rect 15200 14408 15252 14414
rect 15200 14350 15252 14356
rect 16856 14408 16908 14414
rect 16856 14350 16908 14356
rect 12452 13938 12480 14350
rect 15016 14272 15068 14278
rect 15016 14214 15068 14220
rect 14740 14068 14792 14074
rect 14740 14010 14792 14016
rect 12900 14000 12952 14006
rect 12900 13942 12952 13948
rect 12440 13932 12492 13938
rect 12440 13874 12492 13880
rect 12716 13864 12768 13870
rect 12716 13806 12768 13812
rect 11704 13796 11756 13802
rect 11704 13738 11756 13744
rect 12164 13796 12216 13802
rect 12164 13738 12216 13744
rect 11716 13705 11744 13738
rect 11702 13696 11758 13705
rect 11702 13631 11758 13640
rect 11704 12232 11756 12238
rect 11704 12174 11756 12180
rect 11716 11694 11744 12174
rect 11704 11688 11756 11694
rect 11704 11630 11756 11636
rect 11716 11218 11744 11630
rect 12176 11354 12204 13738
rect 12728 13530 12756 13806
rect 12912 13705 12940 13942
rect 13084 13932 13136 13938
rect 13084 13874 13136 13880
rect 13096 13814 13124 13874
rect 14752 13870 14780 14010
rect 13728 13864 13780 13870
rect 13096 13786 13216 13814
rect 13728 13806 13780 13812
rect 14740 13864 14792 13870
rect 14740 13806 14792 13812
rect 13084 13728 13136 13734
rect 12898 13696 12954 13705
rect 13084 13670 13136 13676
rect 12898 13631 12954 13640
rect 12716 13524 12768 13530
rect 12716 13466 12768 13472
rect 12912 13462 12940 13631
rect 12900 13456 12952 13462
rect 12900 13398 12952 13404
rect 13096 13394 13124 13670
rect 13084 13388 13136 13394
rect 13084 13330 13136 13336
rect 13188 13326 13216 13786
rect 13176 13320 13228 13326
rect 13176 13262 13228 13268
rect 12532 13184 12584 13190
rect 12532 13126 12584 13132
rect 13268 13184 13320 13190
rect 13268 13126 13320 13132
rect 12544 12238 12572 13126
rect 12532 12232 12584 12238
rect 12532 12174 12584 12180
rect 13280 12102 13308 13126
rect 13544 12844 13596 12850
rect 13544 12786 13596 12792
rect 13268 12096 13320 12102
rect 13268 12038 13320 12044
rect 12716 11892 12768 11898
rect 12716 11834 12768 11840
rect 12164 11348 12216 11354
rect 12164 11290 12216 11296
rect 11704 11212 11756 11218
rect 11704 11154 11756 11160
rect 11612 11144 11664 11150
rect 11612 11086 11664 11092
rect 12176 9674 12204 11290
rect 12440 9920 12492 9926
rect 12440 9862 12492 9868
rect 11992 9646 12204 9674
rect 11532 9438 11928 9466
rect 11520 9376 11572 9382
rect 11520 9318 11572 9324
rect 11532 6798 11560 9318
rect 11612 8492 11664 8498
rect 11612 8434 11664 8440
rect 11624 8378 11652 8434
rect 11796 8424 11848 8430
rect 11624 8350 11744 8378
rect 11796 8366 11848 8372
rect 11612 8288 11664 8294
rect 11612 8230 11664 8236
rect 11624 8090 11652 8230
rect 11612 8084 11664 8090
rect 11612 8026 11664 8032
rect 11716 7818 11744 8350
rect 11808 7954 11836 8366
rect 11796 7948 11848 7954
rect 11796 7890 11848 7896
rect 11900 7834 11928 9438
rect 11704 7812 11756 7818
rect 11704 7754 11756 7760
rect 11808 7806 11928 7834
rect 11704 7540 11756 7546
rect 11704 7482 11756 7488
rect 11716 7274 11744 7482
rect 11704 7268 11756 7274
rect 11704 7210 11756 7216
rect 11520 6792 11572 6798
rect 11520 6734 11572 6740
rect 11532 5914 11560 6734
rect 11716 6322 11744 7210
rect 11612 6316 11664 6322
rect 11612 6258 11664 6264
rect 11704 6316 11756 6322
rect 11704 6258 11756 6264
rect 11624 6225 11652 6258
rect 11610 6216 11666 6225
rect 11610 6151 11666 6160
rect 11624 6118 11652 6151
rect 11612 6112 11664 6118
rect 11612 6054 11664 6060
rect 11520 5908 11572 5914
rect 11520 5850 11572 5856
rect 11612 5568 11664 5574
rect 11612 5510 11664 5516
rect 11624 5030 11652 5510
rect 11808 5370 11836 7806
rect 11888 7744 11940 7750
rect 11888 7686 11940 7692
rect 11900 7478 11928 7686
rect 11888 7472 11940 7478
rect 11888 7414 11940 7420
rect 11888 7200 11940 7206
rect 11888 7142 11940 7148
rect 11796 5364 11848 5370
rect 11796 5306 11848 5312
rect 11808 5273 11836 5306
rect 11794 5264 11850 5273
rect 11704 5228 11756 5234
rect 11794 5199 11850 5208
rect 11704 5170 11756 5176
rect 11612 5024 11664 5030
rect 11612 4966 11664 4972
rect 11624 4690 11652 4966
rect 11612 4684 11664 4690
rect 11612 4626 11664 4632
rect 11716 4622 11744 5170
rect 11704 4616 11756 4622
rect 11704 4558 11756 4564
rect 11808 4282 11836 5199
rect 11796 4276 11848 4282
rect 11796 4218 11848 4224
rect 11796 4004 11848 4010
rect 11796 3946 11848 3952
rect 11808 3398 11836 3946
rect 11704 3392 11756 3398
rect 11702 3360 11704 3369
rect 11796 3392 11848 3398
rect 11756 3360 11758 3369
rect 11796 3334 11848 3340
rect 11702 3295 11758 3304
rect 11900 3126 11928 7142
rect 11888 3120 11940 3126
rect 11888 3062 11940 3068
rect 11992 2774 12020 9646
rect 12348 8832 12400 8838
rect 12348 8774 12400 8780
rect 12256 8492 12308 8498
rect 12256 8434 12308 8440
rect 12164 7268 12216 7274
rect 12164 7210 12216 7216
rect 12070 6760 12126 6769
rect 12070 6695 12126 6704
rect 12084 6662 12112 6695
rect 12072 6656 12124 6662
rect 12072 6598 12124 6604
rect 12176 6390 12204 7210
rect 12164 6384 12216 6390
rect 12164 6326 12216 6332
rect 12268 6186 12296 8434
rect 12360 7206 12388 8774
rect 12452 7546 12480 9862
rect 12624 9512 12676 9518
rect 12624 9454 12676 9460
rect 12532 9036 12584 9042
rect 12532 8978 12584 8984
rect 12544 8498 12572 8978
rect 12532 8492 12584 8498
rect 12532 8434 12584 8440
rect 12544 7886 12572 8434
rect 12636 8294 12664 9454
rect 12728 8974 12756 11834
rect 12992 10464 13044 10470
rect 12992 10406 13044 10412
rect 12900 9648 12952 9654
rect 12900 9590 12952 9596
rect 12808 9580 12860 9586
rect 12808 9522 12860 9528
rect 12820 9178 12848 9522
rect 12808 9172 12860 9178
rect 12808 9114 12860 9120
rect 12716 8968 12768 8974
rect 12716 8910 12768 8916
rect 12912 8634 12940 9590
rect 12900 8628 12952 8634
rect 12900 8570 12952 8576
rect 12624 8288 12676 8294
rect 12624 8230 12676 8236
rect 12808 8288 12860 8294
rect 12808 8230 12860 8236
rect 12820 7954 12848 8230
rect 12808 7948 12860 7954
rect 12808 7890 12860 7896
rect 12532 7880 12584 7886
rect 12532 7822 12584 7828
rect 12440 7540 12492 7546
rect 12440 7482 12492 7488
rect 12820 7478 12848 7890
rect 12808 7472 12860 7478
rect 12808 7414 12860 7420
rect 12716 7404 12768 7410
rect 12716 7346 12768 7352
rect 12728 7274 12756 7346
rect 12716 7268 12768 7274
rect 12768 7228 12848 7256
rect 12716 7210 12768 7216
rect 12348 7200 12400 7206
rect 12348 7142 12400 7148
rect 12256 6180 12308 6186
rect 12256 6122 12308 6128
rect 12072 6112 12124 6118
rect 12072 6054 12124 6060
rect 12084 5778 12112 6054
rect 12072 5772 12124 5778
rect 12072 5714 12124 5720
rect 12072 5636 12124 5642
rect 12072 5578 12124 5584
rect 12084 5302 12112 5578
rect 12164 5364 12216 5370
rect 12164 5306 12216 5312
rect 12072 5296 12124 5302
rect 12072 5238 12124 5244
rect 12176 5098 12204 5306
rect 12164 5092 12216 5098
rect 12164 5034 12216 5040
rect 12070 4856 12126 4865
rect 12176 4826 12204 5034
rect 12256 5024 12308 5030
rect 12256 4966 12308 4972
rect 12070 4791 12072 4800
rect 12124 4791 12126 4800
rect 12164 4820 12216 4826
rect 12072 4762 12124 4768
rect 12164 4762 12216 4768
rect 12268 4146 12296 4966
rect 12072 4140 12124 4146
rect 12072 4082 12124 4088
rect 12256 4140 12308 4146
rect 12256 4082 12308 4088
rect 12084 3738 12112 4082
rect 12164 4072 12216 4078
rect 12164 4014 12216 4020
rect 12072 3732 12124 3738
rect 12072 3674 12124 3680
rect 12176 3058 12204 4014
rect 12256 4004 12308 4010
rect 12256 3946 12308 3952
rect 12268 3534 12296 3946
rect 12256 3528 12308 3534
rect 12256 3470 12308 3476
rect 12164 3052 12216 3058
rect 12164 2994 12216 3000
rect 12164 2848 12216 2854
rect 12164 2790 12216 2796
rect 11348 2746 11468 2774
rect 11716 2746 12020 2774
rect 11348 2514 11376 2746
rect 11336 2508 11388 2514
rect 11336 2450 11388 2456
rect 11716 2446 11744 2746
rect 11704 2440 11756 2446
rect 11704 2382 11756 2388
rect 10876 2372 10928 2378
rect 10876 2314 10928 2320
rect 10048 2304 10100 2310
rect 10048 2246 10100 2252
rect 10784 2304 10836 2310
rect 10784 2246 10836 2252
rect 8208 1896 8260 1902
rect 8208 1838 8260 1844
rect 10060 1834 10088 2246
rect 10796 2106 10824 2246
rect 10784 2100 10836 2106
rect 10784 2042 10836 2048
rect 10048 1828 10100 1834
rect 10048 1770 10100 1776
rect 12176 1494 12204 2790
rect 12164 1488 12216 1494
rect 12164 1430 12216 1436
rect 12360 800 12388 7142
rect 12532 6928 12584 6934
rect 12532 6870 12584 6876
rect 12544 6458 12572 6870
rect 12820 6458 12848 7228
rect 12900 7200 12952 7206
rect 12900 7142 12952 7148
rect 12532 6452 12584 6458
rect 12532 6394 12584 6400
rect 12808 6452 12860 6458
rect 12808 6394 12860 6400
rect 12912 6390 12940 7142
rect 12716 6384 12768 6390
rect 12716 6326 12768 6332
rect 12900 6384 12952 6390
rect 12900 6326 12952 6332
rect 12624 6180 12676 6186
rect 12624 6122 12676 6128
rect 12440 5160 12492 5166
rect 12440 5102 12492 5108
rect 12452 4282 12480 5102
rect 12532 5024 12584 5030
rect 12532 4966 12584 4972
rect 12544 4554 12572 4966
rect 12532 4548 12584 4554
rect 12532 4490 12584 4496
rect 12530 4448 12586 4457
rect 12530 4383 12586 4392
rect 12440 4276 12492 4282
rect 12440 4218 12492 4224
rect 12438 4176 12494 4185
rect 12438 4111 12494 4120
rect 12452 800 12480 4111
rect 12544 800 12572 4383
rect 12636 800 12664 6122
rect 12728 800 12756 6326
rect 12808 6316 12860 6322
rect 12808 6258 12860 6264
rect 12820 6089 12848 6258
rect 12900 6248 12952 6254
rect 12900 6190 12952 6196
rect 12806 6080 12862 6089
rect 12806 6015 12862 6024
rect 12912 5710 12940 6190
rect 13004 5710 13032 10406
rect 13084 9920 13136 9926
rect 13084 9862 13136 9868
rect 13096 6730 13124 9862
rect 13176 8900 13228 8906
rect 13176 8842 13228 8848
rect 13188 8634 13216 8842
rect 13176 8628 13228 8634
rect 13176 8570 13228 8576
rect 13176 8492 13228 8498
rect 13176 8434 13228 8440
rect 13084 6724 13136 6730
rect 13084 6666 13136 6672
rect 12900 5704 12952 5710
rect 12900 5646 12952 5652
rect 12992 5704 13044 5710
rect 12992 5646 13044 5652
rect 12808 5228 12860 5234
rect 12808 5170 12860 5176
rect 12820 4486 12848 5170
rect 12808 4480 12860 4486
rect 12808 4422 12860 4428
rect 12820 2446 12848 4422
rect 12912 4146 12940 5646
rect 13084 5568 13136 5574
rect 13084 5510 13136 5516
rect 12992 5228 13044 5234
rect 12992 5170 13044 5176
rect 13004 4826 13032 5170
rect 12992 4820 13044 4826
rect 12992 4762 13044 4768
rect 12990 4312 13046 4321
rect 12990 4247 13046 4256
rect 12900 4140 12952 4146
rect 12900 4082 12952 4088
rect 12898 3360 12954 3369
rect 12898 3295 12954 3304
rect 12912 2854 12940 3295
rect 12900 2848 12952 2854
rect 12900 2790 12952 2796
rect 12808 2440 12860 2446
rect 12808 2382 12860 2388
rect 12808 1964 12860 1970
rect 12808 1906 12860 1912
rect 12820 800 12848 1906
rect 13004 800 13032 4247
rect 13096 800 13124 5510
rect 13188 800 13216 8434
rect 13280 4622 13308 12038
rect 13556 11762 13584 12786
rect 13544 11756 13596 11762
rect 13544 11698 13596 11704
rect 13556 11218 13584 11698
rect 13544 11212 13596 11218
rect 13544 11154 13596 11160
rect 13556 10742 13584 11154
rect 13740 11150 13768 13806
rect 14924 13184 14976 13190
rect 14924 13126 14976 13132
rect 14648 12232 14700 12238
rect 14648 12174 14700 12180
rect 14660 11762 14688 12174
rect 14936 11830 14964 13126
rect 15028 12918 15056 14214
rect 15016 12912 15068 12918
rect 15016 12854 15068 12860
rect 15212 12646 15240 14350
rect 16304 14340 16356 14346
rect 16304 14282 16356 14288
rect 15660 14272 15712 14278
rect 15660 14214 15712 14220
rect 15672 13394 15700 14214
rect 15660 13388 15712 13394
rect 15660 13330 15712 13336
rect 15292 13320 15344 13326
rect 15292 13262 15344 13268
rect 15200 12640 15252 12646
rect 15200 12582 15252 12588
rect 14924 11824 14976 11830
rect 14924 11766 14976 11772
rect 14648 11756 14700 11762
rect 14648 11698 14700 11704
rect 15304 11558 15332 13262
rect 15672 12986 15700 13330
rect 16212 13184 16264 13190
rect 16212 13126 16264 13132
rect 15660 12980 15712 12986
rect 15660 12922 15712 12928
rect 15292 11552 15344 11558
rect 15292 11494 15344 11500
rect 13728 11144 13780 11150
rect 13728 11086 13780 11092
rect 13544 10736 13596 10742
rect 13544 10678 13596 10684
rect 15672 10538 15700 12922
rect 16120 12776 16172 12782
rect 16120 12718 16172 12724
rect 16132 11898 16160 12718
rect 16120 11892 16172 11898
rect 16120 11834 16172 11840
rect 16028 11552 16080 11558
rect 16028 11494 16080 11500
rect 16040 11082 16068 11494
rect 16028 11076 16080 11082
rect 16028 11018 16080 11024
rect 15660 10532 15712 10538
rect 15660 10474 15712 10480
rect 16224 9994 16252 13126
rect 16212 9988 16264 9994
rect 16212 9930 16264 9936
rect 14188 9920 14240 9926
rect 14188 9862 14240 9868
rect 14740 9920 14792 9926
rect 14740 9862 14792 9868
rect 15568 9920 15620 9926
rect 15568 9862 15620 9868
rect 13452 9376 13504 9382
rect 13452 9318 13504 9324
rect 13464 8498 13492 9318
rect 13544 8560 13596 8566
rect 13544 8502 13596 8508
rect 13452 8492 13504 8498
rect 13452 8434 13504 8440
rect 13556 8090 13584 8502
rect 13634 8392 13690 8401
rect 13634 8327 13636 8336
rect 13688 8327 13690 8336
rect 13636 8298 13688 8304
rect 13360 8084 13412 8090
rect 13360 8026 13412 8032
rect 13544 8084 13596 8090
rect 13544 8026 13596 8032
rect 13372 7002 13400 8026
rect 13360 6996 13412 7002
rect 13360 6938 13412 6944
rect 13544 6792 13596 6798
rect 13544 6734 13596 6740
rect 14096 6792 14148 6798
rect 14096 6734 14148 6740
rect 13556 6390 13584 6734
rect 13820 6656 13872 6662
rect 13820 6598 13872 6604
rect 13912 6656 13964 6662
rect 13912 6598 13964 6604
rect 13544 6384 13596 6390
rect 13544 6326 13596 6332
rect 13728 6316 13780 6322
rect 13728 6258 13780 6264
rect 13636 6112 13688 6118
rect 13634 6080 13636 6089
rect 13688 6080 13690 6089
rect 13634 6015 13690 6024
rect 13360 5908 13412 5914
rect 13360 5850 13412 5856
rect 13268 4616 13320 4622
rect 13268 4558 13320 4564
rect 13266 3632 13322 3641
rect 13266 3567 13268 3576
rect 13320 3567 13322 3576
rect 13268 3538 13320 3544
rect 13372 800 13400 5850
rect 13740 5574 13768 6258
rect 13832 5914 13860 6598
rect 13820 5908 13872 5914
rect 13820 5850 13872 5856
rect 13728 5568 13780 5574
rect 13728 5510 13780 5516
rect 13634 5264 13690 5273
rect 13634 5199 13636 5208
rect 13688 5199 13690 5208
rect 13636 5170 13688 5176
rect 13544 5160 13596 5166
rect 13544 5102 13596 5108
rect 13556 3738 13584 5102
rect 13740 4690 13768 5510
rect 13728 4684 13780 4690
rect 13728 4626 13780 4632
rect 13924 4570 13952 6598
rect 14108 6458 14136 6734
rect 14096 6452 14148 6458
rect 14096 6394 14148 6400
rect 14200 6390 14228 9862
rect 14280 8356 14332 8362
rect 14280 8298 14332 8304
rect 14292 7886 14320 8298
rect 14280 7880 14332 7886
rect 14280 7822 14332 7828
rect 14292 6866 14320 7822
rect 14752 7818 14780 9862
rect 15580 9518 15608 9862
rect 15568 9512 15620 9518
rect 15568 9454 15620 9460
rect 15200 9376 15252 9382
rect 15200 9318 15252 9324
rect 15108 8628 15160 8634
rect 15108 8570 15160 8576
rect 15014 7848 15070 7857
rect 14740 7812 14792 7818
rect 15014 7783 15070 7792
rect 14740 7754 14792 7760
rect 15028 7750 15056 7783
rect 14372 7744 14424 7750
rect 14372 7686 14424 7692
rect 15016 7744 15068 7750
rect 15016 7686 15068 7692
rect 14280 6860 14332 6866
rect 14280 6802 14332 6808
rect 14188 6384 14240 6390
rect 14188 6326 14240 6332
rect 14186 5808 14242 5817
rect 14096 5772 14148 5778
rect 14292 5778 14320 6802
rect 14186 5743 14242 5752
rect 14280 5772 14332 5778
rect 14096 5714 14148 5720
rect 14108 4826 14136 5714
rect 14200 5710 14228 5743
rect 14280 5714 14332 5720
rect 14188 5704 14240 5710
rect 14188 5646 14240 5652
rect 14096 4820 14148 4826
rect 14096 4762 14148 4768
rect 14384 4729 14412 7686
rect 14648 7200 14700 7206
rect 14646 7168 14648 7177
rect 14700 7168 14702 7177
rect 14646 7103 14702 7112
rect 14924 6996 14976 7002
rect 14924 6938 14976 6944
rect 14740 6724 14792 6730
rect 14740 6666 14792 6672
rect 14556 5296 14608 5302
rect 14556 5238 14608 5244
rect 14370 4720 14426 4729
rect 14370 4655 14426 4664
rect 14568 4622 14596 5238
rect 13648 4542 13952 4570
rect 14556 4616 14608 4622
rect 14556 4558 14608 4564
rect 13544 3732 13596 3738
rect 13544 3674 13596 3680
rect 13556 3233 13584 3674
rect 13542 3224 13598 3233
rect 13542 3159 13598 3168
rect 13556 3058 13584 3159
rect 13648 3058 13676 4542
rect 13820 4480 13872 4486
rect 13820 4422 13872 4428
rect 13728 4140 13780 4146
rect 13728 4082 13780 4088
rect 13740 3194 13768 4082
rect 13728 3188 13780 3194
rect 13728 3130 13780 3136
rect 13726 3088 13782 3097
rect 13544 3052 13596 3058
rect 13544 2994 13596 3000
rect 13636 3052 13688 3058
rect 13726 3023 13782 3032
rect 13636 2994 13688 3000
rect 13452 2644 13504 2650
rect 13452 2586 13504 2592
rect 13464 800 13492 2586
rect 13740 800 13768 3023
rect 13832 800 13860 4422
rect 14096 3596 14148 3602
rect 14096 3538 14148 3544
rect 14108 3194 14136 3538
rect 14096 3188 14148 3194
rect 14096 3130 14148 3136
rect 14372 2848 14424 2854
rect 14372 2790 14424 2796
rect 14462 2816 14518 2825
rect 14384 2446 14412 2790
rect 14462 2751 14518 2760
rect 14372 2440 14424 2446
rect 14372 2382 14424 2388
rect 14096 2032 14148 2038
rect 14096 1974 14148 1980
rect 14108 800 14136 1974
rect 14188 1828 14240 1834
rect 14188 1770 14240 1776
rect 14200 800 14228 1770
rect 14476 800 14504 2751
rect 14556 2100 14608 2106
rect 14556 2042 14608 2048
rect 14568 800 14596 2042
rect 14752 800 14780 6666
rect 14936 6118 14964 6938
rect 15016 6792 15068 6798
rect 15016 6734 15068 6740
rect 15028 6322 15056 6734
rect 15120 6322 15148 8570
rect 15212 7886 15240 9318
rect 15476 8832 15528 8838
rect 15476 8774 15528 8780
rect 15488 8634 15516 8774
rect 15476 8628 15528 8634
rect 15476 8570 15528 8576
rect 16120 8424 16172 8430
rect 16120 8366 16172 8372
rect 15476 8016 15528 8022
rect 15476 7958 15528 7964
rect 15200 7880 15252 7886
rect 15200 7822 15252 7828
rect 15384 7812 15436 7818
rect 15384 7754 15436 7760
rect 15200 7744 15252 7750
rect 15200 7686 15252 7692
rect 15016 6316 15068 6322
rect 15016 6258 15068 6264
rect 15108 6316 15160 6322
rect 15108 6258 15160 6264
rect 14924 6112 14976 6118
rect 14924 6054 14976 6060
rect 14936 5914 14964 6054
rect 14832 5908 14884 5914
rect 14832 5850 14884 5856
rect 14924 5908 14976 5914
rect 14924 5850 14976 5856
rect 14844 5250 14872 5850
rect 14936 5370 14964 5850
rect 14924 5364 14976 5370
rect 14924 5306 14976 5312
rect 14844 5222 15056 5250
rect 14832 1488 14884 1494
rect 14832 1430 14884 1436
rect 14844 800 14872 1430
rect 15028 800 15056 5222
rect 15212 4622 15240 7686
rect 15292 6180 15344 6186
rect 15292 6122 15344 6128
rect 15304 5846 15332 6122
rect 15292 5840 15344 5846
rect 15292 5782 15344 5788
rect 15292 5024 15344 5030
rect 15292 4966 15344 4972
rect 15304 4826 15332 4966
rect 15292 4820 15344 4826
rect 15292 4762 15344 4768
rect 15200 4616 15252 4622
rect 15106 4584 15162 4593
rect 15200 4558 15252 4564
rect 15106 4519 15162 4528
rect 15120 3194 15148 4519
rect 15290 3632 15346 3641
rect 15290 3567 15346 3576
rect 15304 3534 15332 3567
rect 15292 3528 15344 3534
rect 15292 3470 15344 3476
rect 15200 3460 15252 3466
rect 15200 3402 15252 3408
rect 15108 3188 15160 3194
rect 15108 3130 15160 3136
rect 15108 2508 15160 2514
rect 15108 2450 15160 2456
rect 15120 800 15148 2450
rect 15212 1442 15240 3402
rect 15292 2848 15344 2854
rect 15292 2790 15344 2796
rect 15304 2650 15332 2790
rect 15396 2774 15424 7754
rect 15488 7002 15516 7958
rect 16028 7880 16080 7886
rect 16028 7822 16080 7828
rect 15660 7812 15712 7818
rect 15660 7754 15712 7760
rect 15672 7206 15700 7754
rect 15936 7404 15988 7410
rect 15936 7346 15988 7352
rect 15660 7200 15712 7206
rect 15660 7142 15712 7148
rect 15476 6996 15528 7002
rect 15476 6938 15528 6944
rect 15568 6112 15620 6118
rect 15568 6054 15620 6060
rect 15580 5234 15608 6054
rect 15672 5710 15700 7142
rect 15948 6866 15976 7346
rect 15936 6860 15988 6866
rect 15936 6802 15988 6808
rect 15752 6792 15804 6798
rect 15752 6734 15804 6740
rect 15764 5914 15792 6734
rect 15752 5908 15804 5914
rect 15752 5850 15804 5856
rect 15660 5704 15712 5710
rect 15660 5646 15712 5652
rect 15568 5228 15620 5234
rect 15568 5170 15620 5176
rect 15476 5160 15528 5166
rect 15476 5102 15528 5108
rect 15488 4690 15516 5102
rect 15476 4684 15528 4690
rect 15476 4626 15528 4632
rect 15764 4010 15792 5850
rect 15844 5568 15896 5574
rect 15844 5510 15896 5516
rect 15752 4004 15804 4010
rect 15752 3946 15804 3952
rect 15752 3732 15804 3738
rect 15752 3674 15804 3680
rect 15568 3664 15620 3670
rect 15568 3606 15620 3612
rect 15476 3528 15528 3534
rect 15476 3470 15528 3476
rect 15488 3233 15516 3470
rect 15474 3224 15530 3233
rect 15474 3159 15530 3168
rect 15488 3058 15516 3159
rect 15580 3074 15608 3606
rect 15476 3052 15528 3058
rect 15580 3046 15700 3074
rect 15476 2994 15528 3000
rect 15396 2746 15608 2774
rect 15292 2644 15344 2650
rect 15292 2586 15344 2592
rect 15384 2576 15436 2582
rect 15384 2518 15436 2524
rect 15292 2440 15344 2446
rect 15292 2382 15344 2388
rect 15304 1562 15332 2382
rect 15292 1556 15344 1562
rect 15292 1498 15344 1504
rect 15212 1414 15332 1442
rect 15304 800 15332 1414
rect 15396 800 15424 2518
rect 15580 800 15608 2746
rect 15672 800 15700 3046
rect 15764 2774 15792 3674
rect 15856 3534 15884 5510
rect 15934 4856 15990 4865
rect 15934 4791 15936 4800
rect 15988 4791 15990 4800
rect 15936 4762 15988 4768
rect 15936 3936 15988 3942
rect 15936 3878 15988 3884
rect 15844 3528 15896 3534
rect 15844 3470 15896 3476
rect 15764 2746 15884 2774
rect 15856 800 15884 2746
rect 15948 800 15976 3878
rect 16040 2774 16068 7822
rect 16132 6866 16160 8366
rect 16120 6860 16172 6866
rect 16120 6802 16172 6808
rect 16132 5914 16160 6802
rect 16120 5908 16172 5914
rect 16120 5850 16172 5856
rect 16316 4486 16344 14282
rect 16868 13462 16896 14350
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 50294 14172 50602 14181
rect 50294 14170 50300 14172
rect 50356 14170 50380 14172
rect 50436 14170 50460 14172
rect 50516 14170 50540 14172
rect 50596 14170 50602 14172
rect 50356 14118 50358 14170
rect 50538 14118 50540 14170
rect 50294 14116 50300 14118
rect 50356 14116 50380 14118
rect 50436 14116 50460 14118
rect 50516 14116 50540 14118
rect 50596 14116 50602 14118
rect 50294 14107 50602 14116
rect 21548 13864 21600 13870
rect 21548 13806 21600 13812
rect 16856 13456 16908 13462
rect 16856 13398 16908 13404
rect 16868 13326 16896 13398
rect 16396 13320 16448 13326
rect 16672 13320 16724 13326
rect 16448 13280 16528 13308
rect 16396 13262 16448 13268
rect 16396 13184 16448 13190
rect 16396 13126 16448 13132
rect 16408 5370 16436 13126
rect 16500 10266 16528 13280
rect 16672 13262 16724 13268
rect 16856 13320 16908 13326
rect 16856 13262 16908 13268
rect 17316 13320 17368 13326
rect 17316 13262 17368 13268
rect 16580 13184 16632 13190
rect 16580 13126 16632 13132
rect 16592 12986 16620 13126
rect 16580 12980 16632 12986
rect 16580 12922 16632 12928
rect 16684 11529 16712 13262
rect 16948 12232 17000 12238
rect 16948 12174 17000 12180
rect 16960 12102 16988 12174
rect 16856 12096 16908 12102
rect 16856 12038 16908 12044
rect 16948 12096 17000 12102
rect 16948 12038 17000 12044
rect 16868 11830 16896 12038
rect 16856 11824 16908 11830
rect 16856 11766 16908 11772
rect 16670 11520 16726 11529
rect 16670 11455 16726 11464
rect 17328 10674 17356 13262
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 20076 12640 20128 12646
rect 20076 12582 20128 12588
rect 17868 12232 17920 12238
rect 17868 12174 17920 12180
rect 18420 12232 18472 12238
rect 18420 12174 18472 12180
rect 17880 10674 17908 12174
rect 18432 11762 18460 12174
rect 18696 12096 18748 12102
rect 18696 12038 18748 12044
rect 18420 11756 18472 11762
rect 18420 11698 18472 11704
rect 18708 11218 18736 12038
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 19800 11552 19852 11558
rect 19800 11494 19852 11500
rect 19812 11286 19840 11494
rect 19800 11280 19852 11286
rect 19800 11222 19852 11228
rect 18696 11212 18748 11218
rect 18696 11154 18748 11160
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 19156 10736 19208 10742
rect 19156 10678 19208 10684
rect 17316 10668 17368 10674
rect 17316 10610 17368 10616
rect 17868 10668 17920 10674
rect 17868 10610 17920 10616
rect 16948 10532 17000 10538
rect 16948 10474 17000 10480
rect 16488 10260 16540 10266
rect 16488 10202 16540 10208
rect 16500 9722 16528 10202
rect 16580 10056 16632 10062
rect 16580 9998 16632 10004
rect 16488 9716 16540 9722
rect 16488 9658 16540 9664
rect 16592 8974 16620 9998
rect 16960 9518 16988 10474
rect 16948 9512 17000 9518
rect 16948 9454 17000 9460
rect 16580 8968 16632 8974
rect 16580 8910 16632 8916
rect 16592 8090 16620 8910
rect 16672 8832 16724 8838
rect 16672 8774 16724 8780
rect 16684 8430 16712 8774
rect 16672 8424 16724 8430
rect 16672 8366 16724 8372
rect 16580 8084 16632 8090
rect 16580 8026 16632 8032
rect 16960 7546 16988 9454
rect 17328 8430 17356 10610
rect 17776 10600 17828 10606
rect 17776 10542 17828 10548
rect 17316 8424 17368 8430
rect 17316 8366 17368 8372
rect 16948 7540 17000 7546
rect 16948 7482 17000 7488
rect 17328 7410 17356 8366
rect 16856 7404 16908 7410
rect 16856 7346 16908 7352
rect 17132 7404 17184 7410
rect 17132 7346 17184 7352
rect 17316 7404 17368 7410
rect 17316 7346 17368 7352
rect 16672 7200 16724 7206
rect 16672 7142 16724 7148
rect 16684 6798 16712 7142
rect 16868 7002 16896 7346
rect 16856 6996 16908 7002
rect 16856 6938 16908 6944
rect 16672 6792 16724 6798
rect 16672 6734 16724 6740
rect 16672 6656 16724 6662
rect 16672 6598 16724 6604
rect 16580 6180 16632 6186
rect 16580 6122 16632 6128
rect 16396 5364 16448 5370
rect 16396 5306 16448 5312
rect 16592 4978 16620 6122
rect 16684 5370 16712 6598
rect 16948 6452 17000 6458
rect 16948 6394 17000 6400
rect 16856 6112 16908 6118
rect 16856 6054 16908 6060
rect 16672 5364 16724 5370
rect 16672 5306 16724 5312
rect 16500 4950 16620 4978
rect 16500 4622 16528 4950
rect 16684 4842 16712 5306
rect 16592 4814 16712 4842
rect 16488 4616 16540 4622
rect 16488 4558 16540 4564
rect 16304 4480 16356 4486
rect 16304 4422 16356 4428
rect 16488 3936 16540 3942
rect 16488 3878 16540 3884
rect 16210 3632 16266 3641
rect 16210 3567 16266 3576
rect 16224 3534 16252 3567
rect 16212 3528 16264 3534
rect 16212 3470 16264 3476
rect 16304 3460 16356 3466
rect 16304 3402 16356 3408
rect 16120 3188 16172 3194
rect 16120 3130 16172 3136
rect 16132 2922 16160 3130
rect 16316 3126 16344 3402
rect 16304 3120 16356 3126
rect 16304 3062 16356 3068
rect 16120 2916 16172 2922
rect 16120 2858 16172 2864
rect 16040 2746 16160 2774
rect 16132 800 16160 2746
rect 16396 1896 16448 1902
rect 16396 1838 16448 1844
rect 16212 1556 16264 1562
rect 16212 1498 16264 1504
rect 16224 800 16252 1498
rect 16408 800 16436 1838
rect 16500 800 16528 3878
rect 16592 2514 16620 4814
rect 16670 4720 16726 4729
rect 16670 4655 16726 4664
rect 16684 4622 16712 4655
rect 16672 4616 16724 4622
rect 16672 4558 16724 4564
rect 16672 4004 16724 4010
rect 16672 3946 16724 3952
rect 16580 2508 16632 2514
rect 16580 2450 16632 2456
rect 16684 800 16712 3946
rect 16764 3392 16816 3398
rect 16764 3334 16816 3340
rect 16776 800 16804 3334
rect 16868 3058 16896 6054
rect 16960 5556 16988 6394
rect 17040 6112 17092 6118
rect 17040 6054 17092 6060
rect 17052 5681 17080 6054
rect 17038 5672 17094 5681
rect 17038 5607 17094 5616
rect 16960 5528 17080 5556
rect 16856 3052 16908 3058
rect 16856 2994 16908 3000
rect 17052 2938 17080 5528
rect 17144 4826 17172 7346
rect 17500 7336 17552 7342
rect 17500 7278 17552 7284
rect 17224 5840 17276 5846
rect 17224 5782 17276 5788
rect 17132 4820 17184 4826
rect 17132 4762 17184 4768
rect 17236 4706 17264 5782
rect 16960 2910 17080 2938
rect 17144 4678 17264 4706
rect 16960 800 16988 2910
rect 17040 2848 17092 2854
rect 17040 2790 17092 2796
rect 17052 800 17080 2790
rect 17144 1442 17172 4678
rect 17224 4140 17276 4146
rect 17224 4082 17276 4088
rect 17236 3058 17264 4082
rect 17316 3936 17368 3942
rect 17316 3878 17368 3884
rect 17224 3052 17276 3058
rect 17224 2994 17276 3000
rect 17236 2650 17264 2994
rect 17224 2644 17276 2650
rect 17224 2586 17276 2592
rect 17144 1414 17264 1442
rect 17236 800 17264 1414
rect 17328 800 17356 3878
rect 17512 800 17540 7278
rect 17592 7268 17644 7274
rect 17592 7210 17644 7216
rect 17604 4622 17632 7210
rect 17684 5704 17736 5710
rect 17684 5646 17736 5652
rect 17592 4616 17644 4622
rect 17592 4558 17644 4564
rect 17696 4010 17724 5646
rect 17788 4826 17816 10542
rect 17880 10062 17908 10610
rect 17868 10056 17920 10062
rect 17868 9998 17920 10004
rect 18236 9376 18288 9382
rect 18236 9318 18288 9324
rect 17868 8832 17920 8838
rect 17868 8774 17920 8780
rect 17880 7886 17908 8774
rect 18144 8492 18196 8498
rect 18144 8434 18196 8440
rect 18156 7886 18184 8434
rect 17868 7880 17920 7886
rect 17868 7822 17920 7828
rect 18144 7880 18196 7886
rect 18144 7822 18196 7828
rect 17776 4820 17828 4826
rect 17776 4762 17828 4768
rect 17880 4706 17908 7822
rect 18156 7410 18184 7822
rect 18144 7404 18196 7410
rect 18144 7346 18196 7352
rect 18248 6254 18276 9318
rect 18512 8832 18564 8838
rect 18512 8774 18564 8780
rect 18420 6452 18472 6458
rect 18420 6394 18472 6400
rect 18236 6248 18288 6254
rect 18236 6190 18288 6196
rect 18052 5908 18104 5914
rect 18052 5850 18104 5856
rect 18064 5778 18092 5850
rect 18052 5772 18104 5778
rect 18052 5714 18104 5720
rect 18064 5234 18092 5714
rect 18052 5228 18104 5234
rect 18052 5170 18104 5176
rect 17788 4678 17908 4706
rect 17684 4004 17736 4010
rect 17684 3946 17736 3952
rect 17684 2848 17736 2854
rect 17684 2790 17736 2796
rect 17696 2446 17724 2790
rect 17684 2440 17736 2446
rect 17684 2382 17736 2388
rect 17592 2372 17644 2378
rect 17592 2314 17644 2320
rect 17604 800 17632 2314
rect 17788 800 17816 4678
rect 17960 4480 18012 4486
rect 17960 4422 18012 4428
rect 17972 2530 18000 4422
rect 18064 4146 18092 5170
rect 18052 4140 18104 4146
rect 18052 4082 18104 4088
rect 18064 3534 18092 4082
rect 18052 3528 18104 3534
rect 18052 3470 18104 3476
rect 18064 2990 18092 3470
rect 18052 2984 18104 2990
rect 18052 2926 18104 2932
rect 18144 2916 18196 2922
rect 18144 2858 18196 2864
rect 17880 2502 18000 2530
rect 17880 800 17908 2502
rect 18156 1442 18184 2858
rect 18248 2774 18276 6190
rect 18432 4622 18460 6394
rect 18524 6322 18552 8774
rect 18972 8628 19024 8634
rect 18972 8570 19024 8576
rect 18880 7744 18932 7750
rect 18880 7686 18932 7692
rect 18892 6798 18920 7686
rect 18880 6792 18932 6798
rect 18880 6734 18932 6740
rect 18788 6724 18840 6730
rect 18788 6666 18840 6672
rect 18512 6316 18564 6322
rect 18564 6276 18644 6304
rect 18512 6258 18564 6264
rect 18420 4616 18472 4622
rect 18420 4558 18472 4564
rect 18420 2984 18472 2990
rect 18420 2926 18472 2932
rect 18248 2746 18368 2774
rect 18236 2372 18288 2378
rect 18236 2314 18288 2320
rect 18064 1414 18184 1442
rect 18064 800 18092 1414
rect 18248 1170 18276 2314
rect 18156 1142 18276 1170
rect 18156 800 18184 1142
rect 18340 800 18368 2746
rect 18432 2514 18460 2926
rect 18420 2508 18472 2514
rect 18420 2450 18472 2456
rect 18420 2304 18472 2310
rect 18420 2246 18472 2252
rect 18432 800 18460 2246
rect 18616 800 18644 6276
rect 18800 4826 18828 6666
rect 18788 4820 18840 4826
rect 18788 4762 18840 4768
rect 18696 3664 18748 3670
rect 18696 3606 18748 3612
rect 18708 800 18736 3606
rect 18892 800 18920 6734
rect 18984 3534 19012 8570
rect 19168 8430 19196 10678
rect 19248 9988 19300 9994
rect 19248 9930 19300 9936
rect 19260 9654 19288 9930
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 19248 9648 19300 9654
rect 19248 9590 19300 9596
rect 19984 9444 20036 9450
rect 19984 9386 20036 9392
rect 19432 8832 19484 8838
rect 19432 8774 19484 8780
rect 19156 8424 19208 8430
rect 19156 8366 19208 8372
rect 19168 7410 19196 8366
rect 19340 8356 19392 8362
rect 19340 8298 19392 8304
rect 19352 7478 19380 8298
rect 19340 7472 19392 7478
rect 19340 7414 19392 7420
rect 19156 7404 19208 7410
rect 19156 7346 19208 7352
rect 19444 7290 19472 8774
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 19352 7262 19472 7290
rect 19064 6384 19116 6390
rect 19064 6326 19116 6332
rect 19076 5030 19104 6326
rect 19248 6112 19300 6118
rect 19248 6054 19300 6060
rect 19260 5778 19288 6054
rect 19248 5772 19300 5778
rect 19248 5714 19300 5720
rect 19352 5710 19380 7262
rect 19432 6656 19484 6662
rect 19432 6598 19484 6604
rect 19340 5704 19392 5710
rect 19340 5646 19392 5652
rect 19352 5137 19380 5646
rect 19444 5234 19472 6598
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 19996 6322 20024 9386
rect 20088 8294 20116 12582
rect 20904 12368 20956 12374
rect 20904 12310 20956 12316
rect 20812 12300 20864 12306
rect 20812 12242 20864 12248
rect 20536 12164 20588 12170
rect 20536 12106 20588 12112
rect 20548 11898 20576 12106
rect 20536 11892 20588 11898
rect 20536 11834 20588 11840
rect 20444 11756 20496 11762
rect 20444 11698 20496 11704
rect 20456 10810 20484 11698
rect 20824 11694 20852 12242
rect 20916 11762 20944 12310
rect 21272 12232 21324 12238
rect 21324 12192 21404 12220
rect 21272 12174 21324 12180
rect 20904 11756 20956 11762
rect 20904 11698 20956 11704
rect 21088 11756 21140 11762
rect 21088 11698 21140 11704
rect 21272 11756 21324 11762
rect 21272 11698 21324 11704
rect 20812 11688 20864 11694
rect 20812 11630 20864 11636
rect 20628 11280 20680 11286
rect 20628 11222 20680 11228
rect 20444 10804 20496 10810
rect 20444 10746 20496 10752
rect 20640 10674 20668 11222
rect 20824 10810 20852 11630
rect 20916 10810 20944 11698
rect 20812 10804 20864 10810
rect 20812 10746 20864 10752
rect 20904 10804 20956 10810
rect 20904 10746 20956 10752
rect 20168 10668 20220 10674
rect 20168 10610 20220 10616
rect 20628 10668 20680 10674
rect 20628 10610 20680 10616
rect 20180 10266 20208 10610
rect 20536 10532 20588 10538
rect 20536 10474 20588 10480
rect 20444 10464 20496 10470
rect 20444 10406 20496 10412
rect 20168 10260 20220 10266
rect 20168 10202 20220 10208
rect 20456 10062 20484 10406
rect 20444 10056 20496 10062
rect 20444 9998 20496 10004
rect 20444 9512 20496 9518
rect 20444 9454 20496 9460
rect 20456 9178 20484 9454
rect 20444 9172 20496 9178
rect 20444 9114 20496 9120
rect 20168 8968 20220 8974
rect 20168 8910 20220 8916
rect 20076 8288 20128 8294
rect 20076 8230 20128 8236
rect 20088 7886 20116 8230
rect 20076 7880 20128 7886
rect 20076 7822 20128 7828
rect 19984 6316 20036 6322
rect 19984 6258 20036 6264
rect 20180 6202 20208 8910
rect 20352 8900 20404 8906
rect 20352 8842 20404 8848
rect 20364 8634 20392 8842
rect 20548 8634 20576 10474
rect 20720 10464 20772 10470
rect 20720 10406 20772 10412
rect 20628 10056 20680 10062
rect 20628 9998 20680 10004
rect 20352 8628 20404 8634
rect 20352 8570 20404 8576
rect 20536 8628 20588 8634
rect 20536 8570 20588 8576
rect 20260 8492 20312 8498
rect 20260 8434 20312 8440
rect 20444 8492 20496 8498
rect 20444 8434 20496 8440
rect 20272 8265 20300 8434
rect 20258 8256 20314 8265
rect 20258 8191 20314 8200
rect 20272 7002 20300 8191
rect 20352 8016 20404 8022
rect 20352 7958 20404 7964
rect 20364 7750 20392 7958
rect 20352 7744 20404 7750
rect 20352 7686 20404 7692
rect 20260 6996 20312 7002
rect 20260 6938 20312 6944
rect 19996 6174 20208 6202
rect 20260 6180 20312 6186
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 19996 5409 20024 6174
rect 20260 6122 20312 6128
rect 20168 5908 20220 5914
rect 20088 5868 20168 5896
rect 19982 5400 20038 5409
rect 19982 5335 20038 5344
rect 19432 5228 19484 5234
rect 19432 5170 19484 5176
rect 19338 5128 19394 5137
rect 19982 5128 20038 5137
rect 19338 5063 19394 5072
rect 19708 5092 19760 5098
rect 19982 5063 20038 5072
rect 19708 5034 19760 5040
rect 19064 5024 19116 5030
rect 19064 4966 19116 4972
rect 19248 5024 19300 5030
rect 19300 4984 19472 5012
rect 19248 4966 19300 4972
rect 19156 4820 19208 4826
rect 19156 4762 19208 4768
rect 18972 3528 19024 3534
rect 18972 3470 19024 3476
rect 18972 3392 19024 3398
rect 18972 3334 19024 3340
rect 18984 800 19012 3334
rect 19062 2816 19118 2825
rect 19062 2751 19118 2760
rect 19076 2650 19104 2751
rect 19064 2644 19116 2650
rect 19064 2586 19116 2592
rect 19168 800 19196 4762
rect 19340 3936 19392 3942
rect 19338 3904 19340 3913
rect 19392 3904 19394 3913
rect 19338 3839 19394 3848
rect 19444 3754 19472 4984
rect 19616 4616 19668 4622
rect 19614 4584 19616 4593
rect 19668 4584 19670 4593
rect 19614 4519 19670 4528
rect 19720 4486 19748 5034
rect 19800 5024 19852 5030
rect 19798 4992 19800 5001
rect 19852 4992 19854 5001
rect 19798 4927 19854 4936
rect 19708 4480 19760 4486
rect 19708 4422 19760 4428
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 19352 3726 19472 3754
rect 19248 2372 19300 2378
rect 19248 2314 19300 2320
rect 19260 800 19288 2314
rect 19352 1442 19380 3726
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 19432 2916 19484 2922
rect 19432 2858 19484 2864
rect 19444 1578 19472 2858
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 19444 1550 19564 1578
rect 19352 1414 19472 1442
rect 19444 800 19472 1414
rect 19536 800 19564 1550
rect 19996 1442 20024 5063
rect 20088 2825 20116 5868
rect 20168 5850 20220 5856
rect 20272 5642 20300 6122
rect 20260 5636 20312 5642
rect 20260 5578 20312 5584
rect 20364 5522 20392 7686
rect 20456 7546 20484 8434
rect 20444 7540 20496 7546
rect 20444 7482 20496 7488
rect 20456 6361 20484 7482
rect 20536 6724 20588 6730
rect 20536 6666 20588 6672
rect 20442 6352 20498 6361
rect 20548 6322 20576 6666
rect 20442 6287 20498 6296
rect 20536 6316 20588 6322
rect 20536 6258 20588 6264
rect 20444 6112 20496 6118
rect 20444 6054 20496 6060
rect 20456 5817 20484 6054
rect 20442 5808 20498 5817
rect 20442 5743 20498 5752
rect 20444 5568 20496 5574
rect 20180 5494 20392 5522
rect 20442 5536 20444 5545
rect 20496 5536 20498 5545
rect 20074 2816 20130 2825
rect 20074 2751 20130 2760
rect 20180 2446 20208 5494
rect 20442 5471 20498 5480
rect 20258 5400 20314 5409
rect 20258 5335 20314 5344
rect 20272 3738 20300 5335
rect 20548 5250 20576 6258
rect 20640 5370 20668 9998
rect 20732 8974 20760 10406
rect 20824 9926 20852 10746
rect 20904 10671 20956 10677
rect 20904 10613 20956 10619
rect 20812 9920 20864 9926
rect 20812 9862 20864 9868
rect 20812 9580 20864 9586
rect 20812 9522 20864 9528
rect 20720 8968 20772 8974
rect 20720 8910 20772 8916
rect 20720 7200 20772 7206
rect 20720 7142 20772 7148
rect 20732 6882 20760 7142
rect 20824 7002 20852 9522
rect 20812 6996 20864 7002
rect 20812 6938 20864 6944
rect 20732 6854 20852 6882
rect 20720 6656 20772 6662
rect 20720 6598 20772 6604
rect 20628 5364 20680 5370
rect 20628 5306 20680 5312
rect 20732 5302 20760 6598
rect 20824 6322 20852 6854
rect 20812 6316 20864 6322
rect 20812 6258 20864 6264
rect 20824 6225 20852 6258
rect 20810 6216 20866 6225
rect 20810 6151 20866 6160
rect 20812 5704 20864 5710
rect 20812 5646 20864 5652
rect 20720 5296 20772 5302
rect 20548 5222 20668 5250
rect 20720 5238 20772 5244
rect 20824 5234 20852 5646
rect 20444 5160 20496 5166
rect 20444 5102 20496 5108
rect 20456 4672 20484 5102
rect 20536 4684 20588 4690
rect 20456 4644 20536 4672
rect 20352 4480 20404 4486
rect 20352 4422 20404 4428
rect 20260 3732 20312 3738
rect 20260 3674 20312 3680
rect 20260 2576 20312 2582
rect 20260 2518 20312 2524
rect 20168 2440 20220 2446
rect 20168 2382 20220 2388
rect 20076 2304 20128 2310
rect 20076 2246 20128 2252
rect 19720 1414 20024 1442
rect 19720 800 19748 1414
rect 19800 1352 19852 1358
rect 19800 1294 19852 1300
rect 19984 1352 20036 1358
rect 19984 1294 20036 1300
rect 19812 800 19840 1294
rect 19996 800 20024 1294
rect 20088 800 20116 2246
rect 20272 1426 20300 2518
rect 20260 1420 20312 1426
rect 20260 1362 20312 1368
rect 20364 800 20392 4422
rect 20456 4282 20484 4644
rect 20536 4626 20588 4632
rect 20640 4622 20668 5222
rect 20812 5228 20864 5234
rect 20812 5170 20864 5176
rect 20720 5092 20772 5098
rect 20720 5034 20772 5040
rect 20628 4616 20680 4622
rect 20628 4558 20680 4564
rect 20444 4276 20496 4282
rect 20444 4218 20496 4224
rect 20456 4078 20484 4218
rect 20640 4146 20668 4558
rect 20732 4214 20760 5034
rect 20916 4826 20944 10613
rect 20996 10600 21048 10606
rect 20996 10542 21048 10548
rect 21008 10062 21036 10542
rect 20996 10056 21048 10062
rect 20996 9998 21048 10004
rect 20996 6860 21048 6866
rect 20996 6802 21048 6808
rect 20904 4820 20956 4826
rect 20904 4762 20956 4768
rect 21008 4622 21036 6802
rect 21100 5370 21128 11698
rect 21284 10674 21312 11698
rect 21376 11218 21404 12192
rect 21364 11212 21416 11218
rect 21364 11154 21416 11160
rect 21272 10668 21324 10674
rect 21272 10610 21324 10616
rect 21272 8968 21324 8974
rect 21272 8910 21324 8916
rect 21284 8430 21312 8910
rect 21560 8537 21588 13806
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 65654 13628 65962 13637
rect 65654 13626 65660 13628
rect 65716 13626 65740 13628
rect 65796 13626 65820 13628
rect 65876 13626 65900 13628
rect 65956 13626 65962 13628
rect 65716 13574 65718 13626
rect 65898 13574 65900 13626
rect 65654 13572 65660 13574
rect 65716 13572 65740 13574
rect 65796 13572 65820 13574
rect 65876 13572 65900 13574
rect 65956 13572 65962 13574
rect 65654 13563 65962 13572
rect 50294 13084 50602 13093
rect 50294 13082 50300 13084
rect 50356 13082 50380 13084
rect 50436 13082 50460 13084
rect 50516 13082 50540 13084
rect 50596 13082 50602 13084
rect 50356 13030 50358 13082
rect 50538 13030 50540 13082
rect 50294 13028 50300 13030
rect 50356 13028 50380 13030
rect 50436 13028 50460 13030
rect 50516 13028 50540 13030
rect 50596 13028 50602 13030
rect 50294 13019 50602 13028
rect 21732 12844 21784 12850
rect 21732 12786 21784 12792
rect 21744 12238 21772 12786
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 65654 12540 65962 12549
rect 65654 12538 65660 12540
rect 65716 12538 65740 12540
rect 65796 12538 65820 12540
rect 65876 12538 65900 12540
rect 65956 12538 65962 12540
rect 65716 12486 65718 12538
rect 65898 12486 65900 12538
rect 65654 12484 65660 12486
rect 65716 12484 65740 12486
rect 65796 12484 65820 12486
rect 65876 12484 65900 12486
rect 65956 12484 65962 12486
rect 65654 12475 65962 12484
rect 21732 12232 21784 12238
rect 22376 12232 22428 12238
rect 21732 12174 21784 12180
rect 22296 12192 22376 12220
rect 21640 12096 21692 12102
rect 21640 12038 21692 12044
rect 21546 8528 21602 8537
rect 21546 8463 21548 8472
rect 21600 8463 21602 8472
rect 21548 8434 21600 8440
rect 21272 8424 21324 8430
rect 21270 8392 21272 8401
rect 21560 8403 21588 8434
rect 21324 8392 21326 8401
rect 21270 8327 21326 8336
rect 21548 8084 21600 8090
rect 21548 8026 21600 8032
rect 21456 7880 21508 7886
rect 21456 7822 21508 7828
rect 21468 7546 21496 7822
rect 21456 7540 21508 7546
rect 21456 7482 21508 7488
rect 21456 7268 21508 7274
rect 21456 7210 21508 7216
rect 21468 6798 21496 7210
rect 21560 7206 21588 8026
rect 21548 7200 21600 7206
rect 21548 7142 21600 7148
rect 21456 6792 21508 6798
rect 21456 6734 21508 6740
rect 21180 6656 21232 6662
rect 21180 6598 21232 6604
rect 21192 6186 21220 6598
rect 21180 6180 21232 6186
rect 21180 6122 21232 6128
rect 21272 6112 21324 6118
rect 21272 6054 21324 6060
rect 21180 5704 21232 5710
rect 21180 5646 21232 5652
rect 21088 5364 21140 5370
rect 21088 5306 21140 5312
rect 20996 4616 21048 4622
rect 20996 4558 21048 4564
rect 21086 4584 21142 4593
rect 20904 4548 20956 4554
rect 21086 4519 21142 4528
rect 20904 4490 20956 4496
rect 20812 4480 20864 4486
rect 20812 4422 20864 4428
rect 20720 4208 20772 4214
rect 20720 4150 20772 4156
rect 20628 4140 20680 4146
rect 20628 4082 20680 4088
rect 20444 4072 20496 4078
rect 20444 4014 20496 4020
rect 20536 3936 20588 3942
rect 20536 3878 20588 3884
rect 20444 3732 20496 3738
rect 20444 3674 20496 3680
rect 20456 2446 20484 3674
rect 20444 2440 20496 2446
rect 20444 2382 20496 2388
rect 20548 1358 20576 3878
rect 20640 3670 20668 4082
rect 20628 3664 20680 3670
rect 20628 3606 20680 3612
rect 20628 3460 20680 3466
rect 20628 3402 20680 3408
rect 20536 1352 20588 1358
rect 20536 1294 20588 1300
rect 20640 800 20668 3402
rect 20824 3126 20852 4422
rect 20916 3534 20944 4490
rect 20904 3528 20956 3534
rect 20904 3470 20956 3476
rect 20812 3120 20864 3126
rect 20718 3088 20774 3097
rect 20812 3062 20864 3068
rect 20718 3023 20720 3032
rect 20772 3023 20774 3032
rect 20720 2994 20772 3000
rect 20916 2922 20944 3470
rect 20904 2916 20956 2922
rect 20904 2858 20956 2864
rect 21100 2666 21128 4519
rect 20904 2644 20956 2650
rect 20904 2586 20956 2592
rect 21008 2638 21128 2666
rect 20916 800 20944 2586
rect 21008 800 21036 2638
rect 21192 800 21220 5646
rect 21284 5030 21312 6054
rect 21456 5228 21508 5234
rect 21456 5170 21508 5176
rect 21548 5228 21600 5234
rect 21548 5170 21600 5176
rect 21272 5024 21324 5030
rect 21272 4966 21324 4972
rect 21284 4826 21312 4966
rect 21272 4820 21324 4826
rect 21272 4762 21324 4768
rect 21364 4752 21416 4758
rect 21364 4694 21416 4700
rect 21376 3534 21404 4694
rect 21468 4554 21496 5170
rect 21456 4548 21508 4554
rect 21456 4490 21508 4496
rect 21468 4214 21496 4490
rect 21456 4208 21508 4214
rect 21456 4150 21508 4156
rect 21456 4004 21508 4010
rect 21456 3946 21508 3952
rect 21272 3528 21324 3534
rect 21272 3470 21324 3476
rect 21364 3528 21416 3534
rect 21364 3470 21416 3476
rect 21284 3194 21312 3470
rect 21364 3392 21416 3398
rect 21364 3334 21416 3340
rect 21272 3188 21324 3194
rect 21272 3130 21324 3136
rect 21376 3074 21404 3334
rect 21284 3046 21404 3074
rect 21284 2854 21312 3046
rect 21272 2848 21324 2854
rect 21272 2790 21324 2796
rect 21284 800 21312 2790
rect 21468 800 21496 3946
rect 21560 800 21588 5170
rect 21652 4758 21680 12038
rect 21744 11762 21772 12174
rect 21732 11756 21784 11762
rect 21732 11698 21784 11704
rect 22100 11348 22152 11354
rect 22100 11290 22152 11296
rect 22112 10470 22140 11290
rect 22100 10464 22152 10470
rect 22100 10406 22152 10412
rect 22112 10266 22140 10406
rect 22100 10260 22152 10266
rect 22100 10202 22152 10208
rect 21732 9920 21784 9926
rect 21732 9862 21784 9868
rect 21744 9518 21772 9862
rect 21732 9512 21784 9518
rect 21732 9454 21784 9460
rect 21744 8090 21772 9454
rect 22112 9450 22140 10202
rect 22296 9602 22324 12192
rect 22376 12174 22428 12180
rect 22560 12096 22612 12102
rect 22560 12038 22612 12044
rect 22572 11830 22600 12038
rect 50294 11996 50602 12005
rect 50294 11994 50300 11996
rect 50356 11994 50380 11996
rect 50436 11994 50460 11996
rect 50516 11994 50540 11996
rect 50596 11994 50602 11996
rect 50356 11942 50358 11994
rect 50538 11942 50540 11994
rect 50294 11940 50300 11942
rect 50356 11940 50380 11942
rect 50436 11940 50460 11942
rect 50516 11940 50540 11942
rect 50596 11940 50602 11942
rect 50294 11931 50602 11940
rect 22560 11824 22612 11830
rect 22560 11766 22612 11772
rect 22376 11144 22428 11150
rect 22376 11086 22428 11092
rect 22388 10674 22416 11086
rect 22376 10668 22428 10674
rect 22376 10610 22428 10616
rect 22572 10606 22600 11766
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 65654 11452 65962 11461
rect 65654 11450 65660 11452
rect 65716 11450 65740 11452
rect 65796 11450 65820 11452
rect 65876 11450 65900 11452
rect 65956 11450 65962 11452
rect 65716 11398 65718 11450
rect 65898 11398 65900 11450
rect 65654 11396 65660 11398
rect 65716 11396 65740 11398
rect 65796 11396 65820 11398
rect 65876 11396 65900 11398
rect 65956 11396 65962 11398
rect 65654 11387 65962 11396
rect 23204 11348 23256 11354
rect 23204 11290 23256 11296
rect 23112 11280 23164 11286
rect 23112 11222 23164 11228
rect 23020 11144 23072 11150
rect 23020 11086 23072 11092
rect 22652 10668 22704 10674
rect 22652 10610 22704 10616
rect 22560 10600 22612 10606
rect 22560 10542 22612 10548
rect 22560 10192 22612 10198
rect 22560 10134 22612 10140
rect 22204 9574 22324 9602
rect 22572 9586 22600 10134
rect 22664 10062 22692 10610
rect 22652 10056 22704 10062
rect 22652 9998 22704 10004
rect 22560 9580 22612 9586
rect 22100 9444 22152 9450
rect 22100 9386 22152 9392
rect 22100 9172 22152 9178
rect 22100 9114 22152 9120
rect 22112 8906 22140 9114
rect 22100 8900 22152 8906
rect 22100 8842 22152 8848
rect 22112 8498 22140 8842
rect 21916 8492 21968 8498
rect 21916 8434 21968 8440
rect 22100 8492 22152 8498
rect 22100 8434 22152 8440
rect 21732 8084 21784 8090
rect 21732 8026 21784 8032
rect 21928 5778 21956 8434
rect 22008 7404 22060 7410
rect 22008 7346 22060 7352
rect 22020 6934 22048 7346
rect 22008 6928 22060 6934
rect 22008 6870 22060 6876
rect 22100 6724 22152 6730
rect 22100 6666 22152 6672
rect 22112 6458 22140 6666
rect 22100 6452 22152 6458
rect 22100 6394 22152 6400
rect 22112 5778 22140 6394
rect 21916 5772 21968 5778
rect 21916 5714 21968 5720
rect 22100 5772 22152 5778
rect 22100 5714 22152 5720
rect 22098 5536 22154 5545
rect 22098 5471 22154 5480
rect 21824 5024 21876 5030
rect 21824 4966 21876 4972
rect 21640 4752 21692 4758
rect 21640 4694 21692 4700
rect 21640 4140 21692 4146
rect 21640 4082 21692 4088
rect 21652 2854 21680 4082
rect 21732 3936 21784 3942
rect 21732 3878 21784 3884
rect 21744 3534 21772 3878
rect 21836 3738 21864 4966
rect 21916 4820 21968 4826
rect 21916 4762 21968 4768
rect 21928 3942 21956 4762
rect 22112 4622 22140 5471
rect 22100 4616 22152 4622
rect 22100 4558 22152 4564
rect 22100 4140 22152 4146
rect 22100 4082 22152 4088
rect 22008 4072 22060 4078
rect 22112 4049 22140 4082
rect 22008 4014 22060 4020
rect 22098 4040 22154 4049
rect 21916 3936 21968 3942
rect 21916 3878 21968 3884
rect 21824 3732 21876 3738
rect 21824 3674 21876 3680
rect 21824 3596 21876 3602
rect 21824 3538 21876 3544
rect 21732 3528 21784 3534
rect 21732 3470 21784 3476
rect 21836 3210 21864 3538
rect 21744 3182 21864 3210
rect 21640 2848 21692 2854
rect 21640 2790 21692 2796
rect 21744 800 21772 3182
rect 21824 2848 21876 2854
rect 21824 2790 21876 2796
rect 21836 800 21864 2790
rect 22020 800 22048 4014
rect 22204 4010 22232 9574
rect 22560 9522 22612 9528
rect 22572 8786 22600 9522
rect 22664 9382 22692 9998
rect 23032 9722 23060 11086
rect 23020 9716 23072 9722
rect 23020 9658 23072 9664
rect 22928 9512 22980 9518
rect 22928 9454 22980 9460
rect 22652 9376 22704 9382
rect 22652 9318 22704 9324
rect 22940 8906 22968 9454
rect 22928 8900 22980 8906
rect 22928 8842 22980 8848
rect 22744 8832 22796 8838
rect 22572 8758 22692 8786
rect 22744 8774 22796 8780
rect 22558 8256 22614 8265
rect 22558 8191 22614 8200
rect 22284 7744 22336 7750
rect 22284 7686 22336 7692
rect 22296 6322 22324 7686
rect 22572 7342 22600 8191
rect 22560 7336 22612 7342
rect 22560 7278 22612 7284
rect 22468 6792 22520 6798
rect 22468 6734 22520 6740
rect 22480 6322 22508 6734
rect 22284 6316 22336 6322
rect 22284 6258 22336 6264
rect 22468 6316 22520 6322
rect 22468 6258 22520 6264
rect 22284 5024 22336 5030
rect 22284 4966 22336 4972
rect 22098 3975 22154 3984
rect 22192 4004 22244 4010
rect 22192 3946 22244 3952
rect 22192 2984 22244 2990
rect 22192 2926 22244 2932
rect 22204 800 22232 2926
rect 22296 2650 22324 4966
rect 22468 3936 22520 3942
rect 22468 3878 22520 3884
rect 22284 2644 22336 2650
rect 22284 2586 22336 2592
rect 22480 800 22508 3878
rect 22664 2514 22692 8758
rect 22756 8566 22784 8774
rect 22744 8560 22796 8566
rect 22744 8502 22796 8508
rect 22926 8392 22982 8401
rect 22926 8327 22982 8336
rect 22940 6254 22968 8327
rect 23032 7342 23060 9658
rect 23124 7886 23152 11222
rect 23216 10130 23244 11290
rect 23848 11280 23900 11286
rect 23848 11222 23900 11228
rect 23572 11144 23624 11150
rect 23572 11086 23624 11092
rect 23388 10464 23440 10470
rect 23388 10406 23440 10412
rect 23204 10124 23256 10130
rect 23204 10066 23256 10072
rect 23204 9920 23256 9926
rect 23204 9862 23256 9868
rect 23296 9920 23348 9926
rect 23296 9862 23348 9868
rect 23216 9586 23244 9862
rect 23204 9580 23256 9586
rect 23204 9522 23256 9528
rect 23204 9444 23256 9450
rect 23204 9386 23256 9392
rect 23216 9110 23244 9386
rect 23204 9104 23256 9110
rect 23204 9046 23256 9052
rect 23216 8498 23244 9046
rect 23308 8974 23336 9862
rect 23296 8968 23348 8974
rect 23296 8910 23348 8916
rect 23296 8832 23348 8838
rect 23296 8774 23348 8780
rect 23308 8566 23336 8774
rect 23296 8560 23348 8566
rect 23296 8502 23348 8508
rect 23204 8492 23256 8498
rect 23204 8434 23256 8440
rect 23216 7954 23244 8434
rect 23308 8022 23336 8502
rect 23400 8498 23428 10406
rect 23584 10198 23612 11086
rect 23664 11008 23716 11014
rect 23664 10950 23716 10956
rect 23676 10742 23704 10950
rect 23664 10736 23716 10742
rect 23664 10678 23716 10684
rect 23860 10674 23888 11222
rect 24492 11076 24544 11082
rect 24492 11018 24544 11024
rect 23848 10668 23900 10674
rect 23848 10610 23900 10616
rect 23572 10192 23624 10198
rect 23572 10134 23624 10140
rect 24306 8528 24362 8537
rect 23388 8492 23440 8498
rect 24306 8463 24308 8472
rect 23388 8434 23440 8440
rect 24360 8463 24362 8472
rect 24308 8434 24360 8440
rect 23296 8016 23348 8022
rect 23296 7958 23348 7964
rect 23204 7948 23256 7954
rect 23204 7890 23256 7896
rect 23112 7880 23164 7886
rect 23112 7822 23164 7828
rect 23756 7540 23808 7546
rect 23756 7482 23808 7488
rect 23296 7404 23348 7410
rect 23296 7346 23348 7352
rect 23020 7336 23072 7342
rect 23020 7278 23072 7284
rect 23308 6866 23336 7346
rect 23572 7200 23624 7206
rect 23572 7142 23624 7148
rect 23296 6860 23348 6866
rect 23296 6802 23348 6808
rect 23388 6792 23440 6798
rect 23388 6734 23440 6740
rect 23296 6724 23348 6730
rect 23296 6666 23348 6672
rect 22928 6248 22980 6254
rect 22928 6190 22980 6196
rect 23204 6180 23256 6186
rect 23204 6122 23256 6128
rect 23216 5574 23244 6122
rect 23204 5568 23256 5574
rect 23204 5510 23256 5516
rect 23216 5273 23244 5510
rect 23308 5302 23336 6666
rect 23400 5914 23428 6734
rect 23388 5908 23440 5914
rect 23388 5850 23440 5856
rect 23296 5296 23348 5302
rect 23202 5264 23258 5273
rect 22836 5228 22888 5234
rect 23296 5238 23348 5244
rect 23202 5199 23258 5208
rect 22836 5170 22888 5176
rect 22848 3913 22876 5170
rect 23308 4758 23336 5238
rect 23296 4752 23348 4758
rect 23296 4694 23348 4700
rect 23584 4622 23612 7142
rect 23664 6792 23716 6798
rect 23664 6734 23716 6740
rect 23676 6322 23704 6734
rect 23664 6316 23716 6322
rect 23664 6258 23716 6264
rect 23676 5370 23704 6258
rect 23664 5364 23716 5370
rect 23664 5306 23716 5312
rect 23676 4622 23704 5306
rect 23768 5234 23796 7482
rect 24320 5914 24348 8434
rect 24400 7744 24452 7750
rect 24400 7686 24452 7692
rect 24412 7342 24440 7686
rect 24400 7336 24452 7342
rect 24400 7278 24452 7284
rect 24412 7002 24440 7278
rect 24400 6996 24452 7002
rect 24400 6938 24452 6944
rect 24504 6866 24532 11018
rect 50294 10908 50602 10917
rect 50294 10906 50300 10908
rect 50356 10906 50380 10908
rect 50436 10906 50460 10908
rect 50516 10906 50540 10908
rect 50596 10906 50602 10908
rect 50356 10854 50358 10906
rect 50538 10854 50540 10906
rect 50294 10852 50300 10854
rect 50356 10852 50380 10854
rect 50436 10852 50460 10854
rect 50516 10852 50540 10854
rect 50596 10852 50602 10854
rect 50294 10843 50602 10852
rect 26976 10464 27028 10470
rect 26976 10406 27028 10412
rect 24492 6860 24544 6866
rect 24492 6802 24544 6808
rect 24308 5908 24360 5914
rect 24308 5850 24360 5856
rect 23756 5228 23808 5234
rect 23756 5170 23808 5176
rect 23572 4616 23624 4622
rect 23572 4558 23624 4564
rect 23664 4616 23716 4622
rect 24400 4616 24452 4622
rect 23664 4558 23716 4564
rect 24398 4584 24400 4593
rect 24452 4584 24454 4593
rect 24398 4519 24454 4528
rect 24032 3936 24084 3942
rect 22834 3904 22890 3913
rect 24032 3878 24084 3884
rect 24676 3936 24728 3942
rect 24676 3878 24728 3884
rect 22834 3839 22890 3848
rect 22744 3528 22796 3534
rect 22744 3470 22796 3476
rect 22652 2508 22704 2514
rect 22652 2450 22704 2456
rect 22756 800 22784 3470
rect 22848 2446 22876 3839
rect 23572 3528 23624 3534
rect 23572 3470 23624 3476
rect 23020 2848 23072 2854
rect 23020 2790 23072 2796
rect 23296 2848 23348 2854
rect 23296 2790 23348 2796
rect 22836 2440 22888 2446
rect 22836 2382 22888 2388
rect 23032 800 23060 2790
rect 23308 800 23336 2790
rect 23584 800 23612 3470
rect 24044 3466 24072 3878
rect 24032 3460 24084 3466
rect 24032 3402 24084 3408
rect 24688 3398 24716 3878
rect 26056 3528 26108 3534
rect 26056 3470 26108 3476
rect 24676 3392 24728 3398
rect 24676 3334 24728 3340
rect 24952 3392 25004 3398
rect 24952 3334 25004 3340
rect 24124 2848 24176 2854
rect 24124 2790 24176 2796
rect 24676 2848 24728 2854
rect 24676 2790 24728 2796
rect 23848 2576 23900 2582
rect 23848 2518 23900 2524
rect 23860 800 23888 2518
rect 24136 800 24164 2790
rect 24400 2440 24452 2446
rect 24400 2382 24452 2388
rect 24412 800 24440 2382
rect 24688 800 24716 2790
rect 24964 800 24992 3334
rect 25228 2984 25280 2990
rect 25228 2926 25280 2932
rect 25240 800 25268 2926
rect 25780 2848 25832 2854
rect 25780 2790 25832 2796
rect 25504 2304 25556 2310
rect 25504 2246 25556 2252
rect 25516 800 25544 2246
rect 25792 800 25820 2790
rect 26068 800 26096 3470
rect 26422 2952 26478 2961
rect 26422 2887 26478 2896
rect 26436 2854 26464 2887
rect 26332 2848 26384 2854
rect 26332 2790 26384 2796
rect 26424 2848 26476 2854
rect 26424 2790 26476 2796
rect 26344 800 26372 2790
rect 26436 2446 26464 2790
rect 26988 2446 27016 10406
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 65654 10364 65962 10373
rect 65654 10362 65660 10364
rect 65716 10362 65740 10364
rect 65796 10362 65820 10364
rect 65876 10362 65900 10364
rect 65956 10362 65962 10364
rect 65716 10310 65718 10362
rect 65898 10310 65900 10362
rect 65654 10308 65660 10310
rect 65716 10308 65740 10310
rect 65796 10308 65820 10310
rect 65876 10308 65900 10310
rect 65956 10308 65962 10310
rect 65654 10299 65962 10308
rect 50294 9820 50602 9829
rect 50294 9818 50300 9820
rect 50356 9818 50380 9820
rect 50436 9818 50460 9820
rect 50516 9818 50540 9820
rect 50596 9818 50602 9820
rect 50356 9766 50358 9818
rect 50538 9766 50540 9818
rect 50294 9764 50300 9766
rect 50356 9764 50380 9766
rect 50436 9764 50460 9766
rect 50516 9764 50540 9766
rect 50596 9764 50602 9766
rect 50294 9755 50602 9764
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 65654 9276 65962 9285
rect 65654 9274 65660 9276
rect 65716 9274 65740 9276
rect 65796 9274 65820 9276
rect 65876 9274 65900 9276
rect 65956 9274 65962 9276
rect 65716 9222 65718 9274
rect 65898 9222 65900 9274
rect 65654 9220 65660 9222
rect 65716 9220 65740 9222
rect 65796 9220 65820 9222
rect 65876 9220 65900 9222
rect 65956 9220 65962 9222
rect 65654 9211 65962 9220
rect 50294 8732 50602 8741
rect 50294 8730 50300 8732
rect 50356 8730 50380 8732
rect 50436 8730 50460 8732
rect 50516 8730 50540 8732
rect 50596 8730 50602 8732
rect 50356 8678 50358 8730
rect 50538 8678 50540 8730
rect 50294 8676 50300 8678
rect 50356 8676 50380 8678
rect 50436 8676 50460 8678
rect 50516 8676 50540 8678
rect 50596 8676 50602 8678
rect 50294 8667 50602 8676
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 65654 8188 65962 8197
rect 65654 8186 65660 8188
rect 65716 8186 65740 8188
rect 65796 8186 65820 8188
rect 65876 8186 65900 8188
rect 65956 8186 65962 8188
rect 65716 8134 65718 8186
rect 65898 8134 65900 8186
rect 65654 8132 65660 8134
rect 65716 8132 65740 8134
rect 65796 8132 65820 8134
rect 65876 8132 65900 8134
rect 65956 8132 65962 8134
rect 65654 8123 65962 8132
rect 50294 7644 50602 7653
rect 50294 7642 50300 7644
rect 50356 7642 50380 7644
rect 50436 7642 50460 7644
rect 50516 7642 50540 7644
rect 50596 7642 50602 7644
rect 50356 7590 50358 7642
rect 50538 7590 50540 7642
rect 50294 7588 50300 7590
rect 50356 7588 50380 7590
rect 50436 7588 50460 7590
rect 50516 7588 50540 7590
rect 50596 7588 50602 7590
rect 50294 7579 50602 7588
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 65654 7100 65962 7109
rect 65654 7098 65660 7100
rect 65716 7098 65740 7100
rect 65796 7098 65820 7100
rect 65876 7098 65900 7100
rect 65956 7098 65962 7100
rect 65716 7046 65718 7098
rect 65898 7046 65900 7098
rect 65654 7044 65660 7046
rect 65716 7044 65740 7046
rect 65796 7044 65820 7046
rect 65876 7044 65900 7046
rect 65956 7044 65962 7046
rect 65654 7035 65962 7044
rect 50294 6556 50602 6565
rect 50294 6554 50300 6556
rect 50356 6554 50380 6556
rect 50436 6554 50460 6556
rect 50516 6554 50540 6556
rect 50596 6554 50602 6556
rect 50356 6502 50358 6554
rect 50538 6502 50540 6554
rect 50294 6500 50300 6502
rect 50356 6500 50380 6502
rect 50436 6500 50460 6502
rect 50516 6500 50540 6502
rect 50596 6500 50602 6502
rect 50294 6491 50602 6500
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 65654 6012 65962 6021
rect 65654 6010 65660 6012
rect 65716 6010 65740 6012
rect 65796 6010 65820 6012
rect 65876 6010 65900 6012
rect 65956 6010 65962 6012
rect 65716 5958 65718 6010
rect 65898 5958 65900 6010
rect 65654 5956 65660 5958
rect 65716 5956 65740 5958
rect 65796 5956 65820 5958
rect 65876 5956 65900 5958
rect 65956 5956 65962 5958
rect 65654 5947 65962 5956
rect 50294 5468 50602 5477
rect 50294 5466 50300 5468
rect 50356 5466 50380 5468
rect 50436 5466 50460 5468
rect 50516 5466 50540 5468
rect 50596 5466 50602 5468
rect 50356 5414 50358 5466
rect 50538 5414 50540 5466
rect 50294 5412 50300 5414
rect 50356 5412 50380 5414
rect 50436 5412 50460 5414
rect 50516 5412 50540 5414
rect 50596 5412 50602 5414
rect 50294 5403 50602 5412
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 65654 4924 65962 4933
rect 65654 4922 65660 4924
rect 65716 4922 65740 4924
rect 65796 4922 65820 4924
rect 65876 4922 65900 4924
rect 65956 4922 65962 4924
rect 65716 4870 65718 4922
rect 65898 4870 65900 4922
rect 65654 4868 65660 4870
rect 65716 4868 65740 4870
rect 65796 4868 65820 4870
rect 65876 4868 65900 4870
rect 65956 4868 65962 4870
rect 65654 4859 65962 4868
rect 50294 4380 50602 4389
rect 50294 4378 50300 4380
rect 50356 4378 50380 4380
rect 50436 4378 50460 4380
rect 50516 4378 50540 4380
rect 50596 4378 50602 4380
rect 50356 4326 50358 4378
rect 50538 4326 50540 4378
rect 50294 4324 50300 4326
rect 50356 4324 50380 4326
rect 50436 4324 50460 4326
rect 50516 4324 50540 4326
rect 50596 4324 50602 4326
rect 50294 4315 50602 4324
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 65654 3836 65962 3845
rect 65654 3834 65660 3836
rect 65716 3834 65740 3836
rect 65796 3834 65820 3836
rect 65876 3834 65900 3836
rect 65956 3834 65962 3836
rect 65716 3782 65718 3834
rect 65898 3782 65900 3834
rect 65654 3780 65660 3782
rect 65716 3780 65740 3782
rect 65796 3780 65820 3782
rect 65876 3780 65900 3782
rect 65956 3780 65962 3782
rect 65654 3771 65962 3780
rect 51448 3664 51500 3670
rect 51448 3606 51500 3612
rect 27436 3528 27488 3534
rect 27436 3470 27488 3476
rect 27712 3528 27764 3534
rect 27712 3470 27764 3476
rect 28264 3528 28316 3534
rect 28264 3470 28316 3476
rect 29368 3528 29420 3534
rect 29368 3470 29420 3476
rect 30196 3528 30248 3534
rect 30196 3470 30248 3476
rect 31300 3528 31352 3534
rect 31300 3470 31352 3476
rect 32128 3528 32180 3534
rect 32128 3470 32180 3476
rect 32956 3528 33008 3534
rect 32956 3470 33008 3476
rect 39856 3528 39908 3534
rect 39856 3470 39908 3476
rect 40132 3528 40184 3534
rect 40132 3470 40184 3476
rect 40960 3528 41012 3534
rect 40960 3470 41012 3476
rect 41788 3528 41840 3534
rect 41788 3470 41840 3476
rect 42616 3528 42668 3534
rect 42616 3470 42668 3476
rect 43720 3528 43772 3534
rect 43720 3470 43772 3476
rect 45100 3528 45152 3534
rect 45100 3470 45152 3476
rect 45652 3528 45704 3534
rect 45652 3470 45704 3476
rect 46204 3528 46256 3534
rect 46204 3470 46256 3476
rect 47584 3528 47636 3534
rect 47584 3470 47636 3476
rect 47860 3528 47912 3534
rect 47860 3470 47912 3476
rect 49516 3528 49568 3534
rect 49516 3470 49568 3476
rect 50620 3528 50672 3534
rect 50620 3470 50672 3476
rect 51172 3528 51224 3534
rect 51172 3470 51224 3476
rect 27160 2508 27212 2514
rect 27160 2450 27212 2456
rect 26424 2440 26476 2446
rect 26424 2382 26476 2388
rect 26976 2440 27028 2446
rect 26976 2382 27028 2388
rect 26608 2304 26660 2310
rect 26608 2246 26660 2252
rect 26884 2304 26936 2310
rect 26884 2246 26936 2252
rect 26620 800 26648 2246
rect 26896 800 26924 2246
rect 27172 800 27200 2450
rect 27448 800 27476 3470
rect 27724 800 27752 3470
rect 27988 2848 28040 2854
rect 27988 2790 28040 2796
rect 28000 800 28028 2790
rect 28276 800 28304 3470
rect 28540 2848 28592 2854
rect 28540 2790 28592 2796
rect 29092 2848 29144 2854
rect 29092 2790 29144 2796
rect 28552 800 28580 2790
rect 28816 2440 28868 2446
rect 28816 2382 28868 2388
rect 28828 800 28856 2382
rect 29104 800 29132 2790
rect 29380 800 29408 3470
rect 29920 2848 29972 2854
rect 29920 2790 29972 2796
rect 29644 2440 29696 2446
rect 29644 2382 29696 2388
rect 29656 800 29684 2382
rect 29932 800 29960 2790
rect 30208 800 30236 3470
rect 30472 2848 30524 2854
rect 30472 2790 30524 2796
rect 31024 2848 31076 2854
rect 31024 2790 31076 2796
rect 30484 800 30512 2790
rect 30748 2440 30800 2446
rect 30748 2382 30800 2388
rect 30760 800 30788 2382
rect 31036 800 31064 2790
rect 31312 800 31340 3470
rect 31852 2848 31904 2854
rect 31852 2790 31904 2796
rect 31576 2576 31628 2582
rect 31576 2518 31628 2524
rect 31588 800 31616 2518
rect 31864 800 31892 2790
rect 32140 800 32168 3470
rect 32680 2848 32732 2854
rect 32680 2790 32732 2796
rect 32404 2440 32456 2446
rect 32404 2382 32456 2388
rect 32416 800 32444 2382
rect 32692 800 32720 2790
rect 32968 800 32996 3470
rect 37924 2984 37976 2990
rect 37924 2926 37976 2932
rect 39580 2984 39632 2990
rect 39580 2926 39632 2932
rect 33232 2848 33284 2854
rect 33232 2790 33284 2796
rect 33784 2848 33836 2854
rect 33784 2790 33836 2796
rect 34336 2848 34388 2854
rect 34336 2790 34388 2796
rect 34796 2848 34848 2854
rect 34796 2790 34848 2796
rect 35440 2848 35492 2854
rect 35440 2790 35492 2796
rect 36268 2848 36320 2854
rect 36268 2790 36320 2796
rect 36820 2848 36872 2854
rect 36820 2790 36872 2796
rect 37372 2848 37424 2854
rect 37372 2790 37424 2796
rect 33244 800 33272 2790
rect 33508 2576 33560 2582
rect 33508 2518 33560 2524
rect 33520 800 33548 2518
rect 33796 800 33824 2790
rect 34060 2440 34112 2446
rect 34060 2382 34112 2388
rect 34072 800 34100 2382
rect 34348 800 34376 2790
rect 34612 2440 34664 2446
rect 34612 2382 34664 2388
rect 34624 800 34652 2382
rect 34808 1442 34836 2790
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 35164 2440 35216 2446
rect 35164 2382 35216 2388
rect 34808 1414 34928 1442
rect 34900 800 34928 1414
rect 35176 800 35204 2382
rect 35452 800 35480 2790
rect 35716 2440 35768 2446
rect 35716 2382 35768 2388
rect 35992 2440 36044 2446
rect 35992 2382 36044 2388
rect 35728 800 35756 2382
rect 36004 800 36032 2382
rect 36280 800 36308 2790
rect 36544 2440 36596 2446
rect 36544 2382 36596 2388
rect 36556 800 36584 2382
rect 36832 800 36860 2790
rect 37096 2508 37148 2514
rect 37096 2450 37148 2456
rect 37108 800 37136 2450
rect 37384 800 37412 2790
rect 37648 2440 37700 2446
rect 37648 2382 37700 2388
rect 37660 800 37688 2382
rect 37936 800 37964 2926
rect 38476 2916 38528 2922
rect 38476 2858 38528 2864
rect 38200 2508 38252 2514
rect 38200 2450 38252 2456
rect 38212 800 38240 2450
rect 38488 800 38516 2858
rect 39028 2848 39080 2854
rect 39028 2790 39080 2796
rect 38752 2440 38804 2446
rect 38752 2382 38804 2388
rect 38764 800 38792 2382
rect 39040 800 39068 2790
rect 39304 2576 39356 2582
rect 39304 2518 39356 2524
rect 39316 800 39344 2518
rect 39592 800 39620 2926
rect 39868 800 39896 3470
rect 40144 800 40172 3470
rect 40408 2916 40460 2922
rect 40408 2858 40460 2864
rect 40420 800 40448 2858
rect 40684 2508 40736 2514
rect 40684 2450 40736 2456
rect 40696 800 40724 2450
rect 40972 800 41000 3470
rect 41512 2848 41564 2854
rect 41512 2790 41564 2796
rect 41236 2440 41288 2446
rect 41236 2382 41288 2388
rect 41248 800 41276 2382
rect 41524 800 41552 2790
rect 41800 800 41828 3470
rect 42340 2916 42392 2922
rect 42340 2858 42392 2864
rect 42064 2372 42116 2378
rect 42064 2314 42116 2320
rect 42076 800 42104 2314
rect 42352 800 42380 2858
rect 42628 800 42656 3470
rect 43444 2984 43496 2990
rect 43444 2926 43496 2932
rect 42892 2848 42944 2854
rect 42892 2790 42944 2796
rect 42904 800 42932 2790
rect 43168 2576 43220 2582
rect 43168 2518 43220 2524
rect 43180 800 43208 2518
rect 43456 800 43484 2926
rect 43732 800 43760 3470
rect 44272 2916 44324 2922
rect 44272 2858 44324 2864
rect 43996 2508 44048 2514
rect 43996 2450 44048 2456
rect 44008 800 44036 2450
rect 44284 800 44312 2858
rect 44824 2848 44876 2854
rect 44824 2790 44876 2796
rect 44548 2372 44600 2378
rect 44548 2314 44600 2320
rect 44560 800 44588 2314
rect 44836 800 44864 2790
rect 45112 800 45140 3470
rect 45376 2916 45428 2922
rect 45376 2858 45428 2864
rect 45388 800 45416 2858
rect 45664 800 45692 3470
rect 45928 2508 45980 2514
rect 45928 2450 45980 2456
rect 45940 800 45968 2450
rect 46216 800 46244 3470
rect 47308 2984 47360 2990
rect 47308 2926 47360 2932
rect 46756 2848 46808 2854
rect 46756 2790 46808 2796
rect 46480 2440 46532 2446
rect 46480 2382 46532 2388
rect 46492 800 46520 2382
rect 46768 800 46796 2790
rect 47032 2576 47084 2582
rect 47032 2518 47084 2524
rect 47044 800 47072 2518
rect 47320 800 47348 2926
rect 47596 800 47624 3470
rect 47872 800 47900 3470
rect 49240 2984 49292 2990
rect 49240 2926 49292 2932
rect 48136 2916 48188 2922
rect 48136 2858 48188 2864
rect 48148 800 48176 2858
rect 48688 2848 48740 2854
rect 48688 2790 48740 2796
rect 48412 2508 48464 2514
rect 48412 2450 48464 2456
rect 48424 800 48452 2450
rect 48700 800 48728 2790
rect 48964 2440 49016 2446
rect 48964 2382 49016 2388
rect 48976 800 49004 2382
rect 49252 800 49280 2926
rect 49528 800 49556 3470
rect 50294 3292 50602 3301
rect 50294 3290 50300 3292
rect 50356 3290 50380 3292
rect 50436 3290 50460 3292
rect 50516 3290 50540 3292
rect 50596 3290 50602 3292
rect 50356 3238 50358 3290
rect 50538 3238 50540 3290
rect 50294 3236 50300 3238
rect 50356 3236 50380 3238
rect 50436 3236 50460 3238
rect 50516 3236 50540 3238
rect 50596 3236 50602 3238
rect 50294 3227 50602 3236
rect 50068 2916 50120 2922
rect 50068 2858 50120 2864
rect 49792 2372 49844 2378
rect 49792 2314 49844 2320
rect 49804 800 49832 2314
rect 50080 800 50108 2858
rect 50294 2204 50602 2213
rect 50294 2202 50300 2204
rect 50356 2202 50380 2204
rect 50436 2202 50460 2204
rect 50516 2202 50540 2204
rect 50596 2202 50602 2204
rect 50356 2150 50358 2202
rect 50538 2150 50540 2202
rect 50294 2148 50300 2150
rect 50356 2148 50380 2150
rect 50436 2148 50460 2150
rect 50516 2148 50540 2150
rect 50596 2148 50602 2150
rect 50294 2139 50602 2148
rect 50632 1850 50660 3470
rect 50712 2848 50764 2854
rect 50712 2790 50764 2796
rect 50356 1822 50660 1850
rect 50356 800 50384 1822
rect 50724 1442 50752 2790
rect 50896 2576 50948 2582
rect 50896 2518 50948 2524
rect 50632 1414 50752 1442
rect 50632 800 50660 1414
rect 50908 800 50936 2518
rect 51184 800 51212 3470
rect 51460 800 51488 3606
rect 52828 3528 52880 3534
rect 52828 3470 52880 3476
rect 53380 3528 53432 3534
rect 53380 3470 53432 3476
rect 55312 3528 55364 3534
rect 55312 3470 55364 3476
rect 55588 3528 55640 3534
rect 55588 3470 55640 3476
rect 56416 3528 56468 3534
rect 56416 3470 56468 3476
rect 57244 3528 57296 3534
rect 57244 3470 57296 3476
rect 57520 3528 57572 3534
rect 57520 3470 57572 3476
rect 52552 2916 52604 2922
rect 52552 2858 52604 2864
rect 52000 2848 52052 2854
rect 52000 2790 52052 2796
rect 51724 2508 51776 2514
rect 51724 2450 51776 2456
rect 51736 800 51764 2450
rect 52012 800 52040 2790
rect 52276 2440 52328 2446
rect 52276 2382 52328 2388
rect 52288 800 52316 2382
rect 52564 800 52592 2858
rect 52840 800 52868 3470
rect 53104 2848 53156 2854
rect 53104 2790 53156 2796
rect 53116 800 53144 2790
rect 53392 800 53420 3470
rect 55036 2984 55088 2990
rect 55036 2926 55088 2932
rect 53932 2916 53984 2922
rect 53932 2858 53984 2864
rect 53656 2508 53708 2514
rect 53656 2450 53708 2456
rect 53668 800 53696 2450
rect 53944 800 53972 2858
rect 54484 2848 54536 2854
rect 54484 2790 54536 2796
rect 54208 2372 54260 2378
rect 54208 2314 54260 2320
rect 54220 800 54248 2314
rect 54496 800 54524 2790
rect 54760 2576 54812 2582
rect 54760 2518 54812 2524
rect 54772 800 54800 2518
rect 55048 800 55076 2926
rect 55324 800 55352 3470
rect 55600 800 55628 3470
rect 55864 2848 55916 2854
rect 55864 2790 55916 2796
rect 55876 800 55904 2790
rect 56140 2440 56192 2446
rect 56140 2382 56192 2388
rect 56152 800 56180 2382
rect 56428 800 56456 3470
rect 56968 2848 57020 2854
rect 56968 2790 57020 2796
rect 56692 2576 56744 2582
rect 56692 2518 56744 2524
rect 56704 800 56732 2518
rect 56980 800 57008 2790
rect 57256 800 57284 3470
rect 57428 2508 57480 2514
rect 57428 2450 57480 2456
rect 57440 800 57468 2450
rect 57532 800 57560 3470
rect 57612 2916 57664 2922
rect 57612 2858 57664 2864
rect 57624 800 57652 2858
rect 65654 2748 65962 2757
rect 65654 2746 65660 2748
rect 65716 2746 65740 2748
rect 65796 2746 65820 2748
rect 65876 2746 65900 2748
rect 65956 2746 65962 2748
rect 65716 2694 65718 2746
rect 65898 2694 65900 2746
rect 65654 2692 65660 2694
rect 65716 2692 65740 2694
rect 65796 2692 65820 2694
rect 65876 2692 65900 2694
rect 65956 2692 65962 2694
rect 65654 2683 65962 2692
rect 12346 0 12402 800
rect 12438 0 12494 800
rect 12530 0 12586 800
rect 12622 0 12678 800
rect 12714 0 12770 800
rect 12806 0 12862 800
rect 12898 0 12954 800
rect 12990 0 13046 800
rect 13082 0 13138 800
rect 13174 0 13230 800
rect 13266 0 13322 800
rect 13358 0 13414 800
rect 13450 0 13506 800
rect 13542 0 13598 800
rect 13634 0 13690 800
rect 13726 0 13782 800
rect 13818 0 13874 800
rect 13910 0 13966 800
rect 14002 0 14058 800
rect 14094 0 14150 800
rect 14186 0 14242 800
rect 14278 0 14334 800
rect 14370 0 14426 800
rect 14462 0 14518 800
rect 14554 0 14610 800
rect 14646 0 14702 800
rect 14738 0 14794 800
rect 14830 0 14886 800
rect 14922 0 14978 800
rect 15014 0 15070 800
rect 15106 0 15162 800
rect 15198 0 15254 800
rect 15290 0 15346 800
rect 15382 0 15438 800
rect 15474 0 15530 800
rect 15566 0 15622 800
rect 15658 0 15714 800
rect 15750 0 15806 800
rect 15842 0 15898 800
rect 15934 0 15990 800
rect 16026 0 16082 800
rect 16118 0 16174 800
rect 16210 0 16266 800
rect 16302 0 16358 800
rect 16394 0 16450 800
rect 16486 0 16542 800
rect 16578 0 16634 800
rect 16670 0 16726 800
rect 16762 0 16818 800
rect 16854 0 16910 800
rect 16946 0 17002 800
rect 17038 0 17094 800
rect 17130 0 17186 800
rect 17222 0 17278 800
rect 17314 0 17370 800
rect 17406 0 17462 800
rect 17498 0 17554 800
rect 17590 0 17646 800
rect 17682 0 17738 800
rect 17774 0 17830 800
rect 17866 0 17922 800
rect 17958 0 18014 800
rect 18050 0 18106 800
rect 18142 0 18198 800
rect 18234 0 18290 800
rect 18326 0 18382 800
rect 18418 0 18474 800
rect 18510 0 18566 800
rect 18602 0 18658 800
rect 18694 0 18750 800
rect 18786 0 18842 800
rect 18878 0 18934 800
rect 18970 0 19026 800
rect 19062 0 19118 800
rect 19154 0 19210 800
rect 19246 0 19302 800
rect 19338 0 19394 800
rect 19430 0 19486 800
rect 19522 0 19578 800
rect 19614 0 19670 800
rect 19706 0 19762 800
rect 19798 0 19854 800
rect 19890 0 19946 800
rect 19982 0 20038 800
rect 20074 0 20130 800
rect 20166 0 20222 800
rect 20258 0 20314 800
rect 20350 0 20406 800
rect 20442 0 20498 800
rect 20534 0 20590 800
rect 20626 0 20682 800
rect 20718 0 20774 800
rect 20810 0 20866 800
rect 20902 0 20958 800
rect 20994 0 21050 800
rect 21086 0 21142 800
rect 21178 0 21234 800
rect 21270 0 21326 800
rect 21362 0 21418 800
rect 21454 0 21510 800
rect 21546 0 21602 800
rect 21638 0 21694 800
rect 21730 0 21786 800
rect 21822 0 21878 800
rect 21914 0 21970 800
rect 22006 0 22062 800
rect 22098 0 22154 800
rect 22190 0 22246 800
rect 22282 0 22338 800
rect 22374 0 22430 800
rect 22466 0 22522 800
rect 22558 0 22614 800
rect 22650 0 22706 800
rect 22742 0 22798 800
rect 22834 0 22890 800
rect 22926 0 22982 800
rect 23018 0 23074 800
rect 23110 0 23166 800
rect 23202 0 23258 800
rect 23294 0 23350 800
rect 23386 0 23442 800
rect 23478 0 23534 800
rect 23570 0 23626 800
rect 23662 0 23718 800
rect 23754 0 23810 800
rect 23846 0 23902 800
rect 23938 0 23994 800
rect 24030 0 24086 800
rect 24122 0 24178 800
rect 24214 0 24270 800
rect 24306 0 24362 800
rect 24398 0 24454 800
rect 24490 0 24546 800
rect 24582 0 24638 800
rect 24674 0 24730 800
rect 24766 0 24822 800
rect 24858 0 24914 800
rect 24950 0 25006 800
rect 25042 0 25098 800
rect 25134 0 25190 800
rect 25226 0 25282 800
rect 25318 0 25374 800
rect 25410 0 25466 800
rect 25502 0 25558 800
rect 25594 0 25650 800
rect 25686 0 25742 800
rect 25778 0 25834 800
rect 25870 0 25926 800
rect 25962 0 26018 800
rect 26054 0 26110 800
rect 26146 0 26202 800
rect 26238 0 26294 800
rect 26330 0 26386 800
rect 26422 0 26478 800
rect 26514 0 26570 800
rect 26606 0 26662 800
rect 26698 0 26754 800
rect 26790 0 26846 800
rect 26882 0 26938 800
rect 26974 0 27030 800
rect 27066 0 27122 800
rect 27158 0 27214 800
rect 27250 0 27306 800
rect 27342 0 27398 800
rect 27434 0 27490 800
rect 27526 0 27582 800
rect 27618 0 27674 800
rect 27710 0 27766 800
rect 27802 0 27858 800
rect 27894 0 27950 800
rect 27986 0 28042 800
rect 28078 0 28134 800
rect 28170 0 28226 800
rect 28262 0 28318 800
rect 28354 0 28410 800
rect 28446 0 28502 800
rect 28538 0 28594 800
rect 28630 0 28686 800
rect 28722 0 28778 800
rect 28814 0 28870 800
rect 28906 0 28962 800
rect 28998 0 29054 800
rect 29090 0 29146 800
rect 29182 0 29238 800
rect 29274 0 29330 800
rect 29366 0 29422 800
rect 29458 0 29514 800
rect 29550 0 29606 800
rect 29642 0 29698 800
rect 29734 0 29790 800
rect 29826 0 29882 800
rect 29918 0 29974 800
rect 30010 0 30066 800
rect 30102 0 30158 800
rect 30194 0 30250 800
rect 30286 0 30342 800
rect 30378 0 30434 800
rect 30470 0 30526 800
rect 30562 0 30618 800
rect 30654 0 30710 800
rect 30746 0 30802 800
rect 30838 0 30894 800
rect 30930 0 30986 800
rect 31022 0 31078 800
rect 31114 0 31170 800
rect 31206 0 31262 800
rect 31298 0 31354 800
rect 31390 0 31446 800
rect 31482 0 31538 800
rect 31574 0 31630 800
rect 31666 0 31722 800
rect 31758 0 31814 800
rect 31850 0 31906 800
rect 31942 0 31998 800
rect 32034 0 32090 800
rect 32126 0 32182 800
rect 32218 0 32274 800
rect 32310 0 32366 800
rect 32402 0 32458 800
rect 32494 0 32550 800
rect 32586 0 32642 800
rect 32678 0 32734 800
rect 32770 0 32826 800
rect 32862 0 32918 800
rect 32954 0 33010 800
rect 33046 0 33102 800
rect 33138 0 33194 800
rect 33230 0 33286 800
rect 33322 0 33378 800
rect 33414 0 33470 800
rect 33506 0 33562 800
rect 33598 0 33654 800
rect 33690 0 33746 800
rect 33782 0 33838 800
rect 33874 0 33930 800
rect 33966 0 34022 800
rect 34058 0 34114 800
rect 34150 0 34206 800
rect 34242 0 34298 800
rect 34334 0 34390 800
rect 34426 0 34482 800
rect 34518 0 34574 800
rect 34610 0 34666 800
rect 34702 0 34758 800
rect 34794 0 34850 800
rect 34886 0 34942 800
rect 34978 0 35034 800
rect 35070 0 35126 800
rect 35162 0 35218 800
rect 35254 0 35310 800
rect 35346 0 35402 800
rect 35438 0 35494 800
rect 35530 0 35586 800
rect 35622 0 35678 800
rect 35714 0 35770 800
rect 35806 0 35862 800
rect 35898 0 35954 800
rect 35990 0 36046 800
rect 36082 0 36138 800
rect 36174 0 36230 800
rect 36266 0 36322 800
rect 36358 0 36414 800
rect 36450 0 36506 800
rect 36542 0 36598 800
rect 36634 0 36690 800
rect 36726 0 36782 800
rect 36818 0 36874 800
rect 36910 0 36966 800
rect 37002 0 37058 800
rect 37094 0 37150 800
rect 37186 0 37242 800
rect 37278 0 37334 800
rect 37370 0 37426 800
rect 37462 0 37518 800
rect 37554 0 37610 800
rect 37646 0 37702 800
rect 37738 0 37794 800
rect 37830 0 37886 800
rect 37922 0 37978 800
rect 38014 0 38070 800
rect 38106 0 38162 800
rect 38198 0 38254 800
rect 38290 0 38346 800
rect 38382 0 38438 800
rect 38474 0 38530 800
rect 38566 0 38622 800
rect 38658 0 38714 800
rect 38750 0 38806 800
rect 38842 0 38898 800
rect 38934 0 38990 800
rect 39026 0 39082 800
rect 39118 0 39174 800
rect 39210 0 39266 800
rect 39302 0 39358 800
rect 39394 0 39450 800
rect 39486 0 39542 800
rect 39578 0 39634 800
rect 39670 0 39726 800
rect 39762 0 39818 800
rect 39854 0 39910 800
rect 39946 0 40002 800
rect 40038 0 40094 800
rect 40130 0 40186 800
rect 40222 0 40278 800
rect 40314 0 40370 800
rect 40406 0 40462 800
rect 40498 0 40554 800
rect 40590 0 40646 800
rect 40682 0 40738 800
rect 40774 0 40830 800
rect 40866 0 40922 800
rect 40958 0 41014 800
rect 41050 0 41106 800
rect 41142 0 41198 800
rect 41234 0 41290 800
rect 41326 0 41382 800
rect 41418 0 41474 800
rect 41510 0 41566 800
rect 41602 0 41658 800
rect 41694 0 41750 800
rect 41786 0 41842 800
rect 41878 0 41934 800
rect 41970 0 42026 800
rect 42062 0 42118 800
rect 42154 0 42210 800
rect 42246 0 42302 800
rect 42338 0 42394 800
rect 42430 0 42486 800
rect 42522 0 42578 800
rect 42614 0 42670 800
rect 42706 0 42762 800
rect 42798 0 42854 800
rect 42890 0 42946 800
rect 42982 0 43038 800
rect 43074 0 43130 800
rect 43166 0 43222 800
rect 43258 0 43314 800
rect 43350 0 43406 800
rect 43442 0 43498 800
rect 43534 0 43590 800
rect 43626 0 43682 800
rect 43718 0 43774 800
rect 43810 0 43866 800
rect 43902 0 43958 800
rect 43994 0 44050 800
rect 44086 0 44142 800
rect 44178 0 44234 800
rect 44270 0 44326 800
rect 44362 0 44418 800
rect 44454 0 44510 800
rect 44546 0 44602 800
rect 44638 0 44694 800
rect 44730 0 44786 800
rect 44822 0 44878 800
rect 44914 0 44970 800
rect 45006 0 45062 800
rect 45098 0 45154 800
rect 45190 0 45246 800
rect 45282 0 45338 800
rect 45374 0 45430 800
rect 45466 0 45522 800
rect 45558 0 45614 800
rect 45650 0 45706 800
rect 45742 0 45798 800
rect 45834 0 45890 800
rect 45926 0 45982 800
rect 46018 0 46074 800
rect 46110 0 46166 800
rect 46202 0 46258 800
rect 46294 0 46350 800
rect 46386 0 46442 800
rect 46478 0 46534 800
rect 46570 0 46626 800
rect 46662 0 46718 800
rect 46754 0 46810 800
rect 46846 0 46902 800
rect 46938 0 46994 800
rect 47030 0 47086 800
rect 47122 0 47178 800
rect 47214 0 47270 800
rect 47306 0 47362 800
rect 47398 0 47454 800
rect 47490 0 47546 800
rect 47582 0 47638 800
rect 47674 0 47730 800
rect 47766 0 47822 800
rect 47858 0 47914 800
rect 47950 0 48006 800
rect 48042 0 48098 800
rect 48134 0 48190 800
rect 48226 0 48282 800
rect 48318 0 48374 800
rect 48410 0 48466 800
rect 48502 0 48558 800
rect 48594 0 48650 800
rect 48686 0 48742 800
rect 48778 0 48834 800
rect 48870 0 48926 800
rect 48962 0 49018 800
rect 49054 0 49110 800
rect 49146 0 49202 800
rect 49238 0 49294 800
rect 49330 0 49386 800
rect 49422 0 49478 800
rect 49514 0 49570 800
rect 49606 0 49662 800
rect 49698 0 49754 800
rect 49790 0 49846 800
rect 49882 0 49938 800
rect 49974 0 50030 800
rect 50066 0 50122 800
rect 50158 0 50214 800
rect 50250 0 50306 800
rect 50342 0 50398 800
rect 50434 0 50490 800
rect 50526 0 50582 800
rect 50618 0 50674 800
rect 50710 0 50766 800
rect 50802 0 50858 800
rect 50894 0 50950 800
rect 50986 0 51042 800
rect 51078 0 51134 800
rect 51170 0 51226 800
rect 51262 0 51318 800
rect 51354 0 51410 800
rect 51446 0 51502 800
rect 51538 0 51594 800
rect 51630 0 51686 800
rect 51722 0 51778 800
rect 51814 0 51870 800
rect 51906 0 51962 800
rect 51998 0 52054 800
rect 52090 0 52146 800
rect 52182 0 52238 800
rect 52274 0 52330 800
rect 52366 0 52422 800
rect 52458 0 52514 800
rect 52550 0 52606 800
rect 52642 0 52698 800
rect 52734 0 52790 800
rect 52826 0 52882 800
rect 52918 0 52974 800
rect 53010 0 53066 800
rect 53102 0 53158 800
rect 53194 0 53250 800
rect 53286 0 53342 800
rect 53378 0 53434 800
rect 53470 0 53526 800
rect 53562 0 53618 800
rect 53654 0 53710 800
rect 53746 0 53802 800
rect 53838 0 53894 800
rect 53930 0 53986 800
rect 54022 0 54078 800
rect 54114 0 54170 800
rect 54206 0 54262 800
rect 54298 0 54354 800
rect 54390 0 54446 800
rect 54482 0 54538 800
rect 54574 0 54630 800
rect 54666 0 54722 800
rect 54758 0 54814 800
rect 54850 0 54906 800
rect 54942 0 54998 800
rect 55034 0 55090 800
rect 55126 0 55182 800
rect 55218 0 55274 800
rect 55310 0 55366 800
rect 55402 0 55458 800
rect 55494 0 55550 800
rect 55586 0 55642 800
rect 55678 0 55734 800
rect 55770 0 55826 800
rect 55862 0 55918 800
rect 55954 0 56010 800
rect 56046 0 56102 800
rect 56138 0 56194 800
rect 56230 0 56286 800
rect 56322 0 56378 800
rect 56414 0 56470 800
rect 56506 0 56562 800
rect 56598 0 56654 800
rect 56690 0 56746 800
rect 56782 0 56838 800
rect 56874 0 56930 800
rect 56966 0 57022 800
rect 57058 0 57114 800
rect 57150 0 57206 800
rect 57242 0 57298 800
rect 57334 0 57390 800
rect 57426 0 57482 800
rect 57518 0 57574 800
rect 57610 0 57666 800
<< via2 >>
rect 19580 57690 19636 57692
rect 19660 57690 19716 57692
rect 19740 57690 19796 57692
rect 19820 57690 19876 57692
rect 19580 57638 19626 57690
rect 19626 57638 19636 57690
rect 19660 57638 19690 57690
rect 19690 57638 19702 57690
rect 19702 57638 19716 57690
rect 19740 57638 19754 57690
rect 19754 57638 19766 57690
rect 19766 57638 19796 57690
rect 19820 57638 19830 57690
rect 19830 57638 19876 57690
rect 19580 57636 19636 57638
rect 19660 57636 19716 57638
rect 19740 57636 19796 57638
rect 19820 57636 19876 57638
rect 4220 57146 4276 57148
rect 4300 57146 4356 57148
rect 4380 57146 4436 57148
rect 4460 57146 4516 57148
rect 4220 57094 4266 57146
rect 4266 57094 4276 57146
rect 4300 57094 4330 57146
rect 4330 57094 4342 57146
rect 4342 57094 4356 57146
rect 4380 57094 4394 57146
rect 4394 57094 4406 57146
rect 4406 57094 4436 57146
rect 4460 57094 4470 57146
rect 4470 57094 4516 57146
rect 4220 57092 4276 57094
rect 4300 57092 4356 57094
rect 4380 57092 4436 57094
rect 4460 57092 4516 57094
rect 34940 57146 34996 57148
rect 35020 57146 35076 57148
rect 35100 57146 35156 57148
rect 35180 57146 35236 57148
rect 34940 57094 34986 57146
rect 34986 57094 34996 57146
rect 35020 57094 35050 57146
rect 35050 57094 35062 57146
rect 35062 57094 35076 57146
rect 35100 57094 35114 57146
rect 35114 57094 35126 57146
rect 35126 57094 35156 57146
rect 35180 57094 35190 57146
rect 35190 57094 35236 57146
rect 34940 57092 34996 57094
rect 35020 57092 35076 57094
rect 35100 57092 35156 57094
rect 35180 57092 35236 57094
rect 50300 57690 50356 57692
rect 50380 57690 50436 57692
rect 50460 57690 50516 57692
rect 50540 57690 50596 57692
rect 50300 57638 50346 57690
rect 50346 57638 50356 57690
rect 50380 57638 50410 57690
rect 50410 57638 50422 57690
rect 50422 57638 50436 57690
rect 50460 57638 50474 57690
rect 50474 57638 50486 57690
rect 50486 57638 50516 57690
rect 50540 57638 50550 57690
rect 50550 57638 50596 57690
rect 50300 57636 50356 57638
rect 50380 57636 50436 57638
rect 50460 57636 50516 57638
rect 50540 57636 50596 57638
rect 65660 57146 65716 57148
rect 65740 57146 65796 57148
rect 65820 57146 65876 57148
rect 65900 57146 65956 57148
rect 65660 57094 65706 57146
rect 65706 57094 65716 57146
rect 65740 57094 65770 57146
rect 65770 57094 65782 57146
rect 65782 57094 65796 57146
rect 65820 57094 65834 57146
rect 65834 57094 65846 57146
rect 65846 57094 65876 57146
rect 65900 57094 65910 57146
rect 65910 57094 65956 57146
rect 65660 57092 65716 57094
rect 65740 57092 65796 57094
rect 65820 57092 65876 57094
rect 65900 57092 65956 57094
rect 19580 56602 19636 56604
rect 19660 56602 19716 56604
rect 19740 56602 19796 56604
rect 19820 56602 19876 56604
rect 19580 56550 19626 56602
rect 19626 56550 19636 56602
rect 19660 56550 19690 56602
rect 19690 56550 19702 56602
rect 19702 56550 19716 56602
rect 19740 56550 19754 56602
rect 19754 56550 19766 56602
rect 19766 56550 19796 56602
rect 19820 56550 19830 56602
rect 19830 56550 19876 56602
rect 19580 56548 19636 56550
rect 19660 56548 19716 56550
rect 19740 56548 19796 56550
rect 19820 56548 19876 56550
rect 50300 56602 50356 56604
rect 50380 56602 50436 56604
rect 50460 56602 50516 56604
rect 50540 56602 50596 56604
rect 50300 56550 50346 56602
rect 50346 56550 50356 56602
rect 50380 56550 50410 56602
rect 50410 56550 50422 56602
rect 50422 56550 50436 56602
rect 50460 56550 50474 56602
rect 50474 56550 50486 56602
rect 50486 56550 50516 56602
rect 50540 56550 50550 56602
rect 50550 56550 50596 56602
rect 50300 56548 50356 56550
rect 50380 56548 50436 56550
rect 50460 56548 50516 56550
rect 50540 56548 50596 56550
rect 4220 56058 4276 56060
rect 4300 56058 4356 56060
rect 4380 56058 4436 56060
rect 4460 56058 4516 56060
rect 4220 56006 4266 56058
rect 4266 56006 4276 56058
rect 4300 56006 4330 56058
rect 4330 56006 4342 56058
rect 4342 56006 4356 56058
rect 4380 56006 4394 56058
rect 4394 56006 4406 56058
rect 4406 56006 4436 56058
rect 4460 56006 4470 56058
rect 4470 56006 4516 56058
rect 4220 56004 4276 56006
rect 4300 56004 4356 56006
rect 4380 56004 4436 56006
rect 4460 56004 4516 56006
rect 34940 56058 34996 56060
rect 35020 56058 35076 56060
rect 35100 56058 35156 56060
rect 35180 56058 35236 56060
rect 34940 56006 34986 56058
rect 34986 56006 34996 56058
rect 35020 56006 35050 56058
rect 35050 56006 35062 56058
rect 35062 56006 35076 56058
rect 35100 56006 35114 56058
rect 35114 56006 35126 56058
rect 35126 56006 35156 56058
rect 35180 56006 35190 56058
rect 35190 56006 35236 56058
rect 34940 56004 34996 56006
rect 35020 56004 35076 56006
rect 35100 56004 35156 56006
rect 35180 56004 35236 56006
rect 65660 56058 65716 56060
rect 65740 56058 65796 56060
rect 65820 56058 65876 56060
rect 65900 56058 65956 56060
rect 65660 56006 65706 56058
rect 65706 56006 65716 56058
rect 65740 56006 65770 56058
rect 65770 56006 65782 56058
rect 65782 56006 65796 56058
rect 65820 56006 65834 56058
rect 65834 56006 65846 56058
rect 65846 56006 65876 56058
rect 65900 56006 65910 56058
rect 65910 56006 65956 56058
rect 65660 56004 65716 56006
rect 65740 56004 65796 56006
rect 65820 56004 65876 56006
rect 65900 56004 65956 56006
rect 19580 55514 19636 55516
rect 19660 55514 19716 55516
rect 19740 55514 19796 55516
rect 19820 55514 19876 55516
rect 19580 55462 19626 55514
rect 19626 55462 19636 55514
rect 19660 55462 19690 55514
rect 19690 55462 19702 55514
rect 19702 55462 19716 55514
rect 19740 55462 19754 55514
rect 19754 55462 19766 55514
rect 19766 55462 19796 55514
rect 19820 55462 19830 55514
rect 19830 55462 19876 55514
rect 19580 55460 19636 55462
rect 19660 55460 19716 55462
rect 19740 55460 19796 55462
rect 19820 55460 19876 55462
rect 50300 55514 50356 55516
rect 50380 55514 50436 55516
rect 50460 55514 50516 55516
rect 50540 55514 50596 55516
rect 50300 55462 50346 55514
rect 50346 55462 50356 55514
rect 50380 55462 50410 55514
rect 50410 55462 50422 55514
rect 50422 55462 50436 55514
rect 50460 55462 50474 55514
rect 50474 55462 50486 55514
rect 50486 55462 50516 55514
rect 50540 55462 50550 55514
rect 50550 55462 50596 55514
rect 50300 55460 50356 55462
rect 50380 55460 50436 55462
rect 50460 55460 50516 55462
rect 50540 55460 50596 55462
rect 4220 54970 4276 54972
rect 4300 54970 4356 54972
rect 4380 54970 4436 54972
rect 4460 54970 4516 54972
rect 4220 54918 4266 54970
rect 4266 54918 4276 54970
rect 4300 54918 4330 54970
rect 4330 54918 4342 54970
rect 4342 54918 4356 54970
rect 4380 54918 4394 54970
rect 4394 54918 4406 54970
rect 4406 54918 4436 54970
rect 4460 54918 4470 54970
rect 4470 54918 4516 54970
rect 4220 54916 4276 54918
rect 4300 54916 4356 54918
rect 4380 54916 4436 54918
rect 4460 54916 4516 54918
rect 34940 54970 34996 54972
rect 35020 54970 35076 54972
rect 35100 54970 35156 54972
rect 35180 54970 35236 54972
rect 34940 54918 34986 54970
rect 34986 54918 34996 54970
rect 35020 54918 35050 54970
rect 35050 54918 35062 54970
rect 35062 54918 35076 54970
rect 35100 54918 35114 54970
rect 35114 54918 35126 54970
rect 35126 54918 35156 54970
rect 35180 54918 35190 54970
rect 35190 54918 35236 54970
rect 34940 54916 34996 54918
rect 35020 54916 35076 54918
rect 35100 54916 35156 54918
rect 35180 54916 35236 54918
rect 65660 54970 65716 54972
rect 65740 54970 65796 54972
rect 65820 54970 65876 54972
rect 65900 54970 65956 54972
rect 65660 54918 65706 54970
rect 65706 54918 65716 54970
rect 65740 54918 65770 54970
rect 65770 54918 65782 54970
rect 65782 54918 65796 54970
rect 65820 54918 65834 54970
rect 65834 54918 65846 54970
rect 65846 54918 65876 54970
rect 65900 54918 65910 54970
rect 65910 54918 65956 54970
rect 65660 54916 65716 54918
rect 65740 54916 65796 54918
rect 65820 54916 65876 54918
rect 65900 54916 65956 54918
rect 19580 54426 19636 54428
rect 19660 54426 19716 54428
rect 19740 54426 19796 54428
rect 19820 54426 19876 54428
rect 19580 54374 19626 54426
rect 19626 54374 19636 54426
rect 19660 54374 19690 54426
rect 19690 54374 19702 54426
rect 19702 54374 19716 54426
rect 19740 54374 19754 54426
rect 19754 54374 19766 54426
rect 19766 54374 19796 54426
rect 19820 54374 19830 54426
rect 19830 54374 19876 54426
rect 19580 54372 19636 54374
rect 19660 54372 19716 54374
rect 19740 54372 19796 54374
rect 19820 54372 19876 54374
rect 50300 54426 50356 54428
rect 50380 54426 50436 54428
rect 50460 54426 50516 54428
rect 50540 54426 50596 54428
rect 50300 54374 50346 54426
rect 50346 54374 50356 54426
rect 50380 54374 50410 54426
rect 50410 54374 50422 54426
rect 50422 54374 50436 54426
rect 50460 54374 50474 54426
rect 50474 54374 50486 54426
rect 50486 54374 50516 54426
rect 50540 54374 50550 54426
rect 50550 54374 50596 54426
rect 50300 54372 50356 54374
rect 50380 54372 50436 54374
rect 50460 54372 50516 54374
rect 50540 54372 50596 54374
rect 4220 53882 4276 53884
rect 4300 53882 4356 53884
rect 4380 53882 4436 53884
rect 4460 53882 4516 53884
rect 4220 53830 4266 53882
rect 4266 53830 4276 53882
rect 4300 53830 4330 53882
rect 4330 53830 4342 53882
rect 4342 53830 4356 53882
rect 4380 53830 4394 53882
rect 4394 53830 4406 53882
rect 4406 53830 4436 53882
rect 4460 53830 4470 53882
rect 4470 53830 4516 53882
rect 4220 53828 4276 53830
rect 4300 53828 4356 53830
rect 4380 53828 4436 53830
rect 4460 53828 4516 53830
rect 34940 53882 34996 53884
rect 35020 53882 35076 53884
rect 35100 53882 35156 53884
rect 35180 53882 35236 53884
rect 34940 53830 34986 53882
rect 34986 53830 34996 53882
rect 35020 53830 35050 53882
rect 35050 53830 35062 53882
rect 35062 53830 35076 53882
rect 35100 53830 35114 53882
rect 35114 53830 35126 53882
rect 35126 53830 35156 53882
rect 35180 53830 35190 53882
rect 35190 53830 35236 53882
rect 34940 53828 34996 53830
rect 35020 53828 35076 53830
rect 35100 53828 35156 53830
rect 35180 53828 35236 53830
rect 65660 53882 65716 53884
rect 65740 53882 65796 53884
rect 65820 53882 65876 53884
rect 65900 53882 65956 53884
rect 65660 53830 65706 53882
rect 65706 53830 65716 53882
rect 65740 53830 65770 53882
rect 65770 53830 65782 53882
rect 65782 53830 65796 53882
rect 65820 53830 65834 53882
rect 65834 53830 65846 53882
rect 65846 53830 65876 53882
rect 65900 53830 65910 53882
rect 65910 53830 65956 53882
rect 65660 53828 65716 53830
rect 65740 53828 65796 53830
rect 65820 53828 65876 53830
rect 65900 53828 65956 53830
rect 19580 53338 19636 53340
rect 19660 53338 19716 53340
rect 19740 53338 19796 53340
rect 19820 53338 19876 53340
rect 19580 53286 19626 53338
rect 19626 53286 19636 53338
rect 19660 53286 19690 53338
rect 19690 53286 19702 53338
rect 19702 53286 19716 53338
rect 19740 53286 19754 53338
rect 19754 53286 19766 53338
rect 19766 53286 19796 53338
rect 19820 53286 19830 53338
rect 19830 53286 19876 53338
rect 19580 53284 19636 53286
rect 19660 53284 19716 53286
rect 19740 53284 19796 53286
rect 19820 53284 19876 53286
rect 50300 53338 50356 53340
rect 50380 53338 50436 53340
rect 50460 53338 50516 53340
rect 50540 53338 50596 53340
rect 50300 53286 50346 53338
rect 50346 53286 50356 53338
rect 50380 53286 50410 53338
rect 50410 53286 50422 53338
rect 50422 53286 50436 53338
rect 50460 53286 50474 53338
rect 50474 53286 50486 53338
rect 50486 53286 50516 53338
rect 50540 53286 50550 53338
rect 50550 53286 50596 53338
rect 50300 53284 50356 53286
rect 50380 53284 50436 53286
rect 50460 53284 50516 53286
rect 50540 53284 50596 53286
rect 4220 52794 4276 52796
rect 4300 52794 4356 52796
rect 4380 52794 4436 52796
rect 4460 52794 4516 52796
rect 4220 52742 4266 52794
rect 4266 52742 4276 52794
rect 4300 52742 4330 52794
rect 4330 52742 4342 52794
rect 4342 52742 4356 52794
rect 4380 52742 4394 52794
rect 4394 52742 4406 52794
rect 4406 52742 4436 52794
rect 4460 52742 4470 52794
rect 4470 52742 4516 52794
rect 4220 52740 4276 52742
rect 4300 52740 4356 52742
rect 4380 52740 4436 52742
rect 4460 52740 4516 52742
rect 34940 52794 34996 52796
rect 35020 52794 35076 52796
rect 35100 52794 35156 52796
rect 35180 52794 35236 52796
rect 34940 52742 34986 52794
rect 34986 52742 34996 52794
rect 35020 52742 35050 52794
rect 35050 52742 35062 52794
rect 35062 52742 35076 52794
rect 35100 52742 35114 52794
rect 35114 52742 35126 52794
rect 35126 52742 35156 52794
rect 35180 52742 35190 52794
rect 35190 52742 35236 52794
rect 34940 52740 34996 52742
rect 35020 52740 35076 52742
rect 35100 52740 35156 52742
rect 35180 52740 35236 52742
rect 65660 52794 65716 52796
rect 65740 52794 65796 52796
rect 65820 52794 65876 52796
rect 65900 52794 65956 52796
rect 65660 52742 65706 52794
rect 65706 52742 65716 52794
rect 65740 52742 65770 52794
rect 65770 52742 65782 52794
rect 65782 52742 65796 52794
rect 65820 52742 65834 52794
rect 65834 52742 65846 52794
rect 65846 52742 65876 52794
rect 65900 52742 65910 52794
rect 65910 52742 65956 52794
rect 65660 52740 65716 52742
rect 65740 52740 65796 52742
rect 65820 52740 65876 52742
rect 65900 52740 65956 52742
rect 19580 52250 19636 52252
rect 19660 52250 19716 52252
rect 19740 52250 19796 52252
rect 19820 52250 19876 52252
rect 19580 52198 19626 52250
rect 19626 52198 19636 52250
rect 19660 52198 19690 52250
rect 19690 52198 19702 52250
rect 19702 52198 19716 52250
rect 19740 52198 19754 52250
rect 19754 52198 19766 52250
rect 19766 52198 19796 52250
rect 19820 52198 19830 52250
rect 19830 52198 19876 52250
rect 19580 52196 19636 52198
rect 19660 52196 19716 52198
rect 19740 52196 19796 52198
rect 19820 52196 19876 52198
rect 50300 52250 50356 52252
rect 50380 52250 50436 52252
rect 50460 52250 50516 52252
rect 50540 52250 50596 52252
rect 50300 52198 50346 52250
rect 50346 52198 50356 52250
rect 50380 52198 50410 52250
rect 50410 52198 50422 52250
rect 50422 52198 50436 52250
rect 50460 52198 50474 52250
rect 50474 52198 50486 52250
rect 50486 52198 50516 52250
rect 50540 52198 50550 52250
rect 50550 52198 50596 52250
rect 50300 52196 50356 52198
rect 50380 52196 50436 52198
rect 50460 52196 50516 52198
rect 50540 52196 50596 52198
rect 4220 51706 4276 51708
rect 4300 51706 4356 51708
rect 4380 51706 4436 51708
rect 4460 51706 4516 51708
rect 4220 51654 4266 51706
rect 4266 51654 4276 51706
rect 4300 51654 4330 51706
rect 4330 51654 4342 51706
rect 4342 51654 4356 51706
rect 4380 51654 4394 51706
rect 4394 51654 4406 51706
rect 4406 51654 4436 51706
rect 4460 51654 4470 51706
rect 4470 51654 4516 51706
rect 4220 51652 4276 51654
rect 4300 51652 4356 51654
rect 4380 51652 4436 51654
rect 4460 51652 4516 51654
rect 34940 51706 34996 51708
rect 35020 51706 35076 51708
rect 35100 51706 35156 51708
rect 35180 51706 35236 51708
rect 34940 51654 34986 51706
rect 34986 51654 34996 51706
rect 35020 51654 35050 51706
rect 35050 51654 35062 51706
rect 35062 51654 35076 51706
rect 35100 51654 35114 51706
rect 35114 51654 35126 51706
rect 35126 51654 35156 51706
rect 35180 51654 35190 51706
rect 35190 51654 35236 51706
rect 34940 51652 34996 51654
rect 35020 51652 35076 51654
rect 35100 51652 35156 51654
rect 35180 51652 35236 51654
rect 65660 51706 65716 51708
rect 65740 51706 65796 51708
rect 65820 51706 65876 51708
rect 65900 51706 65956 51708
rect 65660 51654 65706 51706
rect 65706 51654 65716 51706
rect 65740 51654 65770 51706
rect 65770 51654 65782 51706
rect 65782 51654 65796 51706
rect 65820 51654 65834 51706
rect 65834 51654 65846 51706
rect 65846 51654 65876 51706
rect 65900 51654 65910 51706
rect 65910 51654 65956 51706
rect 65660 51652 65716 51654
rect 65740 51652 65796 51654
rect 65820 51652 65876 51654
rect 65900 51652 65956 51654
rect 19580 51162 19636 51164
rect 19660 51162 19716 51164
rect 19740 51162 19796 51164
rect 19820 51162 19876 51164
rect 19580 51110 19626 51162
rect 19626 51110 19636 51162
rect 19660 51110 19690 51162
rect 19690 51110 19702 51162
rect 19702 51110 19716 51162
rect 19740 51110 19754 51162
rect 19754 51110 19766 51162
rect 19766 51110 19796 51162
rect 19820 51110 19830 51162
rect 19830 51110 19876 51162
rect 19580 51108 19636 51110
rect 19660 51108 19716 51110
rect 19740 51108 19796 51110
rect 19820 51108 19876 51110
rect 50300 51162 50356 51164
rect 50380 51162 50436 51164
rect 50460 51162 50516 51164
rect 50540 51162 50596 51164
rect 50300 51110 50346 51162
rect 50346 51110 50356 51162
rect 50380 51110 50410 51162
rect 50410 51110 50422 51162
rect 50422 51110 50436 51162
rect 50460 51110 50474 51162
rect 50474 51110 50486 51162
rect 50486 51110 50516 51162
rect 50540 51110 50550 51162
rect 50550 51110 50596 51162
rect 50300 51108 50356 51110
rect 50380 51108 50436 51110
rect 50460 51108 50516 51110
rect 50540 51108 50596 51110
rect 4220 50618 4276 50620
rect 4300 50618 4356 50620
rect 4380 50618 4436 50620
rect 4460 50618 4516 50620
rect 4220 50566 4266 50618
rect 4266 50566 4276 50618
rect 4300 50566 4330 50618
rect 4330 50566 4342 50618
rect 4342 50566 4356 50618
rect 4380 50566 4394 50618
rect 4394 50566 4406 50618
rect 4406 50566 4436 50618
rect 4460 50566 4470 50618
rect 4470 50566 4516 50618
rect 4220 50564 4276 50566
rect 4300 50564 4356 50566
rect 4380 50564 4436 50566
rect 4460 50564 4516 50566
rect 34940 50618 34996 50620
rect 35020 50618 35076 50620
rect 35100 50618 35156 50620
rect 35180 50618 35236 50620
rect 34940 50566 34986 50618
rect 34986 50566 34996 50618
rect 35020 50566 35050 50618
rect 35050 50566 35062 50618
rect 35062 50566 35076 50618
rect 35100 50566 35114 50618
rect 35114 50566 35126 50618
rect 35126 50566 35156 50618
rect 35180 50566 35190 50618
rect 35190 50566 35236 50618
rect 34940 50564 34996 50566
rect 35020 50564 35076 50566
rect 35100 50564 35156 50566
rect 35180 50564 35236 50566
rect 65660 50618 65716 50620
rect 65740 50618 65796 50620
rect 65820 50618 65876 50620
rect 65900 50618 65956 50620
rect 65660 50566 65706 50618
rect 65706 50566 65716 50618
rect 65740 50566 65770 50618
rect 65770 50566 65782 50618
rect 65782 50566 65796 50618
rect 65820 50566 65834 50618
rect 65834 50566 65846 50618
rect 65846 50566 65876 50618
rect 65900 50566 65910 50618
rect 65910 50566 65956 50618
rect 65660 50564 65716 50566
rect 65740 50564 65796 50566
rect 65820 50564 65876 50566
rect 65900 50564 65956 50566
rect 19580 50074 19636 50076
rect 19660 50074 19716 50076
rect 19740 50074 19796 50076
rect 19820 50074 19876 50076
rect 19580 50022 19626 50074
rect 19626 50022 19636 50074
rect 19660 50022 19690 50074
rect 19690 50022 19702 50074
rect 19702 50022 19716 50074
rect 19740 50022 19754 50074
rect 19754 50022 19766 50074
rect 19766 50022 19796 50074
rect 19820 50022 19830 50074
rect 19830 50022 19876 50074
rect 19580 50020 19636 50022
rect 19660 50020 19716 50022
rect 19740 50020 19796 50022
rect 19820 50020 19876 50022
rect 50300 50074 50356 50076
rect 50380 50074 50436 50076
rect 50460 50074 50516 50076
rect 50540 50074 50596 50076
rect 50300 50022 50346 50074
rect 50346 50022 50356 50074
rect 50380 50022 50410 50074
rect 50410 50022 50422 50074
rect 50422 50022 50436 50074
rect 50460 50022 50474 50074
rect 50474 50022 50486 50074
rect 50486 50022 50516 50074
rect 50540 50022 50550 50074
rect 50550 50022 50596 50074
rect 50300 50020 50356 50022
rect 50380 50020 50436 50022
rect 50460 50020 50516 50022
rect 50540 50020 50596 50022
rect 4220 49530 4276 49532
rect 4300 49530 4356 49532
rect 4380 49530 4436 49532
rect 4460 49530 4516 49532
rect 4220 49478 4266 49530
rect 4266 49478 4276 49530
rect 4300 49478 4330 49530
rect 4330 49478 4342 49530
rect 4342 49478 4356 49530
rect 4380 49478 4394 49530
rect 4394 49478 4406 49530
rect 4406 49478 4436 49530
rect 4460 49478 4470 49530
rect 4470 49478 4516 49530
rect 4220 49476 4276 49478
rect 4300 49476 4356 49478
rect 4380 49476 4436 49478
rect 4460 49476 4516 49478
rect 34940 49530 34996 49532
rect 35020 49530 35076 49532
rect 35100 49530 35156 49532
rect 35180 49530 35236 49532
rect 34940 49478 34986 49530
rect 34986 49478 34996 49530
rect 35020 49478 35050 49530
rect 35050 49478 35062 49530
rect 35062 49478 35076 49530
rect 35100 49478 35114 49530
rect 35114 49478 35126 49530
rect 35126 49478 35156 49530
rect 35180 49478 35190 49530
rect 35190 49478 35236 49530
rect 34940 49476 34996 49478
rect 35020 49476 35076 49478
rect 35100 49476 35156 49478
rect 35180 49476 35236 49478
rect 65660 49530 65716 49532
rect 65740 49530 65796 49532
rect 65820 49530 65876 49532
rect 65900 49530 65956 49532
rect 65660 49478 65706 49530
rect 65706 49478 65716 49530
rect 65740 49478 65770 49530
rect 65770 49478 65782 49530
rect 65782 49478 65796 49530
rect 65820 49478 65834 49530
rect 65834 49478 65846 49530
rect 65846 49478 65876 49530
rect 65900 49478 65910 49530
rect 65910 49478 65956 49530
rect 65660 49476 65716 49478
rect 65740 49476 65796 49478
rect 65820 49476 65876 49478
rect 65900 49476 65956 49478
rect 19580 48986 19636 48988
rect 19660 48986 19716 48988
rect 19740 48986 19796 48988
rect 19820 48986 19876 48988
rect 19580 48934 19626 48986
rect 19626 48934 19636 48986
rect 19660 48934 19690 48986
rect 19690 48934 19702 48986
rect 19702 48934 19716 48986
rect 19740 48934 19754 48986
rect 19754 48934 19766 48986
rect 19766 48934 19796 48986
rect 19820 48934 19830 48986
rect 19830 48934 19876 48986
rect 19580 48932 19636 48934
rect 19660 48932 19716 48934
rect 19740 48932 19796 48934
rect 19820 48932 19876 48934
rect 50300 48986 50356 48988
rect 50380 48986 50436 48988
rect 50460 48986 50516 48988
rect 50540 48986 50596 48988
rect 50300 48934 50346 48986
rect 50346 48934 50356 48986
rect 50380 48934 50410 48986
rect 50410 48934 50422 48986
rect 50422 48934 50436 48986
rect 50460 48934 50474 48986
rect 50474 48934 50486 48986
rect 50486 48934 50516 48986
rect 50540 48934 50550 48986
rect 50550 48934 50596 48986
rect 50300 48932 50356 48934
rect 50380 48932 50436 48934
rect 50460 48932 50516 48934
rect 50540 48932 50596 48934
rect 4220 48442 4276 48444
rect 4300 48442 4356 48444
rect 4380 48442 4436 48444
rect 4460 48442 4516 48444
rect 4220 48390 4266 48442
rect 4266 48390 4276 48442
rect 4300 48390 4330 48442
rect 4330 48390 4342 48442
rect 4342 48390 4356 48442
rect 4380 48390 4394 48442
rect 4394 48390 4406 48442
rect 4406 48390 4436 48442
rect 4460 48390 4470 48442
rect 4470 48390 4516 48442
rect 4220 48388 4276 48390
rect 4300 48388 4356 48390
rect 4380 48388 4436 48390
rect 4460 48388 4516 48390
rect 34940 48442 34996 48444
rect 35020 48442 35076 48444
rect 35100 48442 35156 48444
rect 35180 48442 35236 48444
rect 34940 48390 34986 48442
rect 34986 48390 34996 48442
rect 35020 48390 35050 48442
rect 35050 48390 35062 48442
rect 35062 48390 35076 48442
rect 35100 48390 35114 48442
rect 35114 48390 35126 48442
rect 35126 48390 35156 48442
rect 35180 48390 35190 48442
rect 35190 48390 35236 48442
rect 34940 48388 34996 48390
rect 35020 48388 35076 48390
rect 35100 48388 35156 48390
rect 35180 48388 35236 48390
rect 65660 48442 65716 48444
rect 65740 48442 65796 48444
rect 65820 48442 65876 48444
rect 65900 48442 65956 48444
rect 65660 48390 65706 48442
rect 65706 48390 65716 48442
rect 65740 48390 65770 48442
rect 65770 48390 65782 48442
rect 65782 48390 65796 48442
rect 65820 48390 65834 48442
rect 65834 48390 65846 48442
rect 65846 48390 65876 48442
rect 65900 48390 65910 48442
rect 65910 48390 65956 48442
rect 65660 48388 65716 48390
rect 65740 48388 65796 48390
rect 65820 48388 65876 48390
rect 65900 48388 65956 48390
rect 19580 47898 19636 47900
rect 19660 47898 19716 47900
rect 19740 47898 19796 47900
rect 19820 47898 19876 47900
rect 19580 47846 19626 47898
rect 19626 47846 19636 47898
rect 19660 47846 19690 47898
rect 19690 47846 19702 47898
rect 19702 47846 19716 47898
rect 19740 47846 19754 47898
rect 19754 47846 19766 47898
rect 19766 47846 19796 47898
rect 19820 47846 19830 47898
rect 19830 47846 19876 47898
rect 19580 47844 19636 47846
rect 19660 47844 19716 47846
rect 19740 47844 19796 47846
rect 19820 47844 19876 47846
rect 50300 47898 50356 47900
rect 50380 47898 50436 47900
rect 50460 47898 50516 47900
rect 50540 47898 50596 47900
rect 50300 47846 50346 47898
rect 50346 47846 50356 47898
rect 50380 47846 50410 47898
rect 50410 47846 50422 47898
rect 50422 47846 50436 47898
rect 50460 47846 50474 47898
rect 50474 47846 50486 47898
rect 50486 47846 50516 47898
rect 50540 47846 50550 47898
rect 50550 47846 50596 47898
rect 50300 47844 50356 47846
rect 50380 47844 50436 47846
rect 50460 47844 50516 47846
rect 50540 47844 50596 47846
rect 4220 47354 4276 47356
rect 4300 47354 4356 47356
rect 4380 47354 4436 47356
rect 4460 47354 4516 47356
rect 4220 47302 4266 47354
rect 4266 47302 4276 47354
rect 4300 47302 4330 47354
rect 4330 47302 4342 47354
rect 4342 47302 4356 47354
rect 4380 47302 4394 47354
rect 4394 47302 4406 47354
rect 4406 47302 4436 47354
rect 4460 47302 4470 47354
rect 4470 47302 4516 47354
rect 4220 47300 4276 47302
rect 4300 47300 4356 47302
rect 4380 47300 4436 47302
rect 4460 47300 4516 47302
rect 34940 47354 34996 47356
rect 35020 47354 35076 47356
rect 35100 47354 35156 47356
rect 35180 47354 35236 47356
rect 34940 47302 34986 47354
rect 34986 47302 34996 47354
rect 35020 47302 35050 47354
rect 35050 47302 35062 47354
rect 35062 47302 35076 47354
rect 35100 47302 35114 47354
rect 35114 47302 35126 47354
rect 35126 47302 35156 47354
rect 35180 47302 35190 47354
rect 35190 47302 35236 47354
rect 34940 47300 34996 47302
rect 35020 47300 35076 47302
rect 35100 47300 35156 47302
rect 35180 47300 35236 47302
rect 65660 47354 65716 47356
rect 65740 47354 65796 47356
rect 65820 47354 65876 47356
rect 65900 47354 65956 47356
rect 65660 47302 65706 47354
rect 65706 47302 65716 47354
rect 65740 47302 65770 47354
rect 65770 47302 65782 47354
rect 65782 47302 65796 47354
rect 65820 47302 65834 47354
rect 65834 47302 65846 47354
rect 65846 47302 65876 47354
rect 65900 47302 65910 47354
rect 65910 47302 65956 47354
rect 65660 47300 65716 47302
rect 65740 47300 65796 47302
rect 65820 47300 65876 47302
rect 65900 47300 65956 47302
rect 19580 46810 19636 46812
rect 19660 46810 19716 46812
rect 19740 46810 19796 46812
rect 19820 46810 19876 46812
rect 19580 46758 19626 46810
rect 19626 46758 19636 46810
rect 19660 46758 19690 46810
rect 19690 46758 19702 46810
rect 19702 46758 19716 46810
rect 19740 46758 19754 46810
rect 19754 46758 19766 46810
rect 19766 46758 19796 46810
rect 19820 46758 19830 46810
rect 19830 46758 19876 46810
rect 19580 46756 19636 46758
rect 19660 46756 19716 46758
rect 19740 46756 19796 46758
rect 19820 46756 19876 46758
rect 50300 46810 50356 46812
rect 50380 46810 50436 46812
rect 50460 46810 50516 46812
rect 50540 46810 50596 46812
rect 50300 46758 50346 46810
rect 50346 46758 50356 46810
rect 50380 46758 50410 46810
rect 50410 46758 50422 46810
rect 50422 46758 50436 46810
rect 50460 46758 50474 46810
rect 50474 46758 50486 46810
rect 50486 46758 50516 46810
rect 50540 46758 50550 46810
rect 50550 46758 50596 46810
rect 50300 46756 50356 46758
rect 50380 46756 50436 46758
rect 50460 46756 50516 46758
rect 50540 46756 50596 46758
rect 4220 46266 4276 46268
rect 4300 46266 4356 46268
rect 4380 46266 4436 46268
rect 4460 46266 4516 46268
rect 4220 46214 4266 46266
rect 4266 46214 4276 46266
rect 4300 46214 4330 46266
rect 4330 46214 4342 46266
rect 4342 46214 4356 46266
rect 4380 46214 4394 46266
rect 4394 46214 4406 46266
rect 4406 46214 4436 46266
rect 4460 46214 4470 46266
rect 4470 46214 4516 46266
rect 4220 46212 4276 46214
rect 4300 46212 4356 46214
rect 4380 46212 4436 46214
rect 4460 46212 4516 46214
rect 34940 46266 34996 46268
rect 35020 46266 35076 46268
rect 35100 46266 35156 46268
rect 35180 46266 35236 46268
rect 34940 46214 34986 46266
rect 34986 46214 34996 46266
rect 35020 46214 35050 46266
rect 35050 46214 35062 46266
rect 35062 46214 35076 46266
rect 35100 46214 35114 46266
rect 35114 46214 35126 46266
rect 35126 46214 35156 46266
rect 35180 46214 35190 46266
rect 35190 46214 35236 46266
rect 34940 46212 34996 46214
rect 35020 46212 35076 46214
rect 35100 46212 35156 46214
rect 35180 46212 35236 46214
rect 65660 46266 65716 46268
rect 65740 46266 65796 46268
rect 65820 46266 65876 46268
rect 65900 46266 65956 46268
rect 65660 46214 65706 46266
rect 65706 46214 65716 46266
rect 65740 46214 65770 46266
rect 65770 46214 65782 46266
rect 65782 46214 65796 46266
rect 65820 46214 65834 46266
rect 65834 46214 65846 46266
rect 65846 46214 65876 46266
rect 65900 46214 65910 46266
rect 65910 46214 65956 46266
rect 65660 46212 65716 46214
rect 65740 46212 65796 46214
rect 65820 46212 65876 46214
rect 65900 46212 65956 46214
rect 19580 45722 19636 45724
rect 19660 45722 19716 45724
rect 19740 45722 19796 45724
rect 19820 45722 19876 45724
rect 19580 45670 19626 45722
rect 19626 45670 19636 45722
rect 19660 45670 19690 45722
rect 19690 45670 19702 45722
rect 19702 45670 19716 45722
rect 19740 45670 19754 45722
rect 19754 45670 19766 45722
rect 19766 45670 19796 45722
rect 19820 45670 19830 45722
rect 19830 45670 19876 45722
rect 19580 45668 19636 45670
rect 19660 45668 19716 45670
rect 19740 45668 19796 45670
rect 19820 45668 19876 45670
rect 50300 45722 50356 45724
rect 50380 45722 50436 45724
rect 50460 45722 50516 45724
rect 50540 45722 50596 45724
rect 50300 45670 50346 45722
rect 50346 45670 50356 45722
rect 50380 45670 50410 45722
rect 50410 45670 50422 45722
rect 50422 45670 50436 45722
rect 50460 45670 50474 45722
rect 50474 45670 50486 45722
rect 50486 45670 50516 45722
rect 50540 45670 50550 45722
rect 50550 45670 50596 45722
rect 50300 45668 50356 45670
rect 50380 45668 50436 45670
rect 50460 45668 50516 45670
rect 50540 45668 50596 45670
rect 4220 45178 4276 45180
rect 4300 45178 4356 45180
rect 4380 45178 4436 45180
rect 4460 45178 4516 45180
rect 4220 45126 4266 45178
rect 4266 45126 4276 45178
rect 4300 45126 4330 45178
rect 4330 45126 4342 45178
rect 4342 45126 4356 45178
rect 4380 45126 4394 45178
rect 4394 45126 4406 45178
rect 4406 45126 4436 45178
rect 4460 45126 4470 45178
rect 4470 45126 4516 45178
rect 4220 45124 4276 45126
rect 4300 45124 4356 45126
rect 4380 45124 4436 45126
rect 4460 45124 4516 45126
rect 34940 45178 34996 45180
rect 35020 45178 35076 45180
rect 35100 45178 35156 45180
rect 35180 45178 35236 45180
rect 34940 45126 34986 45178
rect 34986 45126 34996 45178
rect 35020 45126 35050 45178
rect 35050 45126 35062 45178
rect 35062 45126 35076 45178
rect 35100 45126 35114 45178
rect 35114 45126 35126 45178
rect 35126 45126 35156 45178
rect 35180 45126 35190 45178
rect 35190 45126 35236 45178
rect 34940 45124 34996 45126
rect 35020 45124 35076 45126
rect 35100 45124 35156 45126
rect 35180 45124 35236 45126
rect 65660 45178 65716 45180
rect 65740 45178 65796 45180
rect 65820 45178 65876 45180
rect 65900 45178 65956 45180
rect 65660 45126 65706 45178
rect 65706 45126 65716 45178
rect 65740 45126 65770 45178
rect 65770 45126 65782 45178
rect 65782 45126 65796 45178
rect 65820 45126 65834 45178
rect 65834 45126 65846 45178
rect 65846 45126 65876 45178
rect 65900 45126 65910 45178
rect 65910 45126 65956 45178
rect 65660 45124 65716 45126
rect 65740 45124 65796 45126
rect 65820 45124 65876 45126
rect 65900 45124 65956 45126
rect 19580 44634 19636 44636
rect 19660 44634 19716 44636
rect 19740 44634 19796 44636
rect 19820 44634 19876 44636
rect 19580 44582 19626 44634
rect 19626 44582 19636 44634
rect 19660 44582 19690 44634
rect 19690 44582 19702 44634
rect 19702 44582 19716 44634
rect 19740 44582 19754 44634
rect 19754 44582 19766 44634
rect 19766 44582 19796 44634
rect 19820 44582 19830 44634
rect 19830 44582 19876 44634
rect 19580 44580 19636 44582
rect 19660 44580 19716 44582
rect 19740 44580 19796 44582
rect 19820 44580 19876 44582
rect 50300 44634 50356 44636
rect 50380 44634 50436 44636
rect 50460 44634 50516 44636
rect 50540 44634 50596 44636
rect 50300 44582 50346 44634
rect 50346 44582 50356 44634
rect 50380 44582 50410 44634
rect 50410 44582 50422 44634
rect 50422 44582 50436 44634
rect 50460 44582 50474 44634
rect 50474 44582 50486 44634
rect 50486 44582 50516 44634
rect 50540 44582 50550 44634
rect 50550 44582 50596 44634
rect 50300 44580 50356 44582
rect 50380 44580 50436 44582
rect 50460 44580 50516 44582
rect 50540 44580 50596 44582
rect 4220 44090 4276 44092
rect 4300 44090 4356 44092
rect 4380 44090 4436 44092
rect 4460 44090 4516 44092
rect 4220 44038 4266 44090
rect 4266 44038 4276 44090
rect 4300 44038 4330 44090
rect 4330 44038 4342 44090
rect 4342 44038 4356 44090
rect 4380 44038 4394 44090
rect 4394 44038 4406 44090
rect 4406 44038 4436 44090
rect 4460 44038 4470 44090
rect 4470 44038 4516 44090
rect 4220 44036 4276 44038
rect 4300 44036 4356 44038
rect 4380 44036 4436 44038
rect 4460 44036 4516 44038
rect 34940 44090 34996 44092
rect 35020 44090 35076 44092
rect 35100 44090 35156 44092
rect 35180 44090 35236 44092
rect 34940 44038 34986 44090
rect 34986 44038 34996 44090
rect 35020 44038 35050 44090
rect 35050 44038 35062 44090
rect 35062 44038 35076 44090
rect 35100 44038 35114 44090
rect 35114 44038 35126 44090
rect 35126 44038 35156 44090
rect 35180 44038 35190 44090
rect 35190 44038 35236 44090
rect 34940 44036 34996 44038
rect 35020 44036 35076 44038
rect 35100 44036 35156 44038
rect 35180 44036 35236 44038
rect 65660 44090 65716 44092
rect 65740 44090 65796 44092
rect 65820 44090 65876 44092
rect 65900 44090 65956 44092
rect 65660 44038 65706 44090
rect 65706 44038 65716 44090
rect 65740 44038 65770 44090
rect 65770 44038 65782 44090
rect 65782 44038 65796 44090
rect 65820 44038 65834 44090
rect 65834 44038 65846 44090
rect 65846 44038 65876 44090
rect 65900 44038 65910 44090
rect 65910 44038 65956 44090
rect 65660 44036 65716 44038
rect 65740 44036 65796 44038
rect 65820 44036 65876 44038
rect 65900 44036 65956 44038
rect 19580 43546 19636 43548
rect 19660 43546 19716 43548
rect 19740 43546 19796 43548
rect 19820 43546 19876 43548
rect 19580 43494 19626 43546
rect 19626 43494 19636 43546
rect 19660 43494 19690 43546
rect 19690 43494 19702 43546
rect 19702 43494 19716 43546
rect 19740 43494 19754 43546
rect 19754 43494 19766 43546
rect 19766 43494 19796 43546
rect 19820 43494 19830 43546
rect 19830 43494 19876 43546
rect 19580 43492 19636 43494
rect 19660 43492 19716 43494
rect 19740 43492 19796 43494
rect 19820 43492 19876 43494
rect 50300 43546 50356 43548
rect 50380 43546 50436 43548
rect 50460 43546 50516 43548
rect 50540 43546 50596 43548
rect 50300 43494 50346 43546
rect 50346 43494 50356 43546
rect 50380 43494 50410 43546
rect 50410 43494 50422 43546
rect 50422 43494 50436 43546
rect 50460 43494 50474 43546
rect 50474 43494 50486 43546
rect 50486 43494 50516 43546
rect 50540 43494 50550 43546
rect 50550 43494 50596 43546
rect 50300 43492 50356 43494
rect 50380 43492 50436 43494
rect 50460 43492 50516 43494
rect 50540 43492 50596 43494
rect 4220 43002 4276 43004
rect 4300 43002 4356 43004
rect 4380 43002 4436 43004
rect 4460 43002 4516 43004
rect 4220 42950 4266 43002
rect 4266 42950 4276 43002
rect 4300 42950 4330 43002
rect 4330 42950 4342 43002
rect 4342 42950 4356 43002
rect 4380 42950 4394 43002
rect 4394 42950 4406 43002
rect 4406 42950 4436 43002
rect 4460 42950 4470 43002
rect 4470 42950 4516 43002
rect 4220 42948 4276 42950
rect 4300 42948 4356 42950
rect 4380 42948 4436 42950
rect 4460 42948 4516 42950
rect 34940 43002 34996 43004
rect 35020 43002 35076 43004
rect 35100 43002 35156 43004
rect 35180 43002 35236 43004
rect 34940 42950 34986 43002
rect 34986 42950 34996 43002
rect 35020 42950 35050 43002
rect 35050 42950 35062 43002
rect 35062 42950 35076 43002
rect 35100 42950 35114 43002
rect 35114 42950 35126 43002
rect 35126 42950 35156 43002
rect 35180 42950 35190 43002
rect 35190 42950 35236 43002
rect 34940 42948 34996 42950
rect 35020 42948 35076 42950
rect 35100 42948 35156 42950
rect 35180 42948 35236 42950
rect 65660 43002 65716 43004
rect 65740 43002 65796 43004
rect 65820 43002 65876 43004
rect 65900 43002 65956 43004
rect 65660 42950 65706 43002
rect 65706 42950 65716 43002
rect 65740 42950 65770 43002
rect 65770 42950 65782 43002
rect 65782 42950 65796 43002
rect 65820 42950 65834 43002
rect 65834 42950 65846 43002
rect 65846 42950 65876 43002
rect 65900 42950 65910 43002
rect 65910 42950 65956 43002
rect 65660 42948 65716 42950
rect 65740 42948 65796 42950
rect 65820 42948 65876 42950
rect 65900 42948 65956 42950
rect 19580 42458 19636 42460
rect 19660 42458 19716 42460
rect 19740 42458 19796 42460
rect 19820 42458 19876 42460
rect 19580 42406 19626 42458
rect 19626 42406 19636 42458
rect 19660 42406 19690 42458
rect 19690 42406 19702 42458
rect 19702 42406 19716 42458
rect 19740 42406 19754 42458
rect 19754 42406 19766 42458
rect 19766 42406 19796 42458
rect 19820 42406 19830 42458
rect 19830 42406 19876 42458
rect 19580 42404 19636 42406
rect 19660 42404 19716 42406
rect 19740 42404 19796 42406
rect 19820 42404 19876 42406
rect 50300 42458 50356 42460
rect 50380 42458 50436 42460
rect 50460 42458 50516 42460
rect 50540 42458 50596 42460
rect 50300 42406 50346 42458
rect 50346 42406 50356 42458
rect 50380 42406 50410 42458
rect 50410 42406 50422 42458
rect 50422 42406 50436 42458
rect 50460 42406 50474 42458
rect 50474 42406 50486 42458
rect 50486 42406 50516 42458
rect 50540 42406 50550 42458
rect 50550 42406 50596 42458
rect 50300 42404 50356 42406
rect 50380 42404 50436 42406
rect 50460 42404 50516 42406
rect 50540 42404 50596 42406
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 34940 41914 34996 41916
rect 35020 41914 35076 41916
rect 35100 41914 35156 41916
rect 35180 41914 35236 41916
rect 34940 41862 34986 41914
rect 34986 41862 34996 41914
rect 35020 41862 35050 41914
rect 35050 41862 35062 41914
rect 35062 41862 35076 41914
rect 35100 41862 35114 41914
rect 35114 41862 35126 41914
rect 35126 41862 35156 41914
rect 35180 41862 35190 41914
rect 35190 41862 35236 41914
rect 34940 41860 34996 41862
rect 35020 41860 35076 41862
rect 35100 41860 35156 41862
rect 35180 41860 35236 41862
rect 65660 41914 65716 41916
rect 65740 41914 65796 41916
rect 65820 41914 65876 41916
rect 65900 41914 65956 41916
rect 65660 41862 65706 41914
rect 65706 41862 65716 41914
rect 65740 41862 65770 41914
rect 65770 41862 65782 41914
rect 65782 41862 65796 41914
rect 65820 41862 65834 41914
rect 65834 41862 65846 41914
rect 65846 41862 65876 41914
rect 65900 41862 65910 41914
rect 65910 41862 65956 41914
rect 65660 41860 65716 41862
rect 65740 41860 65796 41862
rect 65820 41860 65876 41862
rect 65900 41860 65956 41862
rect 19580 41370 19636 41372
rect 19660 41370 19716 41372
rect 19740 41370 19796 41372
rect 19820 41370 19876 41372
rect 19580 41318 19626 41370
rect 19626 41318 19636 41370
rect 19660 41318 19690 41370
rect 19690 41318 19702 41370
rect 19702 41318 19716 41370
rect 19740 41318 19754 41370
rect 19754 41318 19766 41370
rect 19766 41318 19796 41370
rect 19820 41318 19830 41370
rect 19830 41318 19876 41370
rect 19580 41316 19636 41318
rect 19660 41316 19716 41318
rect 19740 41316 19796 41318
rect 19820 41316 19876 41318
rect 50300 41370 50356 41372
rect 50380 41370 50436 41372
rect 50460 41370 50516 41372
rect 50540 41370 50596 41372
rect 50300 41318 50346 41370
rect 50346 41318 50356 41370
rect 50380 41318 50410 41370
rect 50410 41318 50422 41370
rect 50422 41318 50436 41370
rect 50460 41318 50474 41370
rect 50474 41318 50486 41370
rect 50486 41318 50516 41370
rect 50540 41318 50550 41370
rect 50550 41318 50596 41370
rect 50300 41316 50356 41318
rect 50380 41316 50436 41318
rect 50460 41316 50516 41318
rect 50540 41316 50596 41318
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 34940 40826 34996 40828
rect 35020 40826 35076 40828
rect 35100 40826 35156 40828
rect 35180 40826 35236 40828
rect 34940 40774 34986 40826
rect 34986 40774 34996 40826
rect 35020 40774 35050 40826
rect 35050 40774 35062 40826
rect 35062 40774 35076 40826
rect 35100 40774 35114 40826
rect 35114 40774 35126 40826
rect 35126 40774 35156 40826
rect 35180 40774 35190 40826
rect 35190 40774 35236 40826
rect 34940 40772 34996 40774
rect 35020 40772 35076 40774
rect 35100 40772 35156 40774
rect 35180 40772 35236 40774
rect 65660 40826 65716 40828
rect 65740 40826 65796 40828
rect 65820 40826 65876 40828
rect 65900 40826 65956 40828
rect 65660 40774 65706 40826
rect 65706 40774 65716 40826
rect 65740 40774 65770 40826
rect 65770 40774 65782 40826
rect 65782 40774 65796 40826
rect 65820 40774 65834 40826
rect 65834 40774 65846 40826
rect 65846 40774 65876 40826
rect 65900 40774 65910 40826
rect 65910 40774 65956 40826
rect 65660 40772 65716 40774
rect 65740 40772 65796 40774
rect 65820 40772 65876 40774
rect 65900 40772 65956 40774
rect 19580 40282 19636 40284
rect 19660 40282 19716 40284
rect 19740 40282 19796 40284
rect 19820 40282 19876 40284
rect 19580 40230 19626 40282
rect 19626 40230 19636 40282
rect 19660 40230 19690 40282
rect 19690 40230 19702 40282
rect 19702 40230 19716 40282
rect 19740 40230 19754 40282
rect 19754 40230 19766 40282
rect 19766 40230 19796 40282
rect 19820 40230 19830 40282
rect 19830 40230 19876 40282
rect 19580 40228 19636 40230
rect 19660 40228 19716 40230
rect 19740 40228 19796 40230
rect 19820 40228 19876 40230
rect 50300 40282 50356 40284
rect 50380 40282 50436 40284
rect 50460 40282 50516 40284
rect 50540 40282 50596 40284
rect 50300 40230 50346 40282
rect 50346 40230 50356 40282
rect 50380 40230 50410 40282
rect 50410 40230 50422 40282
rect 50422 40230 50436 40282
rect 50460 40230 50474 40282
rect 50474 40230 50486 40282
rect 50486 40230 50516 40282
rect 50540 40230 50550 40282
rect 50550 40230 50596 40282
rect 50300 40228 50356 40230
rect 50380 40228 50436 40230
rect 50460 40228 50516 40230
rect 50540 40228 50596 40230
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 65660 39738 65716 39740
rect 65740 39738 65796 39740
rect 65820 39738 65876 39740
rect 65900 39738 65956 39740
rect 65660 39686 65706 39738
rect 65706 39686 65716 39738
rect 65740 39686 65770 39738
rect 65770 39686 65782 39738
rect 65782 39686 65796 39738
rect 65820 39686 65834 39738
rect 65834 39686 65846 39738
rect 65846 39686 65876 39738
rect 65900 39686 65910 39738
rect 65910 39686 65956 39738
rect 65660 39684 65716 39686
rect 65740 39684 65796 39686
rect 65820 39684 65876 39686
rect 65900 39684 65956 39686
rect 19580 39194 19636 39196
rect 19660 39194 19716 39196
rect 19740 39194 19796 39196
rect 19820 39194 19876 39196
rect 19580 39142 19626 39194
rect 19626 39142 19636 39194
rect 19660 39142 19690 39194
rect 19690 39142 19702 39194
rect 19702 39142 19716 39194
rect 19740 39142 19754 39194
rect 19754 39142 19766 39194
rect 19766 39142 19796 39194
rect 19820 39142 19830 39194
rect 19830 39142 19876 39194
rect 19580 39140 19636 39142
rect 19660 39140 19716 39142
rect 19740 39140 19796 39142
rect 19820 39140 19876 39142
rect 50300 39194 50356 39196
rect 50380 39194 50436 39196
rect 50460 39194 50516 39196
rect 50540 39194 50596 39196
rect 50300 39142 50346 39194
rect 50346 39142 50356 39194
rect 50380 39142 50410 39194
rect 50410 39142 50422 39194
rect 50422 39142 50436 39194
rect 50460 39142 50474 39194
rect 50474 39142 50486 39194
rect 50486 39142 50516 39194
rect 50540 39142 50550 39194
rect 50550 39142 50596 39194
rect 50300 39140 50356 39142
rect 50380 39140 50436 39142
rect 50460 39140 50516 39142
rect 50540 39140 50596 39142
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 65660 38650 65716 38652
rect 65740 38650 65796 38652
rect 65820 38650 65876 38652
rect 65900 38650 65956 38652
rect 65660 38598 65706 38650
rect 65706 38598 65716 38650
rect 65740 38598 65770 38650
rect 65770 38598 65782 38650
rect 65782 38598 65796 38650
rect 65820 38598 65834 38650
rect 65834 38598 65846 38650
rect 65846 38598 65876 38650
rect 65900 38598 65910 38650
rect 65910 38598 65956 38650
rect 65660 38596 65716 38598
rect 65740 38596 65796 38598
rect 65820 38596 65876 38598
rect 65900 38596 65956 38598
rect 19580 38106 19636 38108
rect 19660 38106 19716 38108
rect 19740 38106 19796 38108
rect 19820 38106 19876 38108
rect 19580 38054 19626 38106
rect 19626 38054 19636 38106
rect 19660 38054 19690 38106
rect 19690 38054 19702 38106
rect 19702 38054 19716 38106
rect 19740 38054 19754 38106
rect 19754 38054 19766 38106
rect 19766 38054 19796 38106
rect 19820 38054 19830 38106
rect 19830 38054 19876 38106
rect 19580 38052 19636 38054
rect 19660 38052 19716 38054
rect 19740 38052 19796 38054
rect 19820 38052 19876 38054
rect 50300 38106 50356 38108
rect 50380 38106 50436 38108
rect 50460 38106 50516 38108
rect 50540 38106 50596 38108
rect 50300 38054 50346 38106
rect 50346 38054 50356 38106
rect 50380 38054 50410 38106
rect 50410 38054 50422 38106
rect 50422 38054 50436 38106
rect 50460 38054 50474 38106
rect 50474 38054 50486 38106
rect 50486 38054 50516 38106
rect 50540 38054 50550 38106
rect 50550 38054 50596 38106
rect 50300 38052 50356 38054
rect 50380 38052 50436 38054
rect 50460 38052 50516 38054
rect 50540 38052 50596 38054
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 65660 37562 65716 37564
rect 65740 37562 65796 37564
rect 65820 37562 65876 37564
rect 65900 37562 65956 37564
rect 65660 37510 65706 37562
rect 65706 37510 65716 37562
rect 65740 37510 65770 37562
rect 65770 37510 65782 37562
rect 65782 37510 65796 37562
rect 65820 37510 65834 37562
rect 65834 37510 65846 37562
rect 65846 37510 65876 37562
rect 65900 37510 65910 37562
rect 65910 37510 65956 37562
rect 65660 37508 65716 37510
rect 65740 37508 65796 37510
rect 65820 37508 65876 37510
rect 65900 37508 65956 37510
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 50300 37018 50356 37020
rect 50380 37018 50436 37020
rect 50460 37018 50516 37020
rect 50540 37018 50596 37020
rect 50300 36966 50346 37018
rect 50346 36966 50356 37018
rect 50380 36966 50410 37018
rect 50410 36966 50422 37018
rect 50422 36966 50436 37018
rect 50460 36966 50474 37018
rect 50474 36966 50486 37018
rect 50486 36966 50516 37018
rect 50540 36966 50550 37018
rect 50550 36966 50596 37018
rect 50300 36964 50356 36966
rect 50380 36964 50436 36966
rect 50460 36964 50516 36966
rect 50540 36964 50596 36966
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 65660 36474 65716 36476
rect 65740 36474 65796 36476
rect 65820 36474 65876 36476
rect 65900 36474 65956 36476
rect 65660 36422 65706 36474
rect 65706 36422 65716 36474
rect 65740 36422 65770 36474
rect 65770 36422 65782 36474
rect 65782 36422 65796 36474
rect 65820 36422 65834 36474
rect 65834 36422 65846 36474
rect 65846 36422 65876 36474
rect 65900 36422 65910 36474
rect 65910 36422 65956 36474
rect 65660 36420 65716 36422
rect 65740 36420 65796 36422
rect 65820 36420 65876 36422
rect 65900 36420 65956 36422
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 50300 35930 50356 35932
rect 50380 35930 50436 35932
rect 50460 35930 50516 35932
rect 50540 35930 50596 35932
rect 50300 35878 50346 35930
rect 50346 35878 50356 35930
rect 50380 35878 50410 35930
rect 50410 35878 50422 35930
rect 50422 35878 50436 35930
rect 50460 35878 50474 35930
rect 50474 35878 50486 35930
rect 50486 35878 50516 35930
rect 50540 35878 50550 35930
rect 50550 35878 50596 35930
rect 50300 35876 50356 35878
rect 50380 35876 50436 35878
rect 50460 35876 50516 35878
rect 50540 35876 50596 35878
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 65660 35386 65716 35388
rect 65740 35386 65796 35388
rect 65820 35386 65876 35388
rect 65900 35386 65956 35388
rect 65660 35334 65706 35386
rect 65706 35334 65716 35386
rect 65740 35334 65770 35386
rect 65770 35334 65782 35386
rect 65782 35334 65796 35386
rect 65820 35334 65834 35386
rect 65834 35334 65846 35386
rect 65846 35334 65876 35386
rect 65900 35334 65910 35386
rect 65910 35334 65956 35386
rect 65660 35332 65716 35334
rect 65740 35332 65796 35334
rect 65820 35332 65876 35334
rect 65900 35332 65956 35334
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 50300 34842 50356 34844
rect 50380 34842 50436 34844
rect 50460 34842 50516 34844
rect 50540 34842 50596 34844
rect 50300 34790 50346 34842
rect 50346 34790 50356 34842
rect 50380 34790 50410 34842
rect 50410 34790 50422 34842
rect 50422 34790 50436 34842
rect 50460 34790 50474 34842
rect 50474 34790 50486 34842
rect 50486 34790 50516 34842
rect 50540 34790 50550 34842
rect 50550 34790 50596 34842
rect 50300 34788 50356 34790
rect 50380 34788 50436 34790
rect 50460 34788 50516 34790
rect 50540 34788 50596 34790
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 65660 34298 65716 34300
rect 65740 34298 65796 34300
rect 65820 34298 65876 34300
rect 65900 34298 65956 34300
rect 65660 34246 65706 34298
rect 65706 34246 65716 34298
rect 65740 34246 65770 34298
rect 65770 34246 65782 34298
rect 65782 34246 65796 34298
rect 65820 34246 65834 34298
rect 65834 34246 65846 34298
rect 65846 34246 65876 34298
rect 65900 34246 65910 34298
rect 65910 34246 65956 34298
rect 65660 34244 65716 34246
rect 65740 34244 65796 34246
rect 65820 34244 65876 34246
rect 65900 34244 65956 34246
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 50300 33754 50356 33756
rect 50380 33754 50436 33756
rect 50460 33754 50516 33756
rect 50540 33754 50596 33756
rect 50300 33702 50346 33754
rect 50346 33702 50356 33754
rect 50380 33702 50410 33754
rect 50410 33702 50422 33754
rect 50422 33702 50436 33754
rect 50460 33702 50474 33754
rect 50474 33702 50486 33754
rect 50486 33702 50516 33754
rect 50540 33702 50550 33754
rect 50550 33702 50596 33754
rect 50300 33700 50356 33702
rect 50380 33700 50436 33702
rect 50460 33700 50516 33702
rect 50540 33700 50596 33702
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 65660 33210 65716 33212
rect 65740 33210 65796 33212
rect 65820 33210 65876 33212
rect 65900 33210 65956 33212
rect 65660 33158 65706 33210
rect 65706 33158 65716 33210
rect 65740 33158 65770 33210
rect 65770 33158 65782 33210
rect 65782 33158 65796 33210
rect 65820 33158 65834 33210
rect 65834 33158 65846 33210
rect 65846 33158 65876 33210
rect 65900 33158 65910 33210
rect 65910 33158 65956 33210
rect 65660 33156 65716 33158
rect 65740 33156 65796 33158
rect 65820 33156 65876 33158
rect 65900 33156 65956 33158
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 50300 32666 50356 32668
rect 50380 32666 50436 32668
rect 50460 32666 50516 32668
rect 50540 32666 50596 32668
rect 50300 32614 50346 32666
rect 50346 32614 50356 32666
rect 50380 32614 50410 32666
rect 50410 32614 50422 32666
rect 50422 32614 50436 32666
rect 50460 32614 50474 32666
rect 50474 32614 50486 32666
rect 50486 32614 50516 32666
rect 50540 32614 50550 32666
rect 50550 32614 50596 32666
rect 50300 32612 50356 32614
rect 50380 32612 50436 32614
rect 50460 32612 50516 32614
rect 50540 32612 50596 32614
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 65660 32122 65716 32124
rect 65740 32122 65796 32124
rect 65820 32122 65876 32124
rect 65900 32122 65956 32124
rect 65660 32070 65706 32122
rect 65706 32070 65716 32122
rect 65740 32070 65770 32122
rect 65770 32070 65782 32122
rect 65782 32070 65796 32122
rect 65820 32070 65834 32122
rect 65834 32070 65846 32122
rect 65846 32070 65876 32122
rect 65900 32070 65910 32122
rect 65910 32070 65956 32122
rect 65660 32068 65716 32070
rect 65740 32068 65796 32070
rect 65820 32068 65876 32070
rect 65900 32068 65956 32070
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 50300 31578 50356 31580
rect 50380 31578 50436 31580
rect 50460 31578 50516 31580
rect 50540 31578 50596 31580
rect 50300 31526 50346 31578
rect 50346 31526 50356 31578
rect 50380 31526 50410 31578
rect 50410 31526 50422 31578
rect 50422 31526 50436 31578
rect 50460 31526 50474 31578
rect 50474 31526 50486 31578
rect 50486 31526 50516 31578
rect 50540 31526 50550 31578
rect 50550 31526 50596 31578
rect 50300 31524 50356 31526
rect 50380 31524 50436 31526
rect 50460 31524 50516 31526
rect 50540 31524 50596 31526
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 65660 31034 65716 31036
rect 65740 31034 65796 31036
rect 65820 31034 65876 31036
rect 65900 31034 65956 31036
rect 65660 30982 65706 31034
rect 65706 30982 65716 31034
rect 65740 30982 65770 31034
rect 65770 30982 65782 31034
rect 65782 30982 65796 31034
rect 65820 30982 65834 31034
rect 65834 30982 65846 31034
rect 65846 30982 65876 31034
rect 65900 30982 65910 31034
rect 65910 30982 65956 31034
rect 65660 30980 65716 30982
rect 65740 30980 65796 30982
rect 65820 30980 65876 30982
rect 65900 30980 65956 30982
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 50300 30490 50356 30492
rect 50380 30490 50436 30492
rect 50460 30490 50516 30492
rect 50540 30490 50596 30492
rect 50300 30438 50346 30490
rect 50346 30438 50356 30490
rect 50380 30438 50410 30490
rect 50410 30438 50422 30490
rect 50422 30438 50436 30490
rect 50460 30438 50474 30490
rect 50474 30438 50486 30490
rect 50486 30438 50516 30490
rect 50540 30438 50550 30490
rect 50550 30438 50596 30490
rect 50300 30436 50356 30438
rect 50380 30436 50436 30438
rect 50460 30436 50516 30438
rect 50540 30436 50596 30438
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 65660 29946 65716 29948
rect 65740 29946 65796 29948
rect 65820 29946 65876 29948
rect 65900 29946 65956 29948
rect 65660 29894 65706 29946
rect 65706 29894 65716 29946
rect 65740 29894 65770 29946
rect 65770 29894 65782 29946
rect 65782 29894 65796 29946
rect 65820 29894 65834 29946
rect 65834 29894 65846 29946
rect 65846 29894 65876 29946
rect 65900 29894 65910 29946
rect 65910 29894 65956 29946
rect 65660 29892 65716 29894
rect 65740 29892 65796 29894
rect 65820 29892 65876 29894
rect 65900 29892 65956 29894
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 50300 29402 50356 29404
rect 50380 29402 50436 29404
rect 50460 29402 50516 29404
rect 50540 29402 50596 29404
rect 50300 29350 50346 29402
rect 50346 29350 50356 29402
rect 50380 29350 50410 29402
rect 50410 29350 50422 29402
rect 50422 29350 50436 29402
rect 50460 29350 50474 29402
rect 50474 29350 50486 29402
rect 50486 29350 50516 29402
rect 50540 29350 50550 29402
rect 50550 29350 50596 29402
rect 50300 29348 50356 29350
rect 50380 29348 50436 29350
rect 50460 29348 50516 29350
rect 50540 29348 50596 29350
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 65660 28858 65716 28860
rect 65740 28858 65796 28860
rect 65820 28858 65876 28860
rect 65900 28858 65956 28860
rect 65660 28806 65706 28858
rect 65706 28806 65716 28858
rect 65740 28806 65770 28858
rect 65770 28806 65782 28858
rect 65782 28806 65796 28858
rect 65820 28806 65834 28858
rect 65834 28806 65846 28858
rect 65846 28806 65876 28858
rect 65900 28806 65910 28858
rect 65910 28806 65956 28858
rect 65660 28804 65716 28806
rect 65740 28804 65796 28806
rect 65820 28804 65876 28806
rect 65900 28804 65956 28806
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 50300 28314 50356 28316
rect 50380 28314 50436 28316
rect 50460 28314 50516 28316
rect 50540 28314 50596 28316
rect 50300 28262 50346 28314
rect 50346 28262 50356 28314
rect 50380 28262 50410 28314
rect 50410 28262 50422 28314
rect 50422 28262 50436 28314
rect 50460 28262 50474 28314
rect 50474 28262 50486 28314
rect 50486 28262 50516 28314
rect 50540 28262 50550 28314
rect 50550 28262 50596 28314
rect 50300 28260 50356 28262
rect 50380 28260 50436 28262
rect 50460 28260 50516 28262
rect 50540 28260 50596 28262
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 65660 27770 65716 27772
rect 65740 27770 65796 27772
rect 65820 27770 65876 27772
rect 65900 27770 65956 27772
rect 65660 27718 65706 27770
rect 65706 27718 65716 27770
rect 65740 27718 65770 27770
rect 65770 27718 65782 27770
rect 65782 27718 65796 27770
rect 65820 27718 65834 27770
rect 65834 27718 65846 27770
rect 65846 27718 65876 27770
rect 65900 27718 65910 27770
rect 65910 27718 65956 27770
rect 65660 27716 65716 27718
rect 65740 27716 65796 27718
rect 65820 27716 65876 27718
rect 65900 27716 65956 27718
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 50300 27226 50356 27228
rect 50380 27226 50436 27228
rect 50460 27226 50516 27228
rect 50540 27226 50596 27228
rect 50300 27174 50346 27226
rect 50346 27174 50356 27226
rect 50380 27174 50410 27226
rect 50410 27174 50422 27226
rect 50422 27174 50436 27226
rect 50460 27174 50474 27226
rect 50474 27174 50486 27226
rect 50486 27174 50516 27226
rect 50540 27174 50550 27226
rect 50550 27174 50596 27226
rect 50300 27172 50356 27174
rect 50380 27172 50436 27174
rect 50460 27172 50516 27174
rect 50540 27172 50596 27174
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 65660 26682 65716 26684
rect 65740 26682 65796 26684
rect 65820 26682 65876 26684
rect 65900 26682 65956 26684
rect 65660 26630 65706 26682
rect 65706 26630 65716 26682
rect 65740 26630 65770 26682
rect 65770 26630 65782 26682
rect 65782 26630 65796 26682
rect 65820 26630 65834 26682
rect 65834 26630 65846 26682
rect 65846 26630 65876 26682
rect 65900 26630 65910 26682
rect 65910 26630 65956 26682
rect 65660 26628 65716 26630
rect 65740 26628 65796 26630
rect 65820 26628 65876 26630
rect 65900 26628 65956 26630
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 50300 26138 50356 26140
rect 50380 26138 50436 26140
rect 50460 26138 50516 26140
rect 50540 26138 50596 26140
rect 50300 26086 50346 26138
rect 50346 26086 50356 26138
rect 50380 26086 50410 26138
rect 50410 26086 50422 26138
rect 50422 26086 50436 26138
rect 50460 26086 50474 26138
rect 50474 26086 50486 26138
rect 50486 26086 50516 26138
rect 50540 26086 50550 26138
rect 50550 26086 50596 26138
rect 50300 26084 50356 26086
rect 50380 26084 50436 26086
rect 50460 26084 50516 26086
rect 50540 26084 50596 26086
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 65660 25594 65716 25596
rect 65740 25594 65796 25596
rect 65820 25594 65876 25596
rect 65900 25594 65956 25596
rect 65660 25542 65706 25594
rect 65706 25542 65716 25594
rect 65740 25542 65770 25594
rect 65770 25542 65782 25594
rect 65782 25542 65796 25594
rect 65820 25542 65834 25594
rect 65834 25542 65846 25594
rect 65846 25542 65876 25594
rect 65900 25542 65910 25594
rect 65910 25542 65956 25594
rect 65660 25540 65716 25542
rect 65740 25540 65796 25542
rect 65820 25540 65876 25542
rect 65900 25540 65956 25542
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 50300 25050 50356 25052
rect 50380 25050 50436 25052
rect 50460 25050 50516 25052
rect 50540 25050 50596 25052
rect 50300 24998 50346 25050
rect 50346 24998 50356 25050
rect 50380 24998 50410 25050
rect 50410 24998 50422 25050
rect 50422 24998 50436 25050
rect 50460 24998 50474 25050
rect 50474 24998 50486 25050
rect 50486 24998 50516 25050
rect 50540 24998 50550 25050
rect 50550 24998 50596 25050
rect 50300 24996 50356 24998
rect 50380 24996 50436 24998
rect 50460 24996 50516 24998
rect 50540 24996 50596 24998
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 65660 24506 65716 24508
rect 65740 24506 65796 24508
rect 65820 24506 65876 24508
rect 65900 24506 65956 24508
rect 65660 24454 65706 24506
rect 65706 24454 65716 24506
rect 65740 24454 65770 24506
rect 65770 24454 65782 24506
rect 65782 24454 65796 24506
rect 65820 24454 65834 24506
rect 65834 24454 65846 24506
rect 65846 24454 65876 24506
rect 65900 24454 65910 24506
rect 65910 24454 65956 24506
rect 65660 24452 65716 24454
rect 65740 24452 65796 24454
rect 65820 24452 65876 24454
rect 65900 24452 65956 24454
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 50300 23962 50356 23964
rect 50380 23962 50436 23964
rect 50460 23962 50516 23964
rect 50540 23962 50596 23964
rect 50300 23910 50346 23962
rect 50346 23910 50356 23962
rect 50380 23910 50410 23962
rect 50410 23910 50422 23962
rect 50422 23910 50436 23962
rect 50460 23910 50474 23962
rect 50474 23910 50486 23962
rect 50486 23910 50516 23962
rect 50540 23910 50550 23962
rect 50550 23910 50596 23962
rect 50300 23908 50356 23910
rect 50380 23908 50436 23910
rect 50460 23908 50516 23910
rect 50540 23908 50596 23910
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 65660 23418 65716 23420
rect 65740 23418 65796 23420
rect 65820 23418 65876 23420
rect 65900 23418 65956 23420
rect 65660 23366 65706 23418
rect 65706 23366 65716 23418
rect 65740 23366 65770 23418
rect 65770 23366 65782 23418
rect 65782 23366 65796 23418
rect 65820 23366 65834 23418
rect 65834 23366 65846 23418
rect 65846 23366 65876 23418
rect 65900 23366 65910 23418
rect 65910 23366 65956 23418
rect 65660 23364 65716 23366
rect 65740 23364 65796 23366
rect 65820 23364 65876 23366
rect 65900 23364 65956 23366
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 50300 22874 50356 22876
rect 50380 22874 50436 22876
rect 50460 22874 50516 22876
rect 50540 22874 50596 22876
rect 50300 22822 50346 22874
rect 50346 22822 50356 22874
rect 50380 22822 50410 22874
rect 50410 22822 50422 22874
rect 50422 22822 50436 22874
rect 50460 22822 50474 22874
rect 50474 22822 50486 22874
rect 50486 22822 50516 22874
rect 50540 22822 50550 22874
rect 50550 22822 50596 22874
rect 50300 22820 50356 22822
rect 50380 22820 50436 22822
rect 50460 22820 50516 22822
rect 50540 22820 50596 22822
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 65660 22330 65716 22332
rect 65740 22330 65796 22332
rect 65820 22330 65876 22332
rect 65900 22330 65956 22332
rect 65660 22278 65706 22330
rect 65706 22278 65716 22330
rect 65740 22278 65770 22330
rect 65770 22278 65782 22330
rect 65782 22278 65796 22330
rect 65820 22278 65834 22330
rect 65834 22278 65846 22330
rect 65846 22278 65876 22330
rect 65900 22278 65910 22330
rect 65910 22278 65956 22330
rect 65660 22276 65716 22278
rect 65740 22276 65796 22278
rect 65820 22276 65876 22278
rect 65900 22276 65956 22278
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 50300 21786 50356 21788
rect 50380 21786 50436 21788
rect 50460 21786 50516 21788
rect 50540 21786 50596 21788
rect 50300 21734 50346 21786
rect 50346 21734 50356 21786
rect 50380 21734 50410 21786
rect 50410 21734 50422 21786
rect 50422 21734 50436 21786
rect 50460 21734 50474 21786
rect 50474 21734 50486 21786
rect 50486 21734 50516 21786
rect 50540 21734 50550 21786
rect 50550 21734 50596 21786
rect 50300 21732 50356 21734
rect 50380 21732 50436 21734
rect 50460 21732 50516 21734
rect 50540 21732 50596 21734
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 65660 21242 65716 21244
rect 65740 21242 65796 21244
rect 65820 21242 65876 21244
rect 65900 21242 65956 21244
rect 65660 21190 65706 21242
rect 65706 21190 65716 21242
rect 65740 21190 65770 21242
rect 65770 21190 65782 21242
rect 65782 21190 65796 21242
rect 65820 21190 65834 21242
rect 65834 21190 65846 21242
rect 65846 21190 65876 21242
rect 65900 21190 65910 21242
rect 65910 21190 65956 21242
rect 65660 21188 65716 21190
rect 65740 21188 65796 21190
rect 65820 21188 65876 21190
rect 65900 21188 65956 21190
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 50300 20698 50356 20700
rect 50380 20698 50436 20700
rect 50460 20698 50516 20700
rect 50540 20698 50596 20700
rect 50300 20646 50346 20698
rect 50346 20646 50356 20698
rect 50380 20646 50410 20698
rect 50410 20646 50422 20698
rect 50422 20646 50436 20698
rect 50460 20646 50474 20698
rect 50474 20646 50486 20698
rect 50486 20646 50516 20698
rect 50540 20646 50550 20698
rect 50550 20646 50596 20698
rect 50300 20644 50356 20646
rect 50380 20644 50436 20646
rect 50460 20644 50516 20646
rect 50540 20644 50596 20646
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 65660 20154 65716 20156
rect 65740 20154 65796 20156
rect 65820 20154 65876 20156
rect 65900 20154 65956 20156
rect 65660 20102 65706 20154
rect 65706 20102 65716 20154
rect 65740 20102 65770 20154
rect 65770 20102 65782 20154
rect 65782 20102 65796 20154
rect 65820 20102 65834 20154
rect 65834 20102 65846 20154
rect 65846 20102 65876 20154
rect 65900 20102 65910 20154
rect 65910 20102 65956 20154
rect 65660 20100 65716 20102
rect 65740 20100 65796 20102
rect 65820 20100 65876 20102
rect 65900 20100 65956 20102
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 50300 19610 50356 19612
rect 50380 19610 50436 19612
rect 50460 19610 50516 19612
rect 50540 19610 50596 19612
rect 50300 19558 50346 19610
rect 50346 19558 50356 19610
rect 50380 19558 50410 19610
rect 50410 19558 50422 19610
rect 50422 19558 50436 19610
rect 50460 19558 50474 19610
rect 50474 19558 50486 19610
rect 50486 19558 50516 19610
rect 50540 19558 50550 19610
rect 50550 19558 50596 19610
rect 50300 19556 50356 19558
rect 50380 19556 50436 19558
rect 50460 19556 50516 19558
rect 50540 19556 50596 19558
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 65660 19066 65716 19068
rect 65740 19066 65796 19068
rect 65820 19066 65876 19068
rect 65900 19066 65956 19068
rect 65660 19014 65706 19066
rect 65706 19014 65716 19066
rect 65740 19014 65770 19066
rect 65770 19014 65782 19066
rect 65782 19014 65796 19066
rect 65820 19014 65834 19066
rect 65834 19014 65846 19066
rect 65846 19014 65876 19066
rect 65900 19014 65910 19066
rect 65910 19014 65956 19066
rect 65660 19012 65716 19014
rect 65740 19012 65796 19014
rect 65820 19012 65876 19014
rect 65900 19012 65956 19014
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 50300 18522 50356 18524
rect 50380 18522 50436 18524
rect 50460 18522 50516 18524
rect 50540 18522 50596 18524
rect 50300 18470 50346 18522
rect 50346 18470 50356 18522
rect 50380 18470 50410 18522
rect 50410 18470 50422 18522
rect 50422 18470 50436 18522
rect 50460 18470 50474 18522
rect 50474 18470 50486 18522
rect 50486 18470 50516 18522
rect 50540 18470 50550 18522
rect 50550 18470 50596 18522
rect 50300 18468 50356 18470
rect 50380 18468 50436 18470
rect 50460 18468 50516 18470
rect 50540 18468 50596 18470
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 65660 17978 65716 17980
rect 65740 17978 65796 17980
rect 65820 17978 65876 17980
rect 65900 17978 65956 17980
rect 65660 17926 65706 17978
rect 65706 17926 65716 17978
rect 65740 17926 65770 17978
rect 65770 17926 65782 17978
rect 65782 17926 65796 17978
rect 65820 17926 65834 17978
rect 65834 17926 65846 17978
rect 65846 17926 65876 17978
rect 65900 17926 65910 17978
rect 65910 17926 65956 17978
rect 65660 17924 65716 17926
rect 65740 17924 65796 17926
rect 65820 17924 65876 17926
rect 65900 17924 65956 17926
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 50300 17434 50356 17436
rect 50380 17434 50436 17436
rect 50460 17434 50516 17436
rect 50540 17434 50596 17436
rect 50300 17382 50346 17434
rect 50346 17382 50356 17434
rect 50380 17382 50410 17434
rect 50410 17382 50422 17434
rect 50422 17382 50436 17434
rect 50460 17382 50474 17434
rect 50474 17382 50486 17434
rect 50486 17382 50516 17434
rect 50540 17382 50550 17434
rect 50550 17382 50596 17434
rect 50300 17380 50356 17382
rect 50380 17380 50436 17382
rect 50460 17380 50516 17382
rect 50540 17380 50596 17382
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 65660 16890 65716 16892
rect 65740 16890 65796 16892
rect 65820 16890 65876 16892
rect 65900 16890 65956 16892
rect 65660 16838 65706 16890
rect 65706 16838 65716 16890
rect 65740 16838 65770 16890
rect 65770 16838 65782 16890
rect 65782 16838 65796 16890
rect 65820 16838 65834 16890
rect 65834 16838 65846 16890
rect 65846 16838 65876 16890
rect 65900 16838 65910 16890
rect 65910 16838 65956 16890
rect 65660 16836 65716 16838
rect 65740 16836 65796 16838
rect 65820 16836 65876 16838
rect 65900 16836 65956 16838
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 50300 16346 50356 16348
rect 50380 16346 50436 16348
rect 50460 16346 50516 16348
rect 50540 16346 50596 16348
rect 50300 16294 50346 16346
rect 50346 16294 50356 16346
rect 50380 16294 50410 16346
rect 50410 16294 50422 16346
rect 50422 16294 50436 16346
rect 50460 16294 50474 16346
rect 50474 16294 50486 16346
rect 50486 16294 50516 16346
rect 50540 16294 50550 16346
rect 50550 16294 50596 16346
rect 50300 16292 50356 16294
rect 50380 16292 50436 16294
rect 50460 16292 50516 16294
rect 50540 16292 50596 16294
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 65660 15802 65716 15804
rect 65740 15802 65796 15804
rect 65820 15802 65876 15804
rect 65900 15802 65956 15804
rect 65660 15750 65706 15802
rect 65706 15750 65716 15802
rect 65740 15750 65770 15802
rect 65770 15750 65782 15802
rect 65782 15750 65796 15802
rect 65820 15750 65834 15802
rect 65834 15750 65846 15802
rect 65846 15750 65876 15802
rect 65900 15750 65910 15802
rect 65910 15750 65956 15802
rect 65660 15748 65716 15750
rect 65740 15748 65796 15750
rect 65820 15748 65876 15750
rect 65900 15748 65956 15750
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 50300 15258 50356 15260
rect 50380 15258 50436 15260
rect 50460 15258 50516 15260
rect 50540 15258 50596 15260
rect 50300 15206 50346 15258
rect 50346 15206 50356 15258
rect 50380 15206 50410 15258
rect 50410 15206 50422 15258
rect 50422 15206 50436 15258
rect 50460 15206 50474 15258
rect 50474 15206 50486 15258
rect 50486 15206 50516 15258
rect 50540 15206 50550 15258
rect 50550 15206 50596 15258
rect 50300 15204 50356 15206
rect 50380 15204 50436 15206
rect 50460 15204 50516 15206
rect 50540 15204 50596 15206
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 65660 14714 65716 14716
rect 65740 14714 65796 14716
rect 65820 14714 65876 14716
rect 65900 14714 65956 14716
rect 65660 14662 65706 14714
rect 65706 14662 65716 14714
rect 65740 14662 65770 14714
rect 65770 14662 65782 14714
rect 65782 14662 65796 14714
rect 65820 14662 65834 14714
rect 65834 14662 65846 14714
rect 65846 14662 65876 14714
rect 65900 14662 65910 14714
rect 65910 14662 65956 14714
rect 65660 14660 65716 14662
rect 65740 14660 65796 14662
rect 65820 14660 65876 14662
rect 65900 14660 65956 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 3882 4120 3938 4176
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4250 3612 4252 3632
rect 4252 3612 4304 3632
rect 4304 3612 4306 3632
rect 4250 3576 4306 3612
rect 4526 3304 4582 3360
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 4986 6704 5042 6760
rect 4802 3440 4858 3496
rect 5262 6840 5318 6896
rect 5078 3712 5134 3768
rect 5722 4664 5778 4720
rect 6274 4020 6276 4040
rect 6276 4020 6328 4040
rect 6328 4020 6330 4040
rect 6274 3984 6330 4020
rect 6826 5616 6882 5672
rect 6550 4392 6606 4448
rect 8666 6060 8668 6080
rect 8668 6060 8720 6080
rect 8720 6060 8722 6080
rect 8666 6024 8722 6060
rect 7930 4256 7986 4312
rect 8114 3576 8170 3632
rect 8206 3476 8208 3496
rect 8208 3476 8260 3496
rect 8260 3476 8262 3496
rect 8206 3440 8262 3476
rect 6734 2760 6790 2816
rect 9402 7828 9404 7848
rect 9404 7828 9456 7848
rect 9456 7828 9458 7848
rect 9402 7792 9458 7828
rect 9034 5752 9090 5808
rect 9586 7112 9642 7168
rect 9494 5616 9550 5672
rect 9494 4564 9496 4584
rect 9496 4564 9548 4584
rect 9548 4564 9550 4584
rect 9494 4528 9550 4564
rect 8942 3712 8998 3768
rect 9678 3440 9734 3496
rect 11334 6840 11390 6896
rect 11242 5616 11298 5672
rect 10230 2896 10286 2952
rect 11702 13640 11758 13696
rect 12898 13640 12954 13696
rect 11610 6160 11666 6216
rect 11794 5208 11850 5264
rect 11702 3340 11704 3360
rect 11704 3340 11756 3360
rect 11756 3340 11758 3360
rect 11702 3304 11758 3340
rect 12070 6704 12126 6760
rect 12070 4820 12126 4856
rect 12070 4800 12072 4820
rect 12072 4800 12124 4820
rect 12124 4800 12126 4820
rect 12530 4392 12586 4448
rect 12438 4120 12494 4176
rect 12806 6024 12862 6080
rect 12990 4256 13046 4312
rect 12898 3304 12954 3360
rect 13634 8356 13690 8392
rect 13634 8336 13636 8356
rect 13636 8336 13688 8356
rect 13688 8336 13690 8356
rect 13634 6060 13636 6080
rect 13636 6060 13688 6080
rect 13688 6060 13690 6080
rect 13634 6024 13690 6060
rect 13266 3596 13322 3632
rect 13266 3576 13268 3596
rect 13268 3576 13320 3596
rect 13320 3576 13322 3596
rect 13634 5228 13690 5264
rect 13634 5208 13636 5228
rect 13636 5208 13688 5228
rect 13688 5208 13690 5228
rect 15014 7792 15070 7848
rect 14186 5752 14242 5808
rect 14646 7148 14648 7168
rect 14648 7148 14700 7168
rect 14700 7148 14702 7168
rect 14646 7112 14702 7148
rect 14370 4664 14426 4720
rect 13542 3168 13598 3224
rect 13726 3032 13782 3088
rect 14462 2760 14518 2816
rect 15106 4528 15162 4584
rect 15290 3576 15346 3632
rect 15474 3168 15530 3224
rect 15934 4820 15990 4856
rect 15934 4800 15936 4820
rect 15936 4800 15988 4820
rect 15988 4800 15990 4820
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 50300 14170 50356 14172
rect 50380 14170 50436 14172
rect 50460 14170 50516 14172
rect 50540 14170 50596 14172
rect 50300 14118 50346 14170
rect 50346 14118 50356 14170
rect 50380 14118 50410 14170
rect 50410 14118 50422 14170
rect 50422 14118 50436 14170
rect 50460 14118 50474 14170
rect 50474 14118 50486 14170
rect 50486 14118 50516 14170
rect 50540 14118 50550 14170
rect 50550 14118 50596 14170
rect 50300 14116 50356 14118
rect 50380 14116 50436 14118
rect 50460 14116 50516 14118
rect 50540 14116 50596 14118
rect 16670 11464 16726 11520
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 16210 3576 16266 3632
rect 16670 4664 16726 4720
rect 17038 5616 17094 5672
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 20258 8200 20314 8256
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19982 5344 20038 5400
rect 19338 5072 19394 5128
rect 19982 5072 20038 5128
rect 19062 2760 19118 2816
rect 19338 3884 19340 3904
rect 19340 3884 19392 3904
rect 19392 3884 19394 3904
rect 19338 3848 19394 3884
rect 19614 4564 19616 4584
rect 19616 4564 19668 4584
rect 19668 4564 19670 4584
rect 19614 4528 19670 4564
rect 19798 4972 19800 4992
rect 19800 4972 19852 4992
rect 19852 4972 19854 4992
rect 19798 4936 19854 4972
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 20442 6296 20498 6352
rect 20442 5752 20498 5808
rect 20442 5516 20444 5536
rect 20444 5516 20496 5536
rect 20496 5516 20498 5536
rect 20074 2760 20130 2816
rect 20442 5480 20498 5516
rect 20258 5344 20314 5400
rect 20810 6160 20866 6216
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 65660 13626 65716 13628
rect 65740 13626 65796 13628
rect 65820 13626 65876 13628
rect 65900 13626 65956 13628
rect 65660 13574 65706 13626
rect 65706 13574 65716 13626
rect 65740 13574 65770 13626
rect 65770 13574 65782 13626
rect 65782 13574 65796 13626
rect 65820 13574 65834 13626
rect 65834 13574 65846 13626
rect 65846 13574 65876 13626
rect 65900 13574 65910 13626
rect 65910 13574 65956 13626
rect 65660 13572 65716 13574
rect 65740 13572 65796 13574
rect 65820 13572 65876 13574
rect 65900 13572 65956 13574
rect 50300 13082 50356 13084
rect 50380 13082 50436 13084
rect 50460 13082 50516 13084
rect 50540 13082 50596 13084
rect 50300 13030 50346 13082
rect 50346 13030 50356 13082
rect 50380 13030 50410 13082
rect 50410 13030 50422 13082
rect 50422 13030 50436 13082
rect 50460 13030 50474 13082
rect 50474 13030 50486 13082
rect 50486 13030 50516 13082
rect 50540 13030 50550 13082
rect 50550 13030 50596 13082
rect 50300 13028 50356 13030
rect 50380 13028 50436 13030
rect 50460 13028 50516 13030
rect 50540 13028 50596 13030
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 65660 12538 65716 12540
rect 65740 12538 65796 12540
rect 65820 12538 65876 12540
rect 65900 12538 65956 12540
rect 65660 12486 65706 12538
rect 65706 12486 65716 12538
rect 65740 12486 65770 12538
rect 65770 12486 65782 12538
rect 65782 12486 65796 12538
rect 65820 12486 65834 12538
rect 65834 12486 65846 12538
rect 65846 12486 65876 12538
rect 65900 12486 65910 12538
rect 65910 12486 65956 12538
rect 65660 12484 65716 12486
rect 65740 12484 65796 12486
rect 65820 12484 65876 12486
rect 65900 12484 65956 12486
rect 21546 8492 21602 8528
rect 21546 8472 21548 8492
rect 21548 8472 21600 8492
rect 21600 8472 21602 8492
rect 21270 8372 21272 8392
rect 21272 8372 21324 8392
rect 21324 8372 21326 8392
rect 21270 8336 21326 8372
rect 21086 4528 21142 4584
rect 20718 3052 20774 3088
rect 20718 3032 20720 3052
rect 20720 3032 20772 3052
rect 20772 3032 20774 3052
rect 50300 11994 50356 11996
rect 50380 11994 50436 11996
rect 50460 11994 50516 11996
rect 50540 11994 50596 11996
rect 50300 11942 50346 11994
rect 50346 11942 50356 11994
rect 50380 11942 50410 11994
rect 50410 11942 50422 11994
rect 50422 11942 50436 11994
rect 50460 11942 50474 11994
rect 50474 11942 50486 11994
rect 50486 11942 50516 11994
rect 50540 11942 50550 11994
rect 50550 11942 50596 11994
rect 50300 11940 50356 11942
rect 50380 11940 50436 11942
rect 50460 11940 50516 11942
rect 50540 11940 50596 11942
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 65660 11450 65716 11452
rect 65740 11450 65796 11452
rect 65820 11450 65876 11452
rect 65900 11450 65956 11452
rect 65660 11398 65706 11450
rect 65706 11398 65716 11450
rect 65740 11398 65770 11450
rect 65770 11398 65782 11450
rect 65782 11398 65796 11450
rect 65820 11398 65834 11450
rect 65834 11398 65846 11450
rect 65846 11398 65876 11450
rect 65900 11398 65910 11450
rect 65910 11398 65956 11450
rect 65660 11396 65716 11398
rect 65740 11396 65796 11398
rect 65820 11396 65876 11398
rect 65900 11396 65956 11398
rect 22098 5480 22154 5536
rect 22098 3984 22154 4040
rect 22558 8200 22614 8256
rect 22926 8336 22982 8392
rect 24306 8492 24362 8528
rect 24306 8472 24308 8492
rect 24308 8472 24360 8492
rect 24360 8472 24362 8492
rect 23202 5208 23258 5264
rect 50300 10906 50356 10908
rect 50380 10906 50436 10908
rect 50460 10906 50516 10908
rect 50540 10906 50596 10908
rect 50300 10854 50346 10906
rect 50346 10854 50356 10906
rect 50380 10854 50410 10906
rect 50410 10854 50422 10906
rect 50422 10854 50436 10906
rect 50460 10854 50474 10906
rect 50474 10854 50486 10906
rect 50486 10854 50516 10906
rect 50540 10854 50550 10906
rect 50550 10854 50596 10906
rect 50300 10852 50356 10854
rect 50380 10852 50436 10854
rect 50460 10852 50516 10854
rect 50540 10852 50596 10854
rect 24398 4564 24400 4584
rect 24400 4564 24452 4584
rect 24452 4564 24454 4584
rect 24398 4528 24454 4564
rect 22834 3848 22890 3904
rect 26422 2896 26478 2952
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 65660 10362 65716 10364
rect 65740 10362 65796 10364
rect 65820 10362 65876 10364
rect 65900 10362 65956 10364
rect 65660 10310 65706 10362
rect 65706 10310 65716 10362
rect 65740 10310 65770 10362
rect 65770 10310 65782 10362
rect 65782 10310 65796 10362
rect 65820 10310 65834 10362
rect 65834 10310 65846 10362
rect 65846 10310 65876 10362
rect 65900 10310 65910 10362
rect 65910 10310 65956 10362
rect 65660 10308 65716 10310
rect 65740 10308 65796 10310
rect 65820 10308 65876 10310
rect 65900 10308 65956 10310
rect 50300 9818 50356 9820
rect 50380 9818 50436 9820
rect 50460 9818 50516 9820
rect 50540 9818 50596 9820
rect 50300 9766 50346 9818
rect 50346 9766 50356 9818
rect 50380 9766 50410 9818
rect 50410 9766 50422 9818
rect 50422 9766 50436 9818
rect 50460 9766 50474 9818
rect 50474 9766 50486 9818
rect 50486 9766 50516 9818
rect 50540 9766 50550 9818
rect 50550 9766 50596 9818
rect 50300 9764 50356 9766
rect 50380 9764 50436 9766
rect 50460 9764 50516 9766
rect 50540 9764 50596 9766
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 65660 9274 65716 9276
rect 65740 9274 65796 9276
rect 65820 9274 65876 9276
rect 65900 9274 65956 9276
rect 65660 9222 65706 9274
rect 65706 9222 65716 9274
rect 65740 9222 65770 9274
rect 65770 9222 65782 9274
rect 65782 9222 65796 9274
rect 65820 9222 65834 9274
rect 65834 9222 65846 9274
rect 65846 9222 65876 9274
rect 65900 9222 65910 9274
rect 65910 9222 65956 9274
rect 65660 9220 65716 9222
rect 65740 9220 65796 9222
rect 65820 9220 65876 9222
rect 65900 9220 65956 9222
rect 50300 8730 50356 8732
rect 50380 8730 50436 8732
rect 50460 8730 50516 8732
rect 50540 8730 50596 8732
rect 50300 8678 50346 8730
rect 50346 8678 50356 8730
rect 50380 8678 50410 8730
rect 50410 8678 50422 8730
rect 50422 8678 50436 8730
rect 50460 8678 50474 8730
rect 50474 8678 50486 8730
rect 50486 8678 50516 8730
rect 50540 8678 50550 8730
rect 50550 8678 50596 8730
rect 50300 8676 50356 8678
rect 50380 8676 50436 8678
rect 50460 8676 50516 8678
rect 50540 8676 50596 8678
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 65660 8186 65716 8188
rect 65740 8186 65796 8188
rect 65820 8186 65876 8188
rect 65900 8186 65956 8188
rect 65660 8134 65706 8186
rect 65706 8134 65716 8186
rect 65740 8134 65770 8186
rect 65770 8134 65782 8186
rect 65782 8134 65796 8186
rect 65820 8134 65834 8186
rect 65834 8134 65846 8186
rect 65846 8134 65876 8186
rect 65900 8134 65910 8186
rect 65910 8134 65956 8186
rect 65660 8132 65716 8134
rect 65740 8132 65796 8134
rect 65820 8132 65876 8134
rect 65900 8132 65956 8134
rect 50300 7642 50356 7644
rect 50380 7642 50436 7644
rect 50460 7642 50516 7644
rect 50540 7642 50596 7644
rect 50300 7590 50346 7642
rect 50346 7590 50356 7642
rect 50380 7590 50410 7642
rect 50410 7590 50422 7642
rect 50422 7590 50436 7642
rect 50460 7590 50474 7642
rect 50474 7590 50486 7642
rect 50486 7590 50516 7642
rect 50540 7590 50550 7642
rect 50550 7590 50596 7642
rect 50300 7588 50356 7590
rect 50380 7588 50436 7590
rect 50460 7588 50516 7590
rect 50540 7588 50596 7590
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 65660 7098 65716 7100
rect 65740 7098 65796 7100
rect 65820 7098 65876 7100
rect 65900 7098 65956 7100
rect 65660 7046 65706 7098
rect 65706 7046 65716 7098
rect 65740 7046 65770 7098
rect 65770 7046 65782 7098
rect 65782 7046 65796 7098
rect 65820 7046 65834 7098
rect 65834 7046 65846 7098
rect 65846 7046 65876 7098
rect 65900 7046 65910 7098
rect 65910 7046 65956 7098
rect 65660 7044 65716 7046
rect 65740 7044 65796 7046
rect 65820 7044 65876 7046
rect 65900 7044 65956 7046
rect 50300 6554 50356 6556
rect 50380 6554 50436 6556
rect 50460 6554 50516 6556
rect 50540 6554 50596 6556
rect 50300 6502 50346 6554
rect 50346 6502 50356 6554
rect 50380 6502 50410 6554
rect 50410 6502 50422 6554
rect 50422 6502 50436 6554
rect 50460 6502 50474 6554
rect 50474 6502 50486 6554
rect 50486 6502 50516 6554
rect 50540 6502 50550 6554
rect 50550 6502 50596 6554
rect 50300 6500 50356 6502
rect 50380 6500 50436 6502
rect 50460 6500 50516 6502
rect 50540 6500 50596 6502
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 65660 6010 65716 6012
rect 65740 6010 65796 6012
rect 65820 6010 65876 6012
rect 65900 6010 65956 6012
rect 65660 5958 65706 6010
rect 65706 5958 65716 6010
rect 65740 5958 65770 6010
rect 65770 5958 65782 6010
rect 65782 5958 65796 6010
rect 65820 5958 65834 6010
rect 65834 5958 65846 6010
rect 65846 5958 65876 6010
rect 65900 5958 65910 6010
rect 65910 5958 65956 6010
rect 65660 5956 65716 5958
rect 65740 5956 65796 5958
rect 65820 5956 65876 5958
rect 65900 5956 65956 5958
rect 50300 5466 50356 5468
rect 50380 5466 50436 5468
rect 50460 5466 50516 5468
rect 50540 5466 50596 5468
rect 50300 5414 50346 5466
rect 50346 5414 50356 5466
rect 50380 5414 50410 5466
rect 50410 5414 50422 5466
rect 50422 5414 50436 5466
rect 50460 5414 50474 5466
rect 50474 5414 50486 5466
rect 50486 5414 50516 5466
rect 50540 5414 50550 5466
rect 50550 5414 50596 5466
rect 50300 5412 50356 5414
rect 50380 5412 50436 5414
rect 50460 5412 50516 5414
rect 50540 5412 50596 5414
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 65660 4922 65716 4924
rect 65740 4922 65796 4924
rect 65820 4922 65876 4924
rect 65900 4922 65956 4924
rect 65660 4870 65706 4922
rect 65706 4870 65716 4922
rect 65740 4870 65770 4922
rect 65770 4870 65782 4922
rect 65782 4870 65796 4922
rect 65820 4870 65834 4922
rect 65834 4870 65846 4922
rect 65846 4870 65876 4922
rect 65900 4870 65910 4922
rect 65910 4870 65956 4922
rect 65660 4868 65716 4870
rect 65740 4868 65796 4870
rect 65820 4868 65876 4870
rect 65900 4868 65956 4870
rect 50300 4378 50356 4380
rect 50380 4378 50436 4380
rect 50460 4378 50516 4380
rect 50540 4378 50596 4380
rect 50300 4326 50346 4378
rect 50346 4326 50356 4378
rect 50380 4326 50410 4378
rect 50410 4326 50422 4378
rect 50422 4326 50436 4378
rect 50460 4326 50474 4378
rect 50474 4326 50486 4378
rect 50486 4326 50516 4378
rect 50540 4326 50550 4378
rect 50550 4326 50596 4378
rect 50300 4324 50356 4326
rect 50380 4324 50436 4326
rect 50460 4324 50516 4326
rect 50540 4324 50596 4326
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 65660 3834 65716 3836
rect 65740 3834 65796 3836
rect 65820 3834 65876 3836
rect 65900 3834 65956 3836
rect 65660 3782 65706 3834
rect 65706 3782 65716 3834
rect 65740 3782 65770 3834
rect 65770 3782 65782 3834
rect 65782 3782 65796 3834
rect 65820 3782 65834 3834
rect 65834 3782 65846 3834
rect 65846 3782 65876 3834
rect 65900 3782 65910 3834
rect 65910 3782 65956 3834
rect 65660 3780 65716 3782
rect 65740 3780 65796 3782
rect 65820 3780 65876 3782
rect 65900 3780 65956 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 50300 3290 50356 3292
rect 50380 3290 50436 3292
rect 50460 3290 50516 3292
rect 50540 3290 50596 3292
rect 50300 3238 50346 3290
rect 50346 3238 50356 3290
rect 50380 3238 50410 3290
rect 50410 3238 50422 3290
rect 50422 3238 50436 3290
rect 50460 3238 50474 3290
rect 50474 3238 50486 3290
rect 50486 3238 50516 3290
rect 50540 3238 50550 3290
rect 50550 3238 50596 3290
rect 50300 3236 50356 3238
rect 50380 3236 50436 3238
rect 50460 3236 50516 3238
rect 50540 3236 50596 3238
rect 50300 2202 50356 2204
rect 50380 2202 50436 2204
rect 50460 2202 50516 2204
rect 50540 2202 50596 2204
rect 50300 2150 50346 2202
rect 50346 2150 50356 2202
rect 50380 2150 50410 2202
rect 50410 2150 50422 2202
rect 50422 2150 50436 2202
rect 50460 2150 50474 2202
rect 50474 2150 50486 2202
rect 50486 2150 50516 2202
rect 50540 2150 50550 2202
rect 50550 2150 50596 2202
rect 50300 2148 50356 2150
rect 50380 2148 50436 2150
rect 50460 2148 50516 2150
rect 50540 2148 50596 2150
rect 65660 2746 65716 2748
rect 65740 2746 65796 2748
rect 65820 2746 65876 2748
rect 65900 2746 65956 2748
rect 65660 2694 65706 2746
rect 65706 2694 65716 2746
rect 65740 2694 65770 2746
rect 65770 2694 65782 2746
rect 65782 2694 65796 2746
rect 65820 2694 65834 2746
rect 65834 2694 65846 2746
rect 65846 2694 65876 2746
rect 65900 2694 65910 2746
rect 65910 2694 65956 2746
rect 65660 2692 65716 2694
rect 65740 2692 65796 2694
rect 65820 2692 65876 2694
rect 65900 2692 65956 2694
<< metal3 >>
rect 19570 57696 19886 57697
rect 19570 57632 19576 57696
rect 19640 57632 19656 57696
rect 19720 57632 19736 57696
rect 19800 57632 19816 57696
rect 19880 57632 19886 57696
rect 19570 57631 19886 57632
rect 50290 57696 50606 57697
rect 50290 57632 50296 57696
rect 50360 57632 50376 57696
rect 50440 57632 50456 57696
rect 50520 57632 50536 57696
rect 50600 57632 50606 57696
rect 50290 57631 50606 57632
rect 4210 57152 4526 57153
rect 4210 57088 4216 57152
rect 4280 57088 4296 57152
rect 4360 57088 4376 57152
rect 4440 57088 4456 57152
rect 4520 57088 4526 57152
rect 4210 57087 4526 57088
rect 34930 57152 35246 57153
rect 34930 57088 34936 57152
rect 35000 57088 35016 57152
rect 35080 57088 35096 57152
rect 35160 57088 35176 57152
rect 35240 57088 35246 57152
rect 34930 57087 35246 57088
rect 65650 57152 65966 57153
rect 65650 57088 65656 57152
rect 65720 57088 65736 57152
rect 65800 57088 65816 57152
rect 65880 57088 65896 57152
rect 65960 57088 65966 57152
rect 65650 57087 65966 57088
rect 19570 56608 19886 56609
rect 19570 56544 19576 56608
rect 19640 56544 19656 56608
rect 19720 56544 19736 56608
rect 19800 56544 19816 56608
rect 19880 56544 19886 56608
rect 19570 56543 19886 56544
rect 50290 56608 50606 56609
rect 50290 56544 50296 56608
rect 50360 56544 50376 56608
rect 50440 56544 50456 56608
rect 50520 56544 50536 56608
rect 50600 56544 50606 56608
rect 50290 56543 50606 56544
rect 4210 56064 4526 56065
rect 4210 56000 4216 56064
rect 4280 56000 4296 56064
rect 4360 56000 4376 56064
rect 4440 56000 4456 56064
rect 4520 56000 4526 56064
rect 4210 55999 4526 56000
rect 34930 56064 35246 56065
rect 34930 56000 34936 56064
rect 35000 56000 35016 56064
rect 35080 56000 35096 56064
rect 35160 56000 35176 56064
rect 35240 56000 35246 56064
rect 34930 55999 35246 56000
rect 65650 56064 65966 56065
rect 65650 56000 65656 56064
rect 65720 56000 65736 56064
rect 65800 56000 65816 56064
rect 65880 56000 65896 56064
rect 65960 56000 65966 56064
rect 65650 55999 65966 56000
rect 19570 55520 19886 55521
rect 19570 55456 19576 55520
rect 19640 55456 19656 55520
rect 19720 55456 19736 55520
rect 19800 55456 19816 55520
rect 19880 55456 19886 55520
rect 19570 55455 19886 55456
rect 50290 55520 50606 55521
rect 50290 55456 50296 55520
rect 50360 55456 50376 55520
rect 50440 55456 50456 55520
rect 50520 55456 50536 55520
rect 50600 55456 50606 55520
rect 50290 55455 50606 55456
rect 4210 54976 4526 54977
rect 4210 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4526 54976
rect 4210 54911 4526 54912
rect 34930 54976 35246 54977
rect 34930 54912 34936 54976
rect 35000 54912 35016 54976
rect 35080 54912 35096 54976
rect 35160 54912 35176 54976
rect 35240 54912 35246 54976
rect 34930 54911 35246 54912
rect 65650 54976 65966 54977
rect 65650 54912 65656 54976
rect 65720 54912 65736 54976
rect 65800 54912 65816 54976
rect 65880 54912 65896 54976
rect 65960 54912 65966 54976
rect 65650 54911 65966 54912
rect 19570 54432 19886 54433
rect 19570 54368 19576 54432
rect 19640 54368 19656 54432
rect 19720 54368 19736 54432
rect 19800 54368 19816 54432
rect 19880 54368 19886 54432
rect 19570 54367 19886 54368
rect 50290 54432 50606 54433
rect 50290 54368 50296 54432
rect 50360 54368 50376 54432
rect 50440 54368 50456 54432
rect 50520 54368 50536 54432
rect 50600 54368 50606 54432
rect 50290 54367 50606 54368
rect 4210 53888 4526 53889
rect 4210 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4526 53888
rect 4210 53823 4526 53824
rect 34930 53888 35246 53889
rect 34930 53824 34936 53888
rect 35000 53824 35016 53888
rect 35080 53824 35096 53888
rect 35160 53824 35176 53888
rect 35240 53824 35246 53888
rect 34930 53823 35246 53824
rect 65650 53888 65966 53889
rect 65650 53824 65656 53888
rect 65720 53824 65736 53888
rect 65800 53824 65816 53888
rect 65880 53824 65896 53888
rect 65960 53824 65966 53888
rect 65650 53823 65966 53824
rect 19570 53344 19886 53345
rect 19570 53280 19576 53344
rect 19640 53280 19656 53344
rect 19720 53280 19736 53344
rect 19800 53280 19816 53344
rect 19880 53280 19886 53344
rect 19570 53279 19886 53280
rect 50290 53344 50606 53345
rect 50290 53280 50296 53344
rect 50360 53280 50376 53344
rect 50440 53280 50456 53344
rect 50520 53280 50536 53344
rect 50600 53280 50606 53344
rect 50290 53279 50606 53280
rect 4210 52800 4526 52801
rect 4210 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4526 52800
rect 4210 52735 4526 52736
rect 34930 52800 35246 52801
rect 34930 52736 34936 52800
rect 35000 52736 35016 52800
rect 35080 52736 35096 52800
rect 35160 52736 35176 52800
rect 35240 52736 35246 52800
rect 34930 52735 35246 52736
rect 65650 52800 65966 52801
rect 65650 52736 65656 52800
rect 65720 52736 65736 52800
rect 65800 52736 65816 52800
rect 65880 52736 65896 52800
rect 65960 52736 65966 52800
rect 65650 52735 65966 52736
rect 19570 52256 19886 52257
rect 19570 52192 19576 52256
rect 19640 52192 19656 52256
rect 19720 52192 19736 52256
rect 19800 52192 19816 52256
rect 19880 52192 19886 52256
rect 19570 52191 19886 52192
rect 50290 52256 50606 52257
rect 50290 52192 50296 52256
rect 50360 52192 50376 52256
rect 50440 52192 50456 52256
rect 50520 52192 50536 52256
rect 50600 52192 50606 52256
rect 50290 52191 50606 52192
rect 4210 51712 4526 51713
rect 4210 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4526 51712
rect 4210 51647 4526 51648
rect 34930 51712 35246 51713
rect 34930 51648 34936 51712
rect 35000 51648 35016 51712
rect 35080 51648 35096 51712
rect 35160 51648 35176 51712
rect 35240 51648 35246 51712
rect 34930 51647 35246 51648
rect 65650 51712 65966 51713
rect 65650 51648 65656 51712
rect 65720 51648 65736 51712
rect 65800 51648 65816 51712
rect 65880 51648 65896 51712
rect 65960 51648 65966 51712
rect 65650 51647 65966 51648
rect 19570 51168 19886 51169
rect 19570 51104 19576 51168
rect 19640 51104 19656 51168
rect 19720 51104 19736 51168
rect 19800 51104 19816 51168
rect 19880 51104 19886 51168
rect 19570 51103 19886 51104
rect 50290 51168 50606 51169
rect 50290 51104 50296 51168
rect 50360 51104 50376 51168
rect 50440 51104 50456 51168
rect 50520 51104 50536 51168
rect 50600 51104 50606 51168
rect 50290 51103 50606 51104
rect 4210 50624 4526 50625
rect 4210 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4526 50624
rect 4210 50559 4526 50560
rect 34930 50624 35246 50625
rect 34930 50560 34936 50624
rect 35000 50560 35016 50624
rect 35080 50560 35096 50624
rect 35160 50560 35176 50624
rect 35240 50560 35246 50624
rect 34930 50559 35246 50560
rect 65650 50624 65966 50625
rect 65650 50560 65656 50624
rect 65720 50560 65736 50624
rect 65800 50560 65816 50624
rect 65880 50560 65896 50624
rect 65960 50560 65966 50624
rect 65650 50559 65966 50560
rect 19570 50080 19886 50081
rect 19570 50016 19576 50080
rect 19640 50016 19656 50080
rect 19720 50016 19736 50080
rect 19800 50016 19816 50080
rect 19880 50016 19886 50080
rect 19570 50015 19886 50016
rect 50290 50080 50606 50081
rect 50290 50016 50296 50080
rect 50360 50016 50376 50080
rect 50440 50016 50456 50080
rect 50520 50016 50536 50080
rect 50600 50016 50606 50080
rect 50290 50015 50606 50016
rect 4210 49536 4526 49537
rect 4210 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4526 49536
rect 4210 49471 4526 49472
rect 34930 49536 35246 49537
rect 34930 49472 34936 49536
rect 35000 49472 35016 49536
rect 35080 49472 35096 49536
rect 35160 49472 35176 49536
rect 35240 49472 35246 49536
rect 34930 49471 35246 49472
rect 65650 49536 65966 49537
rect 65650 49472 65656 49536
rect 65720 49472 65736 49536
rect 65800 49472 65816 49536
rect 65880 49472 65896 49536
rect 65960 49472 65966 49536
rect 65650 49471 65966 49472
rect 19570 48992 19886 48993
rect 19570 48928 19576 48992
rect 19640 48928 19656 48992
rect 19720 48928 19736 48992
rect 19800 48928 19816 48992
rect 19880 48928 19886 48992
rect 19570 48927 19886 48928
rect 50290 48992 50606 48993
rect 50290 48928 50296 48992
rect 50360 48928 50376 48992
rect 50440 48928 50456 48992
rect 50520 48928 50536 48992
rect 50600 48928 50606 48992
rect 50290 48927 50606 48928
rect 4210 48448 4526 48449
rect 4210 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4526 48448
rect 4210 48383 4526 48384
rect 34930 48448 35246 48449
rect 34930 48384 34936 48448
rect 35000 48384 35016 48448
rect 35080 48384 35096 48448
rect 35160 48384 35176 48448
rect 35240 48384 35246 48448
rect 34930 48383 35246 48384
rect 65650 48448 65966 48449
rect 65650 48384 65656 48448
rect 65720 48384 65736 48448
rect 65800 48384 65816 48448
rect 65880 48384 65896 48448
rect 65960 48384 65966 48448
rect 65650 48383 65966 48384
rect 19570 47904 19886 47905
rect 19570 47840 19576 47904
rect 19640 47840 19656 47904
rect 19720 47840 19736 47904
rect 19800 47840 19816 47904
rect 19880 47840 19886 47904
rect 19570 47839 19886 47840
rect 50290 47904 50606 47905
rect 50290 47840 50296 47904
rect 50360 47840 50376 47904
rect 50440 47840 50456 47904
rect 50520 47840 50536 47904
rect 50600 47840 50606 47904
rect 50290 47839 50606 47840
rect 4210 47360 4526 47361
rect 4210 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4526 47360
rect 4210 47295 4526 47296
rect 34930 47360 35246 47361
rect 34930 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35246 47360
rect 34930 47295 35246 47296
rect 65650 47360 65966 47361
rect 65650 47296 65656 47360
rect 65720 47296 65736 47360
rect 65800 47296 65816 47360
rect 65880 47296 65896 47360
rect 65960 47296 65966 47360
rect 65650 47295 65966 47296
rect 19570 46816 19886 46817
rect 19570 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19886 46816
rect 19570 46751 19886 46752
rect 50290 46816 50606 46817
rect 50290 46752 50296 46816
rect 50360 46752 50376 46816
rect 50440 46752 50456 46816
rect 50520 46752 50536 46816
rect 50600 46752 50606 46816
rect 50290 46751 50606 46752
rect 4210 46272 4526 46273
rect 4210 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4526 46272
rect 4210 46207 4526 46208
rect 34930 46272 35246 46273
rect 34930 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35246 46272
rect 34930 46207 35246 46208
rect 65650 46272 65966 46273
rect 65650 46208 65656 46272
rect 65720 46208 65736 46272
rect 65800 46208 65816 46272
rect 65880 46208 65896 46272
rect 65960 46208 65966 46272
rect 65650 46207 65966 46208
rect 19570 45728 19886 45729
rect 19570 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19886 45728
rect 19570 45663 19886 45664
rect 50290 45728 50606 45729
rect 50290 45664 50296 45728
rect 50360 45664 50376 45728
rect 50440 45664 50456 45728
rect 50520 45664 50536 45728
rect 50600 45664 50606 45728
rect 50290 45663 50606 45664
rect 4210 45184 4526 45185
rect 4210 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4526 45184
rect 4210 45119 4526 45120
rect 34930 45184 35246 45185
rect 34930 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35246 45184
rect 34930 45119 35246 45120
rect 65650 45184 65966 45185
rect 65650 45120 65656 45184
rect 65720 45120 65736 45184
rect 65800 45120 65816 45184
rect 65880 45120 65896 45184
rect 65960 45120 65966 45184
rect 65650 45119 65966 45120
rect 19570 44640 19886 44641
rect 19570 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19886 44640
rect 19570 44575 19886 44576
rect 50290 44640 50606 44641
rect 50290 44576 50296 44640
rect 50360 44576 50376 44640
rect 50440 44576 50456 44640
rect 50520 44576 50536 44640
rect 50600 44576 50606 44640
rect 50290 44575 50606 44576
rect 4210 44096 4526 44097
rect 4210 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4526 44096
rect 4210 44031 4526 44032
rect 34930 44096 35246 44097
rect 34930 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35246 44096
rect 34930 44031 35246 44032
rect 65650 44096 65966 44097
rect 65650 44032 65656 44096
rect 65720 44032 65736 44096
rect 65800 44032 65816 44096
rect 65880 44032 65896 44096
rect 65960 44032 65966 44096
rect 65650 44031 65966 44032
rect 19570 43552 19886 43553
rect 19570 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19886 43552
rect 19570 43487 19886 43488
rect 50290 43552 50606 43553
rect 50290 43488 50296 43552
rect 50360 43488 50376 43552
rect 50440 43488 50456 43552
rect 50520 43488 50536 43552
rect 50600 43488 50606 43552
rect 50290 43487 50606 43488
rect 4210 43008 4526 43009
rect 4210 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4526 43008
rect 4210 42943 4526 42944
rect 34930 43008 35246 43009
rect 34930 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35246 43008
rect 34930 42943 35246 42944
rect 65650 43008 65966 43009
rect 65650 42944 65656 43008
rect 65720 42944 65736 43008
rect 65800 42944 65816 43008
rect 65880 42944 65896 43008
rect 65960 42944 65966 43008
rect 65650 42943 65966 42944
rect 19570 42464 19886 42465
rect 19570 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19886 42464
rect 19570 42399 19886 42400
rect 50290 42464 50606 42465
rect 50290 42400 50296 42464
rect 50360 42400 50376 42464
rect 50440 42400 50456 42464
rect 50520 42400 50536 42464
rect 50600 42400 50606 42464
rect 50290 42399 50606 42400
rect 4210 41920 4526 41921
rect 4210 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4526 41920
rect 4210 41855 4526 41856
rect 34930 41920 35246 41921
rect 34930 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35246 41920
rect 34930 41855 35246 41856
rect 65650 41920 65966 41921
rect 65650 41856 65656 41920
rect 65720 41856 65736 41920
rect 65800 41856 65816 41920
rect 65880 41856 65896 41920
rect 65960 41856 65966 41920
rect 65650 41855 65966 41856
rect 19570 41376 19886 41377
rect 19570 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19886 41376
rect 19570 41311 19886 41312
rect 50290 41376 50606 41377
rect 50290 41312 50296 41376
rect 50360 41312 50376 41376
rect 50440 41312 50456 41376
rect 50520 41312 50536 41376
rect 50600 41312 50606 41376
rect 50290 41311 50606 41312
rect 4210 40832 4526 40833
rect 4210 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4526 40832
rect 4210 40767 4526 40768
rect 34930 40832 35246 40833
rect 34930 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35246 40832
rect 34930 40767 35246 40768
rect 65650 40832 65966 40833
rect 65650 40768 65656 40832
rect 65720 40768 65736 40832
rect 65800 40768 65816 40832
rect 65880 40768 65896 40832
rect 65960 40768 65966 40832
rect 65650 40767 65966 40768
rect 19570 40288 19886 40289
rect 19570 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19886 40288
rect 19570 40223 19886 40224
rect 50290 40288 50606 40289
rect 50290 40224 50296 40288
rect 50360 40224 50376 40288
rect 50440 40224 50456 40288
rect 50520 40224 50536 40288
rect 50600 40224 50606 40288
rect 50290 40223 50606 40224
rect 4210 39744 4526 39745
rect 4210 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4526 39744
rect 4210 39679 4526 39680
rect 34930 39744 35246 39745
rect 34930 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35246 39744
rect 34930 39679 35246 39680
rect 65650 39744 65966 39745
rect 65650 39680 65656 39744
rect 65720 39680 65736 39744
rect 65800 39680 65816 39744
rect 65880 39680 65896 39744
rect 65960 39680 65966 39744
rect 65650 39679 65966 39680
rect 19570 39200 19886 39201
rect 19570 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19886 39200
rect 19570 39135 19886 39136
rect 50290 39200 50606 39201
rect 50290 39136 50296 39200
rect 50360 39136 50376 39200
rect 50440 39136 50456 39200
rect 50520 39136 50536 39200
rect 50600 39136 50606 39200
rect 50290 39135 50606 39136
rect 4210 38656 4526 38657
rect 4210 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4526 38656
rect 4210 38591 4526 38592
rect 34930 38656 35246 38657
rect 34930 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35246 38656
rect 34930 38591 35246 38592
rect 65650 38656 65966 38657
rect 65650 38592 65656 38656
rect 65720 38592 65736 38656
rect 65800 38592 65816 38656
rect 65880 38592 65896 38656
rect 65960 38592 65966 38656
rect 65650 38591 65966 38592
rect 19570 38112 19886 38113
rect 19570 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19886 38112
rect 19570 38047 19886 38048
rect 50290 38112 50606 38113
rect 50290 38048 50296 38112
rect 50360 38048 50376 38112
rect 50440 38048 50456 38112
rect 50520 38048 50536 38112
rect 50600 38048 50606 38112
rect 50290 38047 50606 38048
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 65650 37568 65966 37569
rect 65650 37504 65656 37568
rect 65720 37504 65736 37568
rect 65800 37504 65816 37568
rect 65880 37504 65896 37568
rect 65960 37504 65966 37568
rect 65650 37503 65966 37504
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 50290 37024 50606 37025
rect 50290 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50606 37024
rect 50290 36959 50606 36960
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 65650 36480 65966 36481
rect 65650 36416 65656 36480
rect 65720 36416 65736 36480
rect 65800 36416 65816 36480
rect 65880 36416 65896 36480
rect 65960 36416 65966 36480
rect 65650 36415 65966 36416
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 50290 35936 50606 35937
rect 50290 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50606 35936
rect 50290 35871 50606 35872
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 65650 35392 65966 35393
rect 65650 35328 65656 35392
rect 65720 35328 65736 35392
rect 65800 35328 65816 35392
rect 65880 35328 65896 35392
rect 65960 35328 65966 35392
rect 65650 35327 65966 35328
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 50290 34848 50606 34849
rect 50290 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50606 34848
rect 50290 34783 50606 34784
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 65650 34304 65966 34305
rect 65650 34240 65656 34304
rect 65720 34240 65736 34304
rect 65800 34240 65816 34304
rect 65880 34240 65896 34304
rect 65960 34240 65966 34304
rect 65650 34239 65966 34240
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 50290 33760 50606 33761
rect 50290 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50606 33760
rect 50290 33695 50606 33696
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 65650 33216 65966 33217
rect 65650 33152 65656 33216
rect 65720 33152 65736 33216
rect 65800 33152 65816 33216
rect 65880 33152 65896 33216
rect 65960 33152 65966 33216
rect 65650 33151 65966 33152
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 19570 32607 19886 32608
rect 50290 32672 50606 32673
rect 50290 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50606 32672
rect 50290 32607 50606 32608
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 65650 32128 65966 32129
rect 65650 32064 65656 32128
rect 65720 32064 65736 32128
rect 65800 32064 65816 32128
rect 65880 32064 65896 32128
rect 65960 32064 65966 32128
rect 65650 32063 65966 32064
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 50290 31584 50606 31585
rect 50290 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50606 31584
rect 50290 31519 50606 31520
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 65650 31040 65966 31041
rect 65650 30976 65656 31040
rect 65720 30976 65736 31040
rect 65800 30976 65816 31040
rect 65880 30976 65896 31040
rect 65960 30976 65966 31040
rect 65650 30975 65966 30976
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 50290 30496 50606 30497
rect 50290 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50606 30496
rect 50290 30431 50606 30432
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 65650 29952 65966 29953
rect 65650 29888 65656 29952
rect 65720 29888 65736 29952
rect 65800 29888 65816 29952
rect 65880 29888 65896 29952
rect 65960 29888 65966 29952
rect 65650 29887 65966 29888
rect 19570 29408 19886 29409
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 50290 29408 50606 29409
rect 50290 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50606 29408
rect 50290 29343 50606 29344
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 65650 28864 65966 28865
rect 65650 28800 65656 28864
rect 65720 28800 65736 28864
rect 65800 28800 65816 28864
rect 65880 28800 65896 28864
rect 65960 28800 65966 28864
rect 65650 28799 65966 28800
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 50290 28320 50606 28321
rect 50290 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50606 28320
rect 50290 28255 50606 28256
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 65650 27776 65966 27777
rect 65650 27712 65656 27776
rect 65720 27712 65736 27776
rect 65800 27712 65816 27776
rect 65880 27712 65896 27776
rect 65960 27712 65966 27776
rect 65650 27711 65966 27712
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 19570 27167 19886 27168
rect 50290 27232 50606 27233
rect 50290 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50606 27232
rect 50290 27167 50606 27168
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 65650 26688 65966 26689
rect 65650 26624 65656 26688
rect 65720 26624 65736 26688
rect 65800 26624 65816 26688
rect 65880 26624 65896 26688
rect 65960 26624 65966 26688
rect 65650 26623 65966 26624
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 50290 26144 50606 26145
rect 50290 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50606 26144
rect 50290 26079 50606 26080
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 65650 25600 65966 25601
rect 65650 25536 65656 25600
rect 65720 25536 65736 25600
rect 65800 25536 65816 25600
rect 65880 25536 65896 25600
rect 65960 25536 65966 25600
rect 65650 25535 65966 25536
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 50290 25056 50606 25057
rect 50290 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50606 25056
rect 50290 24991 50606 24992
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 65650 24512 65966 24513
rect 65650 24448 65656 24512
rect 65720 24448 65736 24512
rect 65800 24448 65816 24512
rect 65880 24448 65896 24512
rect 65960 24448 65966 24512
rect 65650 24447 65966 24448
rect 19570 23968 19886 23969
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 50290 23968 50606 23969
rect 50290 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50606 23968
rect 50290 23903 50606 23904
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 65650 23424 65966 23425
rect 65650 23360 65656 23424
rect 65720 23360 65736 23424
rect 65800 23360 65816 23424
rect 65880 23360 65896 23424
rect 65960 23360 65966 23424
rect 65650 23359 65966 23360
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 50290 22880 50606 22881
rect 50290 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50606 22880
rect 50290 22815 50606 22816
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 65650 22336 65966 22337
rect 65650 22272 65656 22336
rect 65720 22272 65736 22336
rect 65800 22272 65816 22336
rect 65880 22272 65896 22336
rect 65960 22272 65966 22336
rect 65650 22271 65966 22272
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 19570 21727 19886 21728
rect 50290 21792 50606 21793
rect 50290 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50606 21792
rect 50290 21727 50606 21728
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 65650 21248 65966 21249
rect 65650 21184 65656 21248
rect 65720 21184 65736 21248
rect 65800 21184 65816 21248
rect 65880 21184 65896 21248
rect 65960 21184 65966 21248
rect 65650 21183 65966 21184
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 50290 20704 50606 20705
rect 50290 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50606 20704
rect 50290 20639 50606 20640
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 65650 20160 65966 20161
rect 65650 20096 65656 20160
rect 65720 20096 65736 20160
rect 65800 20096 65816 20160
rect 65880 20096 65896 20160
rect 65960 20096 65966 20160
rect 65650 20095 65966 20096
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 50290 19616 50606 19617
rect 50290 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50606 19616
rect 50290 19551 50606 19552
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 65650 19072 65966 19073
rect 65650 19008 65656 19072
rect 65720 19008 65736 19072
rect 65800 19008 65816 19072
rect 65880 19008 65896 19072
rect 65960 19008 65966 19072
rect 65650 19007 65966 19008
rect 19570 18528 19886 18529
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 50290 18528 50606 18529
rect 50290 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50606 18528
rect 50290 18463 50606 18464
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 65650 17984 65966 17985
rect 65650 17920 65656 17984
rect 65720 17920 65736 17984
rect 65800 17920 65816 17984
rect 65880 17920 65896 17984
rect 65960 17920 65966 17984
rect 65650 17919 65966 17920
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 50290 17440 50606 17441
rect 50290 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50606 17440
rect 50290 17375 50606 17376
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 65650 16896 65966 16897
rect 65650 16832 65656 16896
rect 65720 16832 65736 16896
rect 65800 16832 65816 16896
rect 65880 16832 65896 16896
rect 65960 16832 65966 16896
rect 65650 16831 65966 16832
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 50290 16352 50606 16353
rect 50290 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50606 16352
rect 50290 16287 50606 16288
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 65650 15808 65966 15809
rect 65650 15744 65656 15808
rect 65720 15744 65736 15808
rect 65800 15744 65816 15808
rect 65880 15744 65896 15808
rect 65960 15744 65966 15808
rect 65650 15743 65966 15744
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 50290 15264 50606 15265
rect 50290 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50606 15264
rect 50290 15199 50606 15200
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 65650 14720 65966 14721
rect 65650 14656 65656 14720
rect 65720 14656 65736 14720
rect 65800 14656 65816 14720
rect 65880 14656 65896 14720
rect 65960 14656 65966 14720
rect 65650 14655 65966 14656
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 50290 14176 50606 14177
rect 50290 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50606 14176
rect 50290 14111 50606 14112
rect 11697 13698 11763 13701
rect 12893 13698 12959 13701
rect 11697 13696 12959 13698
rect 11697 13640 11702 13696
rect 11758 13640 12898 13696
rect 12954 13640 12959 13696
rect 11697 13638 12959 13640
rect 11697 13635 11763 13638
rect 12893 13635 12959 13638
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 65650 13632 65966 13633
rect 65650 13568 65656 13632
rect 65720 13568 65736 13632
rect 65800 13568 65816 13632
rect 65880 13568 65896 13632
rect 65960 13568 65966 13632
rect 65650 13567 65966 13568
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 50290 13088 50606 13089
rect 50290 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50606 13088
rect 50290 13023 50606 13024
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 65650 12544 65966 12545
rect 65650 12480 65656 12544
rect 65720 12480 65736 12544
rect 65800 12480 65816 12544
rect 65880 12480 65896 12544
rect 65960 12480 65966 12544
rect 65650 12479 65966 12480
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 50290 12000 50606 12001
rect 50290 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50606 12000
rect 50290 11935 50606 11936
rect 16665 11522 16731 11525
rect 16798 11522 16804 11524
rect 16665 11520 16804 11522
rect 16665 11464 16670 11520
rect 16726 11464 16804 11520
rect 16665 11462 16804 11464
rect 16665 11459 16731 11462
rect 16798 11460 16804 11462
rect 16868 11460 16874 11524
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 65650 11456 65966 11457
rect 65650 11392 65656 11456
rect 65720 11392 65736 11456
rect 65800 11392 65816 11456
rect 65880 11392 65896 11456
rect 65960 11392 65966 11456
rect 65650 11391 65966 11392
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 19570 10847 19886 10848
rect 50290 10912 50606 10913
rect 50290 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50606 10912
rect 50290 10847 50606 10848
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 65650 10368 65966 10369
rect 65650 10304 65656 10368
rect 65720 10304 65736 10368
rect 65800 10304 65816 10368
rect 65880 10304 65896 10368
rect 65960 10304 65966 10368
rect 65650 10303 65966 10304
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 50290 9824 50606 9825
rect 50290 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50606 9824
rect 50290 9759 50606 9760
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 65650 9280 65966 9281
rect 65650 9216 65656 9280
rect 65720 9216 65736 9280
rect 65800 9216 65816 9280
rect 65880 9216 65896 9280
rect 65960 9216 65966 9280
rect 65650 9215 65966 9216
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 50290 8736 50606 8737
rect 50290 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50606 8736
rect 50290 8671 50606 8672
rect 21541 8530 21607 8533
rect 24301 8530 24367 8533
rect 21541 8528 24367 8530
rect 21541 8472 21546 8528
rect 21602 8472 24306 8528
rect 24362 8472 24367 8528
rect 21541 8470 24367 8472
rect 21541 8467 21607 8470
rect 24301 8467 24367 8470
rect 6862 8332 6868 8396
rect 6932 8394 6938 8396
rect 13629 8394 13695 8397
rect 6932 8392 13695 8394
rect 6932 8336 13634 8392
rect 13690 8336 13695 8392
rect 6932 8334 13695 8336
rect 6932 8332 6938 8334
rect 13629 8331 13695 8334
rect 21265 8394 21331 8397
rect 22921 8394 22987 8397
rect 21265 8392 22987 8394
rect 21265 8336 21270 8392
rect 21326 8336 22926 8392
rect 22982 8336 22987 8392
rect 21265 8334 22987 8336
rect 21265 8331 21331 8334
rect 22921 8331 22987 8334
rect 20253 8258 20319 8261
rect 22553 8258 22619 8261
rect 20253 8256 22619 8258
rect 20253 8200 20258 8256
rect 20314 8200 22558 8256
rect 22614 8200 22619 8256
rect 20253 8198 22619 8200
rect 20253 8195 20319 8198
rect 22553 8195 22619 8198
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 65650 8192 65966 8193
rect 65650 8128 65656 8192
rect 65720 8128 65736 8192
rect 65800 8128 65816 8192
rect 65880 8128 65896 8192
rect 65960 8128 65966 8192
rect 65650 8127 65966 8128
rect 9397 7850 9463 7853
rect 15009 7850 15075 7853
rect 9397 7848 15075 7850
rect 9397 7792 9402 7848
rect 9458 7792 15014 7848
rect 15070 7792 15075 7848
rect 9397 7790 15075 7792
rect 9397 7787 9463 7790
rect 15009 7787 15075 7790
rect 19570 7648 19886 7649
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 50290 7648 50606 7649
rect 50290 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50606 7648
rect 50290 7583 50606 7584
rect 9581 7170 9647 7173
rect 14641 7170 14707 7173
rect 9581 7168 14707 7170
rect 9581 7112 9586 7168
rect 9642 7112 14646 7168
rect 14702 7112 14707 7168
rect 9581 7110 14707 7112
rect 9581 7107 9647 7110
rect 14641 7107 14707 7110
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 65650 7104 65966 7105
rect 65650 7040 65656 7104
rect 65720 7040 65736 7104
rect 65800 7040 65816 7104
rect 65880 7040 65896 7104
rect 65960 7040 65966 7104
rect 65650 7039 65966 7040
rect 5257 6898 5323 6901
rect 11329 6898 11395 6901
rect 5257 6896 11395 6898
rect 5257 6840 5262 6896
rect 5318 6840 11334 6896
rect 11390 6840 11395 6896
rect 5257 6838 11395 6840
rect 5257 6835 5323 6838
rect 11329 6835 11395 6838
rect 4981 6762 5047 6765
rect 12065 6762 12131 6765
rect 4981 6760 12131 6762
rect 4981 6704 4986 6760
rect 5042 6704 12070 6760
rect 12126 6704 12131 6760
rect 4981 6702 12131 6704
rect 4981 6699 5047 6702
rect 12065 6699 12131 6702
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 50290 6560 50606 6561
rect 50290 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50606 6560
rect 50290 6495 50606 6496
rect 20437 6354 20503 6357
rect 20662 6354 20668 6356
rect 20437 6352 20668 6354
rect 20437 6296 20442 6352
rect 20498 6296 20668 6352
rect 20437 6294 20668 6296
rect 20437 6291 20503 6294
rect 20662 6292 20668 6294
rect 20732 6292 20738 6356
rect 11605 6218 11671 6221
rect 12750 6218 12756 6220
rect 11605 6216 12756 6218
rect 11605 6160 11610 6216
rect 11666 6160 12756 6216
rect 11605 6158 12756 6160
rect 11605 6155 11671 6158
rect 12750 6156 12756 6158
rect 12820 6218 12826 6220
rect 20805 6218 20871 6221
rect 12820 6216 20871 6218
rect 12820 6160 20810 6216
rect 20866 6160 20871 6216
rect 12820 6158 20871 6160
rect 12820 6156 12826 6158
rect 20805 6155 20871 6158
rect 8661 6082 8727 6085
rect 12801 6082 12867 6085
rect 13629 6082 13695 6085
rect 8661 6080 13695 6082
rect 8661 6024 8666 6080
rect 8722 6024 12806 6080
rect 12862 6024 13634 6080
rect 13690 6024 13695 6080
rect 8661 6022 13695 6024
rect 8661 6019 8727 6022
rect 12801 6019 12867 6022
rect 13629 6019 13695 6022
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 65650 6016 65966 6017
rect 65650 5952 65656 6016
rect 65720 5952 65736 6016
rect 65800 5952 65816 6016
rect 65880 5952 65896 6016
rect 65960 5952 65966 6016
rect 65650 5951 65966 5952
rect 9029 5810 9095 5813
rect 14181 5810 14247 5813
rect 20437 5810 20503 5813
rect 9029 5808 20503 5810
rect 9029 5752 9034 5808
rect 9090 5752 14186 5808
rect 14242 5752 20442 5808
rect 20498 5752 20503 5808
rect 9029 5750 20503 5752
rect 9029 5747 9095 5750
rect 14181 5747 14247 5750
rect 20437 5747 20503 5750
rect 6821 5674 6887 5677
rect 9489 5674 9555 5677
rect 6821 5672 9555 5674
rect 6821 5616 6826 5672
rect 6882 5616 9494 5672
rect 9550 5616 9555 5672
rect 6821 5614 9555 5616
rect 6821 5611 6887 5614
rect 9489 5611 9555 5614
rect 11237 5674 11303 5677
rect 13118 5674 13124 5676
rect 11237 5672 13124 5674
rect 11237 5616 11242 5672
rect 11298 5616 13124 5672
rect 11237 5614 13124 5616
rect 11237 5611 11303 5614
rect 13118 5612 13124 5614
rect 13188 5612 13194 5676
rect 17033 5674 17099 5677
rect 17902 5674 17908 5676
rect 17033 5672 17908 5674
rect 17033 5616 17038 5672
rect 17094 5616 17908 5672
rect 17033 5614 17908 5616
rect 17033 5611 17099 5614
rect 17902 5612 17908 5614
rect 17972 5612 17978 5676
rect 20437 5538 20503 5541
rect 22093 5538 22159 5541
rect 20437 5536 22159 5538
rect 20437 5480 20442 5536
rect 20498 5480 22098 5536
rect 22154 5480 22159 5536
rect 20437 5478 22159 5480
rect 20437 5475 20503 5478
rect 22093 5475 22159 5478
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 19570 5407 19886 5408
rect 50290 5472 50606 5473
rect 50290 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50606 5472
rect 50290 5407 50606 5408
rect 19977 5402 20043 5405
rect 20253 5402 20319 5405
rect 19977 5400 20319 5402
rect 19977 5344 19982 5400
rect 20038 5344 20258 5400
rect 20314 5344 20319 5400
rect 19977 5342 20319 5344
rect 19977 5339 20043 5342
rect 20253 5339 20319 5342
rect 11789 5266 11855 5269
rect 13629 5266 13695 5269
rect 23197 5266 23263 5269
rect 11789 5264 23263 5266
rect 11789 5208 11794 5264
rect 11850 5208 13634 5264
rect 13690 5208 23202 5264
rect 23258 5208 23263 5264
rect 11789 5206 23263 5208
rect 11789 5203 11855 5206
rect 13629 5203 13695 5206
rect 23197 5203 23263 5206
rect 19333 5130 19399 5133
rect 19977 5130 20043 5133
rect 19333 5128 20043 5130
rect 19333 5072 19338 5128
rect 19394 5072 19982 5128
rect 20038 5072 20043 5128
rect 19333 5070 20043 5072
rect 19333 5067 19399 5070
rect 19977 5067 20043 5070
rect 19374 4932 19380 4996
rect 19444 4994 19450 4996
rect 19793 4994 19859 4997
rect 19444 4992 19859 4994
rect 19444 4936 19798 4992
rect 19854 4936 19859 4992
rect 19444 4934 19859 4936
rect 19444 4932 19450 4934
rect 19793 4931 19859 4934
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 65650 4928 65966 4929
rect 65650 4864 65656 4928
rect 65720 4864 65736 4928
rect 65800 4864 65816 4928
rect 65880 4864 65896 4928
rect 65960 4864 65966 4928
rect 65650 4863 65966 4864
rect 12065 4858 12131 4861
rect 15929 4858 15995 4861
rect 16798 4858 16804 4860
rect 12065 4856 15762 4858
rect 12065 4800 12070 4856
rect 12126 4800 15762 4856
rect 12065 4798 15762 4800
rect 12065 4795 12131 4798
rect 5717 4722 5783 4725
rect 14365 4722 14431 4725
rect 5717 4720 14431 4722
rect 5717 4664 5722 4720
rect 5778 4664 14370 4720
rect 14426 4664 14431 4720
rect 5717 4662 14431 4664
rect 15702 4722 15762 4798
rect 15929 4856 16804 4858
rect 15929 4800 15934 4856
rect 15990 4800 16804 4856
rect 15929 4798 16804 4800
rect 15929 4795 15995 4798
rect 16798 4796 16804 4798
rect 16868 4796 16874 4860
rect 16665 4722 16731 4725
rect 15702 4720 16731 4722
rect 15702 4664 16670 4720
rect 16726 4664 16731 4720
rect 15702 4662 16731 4664
rect 5717 4659 5783 4662
rect 14365 4659 14431 4662
rect 16665 4659 16731 4662
rect 9489 4586 9555 4589
rect 15101 4586 15167 4589
rect 9489 4584 15167 4586
rect 9489 4528 9494 4584
rect 9550 4528 15106 4584
rect 15162 4528 15167 4584
rect 9489 4526 15167 4528
rect 9489 4523 9555 4526
rect 15101 4523 15167 4526
rect 19609 4586 19675 4589
rect 21081 4586 21147 4589
rect 24393 4586 24459 4589
rect 19609 4584 24459 4586
rect 19609 4528 19614 4584
rect 19670 4528 21086 4584
rect 21142 4528 24398 4584
rect 24454 4528 24459 4584
rect 19609 4526 24459 4528
rect 19609 4523 19675 4526
rect 21081 4523 21147 4526
rect 24393 4523 24459 4526
rect 6545 4450 6611 4453
rect 12525 4450 12591 4453
rect 6545 4448 12591 4450
rect 6545 4392 6550 4448
rect 6606 4392 12530 4448
rect 12586 4392 12591 4448
rect 6545 4390 12591 4392
rect 6545 4387 6611 4390
rect 12525 4387 12591 4390
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 50290 4384 50606 4385
rect 50290 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50606 4384
rect 50290 4319 50606 4320
rect 7925 4314 7991 4317
rect 12985 4314 13051 4317
rect 7925 4312 13051 4314
rect 7925 4256 7930 4312
rect 7986 4256 12990 4312
rect 13046 4256 13051 4312
rect 7925 4254 13051 4256
rect 7925 4251 7991 4254
rect 12985 4251 13051 4254
rect 3877 4178 3943 4181
rect 12433 4178 12499 4181
rect 3877 4176 12499 4178
rect 3877 4120 3882 4176
rect 3938 4120 12438 4176
rect 12494 4120 12499 4176
rect 3877 4118 12499 4120
rect 3877 4115 3943 4118
rect 12433 4115 12499 4118
rect 6269 4042 6335 4045
rect 6862 4042 6868 4044
rect 6269 4040 6868 4042
rect 6269 3984 6274 4040
rect 6330 3984 6868 4040
rect 6269 3982 6868 3984
rect 6269 3979 6335 3982
rect 6862 3980 6868 3982
rect 6932 3980 6938 4044
rect 17902 3980 17908 4044
rect 17972 4042 17978 4044
rect 22093 4042 22159 4045
rect 17972 4040 22159 4042
rect 17972 3984 22098 4040
rect 22154 3984 22159 4040
rect 17972 3982 22159 3984
rect 17972 3980 17978 3982
rect 22093 3979 22159 3982
rect 19333 3906 19399 3909
rect 22829 3906 22895 3909
rect 19333 3904 22895 3906
rect 19333 3848 19338 3904
rect 19394 3848 22834 3904
rect 22890 3848 22895 3904
rect 19333 3846 22895 3848
rect 19333 3843 19399 3846
rect 22829 3843 22895 3846
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 65650 3840 65966 3841
rect 65650 3776 65656 3840
rect 65720 3776 65736 3840
rect 65800 3776 65816 3840
rect 65880 3776 65896 3840
rect 65960 3776 65966 3840
rect 65650 3775 65966 3776
rect 5073 3770 5139 3773
rect 8937 3770 9003 3773
rect 5073 3768 12450 3770
rect 5073 3712 5078 3768
rect 5134 3712 8942 3768
rect 8998 3712 12450 3768
rect 5073 3710 12450 3712
rect 5073 3707 5139 3710
rect 8937 3707 9003 3710
rect 4245 3634 4311 3637
rect 8109 3634 8175 3637
rect 4245 3632 8175 3634
rect 4245 3576 4250 3632
rect 4306 3576 8114 3632
rect 8170 3576 8175 3632
rect 4245 3574 8175 3576
rect 12390 3634 12450 3710
rect 13261 3634 13327 3637
rect 12390 3632 13327 3634
rect 12390 3576 13266 3632
rect 13322 3576 13327 3632
rect 12390 3574 13327 3576
rect 4245 3571 4311 3574
rect 8109 3571 8175 3574
rect 13261 3571 13327 3574
rect 15285 3634 15351 3637
rect 16205 3634 16271 3637
rect 15285 3632 16271 3634
rect 15285 3576 15290 3632
rect 15346 3576 16210 3632
rect 16266 3576 16271 3632
rect 15285 3574 16271 3576
rect 15285 3571 15351 3574
rect 16205 3571 16271 3574
rect 4797 3498 4863 3501
rect 8201 3498 8267 3501
rect 4797 3496 8267 3498
rect 4797 3440 4802 3496
rect 4858 3440 8206 3496
rect 8262 3440 8267 3496
rect 4797 3438 8267 3440
rect 4797 3435 4863 3438
rect 8201 3435 8267 3438
rect 9673 3498 9739 3501
rect 19374 3498 19380 3500
rect 9673 3496 19380 3498
rect 9673 3440 9678 3496
rect 9734 3440 19380 3496
rect 9673 3438 19380 3440
rect 9673 3435 9739 3438
rect 19374 3436 19380 3438
rect 19444 3436 19450 3500
rect 4521 3362 4587 3365
rect 11697 3362 11763 3365
rect 4521 3360 11763 3362
rect 4521 3304 4526 3360
rect 4582 3304 11702 3360
rect 11758 3304 11763 3360
rect 4521 3302 11763 3304
rect 4521 3299 4587 3302
rect 11697 3299 11763 3302
rect 12750 3300 12756 3364
rect 12820 3362 12826 3364
rect 12893 3362 12959 3365
rect 12820 3360 12959 3362
rect 12820 3304 12898 3360
rect 12954 3304 12959 3360
rect 12820 3302 12959 3304
rect 12820 3300 12826 3302
rect 12893 3299 12959 3302
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 50290 3296 50606 3297
rect 50290 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50606 3296
rect 50290 3231 50606 3232
rect 13537 3226 13603 3229
rect 15469 3226 15535 3229
rect 13537 3224 15535 3226
rect 13537 3168 13542 3224
rect 13598 3168 15474 3224
rect 15530 3168 15535 3224
rect 13537 3166 15535 3168
rect 13537 3163 13603 3166
rect 15469 3163 15535 3166
rect 13118 3028 13124 3092
rect 13188 3090 13194 3092
rect 13721 3090 13787 3093
rect 20713 3092 20779 3093
rect 13188 3088 13787 3090
rect 13188 3032 13726 3088
rect 13782 3032 13787 3088
rect 13188 3030 13787 3032
rect 13188 3028 13194 3030
rect 13721 3027 13787 3030
rect 20662 3028 20668 3092
rect 20732 3090 20779 3092
rect 20732 3088 20824 3090
rect 20774 3032 20824 3088
rect 20732 3030 20824 3032
rect 20732 3028 20779 3030
rect 20713 3027 20779 3028
rect 10225 2954 10291 2957
rect 26417 2954 26483 2957
rect 10225 2952 26483 2954
rect 10225 2896 10230 2952
rect 10286 2896 26422 2952
rect 26478 2896 26483 2952
rect 10225 2894 26483 2896
rect 10225 2891 10291 2894
rect 26417 2891 26483 2894
rect 6729 2818 6795 2821
rect 14457 2818 14523 2821
rect 6729 2816 14523 2818
rect 6729 2760 6734 2816
rect 6790 2760 14462 2816
rect 14518 2760 14523 2816
rect 6729 2758 14523 2760
rect 6729 2755 6795 2758
rect 14457 2755 14523 2758
rect 19057 2818 19123 2821
rect 20069 2818 20135 2821
rect 19057 2816 20135 2818
rect 19057 2760 19062 2816
rect 19118 2760 20074 2816
rect 20130 2760 20135 2816
rect 19057 2758 20135 2760
rect 19057 2755 19123 2758
rect 20069 2755 20135 2758
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 65650 2752 65966 2753
rect 65650 2688 65656 2752
rect 65720 2688 65736 2752
rect 65800 2688 65816 2752
rect 65880 2688 65896 2752
rect 65960 2688 65966 2752
rect 65650 2687 65966 2688
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
rect 50290 2208 50606 2209
rect 50290 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50606 2208
rect 50290 2143 50606 2144
<< via3 >>
rect 19576 57692 19640 57696
rect 19576 57636 19580 57692
rect 19580 57636 19636 57692
rect 19636 57636 19640 57692
rect 19576 57632 19640 57636
rect 19656 57692 19720 57696
rect 19656 57636 19660 57692
rect 19660 57636 19716 57692
rect 19716 57636 19720 57692
rect 19656 57632 19720 57636
rect 19736 57692 19800 57696
rect 19736 57636 19740 57692
rect 19740 57636 19796 57692
rect 19796 57636 19800 57692
rect 19736 57632 19800 57636
rect 19816 57692 19880 57696
rect 19816 57636 19820 57692
rect 19820 57636 19876 57692
rect 19876 57636 19880 57692
rect 19816 57632 19880 57636
rect 50296 57692 50360 57696
rect 50296 57636 50300 57692
rect 50300 57636 50356 57692
rect 50356 57636 50360 57692
rect 50296 57632 50360 57636
rect 50376 57692 50440 57696
rect 50376 57636 50380 57692
rect 50380 57636 50436 57692
rect 50436 57636 50440 57692
rect 50376 57632 50440 57636
rect 50456 57692 50520 57696
rect 50456 57636 50460 57692
rect 50460 57636 50516 57692
rect 50516 57636 50520 57692
rect 50456 57632 50520 57636
rect 50536 57692 50600 57696
rect 50536 57636 50540 57692
rect 50540 57636 50596 57692
rect 50596 57636 50600 57692
rect 50536 57632 50600 57636
rect 4216 57148 4280 57152
rect 4216 57092 4220 57148
rect 4220 57092 4276 57148
rect 4276 57092 4280 57148
rect 4216 57088 4280 57092
rect 4296 57148 4360 57152
rect 4296 57092 4300 57148
rect 4300 57092 4356 57148
rect 4356 57092 4360 57148
rect 4296 57088 4360 57092
rect 4376 57148 4440 57152
rect 4376 57092 4380 57148
rect 4380 57092 4436 57148
rect 4436 57092 4440 57148
rect 4376 57088 4440 57092
rect 4456 57148 4520 57152
rect 4456 57092 4460 57148
rect 4460 57092 4516 57148
rect 4516 57092 4520 57148
rect 4456 57088 4520 57092
rect 34936 57148 35000 57152
rect 34936 57092 34940 57148
rect 34940 57092 34996 57148
rect 34996 57092 35000 57148
rect 34936 57088 35000 57092
rect 35016 57148 35080 57152
rect 35016 57092 35020 57148
rect 35020 57092 35076 57148
rect 35076 57092 35080 57148
rect 35016 57088 35080 57092
rect 35096 57148 35160 57152
rect 35096 57092 35100 57148
rect 35100 57092 35156 57148
rect 35156 57092 35160 57148
rect 35096 57088 35160 57092
rect 35176 57148 35240 57152
rect 35176 57092 35180 57148
rect 35180 57092 35236 57148
rect 35236 57092 35240 57148
rect 35176 57088 35240 57092
rect 65656 57148 65720 57152
rect 65656 57092 65660 57148
rect 65660 57092 65716 57148
rect 65716 57092 65720 57148
rect 65656 57088 65720 57092
rect 65736 57148 65800 57152
rect 65736 57092 65740 57148
rect 65740 57092 65796 57148
rect 65796 57092 65800 57148
rect 65736 57088 65800 57092
rect 65816 57148 65880 57152
rect 65816 57092 65820 57148
rect 65820 57092 65876 57148
rect 65876 57092 65880 57148
rect 65816 57088 65880 57092
rect 65896 57148 65960 57152
rect 65896 57092 65900 57148
rect 65900 57092 65956 57148
rect 65956 57092 65960 57148
rect 65896 57088 65960 57092
rect 19576 56604 19640 56608
rect 19576 56548 19580 56604
rect 19580 56548 19636 56604
rect 19636 56548 19640 56604
rect 19576 56544 19640 56548
rect 19656 56604 19720 56608
rect 19656 56548 19660 56604
rect 19660 56548 19716 56604
rect 19716 56548 19720 56604
rect 19656 56544 19720 56548
rect 19736 56604 19800 56608
rect 19736 56548 19740 56604
rect 19740 56548 19796 56604
rect 19796 56548 19800 56604
rect 19736 56544 19800 56548
rect 19816 56604 19880 56608
rect 19816 56548 19820 56604
rect 19820 56548 19876 56604
rect 19876 56548 19880 56604
rect 19816 56544 19880 56548
rect 50296 56604 50360 56608
rect 50296 56548 50300 56604
rect 50300 56548 50356 56604
rect 50356 56548 50360 56604
rect 50296 56544 50360 56548
rect 50376 56604 50440 56608
rect 50376 56548 50380 56604
rect 50380 56548 50436 56604
rect 50436 56548 50440 56604
rect 50376 56544 50440 56548
rect 50456 56604 50520 56608
rect 50456 56548 50460 56604
rect 50460 56548 50516 56604
rect 50516 56548 50520 56604
rect 50456 56544 50520 56548
rect 50536 56604 50600 56608
rect 50536 56548 50540 56604
rect 50540 56548 50596 56604
rect 50596 56548 50600 56604
rect 50536 56544 50600 56548
rect 4216 56060 4280 56064
rect 4216 56004 4220 56060
rect 4220 56004 4276 56060
rect 4276 56004 4280 56060
rect 4216 56000 4280 56004
rect 4296 56060 4360 56064
rect 4296 56004 4300 56060
rect 4300 56004 4356 56060
rect 4356 56004 4360 56060
rect 4296 56000 4360 56004
rect 4376 56060 4440 56064
rect 4376 56004 4380 56060
rect 4380 56004 4436 56060
rect 4436 56004 4440 56060
rect 4376 56000 4440 56004
rect 4456 56060 4520 56064
rect 4456 56004 4460 56060
rect 4460 56004 4516 56060
rect 4516 56004 4520 56060
rect 4456 56000 4520 56004
rect 34936 56060 35000 56064
rect 34936 56004 34940 56060
rect 34940 56004 34996 56060
rect 34996 56004 35000 56060
rect 34936 56000 35000 56004
rect 35016 56060 35080 56064
rect 35016 56004 35020 56060
rect 35020 56004 35076 56060
rect 35076 56004 35080 56060
rect 35016 56000 35080 56004
rect 35096 56060 35160 56064
rect 35096 56004 35100 56060
rect 35100 56004 35156 56060
rect 35156 56004 35160 56060
rect 35096 56000 35160 56004
rect 35176 56060 35240 56064
rect 35176 56004 35180 56060
rect 35180 56004 35236 56060
rect 35236 56004 35240 56060
rect 35176 56000 35240 56004
rect 65656 56060 65720 56064
rect 65656 56004 65660 56060
rect 65660 56004 65716 56060
rect 65716 56004 65720 56060
rect 65656 56000 65720 56004
rect 65736 56060 65800 56064
rect 65736 56004 65740 56060
rect 65740 56004 65796 56060
rect 65796 56004 65800 56060
rect 65736 56000 65800 56004
rect 65816 56060 65880 56064
rect 65816 56004 65820 56060
rect 65820 56004 65876 56060
rect 65876 56004 65880 56060
rect 65816 56000 65880 56004
rect 65896 56060 65960 56064
rect 65896 56004 65900 56060
rect 65900 56004 65956 56060
rect 65956 56004 65960 56060
rect 65896 56000 65960 56004
rect 19576 55516 19640 55520
rect 19576 55460 19580 55516
rect 19580 55460 19636 55516
rect 19636 55460 19640 55516
rect 19576 55456 19640 55460
rect 19656 55516 19720 55520
rect 19656 55460 19660 55516
rect 19660 55460 19716 55516
rect 19716 55460 19720 55516
rect 19656 55456 19720 55460
rect 19736 55516 19800 55520
rect 19736 55460 19740 55516
rect 19740 55460 19796 55516
rect 19796 55460 19800 55516
rect 19736 55456 19800 55460
rect 19816 55516 19880 55520
rect 19816 55460 19820 55516
rect 19820 55460 19876 55516
rect 19876 55460 19880 55516
rect 19816 55456 19880 55460
rect 50296 55516 50360 55520
rect 50296 55460 50300 55516
rect 50300 55460 50356 55516
rect 50356 55460 50360 55516
rect 50296 55456 50360 55460
rect 50376 55516 50440 55520
rect 50376 55460 50380 55516
rect 50380 55460 50436 55516
rect 50436 55460 50440 55516
rect 50376 55456 50440 55460
rect 50456 55516 50520 55520
rect 50456 55460 50460 55516
rect 50460 55460 50516 55516
rect 50516 55460 50520 55516
rect 50456 55456 50520 55460
rect 50536 55516 50600 55520
rect 50536 55460 50540 55516
rect 50540 55460 50596 55516
rect 50596 55460 50600 55516
rect 50536 55456 50600 55460
rect 4216 54972 4280 54976
rect 4216 54916 4220 54972
rect 4220 54916 4276 54972
rect 4276 54916 4280 54972
rect 4216 54912 4280 54916
rect 4296 54972 4360 54976
rect 4296 54916 4300 54972
rect 4300 54916 4356 54972
rect 4356 54916 4360 54972
rect 4296 54912 4360 54916
rect 4376 54972 4440 54976
rect 4376 54916 4380 54972
rect 4380 54916 4436 54972
rect 4436 54916 4440 54972
rect 4376 54912 4440 54916
rect 4456 54972 4520 54976
rect 4456 54916 4460 54972
rect 4460 54916 4516 54972
rect 4516 54916 4520 54972
rect 4456 54912 4520 54916
rect 34936 54972 35000 54976
rect 34936 54916 34940 54972
rect 34940 54916 34996 54972
rect 34996 54916 35000 54972
rect 34936 54912 35000 54916
rect 35016 54972 35080 54976
rect 35016 54916 35020 54972
rect 35020 54916 35076 54972
rect 35076 54916 35080 54972
rect 35016 54912 35080 54916
rect 35096 54972 35160 54976
rect 35096 54916 35100 54972
rect 35100 54916 35156 54972
rect 35156 54916 35160 54972
rect 35096 54912 35160 54916
rect 35176 54972 35240 54976
rect 35176 54916 35180 54972
rect 35180 54916 35236 54972
rect 35236 54916 35240 54972
rect 35176 54912 35240 54916
rect 65656 54972 65720 54976
rect 65656 54916 65660 54972
rect 65660 54916 65716 54972
rect 65716 54916 65720 54972
rect 65656 54912 65720 54916
rect 65736 54972 65800 54976
rect 65736 54916 65740 54972
rect 65740 54916 65796 54972
rect 65796 54916 65800 54972
rect 65736 54912 65800 54916
rect 65816 54972 65880 54976
rect 65816 54916 65820 54972
rect 65820 54916 65876 54972
rect 65876 54916 65880 54972
rect 65816 54912 65880 54916
rect 65896 54972 65960 54976
rect 65896 54916 65900 54972
rect 65900 54916 65956 54972
rect 65956 54916 65960 54972
rect 65896 54912 65960 54916
rect 19576 54428 19640 54432
rect 19576 54372 19580 54428
rect 19580 54372 19636 54428
rect 19636 54372 19640 54428
rect 19576 54368 19640 54372
rect 19656 54428 19720 54432
rect 19656 54372 19660 54428
rect 19660 54372 19716 54428
rect 19716 54372 19720 54428
rect 19656 54368 19720 54372
rect 19736 54428 19800 54432
rect 19736 54372 19740 54428
rect 19740 54372 19796 54428
rect 19796 54372 19800 54428
rect 19736 54368 19800 54372
rect 19816 54428 19880 54432
rect 19816 54372 19820 54428
rect 19820 54372 19876 54428
rect 19876 54372 19880 54428
rect 19816 54368 19880 54372
rect 50296 54428 50360 54432
rect 50296 54372 50300 54428
rect 50300 54372 50356 54428
rect 50356 54372 50360 54428
rect 50296 54368 50360 54372
rect 50376 54428 50440 54432
rect 50376 54372 50380 54428
rect 50380 54372 50436 54428
rect 50436 54372 50440 54428
rect 50376 54368 50440 54372
rect 50456 54428 50520 54432
rect 50456 54372 50460 54428
rect 50460 54372 50516 54428
rect 50516 54372 50520 54428
rect 50456 54368 50520 54372
rect 50536 54428 50600 54432
rect 50536 54372 50540 54428
rect 50540 54372 50596 54428
rect 50596 54372 50600 54428
rect 50536 54368 50600 54372
rect 4216 53884 4280 53888
rect 4216 53828 4220 53884
rect 4220 53828 4276 53884
rect 4276 53828 4280 53884
rect 4216 53824 4280 53828
rect 4296 53884 4360 53888
rect 4296 53828 4300 53884
rect 4300 53828 4356 53884
rect 4356 53828 4360 53884
rect 4296 53824 4360 53828
rect 4376 53884 4440 53888
rect 4376 53828 4380 53884
rect 4380 53828 4436 53884
rect 4436 53828 4440 53884
rect 4376 53824 4440 53828
rect 4456 53884 4520 53888
rect 4456 53828 4460 53884
rect 4460 53828 4516 53884
rect 4516 53828 4520 53884
rect 4456 53824 4520 53828
rect 34936 53884 35000 53888
rect 34936 53828 34940 53884
rect 34940 53828 34996 53884
rect 34996 53828 35000 53884
rect 34936 53824 35000 53828
rect 35016 53884 35080 53888
rect 35016 53828 35020 53884
rect 35020 53828 35076 53884
rect 35076 53828 35080 53884
rect 35016 53824 35080 53828
rect 35096 53884 35160 53888
rect 35096 53828 35100 53884
rect 35100 53828 35156 53884
rect 35156 53828 35160 53884
rect 35096 53824 35160 53828
rect 35176 53884 35240 53888
rect 35176 53828 35180 53884
rect 35180 53828 35236 53884
rect 35236 53828 35240 53884
rect 35176 53824 35240 53828
rect 65656 53884 65720 53888
rect 65656 53828 65660 53884
rect 65660 53828 65716 53884
rect 65716 53828 65720 53884
rect 65656 53824 65720 53828
rect 65736 53884 65800 53888
rect 65736 53828 65740 53884
rect 65740 53828 65796 53884
rect 65796 53828 65800 53884
rect 65736 53824 65800 53828
rect 65816 53884 65880 53888
rect 65816 53828 65820 53884
rect 65820 53828 65876 53884
rect 65876 53828 65880 53884
rect 65816 53824 65880 53828
rect 65896 53884 65960 53888
rect 65896 53828 65900 53884
rect 65900 53828 65956 53884
rect 65956 53828 65960 53884
rect 65896 53824 65960 53828
rect 19576 53340 19640 53344
rect 19576 53284 19580 53340
rect 19580 53284 19636 53340
rect 19636 53284 19640 53340
rect 19576 53280 19640 53284
rect 19656 53340 19720 53344
rect 19656 53284 19660 53340
rect 19660 53284 19716 53340
rect 19716 53284 19720 53340
rect 19656 53280 19720 53284
rect 19736 53340 19800 53344
rect 19736 53284 19740 53340
rect 19740 53284 19796 53340
rect 19796 53284 19800 53340
rect 19736 53280 19800 53284
rect 19816 53340 19880 53344
rect 19816 53284 19820 53340
rect 19820 53284 19876 53340
rect 19876 53284 19880 53340
rect 19816 53280 19880 53284
rect 50296 53340 50360 53344
rect 50296 53284 50300 53340
rect 50300 53284 50356 53340
rect 50356 53284 50360 53340
rect 50296 53280 50360 53284
rect 50376 53340 50440 53344
rect 50376 53284 50380 53340
rect 50380 53284 50436 53340
rect 50436 53284 50440 53340
rect 50376 53280 50440 53284
rect 50456 53340 50520 53344
rect 50456 53284 50460 53340
rect 50460 53284 50516 53340
rect 50516 53284 50520 53340
rect 50456 53280 50520 53284
rect 50536 53340 50600 53344
rect 50536 53284 50540 53340
rect 50540 53284 50596 53340
rect 50596 53284 50600 53340
rect 50536 53280 50600 53284
rect 4216 52796 4280 52800
rect 4216 52740 4220 52796
rect 4220 52740 4276 52796
rect 4276 52740 4280 52796
rect 4216 52736 4280 52740
rect 4296 52796 4360 52800
rect 4296 52740 4300 52796
rect 4300 52740 4356 52796
rect 4356 52740 4360 52796
rect 4296 52736 4360 52740
rect 4376 52796 4440 52800
rect 4376 52740 4380 52796
rect 4380 52740 4436 52796
rect 4436 52740 4440 52796
rect 4376 52736 4440 52740
rect 4456 52796 4520 52800
rect 4456 52740 4460 52796
rect 4460 52740 4516 52796
rect 4516 52740 4520 52796
rect 4456 52736 4520 52740
rect 34936 52796 35000 52800
rect 34936 52740 34940 52796
rect 34940 52740 34996 52796
rect 34996 52740 35000 52796
rect 34936 52736 35000 52740
rect 35016 52796 35080 52800
rect 35016 52740 35020 52796
rect 35020 52740 35076 52796
rect 35076 52740 35080 52796
rect 35016 52736 35080 52740
rect 35096 52796 35160 52800
rect 35096 52740 35100 52796
rect 35100 52740 35156 52796
rect 35156 52740 35160 52796
rect 35096 52736 35160 52740
rect 35176 52796 35240 52800
rect 35176 52740 35180 52796
rect 35180 52740 35236 52796
rect 35236 52740 35240 52796
rect 35176 52736 35240 52740
rect 65656 52796 65720 52800
rect 65656 52740 65660 52796
rect 65660 52740 65716 52796
rect 65716 52740 65720 52796
rect 65656 52736 65720 52740
rect 65736 52796 65800 52800
rect 65736 52740 65740 52796
rect 65740 52740 65796 52796
rect 65796 52740 65800 52796
rect 65736 52736 65800 52740
rect 65816 52796 65880 52800
rect 65816 52740 65820 52796
rect 65820 52740 65876 52796
rect 65876 52740 65880 52796
rect 65816 52736 65880 52740
rect 65896 52796 65960 52800
rect 65896 52740 65900 52796
rect 65900 52740 65956 52796
rect 65956 52740 65960 52796
rect 65896 52736 65960 52740
rect 19576 52252 19640 52256
rect 19576 52196 19580 52252
rect 19580 52196 19636 52252
rect 19636 52196 19640 52252
rect 19576 52192 19640 52196
rect 19656 52252 19720 52256
rect 19656 52196 19660 52252
rect 19660 52196 19716 52252
rect 19716 52196 19720 52252
rect 19656 52192 19720 52196
rect 19736 52252 19800 52256
rect 19736 52196 19740 52252
rect 19740 52196 19796 52252
rect 19796 52196 19800 52252
rect 19736 52192 19800 52196
rect 19816 52252 19880 52256
rect 19816 52196 19820 52252
rect 19820 52196 19876 52252
rect 19876 52196 19880 52252
rect 19816 52192 19880 52196
rect 50296 52252 50360 52256
rect 50296 52196 50300 52252
rect 50300 52196 50356 52252
rect 50356 52196 50360 52252
rect 50296 52192 50360 52196
rect 50376 52252 50440 52256
rect 50376 52196 50380 52252
rect 50380 52196 50436 52252
rect 50436 52196 50440 52252
rect 50376 52192 50440 52196
rect 50456 52252 50520 52256
rect 50456 52196 50460 52252
rect 50460 52196 50516 52252
rect 50516 52196 50520 52252
rect 50456 52192 50520 52196
rect 50536 52252 50600 52256
rect 50536 52196 50540 52252
rect 50540 52196 50596 52252
rect 50596 52196 50600 52252
rect 50536 52192 50600 52196
rect 4216 51708 4280 51712
rect 4216 51652 4220 51708
rect 4220 51652 4276 51708
rect 4276 51652 4280 51708
rect 4216 51648 4280 51652
rect 4296 51708 4360 51712
rect 4296 51652 4300 51708
rect 4300 51652 4356 51708
rect 4356 51652 4360 51708
rect 4296 51648 4360 51652
rect 4376 51708 4440 51712
rect 4376 51652 4380 51708
rect 4380 51652 4436 51708
rect 4436 51652 4440 51708
rect 4376 51648 4440 51652
rect 4456 51708 4520 51712
rect 4456 51652 4460 51708
rect 4460 51652 4516 51708
rect 4516 51652 4520 51708
rect 4456 51648 4520 51652
rect 34936 51708 35000 51712
rect 34936 51652 34940 51708
rect 34940 51652 34996 51708
rect 34996 51652 35000 51708
rect 34936 51648 35000 51652
rect 35016 51708 35080 51712
rect 35016 51652 35020 51708
rect 35020 51652 35076 51708
rect 35076 51652 35080 51708
rect 35016 51648 35080 51652
rect 35096 51708 35160 51712
rect 35096 51652 35100 51708
rect 35100 51652 35156 51708
rect 35156 51652 35160 51708
rect 35096 51648 35160 51652
rect 35176 51708 35240 51712
rect 35176 51652 35180 51708
rect 35180 51652 35236 51708
rect 35236 51652 35240 51708
rect 35176 51648 35240 51652
rect 65656 51708 65720 51712
rect 65656 51652 65660 51708
rect 65660 51652 65716 51708
rect 65716 51652 65720 51708
rect 65656 51648 65720 51652
rect 65736 51708 65800 51712
rect 65736 51652 65740 51708
rect 65740 51652 65796 51708
rect 65796 51652 65800 51708
rect 65736 51648 65800 51652
rect 65816 51708 65880 51712
rect 65816 51652 65820 51708
rect 65820 51652 65876 51708
rect 65876 51652 65880 51708
rect 65816 51648 65880 51652
rect 65896 51708 65960 51712
rect 65896 51652 65900 51708
rect 65900 51652 65956 51708
rect 65956 51652 65960 51708
rect 65896 51648 65960 51652
rect 19576 51164 19640 51168
rect 19576 51108 19580 51164
rect 19580 51108 19636 51164
rect 19636 51108 19640 51164
rect 19576 51104 19640 51108
rect 19656 51164 19720 51168
rect 19656 51108 19660 51164
rect 19660 51108 19716 51164
rect 19716 51108 19720 51164
rect 19656 51104 19720 51108
rect 19736 51164 19800 51168
rect 19736 51108 19740 51164
rect 19740 51108 19796 51164
rect 19796 51108 19800 51164
rect 19736 51104 19800 51108
rect 19816 51164 19880 51168
rect 19816 51108 19820 51164
rect 19820 51108 19876 51164
rect 19876 51108 19880 51164
rect 19816 51104 19880 51108
rect 50296 51164 50360 51168
rect 50296 51108 50300 51164
rect 50300 51108 50356 51164
rect 50356 51108 50360 51164
rect 50296 51104 50360 51108
rect 50376 51164 50440 51168
rect 50376 51108 50380 51164
rect 50380 51108 50436 51164
rect 50436 51108 50440 51164
rect 50376 51104 50440 51108
rect 50456 51164 50520 51168
rect 50456 51108 50460 51164
rect 50460 51108 50516 51164
rect 50516 51108 50520 51164
rect 50456 51104 50520 51108
rect 50536 51164 50600 51168
rect 50536 51108 50540 51164
rect 50540 51108 50596 51164
rect 50596 51108 50600 51164
rect 50536 51104 50600 51108
rect 4216 50620 4280 50624
rect 4216 50564 4220 50620
rect 4220 50564 4276 50620
rect 4276 50564 4280 50620
rect 4216 50560 4280 50564
rect 4296 50620 4360 50624
rect 4296 50564 4300 50620
rect 4300 50564 4356 50620
rect 4356 50564 4360 50620
rect 4296 50560 4360 50564
rect 4376 50620 4440 50624
rect 4376 50564 4380 50620
rect 4380 50564 4436 50620
rect 4436 50564 4440 50620
rect 4376 50560 4440 50564
rect 4456 50620 4520 50624
rect 4456 50564 4460 50620
rect 4460 50564 4516 50620
rect 4516 50564 4520 50620
rect 4456 50560 4520 50564
rect 34936 50620 35000 50624
rect 34936 50564 34940 50620
rect 34940 50564 34996 50620
rect 34996 50564 35000 50620
rect 34936 50560 35000 50564
rect 35016 50620 35080 50624
rect 35016 50564 35020 50620
rect 35020 50564 35076 50620
rect 35076 50564 35080 50620
rect 35016 50560 35080 50564
rect 35096 50620 35160 50624
rect 35096 50564 35100 50620
rect 35100 50564 35156 50620
rect 35156 50564 35160 50620
rect 35096 50560 35160 50564
rect 35176 50620 35240 50624
rect 35176 50564 35180 50620
rect 35180 50564 35236 50620
rect 35236 50564 35240 50620
rect 35176 50560 35240 50564
rect 65656 50620 65720 50624
rect 65656 50564 65660 50620
rect 65660 50564 65716 50620
rect 65716 50564 65720 50620
rect 65656 50560 65720 50564
rect 65736 50620 65800 50624
rect 65736 50564 65740 50620
rect 65740 50564 65796 50620
rect 65796 50564 65800 50620
rect 65736 50560 65800 50564
rect 65816 50620 65880 50624
rect 65816 50564 65820 50620
rect 65820 50564 65876 50620
rect 65876 50564 65880 50620
rect 65816 50560 65880 50564
rect 65896 50620 65960 50624
rect 65896 50564 65900 50620
rect 65900 50564 65956 50620
rect 65956 50564 65960 50620
rect 65896 50560 65960 50564
rect 19576 50076 19640 50080
rect 19576 50020 19580 50076
rect 19580 50020 19636 50076
rect 19636 50020 19640 50076
rect 19576 50016 19640 50020
rect 19656 50076 19720 50080
rect 19656 50020 19660 50076
rect 19660 50020 19716 50076
rect 19716 50020 19720 50076
rect 19656 50016 19720 50020
rect 19736 50076 19800 50080
rect 19736 50020 19740 50076
rect 19740 50020 19796 50076
rect 19796 50020 19800 50076
rect 19736 50016 19800 50020
rect 19816 50076 19880 50080
rect 19816 50020 19820 50076
rect 19820 50020 19876 50076
rect 19876 50020 19880 50076
rect 19816 50016 19880 50020
rect 50296 50076 50360 50080
rect 50296 50020 50300 50076
rect 50300 50020 50356 50076
rect 50356 50020 50360 50076
rect 50296 50016 50360 50020
rect 50376 50076 50440 50080
rect 50376 50020 50380 50076
rect 50380 50020 50436 50076
rect 50436 50020 50440 50076
rect 50376 50016 50440 50020
rect 50456 50076 50520 50080
rect 50456 50020 50460 50076
rect 50460 50020 50516 50076
rect 50516 50020 50520 50076
rect 50456 50016 50520 50020
rect 50536 50076 50600 50080
rect 50536 50020 50540 50076
rect 50540 50020 50596 50076
rect 50596 50020 50600 50076
rect 50536 50016 50600 50020
rect 4216 49532 4280 49536
rect 4216 49476 4220 49532
rect 4220 49476 4276 49532
rect 4276 49476 4280 49532
rect 4216 49472 4280 49476
rect 4296 49532 4360 49536
rect 4296 49476 4300 49532
rect 4300 49476 4356 49532
rect 4356 49476 4360 49532
rect 4296 49472 4360 49476
rect 4376 49532 4440 49536
rect 4376 49476 4380 49532
rect 4380 49476 4436 49532
rect 4436 49476 4440 49532
rect 4376 49472 4440 49476
rect 4456 49532 4520 49536
rect 4456 49476 4460 49532
rect 4460 49476 4516 49532
rect 4516 49476 4520 49532
rect 4456 49472 4520 49476
rect 34936 49532 35000 49536
rect 34936 49476 34940 49532
rect 34940 49476 34996 49532
rect 34996 49476 35000 49532
rect 34936 49472 35000 49476
rect 35016 49532 35080 49536
rect 35016 49476 35020 49532
rect 35020 49476 35076 49532
rect 35076 49476 35080 49532
rect 35016 49472 35080 49476
rect 35096 49532 35160 49536
rect 35096 49476 35100 49532
rect 35100 49476 35156 49532
rect 35156 49476 35160 49532
rect 35096 49472 35160 49476
rect 35176 49532 35240 49536
rect 35176 49476 35180 49532
rect 35180 49476 35236 49532
rect 35236 49476 35240 49532
rect 35176 49472 35240 49476
rect 65656 49532 65720 49536
rect 65656 49476 65660 49532
rect 65660 49476 65716 49532
rect 65716 49476 65720 49532
rect 65656 49472 65720 49476
rect 65736 49532 65800 49536
rect 65736 49476 65740 49532
rect 65740 49476 65796 49532
rect 65796 49476 65800 49532
rect 65736 49472 65800 49476
rect 65816 49532 65880 49536
rect 65816 49476 65820 49532
rect 65820 49476 65876 49532
rect 65876 49476 65880 49532
rect 65816 49472 65880 49476
rect 65896 49532 65960 49536
rect 65896 49476 65900 49532
rect 65900 49476 65956 49532
rect 65956 49476 65960 49532
rect 65896 49472 65960 49476
rect 19576 48988 19640 48992
rect 19576 48932 19580 48988
rect 19580 48932 19636 48988
rect 19636 48932 19640 48988
rect 19576 48928 19640 48932
rect 19656 48988 19720 48992
rect 19656 48932 19660 48988
rect 19660 48932 19716 48988
rect 19716 48932 19720 48988
rect 19656 48928 19720 48932
rect 19736 48988 19800 48992
rect 19736 48932 19740 48988
rect 19740 48932 19796 48988
rect 19796 48932 19800 48988
rect 19736 48928 19800 48932
rect 19816 48988 19880 48992
rect 19816 48932 19820 48988
rect 19820 48932 19876 48988
rect 19876 48932 19880 48988
rect 19816 48928 19880 48932
rect 50296 48988 50360 48992
rect 50296 48932 50300 48988
rect 50300 48932 50356 48988
rect 50356 48932 50360 48988
rect 50296 48928 50360 48932
rect 50376 48988 50440 48992
rect 50376 48932 50380 48988
rect 50380 48932 50436 48988
rect 50436 48932 50440 48988
rect 50376 48928 50440 48932
rect 50456 48988 50520 48992
rect 50456 48932 50460 48988
rect 50460 48932 50516 48988
rect 50516 48932 50520 48988
rect 50456 48928 50520 48932
rect 50536 48988 50600 48992
rect 50536 48932 50540 48988
rect 50540 48932 50596 48988
rect 50596 48932 50600 48988
rect 50536 48928 50600 48932
rect 4216 48444 4280 48448
rect 4216 48388 4220 48444
rect 4220 48388 4276 48444
rect 4276 48388 4280 48444
rect 4216 48384 4280 48388
rect 4296 48444 4360 48448
rect 4296 48388 4300 48444
rect 4300 48388 4356 48444
rect 4356 48388 4360 48444
rect 4296 48384 4360 48388
rect 4376 48444 4440 48448
rect 4376 48388 4380 48444
rect 4380 48388 4436 48444
rect 4436 48388 4440 48444
rect 4376 48384 4440 48388
rect 4456 48444 4520 48448
rect 4456 48388 4460 48444
rect 4460 48388 4516 48444
rect 4516 48388 4520 48444
rect 4456 48384 4520 48388
rect 34936 48444 35000 48448
rect 34936 48388 34940 48444
rect 34940 48388 34996 48444
rect 34996 48388 35000 48444
rect 34936 48384 35000 48388
rect 35016 48444 35080 48448
rect 35016 48388 35020 48444
rect 35020 48388 35076 48444
rect 35076 48388 35080 48444
rect 35016 48384 35080 48388
rect 35096 48444 35160 48448
rect 35096 48388 35100 48444
rect 35100 48388 35156 48444
rect 35156 48388 35160 48444
rect 35096 48384 35160 48388
rect 35176 48444 35240 48448
rect 35176 48388 35180 48444
rect 35180 48388 35236 48444
rect 35236 48388 35240 48444
rect 35176 48384 35240 48388
rect 65656 48444 65720 48448
rect 65656 48388 65660 48444
rect 65660 48388 65716 48444
rect 65716 48388 65720 48444
rect 65656 48384 65720 48388
rect 65736 48444 65800 48448
rect 65736 48388 65740 48444
rect 65740 48388 65796 48444
rect 65796 48388 65800 48444
rect 65736 48384 65800 48388
rect 65816 48444 65880 48448
rect 65816 48388 65820 48444
rect 65820 48388 65876 48444
rect 65876 48388 65880 48444
rect 65816 48384 65880 48388
rect 65896 48444 65960 48448
rect 65896 48388 65900 48444
rect 65900 48388 65956 48444
rect 65956 48388 65960 48444
rect 65896 48384 65960 48388
rect 19576 47900 19640 47904
rect 19576 47844 19580 47900
rect 19580 47844 19636 47900
rect 19636 47844 19640 47900
rect 19576 47840 19640 47844
rect 19656 47900 19720 47904
rect 19656 47844 19660 47900
rect 19660 47844 19716 47900
rect 19716 47844 19720 47900
rect 19656 47840 19720 47844
rect 19736 47900 19800 47904
rect 19736 47844 19740 47900
rect 19740 47844 19796 47900
rect 19796 47844 19800 47900
rect 19736 47840 19800 47844
rect 19816 47900 19880 47904
rect 19816 47844 19820 47900
rect 19820 47844 19876 47900
rect 19876 47844 19880 47900
rect 19816 47840 19880 47844
rect 50296 47900 50360 47904
rect 50296 47844 50300 47900
rect 50300 47844 50356 47900
rect 50356 47844 50360 47900
rect 50296 47840 50360 47844
rect 50376 47900 50440 47904
rect 50376 47844 50380 47900
rect 50380 47844 50436 47900
rect 50436 47844 50440 47900
rect 50376 47840 50440 47844
rect 50456 47900 50520 47904
rect 50456 47844 50460 47900
rect 50460 47844 50516 47900
rect 50516 47844 50520 47900
rect 50456 47840 50520 47844
rect 50536 47900 50600 47904
rect 50536 47844 50540 47900
rect 50540 47844 50596 47900
rect 50596 47844 50600 47900
rect 50536 47840 50600 47844
rect 4216 47356 4280 47360
rect 4216 47300 4220 47356
rect 4220 47300 4276 47356
rect 4276 47300 4280 47356
rect 4216 47296 4280 47300
rect 4296 47356 4360 47360
rect 4296 47300 4300 47356
rect 4300 47300 4356 47356
rect 4356 47300 4360 47356
rect 4296 47296 4360 47300
rect 4376 47356 4440 47360
rect 4376 47300 4380 47356
rect 4380 47300 4436 47356
rect 4436 47300 4440 47356
rect 4376 47296 4440 47300
rect 4456 47356 4520 47360
rect 4456 47300 4460 47356
rect 4460 47300 4516 47356
rect 4516 47300 4520 47356
rect 4456 47296 4520 47300
rect 34936 47356 35000 47360
rect 34936 47300 34940 47356
rect 34940 47300 34996 47356
rect 34996 47300 35000 47356
rect 34936 47296 35000 47300
rect 35016 47356 35080 47360
rect 35016 47300 35020 47356
rect 35020 47300 35076 47356
rect 35076 47300 35080 47356
rect 35016 47296 35080 47300
rect 35096 47356 35160 47360
rect 35096 47300 35100 47356
rect 35100 47300 35156 47356
rect 35156 47300 35160 47356
rect 35096 47296 35160 47300
rect 35176 47356 35240 47360
rect 35176 47300 35180 47356
rect 35180 47300 35236 47356
rect 35236 47300 35240 47356
rect 35176 47296 35240 47300
rect 65656 47356 65720 47360
rect 65656 47300 65660 47356
rect 65660 47300 65716 47356
rect 65716 47300 65720 47356
rect 65656 47296 65720 47300
rect 65736 47356 65800 47360
rect 65736 47300 65740 47356
rect 65740 47300 65796 47356
rect 65796 47300 65800 47356
rect 65736 47296 65800 47300
rect 65816 47356 65880 47360
rect 65816 47300 65820 47356
rect 65820 47300 65876 47356
rect 65876 47300 65880 47356
rect 65816 47296 65880 47300
rect 65896 47356 65960 47360
rect 65896 47300 65900 47356
rect 65900 47300 65956 47356
rect 65956 47300 65960 47356
rect 65896 47296 65960 47300
rect 19576 46812 19640 46816
rect 19576 46756 19580 46812
rect 19580 46756 19636 46812
rect 19636 46756 19640 46812
rect 19576 46752 19640 46756
rect 19656 46812 19720 46816
rect 19656 46756 19660 46812
rect 19660 46756 19716 46812
rect 19716 46756 19720 46812
rect 19656 46752 19720 46756
rect 19736 46812 19800 46816
rect 19736 46756 19740 46812
rect 19740 46756 19796 46812
rect 19796 46756 19800 46812
rect 19736 46752 19800 46756
rect 19816 46812 19880 46816
rect 19816 46756 19820 46812
rect 19820 46756 19876 46812
rect 19876 46756 19880 46812
rect 19816 46752 19880 46756
rect 50296 46812 50360 46816
rect 50296 46756 50300 46812
rect 50300 46756 50356 46812
rect 50356 46756 50360 46812
rect 50296 46752 50360 46756
rect 50376 46812 50440 46816
rect 50376 46756 50380 46812
rect 50380 46756 50436 46812
rect 50436 46756 50440 46812
rect 50376 46752 50440 46756
rect 50456 46812 50520 46816
rect 50456 46756 50460 46812
rect 50460 46756 50516 46812
rect 50516 46756 50520 46812
rect 50456 46752 50520 46756
rect 50536 46812 50600 46816
rect 50536 46756 50540 46812
rect 50540 46756 50596 46812
rect 50596 46756 50600 46812
rect 50536 46752 50600 46756
rect 4216 46268 4280 46272
rect 4216 46212 4220 46268
rect 4220 46212 4276 46268
rect 4276 46212 4280 46268
rect 4216 46208 4280 46212
rect 4296 46268 4360 46272
rect 4296 46212 4300 46268
rect 4300 46212 4356 46268
rect 4356 46212 4360 46268
rect 4296 46208 4360 46212
rect 4376 46268 4440 46272
rect 4376 46212 4380 46268
rect 4380 46212 4436 46268
rect 4436 46212 4440 46268
rect 4376 46208 4440 46212
rect 4456 46268 4520 46272
rect 4456 46212 4460 46268
rect 4460 46212 4516 46268
rect 4516 46212 4520 46268
rect 4456 46208 4520 46212
rect 34936 46268 35000 46272
rect 34936 46212 34940 46268
rect 34940 46212 34996 46268
rect 34996 46212 35000 46268
rect 34936 46208 35000 46212
rect 35016 46268 35080 46272
rect 35016 46212 35020 46268
rect 35020 46212 35076 46268
rect 35076 46212 35080 46268
rect 35016 46208 35080 46212
rect 35096 46268 35160 46272
rect 35096 46212 35100 46268
rect 35100 46212 35156 46268
rect 35156 46212 35160 46268
rect 35096 46208 35160 46212
rect 35176 46268 35240 46272
rect 35176 46212 35180 46268
rect 35180 46212 35236 46268
rect 35236 46212 35240 46268
rect 35176 46208 35240 46212
rect 65656 46268 65720 46272
rect 65656 46212 65660 46268
rect 65660 46212 65716 46268
rect 65716 46212 65720 46268
rect 65656 46208 65720 46212
rect 65736 46268 65800 46272
rect 65736 46212 65740 46268
rect 65740 46212 65796 46268
rect 65796 46212 65800 46268
rect 65736 46208 65800 46212
rect 65816 46268 65880 46272
rect 65816 46212 65820 46268
rect 65820 46212 65876 46268
rect 65876 46212 65880 46268
rect 65816 46208 65880 46212
rect 65896 46268 65960 46272
rect 65896 46212 65900 46268
rect 65900 46212 65956 46268
rect 65956 46212 65960 46268
rect 65896 46208 65960 46212
rect 19576 45724 19640 45728
rect 19576 45668 19580 45724
rect 19580 45668 19636 45724
rect 19636 45668 19640 45724
rect 19576 45664 19640 45668
rect 19656 45724 19720 45728
rect 19656 45668 19660 45724
rect 19660 45668 19716 45724
rect 19716 45668 19720 45724
rect 19656 45664 19720 45668
rect 19736 45724 19800 45728
rect 19736 45668 19740 45724
rect 19740 45668 19796 45724
rect 19796 45668 19800 45724
rect 19736 45664 19800 45668
rect 19816 45724 19880 45728
rect 19816 45668 19820 45724
rect 19820 45668 19876 45724
rect 19876 45668 19880 45724
rect 19816 45664 19880 45668
rect 50296 45724 50360 45728
rect 50296 45668 50300 45724
rect 50300 45668 50356 45724
rect 50356 45668 50360 45724
rect 50296 45664 50360 45668
rect 50376 45724 50440 45728
rect 50376 45668 50380 45724
rect 50380 45668 50436 45724
rect 50436 45668 50440 45724
rect 50376 45664 50440 45668
rect 50456 45724 50520 45728
rect 50456 45668 50460 45724
rect 50460 45668 50516 45724
rect 50516 45668 50520 45724
rect 50456 45664 50520 45668
rect 50536 45724 50600 45728
rect 50536 45668 50540 45724
rect 50540 45668 50596 45724
rect 50596 45668 50600 45724
rect 50536 45664 50600 45668
rect 4216 45180 4280 45184
rect 4216 45124 4220 45180
rect 4220 45124 4276 45180
rect 4276 45124 4280 45180
rect 4216 45120 4280 45124
rect 4296 45180 4360 45184
rect 4296 45124 4300 45180
rect 4300 45124 4356 45180
rect 4356 45124 4360 45180
rect 4296 45120 4360 45124
rect 4376 45180 4440 45184
rect 4376 45124 4380 45180
rect 4380 45124 4436 45180
rect 4436 45124 4440 45180
rect 4376 45120 4440 45124
rect 4456 45180 4520 45184
rect 4456 45124 4460 45180
rect 4460 45124 4516 45180
rect 4516 45124 4520 45180
rect 4456 45120 4520 45124
rect 34936 45180 35000 45184
rect 34936 45124 34940 45180
rect 34940 45124 34996 45180
rect 34996 45124 35000 45180
rect 34936 45120 35000 45124
rect 35016 45180 35080 45184
rect 35016 45124 35020 45180
rect 35020 45124 35076 45180
rect 35076 45124 35080 45180
rect 35016 45120 35080 45124
rect 35096 45180 35160 45184
rect 35096 45124 35100 45180
rect 35100 45124 35156 45180
rect 35156 45124 35160 45180
rect 35096 45120 35160 45124
rect 35176 45180 35240 45184
rect 35176 45124 35180 45180
rect 35180 45124 35236 45180
rect 35236 45124 35240 45180
rect 35176 45120 35240 45124
rect 65656 45180 65720 45184
rect 65656 45124 65660 45180
rect 65660 45124 65716 45180
rect 65716 45124 65720 45180
rect 65656 45120 65720 45124
rect 65736 45180 65800 45184
rect 65736 45124 65740 45180
rect 65740 45124 65796 45180
rect 65796 45124 65800 45180
rect 65736 45120 65800 45124
rect 65816 45180 65880 45184
rect 65816 45124 65820 45180
rect 65820 45124 65876 45180
rect 65876 45124 65880 45180
rect 65816 45120 65880 45124
rect 65896 45180 65960 45184
rect 65896 45124 65900 45180
rect 65900 45124 65956 45180
rect 65956 45124 65960 45180
rect 65896 45120 65960 45124
rect 19576 44636 19640 44640
rect 19576 44580 19580 44636
rect 19580 44580 19636 44636
rect 19636 44580 19640 44636
rect 19576 44576 19640 44580
rect 19656 44636 19720 44640
rect 19656 44580 19660 44636
rect 19660 44580 19716 44636
rect 19716 44580 19720 44636
rect 19656 44576 19720 44580
rect 19736 44636 19800 44640
rect 19736 44580 19740 44636
rect 19740 44580 19796 44636
rect 19796 44580 19800 44636
rect 19736 44576 19800 44580
rect 19816 44636 19880 44640
rect 19816 44580 19820 44636
rect 19820 44580 19876 44636
rect 19876 44580 19880 44636
rect 19816 44576 19880 44580
rect 50296 44636 50360 44640
rect 50296 44580 50300 44636
rect 50300 44580 50356 44636
rect 50356 44580 50360 44636
rect 50296 44576 50360 44580
rect 50376 44636 50440 44640
rect 50376 44580 50380 44636
rect 50380 44580 50436 44636
rect 50436 44580 50440 44636
rect 50376 44576 50440 44580
rect 50456 44636 50520 44640
rect 50456 44580 50460 44636
rect 50460 44580 50516 44636
rect 50516 44580 50520 44636
rect 50456 44576 50520 44580
rect 50536 44636 50600 44640
rect 50536 44580 50540 44636
rect 50540 44580 50596 44636
rect 50596 44580 50600 44636
rect 50536 44576 50600 44580
rect 4216 44092 4280 44096
rect 4216 44036 4220 44092
rect 4220 44036 4276 44092
rect 4276 44036 4280 44092
rect 4216 44032 4280 44036
rect 4296 44092 4360 44096
rect 4296 44036 4300 44092
rect 4300 44036 4356 44092
rect 4356 44036 4360 44092
rect 4296 44032 4360 44036
rect 4376 44092 4440 44096
rect 4376 44036 4380 44092
rect 4380 44036 4436 44092
rect 4436 44036 4440 44092
rect 4376 44032 4440 44036
rect 4456 44092 4520 44096
rect 4456 44036 4460 44092
rect 4460 44036 4516 44092
rect 4516 44036 4520 44092
rect 4456 44032 4520 44036
rect 34936 44092 35000 44096
rect 34936 44036 34940 44092
rect 34940 44036 34996 44092
rect 34996 44036 35000 44092
rect 34936 44032 35000 44036
rect 35016 44092 35080 44096
rect 35016 44036 35020 44092
rect 35020 44036 35076 44092
rect 35076 44036 35080 44092
rect 35016 44032 35080 44036
rect 35096 44092 35160 44096
rect 35096 44036 35100 44092
rect 35100 44036 35156 44092
rect 35156 44036 35160 44092
rect 35096 44032 35160 44036
rect 35176 44092 35240 44096
rect 35176 44036 35180 44092
rect 35180 44036 35236 44092
rect 35236 44036 35240 44092
rect 35176 44032 35240 44036
rect 65656 44092 65720 44096
rect 65656 44036 65660 44092
rect 65660 44036 65716 44092
rect 65716 44036 65720 44092
rect 65656 44032 65720 44036
rect 65736 44092 65800 44096
rect 65736 44036 65740 44092
rect 65740 44036 65796 44092
rect 65796 44036 65800 44092
rect 65736 44032 65800 44036
rect 65816 44092 65880 44096
rect 65816 44036 65820 44092
rect 65820 44036 65876 44092
rect 65876 44036 65880 44092
rect 65816 44032 65880 44036
rect 65896 44092 65960 44096
rect 65896 44036 65900 44092
rect 65900 44036 65956 44092
rect 65956 44036 65960 44092
rect 65896 44032 65960 44036
rect 19576 43548 19640 43552
rect 19576 43492 19580 43548
rect 19580 43492 19636 43548
rect 19636 43492 19640 43548
rect 19576 43488 19640 43492
rect 19656 43548 19720 43552
rect 19656 43492 19660 43548
rect 19660 43492 19716 43548
rect 19716 43492 19720 43548
rect 19656 43488 19720 43492
rect 19736 43548 19800 43552
rect 19736 43492 19740 43548
rect 19740 43492 19796 43548
rect 19796 43492 19800 43548
rect 19736 43488 19800 43492
rect 19816 43548 19880 43552
rect 19816 43492 19820 43548
rect 19820 43492 19876 43548
rect 19876 43492 19880 43548
rect 19816 43488 19880 43492
rect 50296 43548 50360 43552
rect 50296 43492 50300 43548
rect 50300 43492 50356 43548
rect 50356 43492 50360 43548
rect 50296 43488 50360 43492
rect 50376 43548 50440 43552
rect 50376 43492 50380 43548
rect 50380 43492 50436 43548
rect 50436 43492 50440 43548
rect 50376 43488 50440 43492
rect 50456 43548 50520 43552
rect 50456 43492 50460 43548
rect 50460 43492 50516 43548
rect 50516 43492 50520 43548
rect 50456 43488 50520 43492
rect 50536 43548 50600 43552
rect 50536 43492 50540 43548
rect 50540 43492 50596 43548
rect 50596 43492 50600 43548
rect 50536 43488 50600 43492
rect 4216 43004 4280 43008
rect 4216 42948 4220 43004
rect 4220 42948 4276 43004
rect 4276 42948 4280 43004
rect 4216 42944 4280 42948
rect 4296 43004 4360 43008
rect 4296 42948 4300 43004
rect 4300 42948 4356 43004
rect 4356 42948 4360 43004
rect 4296 42944 4360 42948
rect 4376 43004 4440 43008
rect 4376 42948 4380 43004
rect 4380 42948 4436 43004
rect 4436 42948 4440 43004
rect 4376 42944 4440 42948
rect 4456 43004 4520 43008
rect 4456 42948 4460 43004
rect 4460 42948 4516 43004
rect 4516 42948 4520 43004
rect 4456 42944 4520 42948
rect 34936 43004 35000 43008
rect 34936 42948 34940 43004
rect 34940 42948 34996 43004
rect 34996 42948 35000 43004
rect 34936 42944 35000 42948
rect 35016 43004 35080 43008
rect 35016 42948 35020 43004
rect 35020 42948 35076 43004
rect 35076 42948 35080 43004
rect 35016 42944 35080 42948
rect 35096 43004 35160 43008
rect 35096 42948 35100 43004
rect 35100 42948 35156 43004
rect 35156 42948 35160 43004
rect 35096 42944 35160 42948
rect 35176 43004 35240 43008
rect 35176 42948 35180 43004
rect 35180 42948 35236 43004
rect 35236 42948 35240 43004
rect 35176 42944 35240 42948
rect 65656 43004 65720 43008
rect 65656 42948 65660 43004
rect 65660 42948 65716 43004
rect 65716 42948 65720 43004
rect 65656 42944 65720 42948
rect 65736 43004 65800 43008
rect 65736 42948 65740 43004
rect 65740 42948 65796 43004
rect 65796 42948 65800 43004
rect 65736 42944 65800 42948
rect 65816 43004 65880 43008
rect 65816 42948 65820 43004
rect 65820 42948 65876 43004
rect 65876 42948 65880 43004
rect 65816 42944 65880 42948
rect 65896 43004 65960 43008
rect 65896 42948 65900 43004
rect 65900 42948 65956 43004
rect 65956 42948 65960 43004
rect 65896 42944 65960 42948
rect 19576 42460 19640 42464
rect 19576 42404 19580 42460
rect 19580 42404 19636 42460
rect 19636 42404 19640 42460
rect 19576 42400 19640 42404
rect 19656 42460 19720 42464
rect 19656 42404 19660 42460
rect 19660 42404 19716 42460
rect 19716 42404 19720 42460
rect 19656 42400 19720 42404
rect 19736 42460 19800 42464
rect 19736 42404 19740 42460
rect 19740 42404 19796 42460
rect 19796 42404 19800 42460
rect 19736 42400 19800 42404
rect 19816 42460 19880 42464
rect 19816 42404 19820 42460
rect 19820 42404 19876 42460
rect 19876 42404 19880 42460
rect 19816 42400 19880 42404
rect 50296 42460 50360 42464
rect 50296 42404 50300 42460
rect 50300 42404 50356 42460
rect 50356 42404 50360 42460
rect 50296 42400 50360 42404
rect 50376 42460 50440 42464
rect 50376 42404 50380 42460
rect 50380 42404 50436 42460
rect 50436 42404 50440 42460
rect 50376 42400 50440 42404
rect 50456 42460 50520 42464
rect 50456 42404 50460 42460
rect 50460 42404 50516 42460
rect 50516 42404 50520 42460
rect 50456 42400 50520 42404
rect 50536 42460 50600 42464
rect 50536 42404 50540 42460
rect 50540 42404 50596 42460
rect 50596 42404 50600 42460
rect 50536 42400 50600 42404
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 34936 41916 35000 41920
rect 34936 41860 34940 41916
rect 34940 41860 34996 41916
rect 34996 41860 35000 41916
rect 34936 41856 35000 41860
rect 35016 41916 35080 41920
rect 35016 41860 35020 41916
rect 35020 41860 35076 41916
rect 35076 41860 35080 41916
rect 35016 41856 35080 41860
rect 35096 41916 35160 41920
rect 35096 41860 35100 41916
rect 35100 41860 35156 41916
rect 35156 41860 35160 41916
rect 35096 41856 35160 41860
rect 35176 41916 35240 41920
rect 35176 41860 35180 41916
rect 35180 41860 35236 41916
rect 35236 41860 35240 41916
rect 35176 41856 35240 41860
rect 65656 41916 65720 41920
rect 65656 41860 65660 41916
rect 65660 41860 65716 41916
rect 65716 41860 65720 41916
rect 65656 41856 65720 41860
rect 65736 41916 65800 41920
rect 65736 41860 65740 41916
rect 65740 41860 65796 41916
rect 65796 41860 65800 41916
rect 65736 41856 65800 41860
rect 65816 41916 65880 41920
rect 65816 41860 65820 41916
rect 65820 41860 65876 41916
rect 65876 41860 65880 41916
rect 65816 41856 65880 41860
rect 65896 41916 65960 41920
rect 65896 41860 65900 41916
rect 65900 41860 65956 41916
rect 65956 41860 65960 41916
rect 65896 41856 65960 41860
rect 19576 41372 19640 41376
rect 19576 41316 19580 41372
rect 19580 41316 19636 41372
rect 19636 41316 19640 41372
rect 19576 41312 19640 41316
rect 19656 41372 19720 41376
rect 19656 41316 19660 41372
rect 19660 41316 19716 41372
rect 19716 41316 19720 41372
rect 19656 41312 19720 41316
rect 19736 41372 19800 41376
rect 19736 41316 19740 41372
rect 19740 41316 19796 41372
rect 19796 41316 19800 41372
rect 19736 41312 19800 41316
rect 19816 41372 19880 41376
rect 19816 41316 19820 41372
rect 19820 41316 19876 41372
rect 19876 41316 19880 41372
rect 19816 41312 19880 41316
rect 50296 41372 50360 41376
rect 50296 41316 50300 41372
rect 50300 41316 50356 41372
rect 50356 41316 50360 41372
rect 50296 41312 50360 41316
rect 50376 41372 50440 41376
rect 50376 41316 50380 41372
rect 50380 41316 50436 41372
rect 50436 41316 50440 41372
rect 50376 41312 50440 41316
rect 50456 41372 50520 41376
rect 50456 41316 50460 41372
rect 50460 41316 50516 41372
rect 50516 41316 50520 41372
rect 50456 41312 50520 41316
rect 50536 41372 50600 41376
rect 50536 41316 50540 41372
rect 50540 41316 50596 41372
rect 50596 41316 50600 41372
rect 50536 41312 50600 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 34936 40828 35000 40832
rect 34936 40772 34940 40828
rect 34940 40772 34996 40828
rect 34996 40772 35000 40828
rect 34936 40768 35000 40772
rect 35016 40828 35080 40832
rect 35016 40772 35020 40828
rect 35020 40772 35076 40828
rect 35076 40772 35080 40828
rect 35016 40768 35080 40772
rect 35096 40828 35160 40832
rect 35096 40772 35100 40828
rect 35100 40772 35156 40828
rect 35156 40772 35160 40828
rect 35096 40768 35160 40772
rect 35176 40828 35240 40832
rect 35176 40772 35180 40828
rect 35180 40772 35236 40828
rect 35236 40772 35240 40828
rect 35176 40768 35240 40772
rect 65656 40828 65720 40832
rect 65656 40772 65660 40828
rect 65660 40772 65716 40828
rect 65716 40772 65720 40828
rect 65656 40768 65720 40772
rect 65736 40828 65800 40832
rect 65736 40772 65740 40828
rect 65740 40772 65796 40828
rect 65796 40772 65800 40828
rect 65736 40768 65800 40772
rect 65816 40828 65880 40832
rect 65816 40772 65820 40828
rect 65820 40772 65876 40828
rect 65876 40772 65880 40828
rect 65816 40768 65880 40772
rect 65896 40828 65960 40832
rect 65896 40772 65900 40828
rect 65900 40772 65956 40828
rect 65956 40772 65960 40828
rect 65896 40768 65960 40772
rect 19576 40284 19640 40288
rect 19576 40228 19580 40284
rect 19580 40228 19636 40284
rect 19636 40228 19640 40284
rect 19576 40224 19640 40228
rect 19656 40284 19720 40288
rect 19656 40228 19660 40284
rect 19660 40228 19716 40284
rect 19716 40228 19720 40284
rect 19656 40224 19720 40228
rect 19736 40284 19800 40288
rect 19736 40228 19740 40284
rect 19740 40228 19796 40284
rect 19796 40228 19800 40284
rect 19736 40224 19800 40228
rect 19816 40284 19880 40288
rect 19816 40228 19820 40284
rect 19820 40228 19876 40284
rect 19876 40228 19880 40284
rect 19816 40224 19880 40228
rect 50296 40284 50360 40288
rect 50296 40228 50300 40284
rect 50300 40228 50356 40284
rect 50356 40228 50360 40284
rect 50296 40224 50360 40228
rect 50376 40284 50440 40288
rect 50376 40228 50380 40284
rect 50380 40228 50436 40284
rect 50436 40228 50440 40284
rect 50376 40224 50440 40228
rect 50456 40284 50520 40288
rect 50456 40228 50460 40284
rect 50460 40228 50516 40284
rect 50516 40228 50520 40284
rect 50456 40224 50520 40228
rect 50536 40284 50600 40288
rect 50536 40228 50540 40284
rect 50540 40228 50596 40284
rect 50596 40228 50600 40284
rect 50536 40224 50600 40228
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 65656 39740 65720 39744
rect 65656 39684 65660 39740
rect 65660 39684 65716 39740
rect 65716 39684 65720 39740
rect 65656 39680 65720 39684
rect 65736 39740 65800 39744
rect 65736 39684 65740 39740
rect 65740 39684 65796 39740
rect 65796 39684 65800 39740
rect 65736 39680 65800 39684
rect 65816 39740 65880 39744
rect 65816 39684 65820 39740
rect 65820 39684 65876 39740
rect 65876 39684 65880 39740
rect 65816 39680 65880 39684
rect 65896 39740 65960 39744
rect 65896 39684 65900 39740
rect 65900 39684 65956 39740
rect 65956 39684 65960 39740
rect 65896 39680 65960 39684
rect 19576 39196 19640 39200
rect 19576 39140 19580 39196
rect 19580 39140 19636 39196
rect 19636 39140 19640 39196
rect 19576 39136 19640 39140
rect 19656 39196 19720 39200
rect 19656 39140 19660 39196
rect 19660 39140 19716 39196
rect 19716 39140 19720 39196
rect 19656 39136 19720 39140
rect 19736 39196 19800 39200
rect 19736 39140 19740 39196
rect 19740 39140 19796 39196
rect 19796 39140 19800 39196
rect 19736 39136 19800 39140
rect 19816 39196 19880 39200
rect 19816 39140 19820 39196
rect 19820 39140 19876 39196
rect 19876 39140 19880 39196
rect 19816 39136 19880 39140
rect 50296 39196 50360 39200
rect 50296 39140 50300 39196
rect 50300 39140 50356 39196
rect 50356 39140 50360 39196
rect 50296 39136 50360 39140
rect 50376 39196 50440 39200
rect 50376 39140 50380 39196
rect 50380 39140 50436 39196
rect 50436 39140 50440 39196
rect 50376 39136 50440 39140
rect 50456 39196 50520 39200
rect 50456 39140 50460 39196
rect 50460 39140 50516 39196
rect 50516 39140 50520 39196
rect 50456 39136 50520 39140
rect 50536 39196 50600 39200
rect 50536 39140 50540 39196
rect 50540 39140 50596 39196
rect 50596 39140 50600 39196
rect 50536 39136 50600 39140
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 65656 38652 65720 38656
rect 65656 38596 65660 38652
rect 65660 38596 65716 38652
rect 65716 38596 65720 38652
rect 65656 38592 65720 38596
rect 65736 38652 65800 38656
rect 65736 38596 65740 38652
rect 65740 38596 65796 38652
rect 65796 38596 65800 38652
rect 65736 38592 65800 38596
rect 65816 38652 65880 38656
rect 65816 38596 65820 38652
rect 65820 38596 65876 38652
rect 65876 38596 65880 38652
rect 65816 38592 65880 38596
rect 65896 38652 65960 38656
rect 65896 38596 65900 38652
rect 65900 38596 65956 38652
rect 65956 38596 65960 38652
rect 65896 38592 65960 38596
rect 19576 38108 19640 38112
rect 19576 38052 19580 38108
rect 19580 38052 19636 38108
rect 19636 38052 19640 38108
rect 19576 38048 19640 38052
rect 19656 38108 19720 38112
rect 19656 38052 19660 38108
rect 19660 38052 19716 38108
rect 19716 38052 19720 38108
rect 19656 38048 19720 38052
rect 19736 38108 19800 38112
rect 19736 38052 19740 38108
rect 19740 38052 19796 38108
rect 19796 38052 19800 38108
rect 19736 38048 19800 38052
rect 19816 38108 19880 38112
rect 19816 38052 19820 38108
rect 19820 38052 19876 38108
rect 19876 38052 19880 38108
rect 19816 38048 19880 38052
rect 50296 38108 50360 38112
rect 50296 38052 50300 38108
rect 50300 38052 50356 38108
rect 50356 38052 50360 38108
rect 50296 38048 50360 38052
rect 50376 38108 50440 38112
rect 50376 38052 50380 38108
rect 50380 38052 50436 38108
rect 50436 38052 50440 38108
rect 50376 38048 50440 38052
rect 50456 38108 50520 38112
rect 50456 38052 50460 38108
rect 50460 38052 50516 38108
rect 50516 38052 50520 38108
rect 50456 38048 50520 38052
rect 50536 38108 50600 38112
rect 50536 38052 50540 38108
rect 50540 38052 50596 38108
rect 50596 38052 50600 38108
rect 50536 38048 50600 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 65656 37564 65720 37568
rect 65656 37508 65660 37564
rect 65660 37508 65716 37564
rect 65716 37508 65720 37564
rect 65656 37504 65720 37508
rect 65736 37564 65800 37568
rect 65736 37508 65740 37564
rect 65740 37508 65796 37564
rect 65796 37508 65800 37564
rect 65736 37504 65800 37508
rect 65816 37564 65880 37568
rect 65816 37508 65820 37564
rect 65820 37508 65876 37564
rect 65876 37508 65880 37564
rect 65816 37504 65880 37508
rect 65896 37564 65960 37568
rect 65896 37508 65900 37564
rect 65900 37508 65956 37564
rect 65956 37508 65960 37564
rect 65896 37504 65960 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 50296 37020 50360 37024
rect 50296 36964 50300 37020
rect 50300 36964 50356 37020
rect 50356 36964 50360 37020
rect 50296 36960 50360 36964
rect 50376 37020 50440 37024
rect 50376 36964 50380 37020
rect 50380 36964 50436 37020
rect 50436 36964 50440 37020
rect 50376 36960 50440 36964
rect 50456 37020 50520 37024
rect 50456 36964 50460 37020
rect 50460 36964 50516 37020
rect 50516 36964 50520 37020
rect 50456 36960 50520 36964
rect 50536 37020 50600 37024
rect 50536 36964 50540 37020
rect 50540 36964 50596 37020
rect 50596 36964 50600 37020
rect 50536 36960 50600 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 65656 36476 65720 36480
rect 65656 36420 65660 36476
rect 65660 36420 65716 36476
rect 65716 36420 65720 36476
rect 65656 36416 65720 36420
rect 65736 36476 65800 36480
rect 65736 36420 65740 36476
rect 65740 36420 65796 36476
rect 65796 36420 65800 36476
rect 65736 36416 65800 36420
rect 65816 36476 65880 36480
rect 65816 36420 65820 36476
rect 65820 36420 65876 36476
rect 65876 36420 65880 36476
rect 65816 36416 65880 36420
rect 65896 36476 65960 36480
rect 65896 36420 65900 36476
rect 65900 36420 65956 36476
rect 65956 36420 65960 36476
rect 65896 36416 65960 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 50296 35932 50360 35936
rect 50296 35876 50300 35932
rect 50300 35876 50356 35932
rect 50356 35876 50360 35932
rect 50296 35872 50360 35876
rect 50376 35932 50440 35936
rect 50376 35876 50380 35932
rect 50380 35876 50436 35932
rect 50436 35876 50440 35932
rect 50376 35872 50440 35876
rect 50456 35932 50520 35936
rect 50456 35876 50460 35932
rect 50460 35876 50516 35932
rect 50516 35876 50520 35932
rect 50456 35872 50520 35876
rect 50536 35932 50600 35936
rect 50536 35876 50540 35932
rect 50540 35876 50596 35932
rect 50596 35876 50600 35932
rect 50536 35872 50600 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 65656 35388 65720 35392
rect 65656 35332 65660 35388
rect 65660 35332 65716 35388
rect 65716 35332 65720 35388
rect 65656 35328 65720 35332
rect 65736 35388 65800 35392
rect 65736 35332 65740 35388
rect 65740 35332 65796 35388
rect 65796 35332 65800 35388
rect 65736 35328 65800 35332
rect 65816 35388 65880 35392
rect 65816 35332 65820 35388
rect 65820 35332 65876 35388
rect 65876 35332 65880 35388
rect 65816 35328 65880 35332
rect 65896 35388 65960 35392
rect 65896 35332 65900 35388
rect 65900 35332 65956 35388
rect 65956 35332 65960 35388
rect 65896 35328 65960 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 50296 34844 50360 34848
rect 50296 34788 50300 34844
rect 50300 34788 50356 34844
rect 50356 34788 50360 34844
rect 50296 34784 50360 34788
rect 50376 34844 50440 34848
rect 50376 34788 50380 34844
rect 50380 34788 50436 34844
rect 50436 34788 50440 34844
rect 50376 34784 50440 34788
rect 50456 34844 50520 34848
rect 50456 34788 50460 34844
rect 50460 34788 50516 34844
rect 50516 34788 50520 34844
rect 50456 34784 50520 34788
rect 50536 34844 50600 34848
rect 50536 34788 50540 34844
rect 50540 34788 50596 34844
rect 50596 34788 50600 34844
rect 50536 34784 50600 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 65656 34300 65720 34304
rect 65656 34244 65660 34300
rect 65660 34244 65716 34300
rect 65716 34244 65720 34300
rect 65656 34240 65720 34244
rect 65736 34300 65800 34304
rect 65736 34244 65740 34300
rect 65740 34244 65796 34300
rect 65796 34244 65800 34300
rect 65736 34240 65800 34244
rect 65816 34300 65880 34304
rect 65816 34244 65820 34300
rect 65820 34244 65876 34300
rect 65876 34244 65880 34300
rect 65816 34240 65880 34244
rect 65896 34300 65960 34304
rect 65896 34244 65900 34300
rect 65900 34244 65956 34300
rect 65956 34244 65960 34300
rect 65896 34240 65960 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 50296 33756 50360 33760
rect 50296 33700 50300 33756
rect 50300 33700 50356 33756
rect 50356 33700 50360 33756
rect 50296 33696 50360 33700
rect 50376 33756 50440 33760
rect 50376 33700 50380 33756
rect 50380 33700 50436 33756
rect 50436 33700 50440 33756
rect 50376 33696 50440 33700
rect 50456 33756 50520 33760
rect 50456 33700 50460 33756
rect 50460 33700 50516 33756
rect 50516 33700 50520 33756
rect 50456 33696 50520 33700
rect 50536 33756 50600 33760
rect 50536 33700 50540 33756
rect 50540 33700 50596 33756
rect 50596 33700 50600 33756
rect 50536 33696 50600 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 65656 33212 65720 33216
rect 65656 33156 65660 33212
rect 65660 33156 65716 33212
rect 65716 33156 65720 33212
rect 65656 33152 65720 33156
rect 65736 33212 65800 33216
rect 65736 33156 65740 33212
rect 65740 33156 65796 33212
rect 65796 33156 65800 33212
rect 65736 33152 65800 33156
rect 65816 33212 65880 33216
rect 65816 33156 65820 33212
rect 65820 33156 65876 33212
rect 65876 33156 65880 33212
rect 65816 33152 65880 33156
rect 65896 33212 65960 33216
rect 65896 33156 65900 33212
rect 65900 33156 65956 33212
rect 65956 33156 65960 33212
rect 65896 33152 65960 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 50296 32668 50360 32672
rect 50296 32612 50300 32668
rect 50300 32612 50356 32668
rect 50356 32612 50360 32668
rect 50296 32608 50360 32612
rect 50376 32668 50440 32672
rect 50376 32612 50380 32668
rect 50380 32612 50436 32668
rect 50436 32612 50440 32668
rect 50376 32608 50440 32612
rect 50456 32668 50520 32672
rect 50456 32612 50460 32668
rect 50460 32612 50516 32668
rect 50516 32612 50520 32668
rect 50456 32608 50520 32612
rect 50536 32668 50600 32672
rect 50536 32612 50540 32668
rect 50540 32612 50596 32668
rect 50596 32612 50600 32668
rect 50536 32608 50600 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 65656 32124 65720 32128
rect 65656 32068 65660 32124
rect 65660 32068 65716 32124
rect 65716 32068 65720 32124
rect 65656 32064 65720 32068
rect 65736 32124 65800 32128
rect 65736 32068 65740 32124
rect 65740 32068 65796 32124
rect 65796 32068 65800 32124
rect 65736 32064 65800 32068
rect 65816 32124 65880 32128
rect 65816 32068 65820 32124
rect 65820 32068 65876 32124
rect 65876 32068 65880 32124
rect 65816 32064 65880 32068
rect 65896 32124 65960 32128
rect 65896 32068 65900 32124
rect 65900 32068 65956 32124
rect 65956 32068 65960 32124
rect 65896 32064 65960 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 50296 31580 50360 31584
rect 50296 31524 50300 31580
rect 50300 31524 50356 31580
rect 50356 31524 50360 31580
rect 50296 31520 50360 31524
rect 50376 31580 50440 31584
rect 50376 31524 50380 31580
rect 50380 31524 50436 31580
rect 50436 31524 50440 31580
rect 50376 31520 50440 31524
rect 50456 31580 50520 31584
rect 50456 31524 50460 31580
rect 50460 31524 50516 31580
rect 50516 31524 50520 31580
rect 50456 31520 50520 31524
rect 50536 31580 50600 31584
rect 50536 31524 50540 31580
rect 50540 31524 50596 31580
rect 50596 31524 50600 31580
rect 50536 31520 50600 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 65656 31036 65720 31040
rect 65656 30980 65660 31036
rect 65660 30980 65716 31036
rect 65716 30980 65720 31036
rect 65656 30976 65720 30980
rect 65736 31036 65800 31040
rect 65736 30980 65740 31036
rect 65740 30980 65796 31036
rect 65796 30980 65800 31036
rect 65736 30976 65800 30980
rect 65816 31036 65880 31040
rect 65816 30980 65820 31036
rect 65820 30980 65876 31036
rect 65876 30980 65880 31036
rect 65816 30976 65880 30980
rect 65896 31036 65960 31040
rect 65896 30980 65900 31036
rect 65900 30980 65956 31036
rect 65956 30980 65960 31036
rect 65896 30976 65960 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 50296 30492 50360 30496
rect 50296 30436 50300 30492
rect 50300 30436 50356 30492
rect 50356 30436 50360 30492
rect 50296 30432 50360 30436
rect 50376 30492 50440 30496
rect 50376 30436 50380 30492
rect 50380 30436 50436 30492
rect 50436 30436 50440 30492
rect 50376 30432 50440 30436
rect 50456 30492 50520 30496
rect 50456 30436 50460 30492
rect 50460 30436 50516 30492
rect 50516 30436 50520 30492
rect 50456 30432 50520 30436
rect 50536 30492 50600 30496
rect 50536 30436 50540 30492
rect 50540 30436 50596 30492
rect 50596 30436 50600 30492
rect 50536 30432 50600 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 65656 29948 65720 29952
rect 65656 29892 65660 29948
rect 65660 29892 65716 29948
rect 65716 29892 65720 29948
rect 65656 29888 65720 29892
rect 65736 29948 65800 29952
rect 65736 29892 65740 29948
rect 65740 29892 65796 29948
rect 65796 29892 65800 29948
rect 65736 29888 65800 29892
rect 65816 29948 65880 29952
rect 65816 29892 65820 29948
rect 65820 29892 65876 29948
rect 65876 29892 65880 29948
rect 65816 29888 65880 29892
rect 65896 29948 65960 29952
rect 65896 29892 65900 29948
rect 65900 29892 65956 29948
rect 65956 29892 65960 29948
rect 65896 29888 65960 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 50296 29404 50360 29408
rect 50296 29348 50300 29404
rect 50300 29348 50356 29404
rect 50356 29348 50360 29404
rect 50296 29344 50360 29348
rect 50376 29404 50440 29408
rect 50376 29348 50380 29404
rect 50380 29348 50436 29404
rect 50436 29348 50440 29404
rect 50376 29344 50440 29348
rect 50456 29404 50520 29408
rect 50456 29348 50460 29404
rect 50460 29348 50516 29404
rect 50516 29348 50520 29404
rect 50456 29344 50520 29348
rect 50536 29404 50600 29408
rect 50536 29348 50540 29404
rect 50540 29348 50596 29404
rect 50596 29348 50600 29404
rect 50536 29344 50600 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 65656 28860 65720 28864
rect 65656 28804 65660 28860
rect 65660 28804 65716 28860
rect 65716 28804 65720 28860
rect 65656 28800 65720 28804
rect 65736 28860 65800 28864
rect 65736 28804 65740 28860
rect 65740 28804 65796 28860
rect 65796 28804 65800 28860
rect 65736 28800 65800 28804
rect 65816 28860 65880 28864
rect 65816 28804 65820 28860
rect 65820 28804 65876 28860
rect 65876 28804 65880 28860
rect 65816 28800 65880 28804
rect 65896 28860 65960 28864
rect 65896 28804 65900 28860
rect 65900 28804 65956 28860
rect 65956 28804 65960 28860
rect 65896 28800 65960 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 50296 28316 50360 28320
rect 50296 28260 50300 28316
rect 50300 28260 50356 28316
rect 50356 28260 50360 28316
rect 50296 28256 50360 28260
rect 50376 28316 50440 28320
rect 50376 28260 50380 28316
rect 50380 28260 50436 28316
rect 50436 28260 50440 28316
rect 50376 28256 50440 28260
rect 50456 28316 50520 28320
rect 50456 28260 50460 28316
rect 50460 28260 50516 28316
rect 50516 28260 50520 28316
rect 50456 28256 50520 28260
rect 50536 28316 50600 28320
rect 50536 28260 50540 28316
rect 50540 28260 50596 28316
rect 50596 28260 50600 28316
rect 50536 28256 50600 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 65656 27772 65720 27776
rect 65656 27716 65660 27772
rect 65660 27716 65716 27772
rect 65716 27716 65720 27772
rect 65656 27712 65720 27716
rect 65736 27772 65800 27776
rect 65736 27716 65740 27772
rect 65740 27716 65796 27772
rect 65796 27716 65800 27772
rect 65736 27712 65800 27716
rect 65816 27772 65880 27776
rect 65816 27716 65820 27772
rect 65820 27716 65876 27772
rect 65876 27716 65880 27772
rect 65816 27712 65880 27716
rect 65896 27772 65960 27776
rect 65896 27716 65900 27772
rect 65900 27716 65956 27772
rect 65956 27716 65960 27772
rect 65896 27712 65960 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 50296 27228 50360 27232
rect 50296 27172 50300 27228
rect 50300 27172 50356 27228
rect 50356 27172 50360 27228
rect 50296 27168 50360 27172
rect 50376 27228 50440 27232
rect 50376 27172 50380 27228
rect 50380 27172 50436 27228
rect 50436 27172 50440 27228
rect 50376 27168 50440 27172
rect 50456 27228 50520 27232
rect 50456 27172 50460 27228
rect 50460 27172 50516 27228
rect 50516 27172 50520 27228
rect 50456 27168 50520 27172
rect 50536 27228 50600 27232
rect 50536 27172 50540 27228
rect 50540 27172 50596 27228
rect 50596 27172 50600 27228
rect 50536 27168 50600 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 65656 26684 65720 26688
rect 65656 26628 65660 26684
rect 65660 26628 65716 26684
rect 65716 26628 65720 26684
rect 65656 26624 65720 26628
rect 65736 26684 65800 26688
rect 65736 26628 65740 26684
rect 65740 26628 65796 26684
rect 65796 26628 65800 26684
rect 65736 26624 65800 26628
rect 65816 26684 65880 26688
rect 65816 26628 65820 26684
rect 65820 26628 65876 26684
rect 65876 26628 65880 26684
rect 65816 26624 65880 26628
rect 65896 26684 65960 26688
rect 65896 26628 65900 26684
rect 65900 26628 65956 26684
rect 65956 26628 65960 26684
rect 65896 26624 65960 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 50296 26140 50360 26144
rect 50296 26084 50300 26140
rect 50300 26084 50356 26140
rect 50356 26084 50360 26140
rect 50296 26080 50360 26084
rect 50376 26140 50440 26144
rect 50376 26084 50380 26140
rect 50380 26084 50436 26140
rect 50436 26084 50440 26140
rect 50376 26080 50440 26084
rect 50456 26140 50520 26144
rect 50456 26084 50460 26140
rect 50460 26084 50516 26140
rect 50516 26084 50520 26140
rect 50456 26080 50520 26084
rect 50536 26140 50600 26144
rect 50536 26084 50540 26140
rect 50540 26084 50596 26140
rect 50596 26084 50600 26140
rect 50536 26080 50600 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 65656 25596 65720 25600
rect 65656 25540 65660 25596
rect 65660 25540 65716 25596
rect 65716 25540 65720 25596
rect 65656 25536 65720 25540
rect 65736 25596 65800 25600
rect 65736 25540 65740 25596
rect 65740 25540 65796 25596
rect 65796 25540 65800 25596
rect 65736 25536 65800 25540
rect 65816 25596 65880 25600
rect 65816 25540 65820 25596
rect 65820 25540 65876 25596
rect 65876 25540 65880 25596
rect 65816 25536 65880 25540
rect 65896 25596 65960 25600
rect 65896 25540 65900 25596
rect 65900 25540 65956 25596
rect 65956 25540 65960 25596
rect 65896 25536 65960 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 50296 25052 50360 25056
rect 50296 24996 50300 25052
rect 50300 24996 50356 25052
rect 50356 24996 50360 25052
rect 50296 24992 50360 24996
rect 50376 25052 50440 25056
rect 50376 24996 50380 25052
rect 50380 24996 50436 25052
rect 50436 24996 50440 25052
rect 50376 24992 50440 24996
rect 50456 25052 50520 25056
rect 50456 24996 50460 25052
rect 50460 24996 50516 25052
rect 50516 24996 50520 25052
rect 50456 24992 50520 24996
rect 50536 25052 50600 25056
rect 50536 24996 50540 25052
rect 50540 24996 50596 25052
rect 50596 24996 50600 25052
rect 50536 24992 50600 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 65656 24508 65720 24512
rect 65656 24452 65660 24508
rect 65660 24452 65716 24508
rect 65716 24452 65720 24508
rect 65656 24448 65720 24452
rect 65736 24508 65800 24512
rect 65736 24452 65740 24508
rect 65740 24452 65796 24508
rect 65796 24452 65800 24508
rect 65736 24448 65800 24452
rect 65816 24508 65880 24512
rect 65816 24452 65820 24508
rect 65820 24452 65876 24508
rect 65876 24452 65880 24508
rect 65816 24448 65880 24452
rect 65896 24508 65960 24512
rect 65896 24452 65900 24508
rect 65900 24452 65956 24508
rect 65956 24452 65960 24508
rect 65896 24448 65960 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 50296 23964 50360 23968
rect 50296 23908 50300 23964
rect 50300 23908 50356 23964
rect 50356 23908 50360 23964
rect 50296 23904 50360 23908
rect 50376 23964 50440 23968
rect 50376 23908 50380 23964
rect 50380 23908 50436 23964
rect 50436 23908 50440 23964
rect 50376 23904 50440 23908
rect 50456 23964 50520 23968
rect 50456 23908 50460 23964
rect 50460 23908 50516 23964
rect 50516 23908 50520 23964
rect 50456 23904 50520 23908
rect 50536 23964 50600 23968
rect 50536 23908 50540 23964
rect 50540 23908 50596 23964
rect 50596 23908 50600 23964
rect 50536 23904 50600 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 65656 23420 65720 23424
rect 65656 23364 65660 23420
rect 65660 23364 65716 23420
rect 65716 23364 65720 23420
rect 65656 23360 65720 23364
rect 65736 23420 65800 23424
rect 65736 23364 65740 23420
rect 65740 23364 65796 23420
rect 65796 23364 65800 23420
rect 65736 23360 65800 23364
rect 65816 23420 65880 23424
rect 65816 23364 65820 23420
rect 65820 23364 65876 23420
rect 65876 23364 65880 23420
rect 65816 23360 65880 23364
rect 65896 23420 65960 23424
rect 65896 23364 65900 23420
rect 65900 23364 65956 23420
rect 65956 23364 65960 23420
rect 65896 23360 65960 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 50296 22876 50360 22880
rect 50296 22820 50300 22876
rect 50300 22820 50356 22876
rect 50356 22820 50360 22876
rect 50296 22816 50360 22820
rect 50376 22876 50440 22880
rect 50376 22820 50380 22876
rect 50380 22820 50436 22876
rect 50436 22820 50440 22876
rect 50376 22816 50440 22820
rect 50456 22876 50520 22880
rect 50456 22820 50460 22876
rect 50460 22820 50516 22876
rect 50516 22820 50520 22876
rect 50456 22816 50520 22820
rect 50536 22876 50600 22880
rect 50536 22820 50540 22876
rect 50540 22820 50596 22876
rect 50596 22820 50600 22876
rect 50536 22816 50600 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 65656 22332 65720 22336
rect 65656 22276 65660 22332
rect 65660 22276 65716 22332
rect 65716 22276 65720 22332
rect 65656 22272 65720 22276
rect 65736 22332 65800 22336
rect 65736 22276 65740 22332
rect 65740 22276 65796 22332
rect 65796 22276 65800 22332
rect 65736 22272 65800 22276
rect 65816 22332 65880 22336
rect 65816 22276 65820 22332
rect 65820 22276 65876 22332
rect 65876 22276 65880 22332
rect 65816 22272 65880 22276
rect 65896 22332 65960 22336
rect 65896 22276 65900 22332
rect 65900 22276 65956 22332
rect 65956 22276 65960 22332
rect 65896 22272 65960 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 50296 21788 50360 21792
rect 50296 21732 50300 21788
rect 50300 21732 50356 21788
rect 50356 21732 50360 21788
rect 50296 21728 50360 21732
rect 50376 21788 50440 21792
rect 50376 21732 50380 21788
rect 50380 21732 50436 21788
rect 50436 21732 50440 21788
rect 50376 21728 50440 21732
rect 50456 21788 50520 21792
rect 50456 21732 50460 21788
rect 50460 21732 50516 21788
rect 50516 21732 50520 21788
rect 50456 21728 50520 21732
rect 50536 21788 50600 21792
rect 50536 21732 50540 21788
rect 50540 21732 50596 21788
rect 50596 21732 50600 21788
rect 50536 21728 50600 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 65656 21244 65720 21248
rect 65656 21188 65660 21244
rect 65660 21188 65716 21244
rect 65716 21188 65720 21244
rect 65656 21184 65720 21188
rect 65736 21244 65800 21248
rect 65736 21188 65740 21244
rect 65740 21188 65796 21244
rect 65796 21188 65800 21244
rect 65736 21184 65800 21188
rect 65816 21244 65880 21248
rect 65816 21188 65820 21244
rect 65820 21188 65876 21244
rect 65876 21188 65880 21244
rect 65816 21184 65880 21188
rect 65896 21244 65960 21248
rect 65896 21188 65900 21244
rect 65900 21188 65956 21244
rect 65956 21188 65960 21244
rect 65896 21184 65960 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 50296 20700 50360 20704
rect 50296 20644 50300 20700
rect 50300 20644 50356 20700
rect 50356 20644 50360 20700
rect 50296 20640 50360 20644
rect 50376 20700 50440 20704
rect 50376 20644 50380 20700
rect 50380 20644 50436 20700
rect 50436 20644 50440 20700
rect 50376 20640 50440 20644
rect 50456 20700 50520 20704
rect 50456 20644 50460 20700
rect 50460 20644 50516 20700
rect 50516 20644 50520 20700
rect 50456 20640 50520 20644
rect 50536 20700 50600 20704
rect 50536 20644 50540 20700
rect 50540 20644 50596 20700
rect 50596 20644 50600 20700
rect 50536 20640 50600 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 65656 20156 65720 20160
rect 65656 20100 65660 20156
rect 65660 20100 65716 20156
rect 65716 20100 65720 20156
rect 65656 20096 65720 20100
rect 65736 20156 65800 20160
rect 65736 20100 65740 20156
rect 65740 20100 65796 20156
rect 65796 20100 65800 20156
rect 65736 20096 65800 20100
rect 65816 20156 65880 20160
rect 65816 20100 65820 20156
rect 65820 20100 65876 20156
rect 65876 20100 65880 20156
rect 65816 20096 65880 20100
rect 65896 20156 65960 20160
rect 65896 20100 65900 20156
rect 65900 20100 65956 20156
rect 65956 20100 65960 20156
rect 65896 20096 65960 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 50296 19612 50360 19616
rect 50296 19556 50300 19612
rect 50300 19556 50356 19612
rect 50356 19556 50360 19612
rect 50296 19552 50360 19556
rect 50376 19612 50440 19616
rect 50376 19556 50380 19612
rect 50380 19556 50436 19612
rect 50436 19556 50440 19612
rect 50376 19552 50440 19556
rect 50456 19612 50520 19616
rect 50456 19556 50460 19612
rect 50460 19556 50516 19612
rect 50516 19556 50520 19612
rect 50456 19552 50520 19556
rect 50536 19612 50600 19616
rect 50536 19556 50540 19612
rect 50540 19556 50596 19612
rect 50596 19556 50600 19612
rect 50536 19552 50600 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 65656 19068 65720 19072
rect 65656 19012 65660 19068
rect 65660 19012 65716 19068
rect 65716 19012 65720 19068
rect 65656 19008 65720 19012
rect 65736 19068 65800 19072
rect 65736 19012 65740 19068
rect 65740 19012 65796 19068
rect 65796 19012 65800 19068
rect 65736 19008 65800 19012
rect 65816 19068 65880 19072
rect 65816 19012 65820 19068
rect 65820 19012 65876 19068
rect 65876 19012 65880 19068
rect 65816 19008 65880 19012
rect 65896 19068 65960 19072
rect 65896 19012 65900 19068
rect 65900 19012 65956 19068
rect 65956 19012 65960 19068
rect 65896 19008 65960 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 50296 18524 50360 18528
rect 50296 18468 50300 18524
rect 50300 18468 50356 18524
rect 50356 18468 50360 18524
rect 50296 18464 50360 18468
rect 50376 18524 50440 18528
rect 50376 18468 50380 18524
rect 50380 18468 50436 18524
rect 50436 18468 50440 18524
rect 50376 18464 50440 18468
rect 50456 18524 50520 18528
rect 50456 18468 50460 18524
rect 50460 18468 50516 18524
rect 50516 18468 50520 18524
rect 50456 18464 50520 18468
rect 50536 18524 50600 18528
rect 50536 18468 50540 18524
rect 50540 18468 50596 18524
rect 50596 18468 50600 18524
rect 50536 18464 50600 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 65656 17980 65720 17984
rect 65656 17924 65660 17980
rect 65660 17924 65716 17980
rect 65716 17924 65720 17980
rect 65656 17920 65720 17924
rect 65736 17980 65800 17984
rect 65736 17924 65740 17980
rect 65740 17924 65796 17980
rect 65796 17924 65800 17980
rect 65736 17920 65800 17924
rect 65816 17980 65880 17984
rect 65816 17924 65820 17980
rect 65820 17924 65876 17980
rect 65876 17924 65880 17980
rect 65816 17920 65880 17924
rect 65896 17980 65960 17984
rect 65896 17924 65900 17980
rect 65900 17924 65956 17980
rect 65956 17924 65960 17980
rect 65896 17920 65960 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 50296 17436 50360 17440
rect 50296 17380 50300 17436
rect 50300 17380 50356 17436
rect 50356 17380 50360 17436
rect 50296 17376 50360 17380
rect 50376 17436 50440 17440
rect 50376 17380 50380 17436
rect 50380 17380 50436 17436
rect 50436 17380 50440 17436
rect 50376 17376 50440 17380
rect 50456 17436 50520 17440
rect 50456 17380 50460 17436
rect 50460 17380 50516 17436
rect 50516 17380 50520 17436
rect 50456 17376 50520 17380
rect 50536 17436 50600 17440
rect 50536 17380 50540 17436
rect 50540 17380 50596 17436
rect 50596 17380 50600 17436
rect 50536 17376 50600 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 65656 16892 65720 16896
rect 65656 16836 65660 16892
rect 65660 16836 65716 16892
rect 65716 16836 65720 16892
rect 65656 16832 65720 16836
rect 65736 16892 65800 16896
rect 65736 16836 65740 16892
rect 65740 16836 65796 16892
rect 65796 16836 65800 16892
rect 65736 16832 65800 16836
rect 65816 16892 65880 16896
rect 65816 16836 65820 16892
rect 65820 16836 65876 16892
rect 65876 16836 65880 16892
rect 65816 16832 65880 16836
rect 65896 16892 65960 16896
rect 65896 16836 65900 16892
rect 65900 16836 65956 16892
rect 65956 16836 65960 16892
rect 65896 16832 65960 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 50296 16348 50360 16352
rect 50296 16292 50300 16348
rect 50300 16292 50356 16348
rect 50356 16292 50360 16348
rect 50296 16288 50360 16292
rect 50376 16348 50440 16352
rect 50376 16292 50380 16348
rect 50380 16292 50436 16348
rect 50436 16292 50440 16348
rect 50376 16288 50440 16292
rect 50456 16348 50520 16352
rect 50456 16292 50460 16348
rect 50460 16292 50516 16348
rect 50516 16292 50520 16348
rect 50456 16288 50520 16292
rect 50536 16348 50600 16352
rect 50536 16292 50540 16348
rect 50540 16292 50596 16348
rect 50596 16292 50600 16348
rect 50536 16288 50600 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 65656 15804 65720 15808
rect 65656 15748 65660 15804
rect 65660 15748 65716 15804
rect 65716 15748 65720 15804
rect 65656 15744 65720 15748
rect 65736 15804 65800 15808
rect 65736 15748 65740 15804
rect 65740 15748 65796 15804
rect 65796 15748 65800 15804
rect 65736 15744 65800 15748
rect 65816 15804 65880 15808
rect 65816 15748 65820 15804
rect 65820 15748 65876 15804
rect 65876 15748 65880 15804
rect 65816 15744 65880 15748
rect 65896 15804 65960 15808
rect 65896 15748 65900 15804
rect 65900 15748 65956 15804
rect 65956 15748 65960 15804
rect 65896 15744 65960 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 50296 15260 50360 15264
rect 50296 15204 50300 15260
rect 50300 15204 50356 15260
rect 50356 15204 50360 15260
rect 50296 15200 50360 15204
rect 50376 15260 50440 15264
rect 50376 15204 50380 15260
rect 50380 15204 50436 15260
rect 50436 15204 50440 15260
rect 50376 15200 50440 15204
rect 50456 15260 50520 15264
rect 50456 15204 50460 15260
rect 50460 15204 50516 15260
rect 50516 15204 50520 15260
rect 50456 15200 50520 15204
rect 50536 15260 50600 15264
rect 50536 15204 50540 15260
rect 50540 15204 50596 15260
rect 50596 15204 50600 15260
rect 50536 15200 50600 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 65656 14716 65720 14720
rect 65656 14660 65660 14716
rect 65660 14660 65716 14716
rect 65716 14660 65720 14716
rect 65656 14656 65720 14660
rect 65736 14716 65800 14720
rect 65736 14660 65740 14716
rect 65740 14660 65796 14716
rect 65796 14660 65800 14716
rect 65736 14656 65800 14660
rect 65816 14716 65880 14720
rect 65816 14660 65820 14716
rect 65820 14660 65876 14716
rect 65876 14660 65880 14716
rect 65816 14656 65880 14660
rect 65896 14716 65960 14720
rect 65896 14660 65900 14716
rect 65900 14660 65956 14716
rect 65956 14660 65960 14716
rect 65896 14656 65960 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 50296 14172 50360 14176
rect 50296 14116 50300 14172
rect 50300 14116 50356 14172
rect 50356 14116 50360 14172
rect 50296 14112 50360 14116
rect 50376 14172 50440 14176
rect 50376 14116 50380 14172
rect 50380 14116 50436 14172
rect 50436 14116 50440 14172
rect 50376 14112 50440 14116
rect 50456 14172 50520 14176
rect 50456 14116 50460 14172
rect 50460 14116 50516 14172
rect 50516 14116 50520 14172
rect 50456 14112 50520 14116
rect 50536 14172 50600 14176
rect 50536 14116 50540 14172
rect 50540 14116 50596 14172
rect 50596 14116 50600 14172
rect 50536 14112 50600 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 65656 13628 65720 13632
rect 65656 13572 65660 13628
rect 65660 13572 65716 13628
rect 65716 13572 65720 13628
rect 65656 13568 65720 13572
rect 65736 13628 65800 13632
rect 65736 13572 65740 13628
rect 65740 13572 65796 13628
rect 65796 13572 65800 13628
rect 65736 13568 65800 13572
rect 65816 13628 65880 13632
rect 65816 13572 65820 13628
rect 65820 13572 65876 13628
rect 65876 13572 65880 13628
rect 65816 13568 65880 13572
rect 65896 13628 65960 13632
rect 65896 13572 65900 13628
rect 65900 13572 65956 13628
rect 65956 13572 65960 13628
rect 65896 13568 65960 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 50296 13084 50360 13088
rect 50296 13028 50300 13084
rect 50300 13028 50356 13084
rect 50356 13028 50360 13084
rect 50296 13024 50360 13028
rect 50376 13084 50440 13088
rect 50376 13028 50380 13084
rect 50380 13028 50436 13084
rect 50436 13028 50440 13084
rect 50376 13024 50440 13028
rect 50456 13084 50520 13088
rect 50456 13028 50460 13084
rect 50460 13028 50516 13084
rect 50516 13028 50520 13084
rect 50456 13024 50520 13028
rect 50536 13084 50600 13088
rect 50536 13028 50540 13084
rect 50540 13028 50596 13084
rect 50596 13028 50600 13084
rect 50536 13024 50600 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 65656 12540 65720 12544
rect 65656 12484 65660 12540
rect 65660 12484 65716 12540
rect 65716 12484 65720 12540
rect 65656 12480 65720 12484
rect 65736 12540 65800 12544
rect 65736 12484 65740 12540
rect 65740 12484 65796 12540
rect 65796 12484 65800 12540
rect 65736 12480 65800 12484
rect 65816 12540 65880 12544
rect 65816 12484 65820 12540
rect 65820 12484 65876 12540
rect 65876 12484 65880 12540
rect 65816 12480 65880 12484
rect 65896 12540 65960 12544
rect 65896 12484 65900 12540
rect 65900 12484 65956 12540
rect 65956 12484 65960 12540
rect 65896 12480 65960 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 50296 11996 50360 12000
rect 50296 11940 50300 11996
rect 50300 11940 50356 11996
rect 50356 11940 50360 11996
rect 50296 11936 50360 11940
rect 50376 11996 50440 12000
rect 50376 11940 50380 11996
rect 50380 11940 50436 11996
rect 50436 11940 50440 11996
rect 50376 11936 50440 11940
rect 50456 11996 50520 12000
rect 50456 11940 50460 11996
rect 50460 11940 50516 11996
rect 50516 11940 50520 11996
rect 50456 11936 50520 11940
rect 50536 11996 50600 12000
rect 50536 11940 50540 11996
rect 50540 11940 50596 11996
rect 50596 11940 50600 11996
rect 50536 11936 50600 11940
rect 16804 11460 16868 11524
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 65656 11452 65720 11456
rect 65656 11396 65660 11452
rect 65660 11396 65716 11452
rect 65716 11396 65720 11452
rect 65656 11392 65720 11396
rect 65736 11452 65800 11456
rect 65736 11396 65740 11452
rect 65740 11396 65796 11452
rect 65796 11396 65800 11452
rect 65736 11392 65800 11396
rect 65816 11452 65880 11456
rect 65816 11396 65820 11452
rect 65820 11396 65876 11452
rect 65876 11396 65880 11452
rect 65816 11392 65880 11396
rect 65896 11452 65960 11456
rect 65896 11396 65900 11452
rect 65900 11396 65956 11452
rect 65956 11396 65960 11452
rect 65896 11392 65960 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 50296 10908 50360 10912
rect 50296 10852 50300 10908
rect 50300 10852 50356 10908
rect 50356 10852 50360 10908
rect 50296 10848 50360 10852
rect 50376 10908 50440 10912
rect 50376 10852 50380 10908
rect 50380 10852 50436 10908
rect 50436 10852 50440 10908
rect 50376 10848 50440 10852
rect 50456 10908 50520 10912
rect 50456 10852 50460 10908
rect 50460 10852 50516 10908
rect 50516 10852 50520 10908
rect 50456 10848 50520 10852
rect 50536 10908 50600 10912
rect 50536 10852 50540 10908
rect 50540 10852 50596 10908
rect 50596 10852 50600 10908
rect 50536 10848 50600 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 65656 10364 65720 10368
rect 65656 10308 65660 10364
rect 65660 10308 65716 10364
rect 65716 10308 65720 10364
rect 65656 10304 65720 10308
rect 65736 10364 65800 10368
rect 65736 10308 65740 10364
rect 65740 10308 65796 10364
rect 65796 10308 65800 10364
rect 65736 10304 65800 10308
rect 65816 10364 65880 10368
rect 65816 10308 65820 10364
rect 65820 10308 65876 10364
rect 65876 10308 65880 10364
rect 65816 10304 65880 10308
rect 65896 10364 65960 10368
rect 65896 10308 65900 10364
rect 65900 10308 65956 10364
rect 65956 10308 65960 10364
rect 65896 10304 65960 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 50296 9820 50360 9824
rect 50296 9764 50300 9820
rect 50300 9764 50356 9820
rect 50356 9764 50360 9820
rect 50296 9760 50360 9764
rect 50376 9820 50440 9824
rect 50376 9764 50380 9820
rect 50380 9764 50436 9820
rect 50436 9764 50440 9820
rect 50376 9760 50440 9764
rect 50456 9820 50520 9824
rect 50456 9764 50460 9820
rect 50460 9764 50516 9820
rect 50516 9764 50520 9820
rect 50456 9760 50520 9764
rect 50536 9820 50600 9824
rect 50536 9764 50540 9820
rect 50540 9764 50596 9820
rect 50596 9764 50600 9820
rect 50536 9760 50600 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 65656 9276 65720 9280
rect 65656 9220 65660 9276
rect 65660 9220 65716 9276
rect 65716 9220 65720 9276
rect 65656 9216 65720 9220
rect 65736 9276 65800 9280
rect 65736 9220 65740 9276
rect 65740 9220 65796 9276
rect 65796 9220 65800 9276
rect 65736 9216 65800 9220
rect 65816 9276 65880 9280
rect 65816 9220 65820 9276
rect 65820 9220 65876 9276
rect 65876 9220 65880 9276
rect 65816 9216 65880 9220
rect 65896 9276 65960 9280
rect 65896 9220 65900 9276
rect 65900 9220 65956 9276
rect 65956 9220 65960 9276
rect 65896 9216 65960 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 50296 8732 50360 8736
rect 50296 8676 50300 8732
rect 50300 8676 50356 8732
rect 50356 8676 50360 8732
rect 50296 8672 50360 8676
rect 50376 8732 50440 8736
rect 50376 8676 50380 8732
rect 50380 8676 50436 8732
rect 50436 8676 50440 8732
rect 50376 8672 50440 8676
rect 50456 8732 50520 8736
rect 50456 8676 50460 8732
rect 50460 8676 50516 8732
rect 50516 8676 50520 8732
rect 50456 8672 50520 8676
rect 50536 8732 50600 8736
rect 50536 8676 50540 8732
rect 50540 8676 50596 8732
rect 50596 8676 50600 8732
rect 50536 8672 50600 8676
rect 6868 8332 6932 8396
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 65656 8188 65720 8192
rect 65656 8132 65660 8188
rect 65660 8132 65716 8188
rect 65716 8132 65720 8188
rect 65656 8128 65720 8132
rect 65736 8188 65800 8192
rect 65736 8132 65740 8188
rect 65740 8132 65796 8188
rect 65796 8132 65800 8188
rect 65736 8128 65800 8132
rect 65816 8188 65880 8192
rect 65816 8132 65820 8188
rect 65820 8132 65876 8188
rect 65876 8132 65880 8188
rect 65816 8128 65880 8132
rect 65896 8188 65960 8192
rect 65896 8132 65900 8188
rect 65900 8132 65956 8188
rect 65956 8132 65960 8188
rect 65896 8128 65960 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 50296 7644 50360 7648
rect 50296 7588 50300 7644
rect 50300 7588 50356 7644
rect 50356 7588 50360 7644
rect 50296 7584 50360 7588
rect 50376 7644 50440 7648
rect 50376 7588 50380 7644
rect 50380 7588 50436 7644
rect 50436 7588 50440 7644
rect 50376 7584 50440 7588
rect 50456 7644 50520 7648
rect 50456 7588 50460 7644
rect 50460 7588 50516 7644
rect 50516 7588 50520 7644
rect 50456 7584 50520 7588
rect 50536 7644 50600 7648
rect 50536 7588 50540 7644
rect 50540 7588 50596 7644
rect 50596 7588 50600 7644
rect 50536 7584 50600 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 65656 7100 65720 7104
rect 65656 7044 65660 7100
rect 65660 7044 65716 7100
rect 65716 7044 65720 7100
rect 65656 7040 65720 7044
rect 65736 7100 65800 7104
rect 65736 7044 65740 7100
rect 65740 7044 65796 7100
rect 65796 7044 65800 7100
rect 65736 7040 65800 7044
rect 65816 7100 65880 7104
rect 65816 7044 65820 7100
rect 65820 7044 65876 7100
rect 65876 7044 65880 7100
rect 65816 7040 65880 7044
rect 65896 7100 65960 7104
rect 65896 7044 65900 7100
rect 65900 7044 65956 7100
rect 65956 7044 65960 7100
rect 65896 7040 65960 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 50296 6556 50360 6560
rect 50296 6500 50300 6556
rect 50300 6500 50356 6556
rect 50356 6500 50360 6556
rect 50296 6496 50360 6500
rect 50376 6556 50440 6560
rect 50376 6500 50380 6556
rect 50380 6500 50436 6556
rect 50436 6500 50440 6556
rect 50376 6496 50440 6500
rect 50456 6556 50520 6560
rect 50456 6500 50460 6556
rect 50460 6500 50516 6556
rect 50516 6500 50520 6556
rect 50456 6496 50520 6500
rect 50536 6556 50600 6560
rect 50536 6500 50540 6556
rect 50540 6500 50596 6556
rect 50596 6500 50600 6556
rect 50536 6496 50600 6500
rect 20668 6292 20732 6356
rect 12756 6156 12820 6220
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 65656 6012 65720 6016
rect 65656 5956 65660 6012
rect 65660 5956 65716 6012
rect 65716 5956 65720 6012
rect 65656 5952 65720 5956
rect 65736 6012 65800 6016
rect 65736 5956 65740 6012
rect 65740 5956 65796 6012
rect 65796 5956 65800 6012
rect 65736 5952 65800 5956
rect 65816 6012 65880 6016
rect 65816 5956 65820 6012
rect 65820 5956 65876 6012
rect 65876 5956 65880 6012
rect 65816 5952 65880 5956
rect 65896 6012 65960 6016
rect 65896 5956 65900 6012
rect 65900 5956 65956 6012
rect 65956 5956 65960 6012
rect 65896 5952 65960 5956
rect 13124 5612 13188 5676
rect 17908 5612 17972 5676
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 50296 5468 50360 5472
rect 50296 5412 50300 5468
rect 50300 5412 50356 5468
rect 50356 5412 50360 5468
rect 50296 5408 50360 5412
rect 50376 5468 50440 5472
rect 50376 5412 50380 5468
rect 50380 5412 50436 5468
rect 50436 5412 50440 5468
rect 50376 5408 50440 5412
rect 50456 5468 50520 5472
rect 50456 5412 50460 5468
rect 50460 5412 50516 5468
rect 50516 5412 50520 5468
rect 50456 5408 50520 5412
rect 50536 5468 50600 5472
rect 50536 5412 50540 5468
rect 50540 5412 50596 5468
rect 50596 5412 50600 5468
rect 50536 5408 50600 5412
rect 19380 4932 19444 4996
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 65656 4924 65720 4928
rect 65656 4868 65660 4924
rect 65660 4868 65716 4924
rect 65716 4868 65720 4924
rect 65656 4864 65720 4868
rect 65736 4924 65800 4928
rect 65736 4868 65740 4924
rect 65740 4868 65796 4924
rect 65796 4868 65800 4924
rect 65736 4864 65800 4868
rect 65816 4924 65880 4928
rect 65816 4868 65820 4924
rect 65820 4868 65876 4924
rect 65876 4868 65880 4924
rect 65816 4864 65880 4868
rect 65896 4924 65960 4928
rect 65896 4868 65900 4924
rect 65900 4868 65956 4924
rect 65956 4868 65960 4924
rect 65896 4864 65960 4868
rect 16804 4796 16868 4860
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 50296 4380 50360 4384
rect 50296 4324 50300 4380
rect 50300 4324 50356 4380
rect 50356 4324 50360 4380
rect 50296 4320 50360 4324
rect 50376 4380 50440 4384
rect 50376 4324 50380 4380
rect 50380 4324 50436 4380
rect 50436 4324 50440 4380
rect 50376 4320 50440 4324
rect 50456 4380 50520 4384
rect 50456 4324 50460 4380
rect 50460 4324 50516 4380
rect 50516 4324 50520 4380
rect 50456 4320 50520 4324
rect 50536 4380 50600 4384
rect 50536 4324 50540 4380
rect 50540 4324 50596 4380
rect 50596 4324 50600 4380
rect 50536 4320 50600 4324
rect 6868 3980 6932 4044
rect 17908 3980 17972 4044
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 65656 3836 65720 3840
rect 65656 3780 65660 3836
rect 65660 3780 65716 3836
rect 65716 3780 65720 3836
rect 65656 3776 65720 3780
rect 65736 3836 65800 3840
rect 65736 3780 65740 3836
rect 65740 3780 65796 3836
rect 65796 3780 65800 3836
rect 65736 3776 65800 3780
rect 65816 3836 65880 3840
rect 65816 3780 65820 3836
rect 65820 3780 65876 3836
rect 65876 3780 65880 3836
rect 65816 3776 65880 3780
rect 65896 3836 65960 3840
rect 65896 3780 65900 3836
rect 65900 3780 65956 3836
rect 65956 3780 65960 3836
rect 65896 3776 65960 3780
rect 19380 3436 19444 3500
rect 12756 3300 12820 3364
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 50296 3292 50360 3296
rect 50296 3236 50300 3292
rect 50300 3236 50356 3292
rect 50356 3236 50360 3292
rect 50296 3232 50360 3236
rect 50376 3292 50440 3296
rect 50376 3236 50380 3292
rect 50380 3236 50436 3292
rect 50436 3236 50440 3292
rect 50376 3232 50440 3236
rect 50456 3292 50520 3296
rect 50456 3236 50460 3292
rect 50460 3236 50516 3292
rect 50516 3236 50520 3292
rect 50456 3232 50520 3236
rect 50536 3292 50600 3296
rect 50536 3236 50540 3292
rect 50540 3236 50596 3292
rect 50596 3236 50600 3292
rect 50536 3232 50600 3236
rect 13124 3028 13188 3092
rect 20668 3088 20732 3092
rect 20668 3032 20718 3088
rect 20718 3032 20732 3088
rect 20668 3028 20732 3032
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 65656 2748 65720 2752
rect 65656 2692 65660 2748
rect 65660 2692 65716 2748
rect 65716 2692 65720 2748
rect 65656 2688 65720 2692
rect 65736 2748 65800 2752
rect 65736 2692 65740 2748
rect 65740 2692 65796 2748
rect 65796 2692 65800 2748
rect 65736 2688 65800 2692
rect 65816 2748 65880 2752
rect 65816 2692 65820 2748
rect 65820 2692 65876 2748
rect 65876 2692 65880 2748
rect 65816 2688 65880 2692
rect 65896 2748 65960 2752
rect 65896 2692 65900 2748
rect 65900 2692 65956 2748
rect 65956 2692 65960 2748
rect 65896 2688 65960 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
rect 50296 2204 50360 2208
rect 50296 2148 50300 2204
rect 50300 2148 50356 2204
rect 50356 2148 50360 2204
rect 50296 2144 50360 2148
rect 50376 2204 50440 2208
rect 50376 2148 50380 2204
rect 50380 2148 50436 2204
rect 50436 2148 50440 2204
rect 50376 2144 50440 2148
rect 50456 2204 50520 2208
rect 50456 2148 50460 2204
rect 50460 2148 50516 2204
rect 50516 2148 50520 2204
rect 50456 2144 50520 2148
rect 50536 2204 50600 2208
rect 50536 2148 50540 2204
rect 50540 2148 50596 2204
rect 50596 2148 50600 2204
rect 50536 2144 50600 2148
<< metal4 >>
rect 4208 57152 4528 57712
rect 4208 57088 4216 57152
rect 4280 57088 4296 57152
rect 4360 57088 4376 57152
rect 4440 57088 4456 57152
rect 4520 57088 4528 57152
rect 4208 56064 4528 57088
rect 4208 56000 4216 56064
rect 4280 56000 4296 56064
rect 4360 56000 4376 56064
rect 4440 56000 4456 56064
rect 4520 56000 4528 56064
rect 4208 54976 4528 56000
rect 4208 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4528 54976
rect 4208 53888 4528 54912
rect 4208 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4528 53888
rect 4208 52800 4528 53824
rect 4208 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4528 52800
rect 4208 51712 4528 52736
rect 4208 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4528 51712
rect 4208 50624 4528 51648
rect 4208 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4528 50624
rect 4208 49536 4528 50560
rect 4208 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4528 49536
rect 4208 48448 4528 49472
rect 4208 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4528 48448
rect 4208 47360 4528 48384
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 46272 4528 47296
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 45184 4528 46208
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 44096 4528 45120
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 43008 4528 44032
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 41920 4528 42944
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 19568 57696 19888 57712
rect 19568 57632 19576 57696
rect 19640 57632 19656 57696
rect 19720 57632 19736 57696
rect 19800 57632 19816 57696
rect 19880 57632 19888 57696
rect 19568 56608 19888 57632
rect 19568 56544 19576 56608
rect 19640 56544 19656 56608
rect 19720 56544 19736 56608
rect 19800 56544 19816 56608
rect 19880 56544 19888 56608
rect 19568 55520 19888 56544
rect 19568 55456 19576 55520
rect 19640 55456 19656 55520
rect 19720 55456 19736 55520
rect 19800 55456 19816 55520
rect 19880 55456 19888 55520
rect 19568 54432 19888 55456
rect 19568 54368 19576 54432
rect 19640 54368 19656 54432
rect 19720 54368 19736 54432
rect 19800 54368 19816 54432
rect 19880 54368 19888 54432
rect 19568 53344 19888 54368
rect 19568 53280 19576 53344
rect 19640 53280 19656 53344
rect 19720 53280 19736 53344
rect 19800 53280 19816 53344
rect 19880 53280 19888 53344
rect 19568 52256 19888 53280
rect 19568 52192 19576 52256
rect 19640 52192 19656 52256
rect 19720 52192 19736 52256
rect 19800 52192 19816 52256
rect 19880 52192 19888 52256
rect 19568 51168 19888 52192
rect 19568 51104 19576 51168
rect 19640 51104 19656 51168
rect 19720 51104 19736 51168
rect 19800 51104 19816 51168
rect 19880 51104 19888 51168
rect 19568 50080 19888 51104
rect 19568 50016 19576 50080
rect 19640 50016 19656 50080
rect 19720 50016 19736 50080
rect 19800 50016 19816 50080
rect 19880 50016 19888 50080
rect 19568 48992 19888 50016
rect 19568 48928 19576 48992
rect 19640 48928 19656 48992
rect 19720 48928 19736 48992
rect 19800 48928 19816 48992
rect 19880 48928 19888 48992
rect 19568 47904 19888 48928
rect 19568 47840 19576 47904
rect 19640 47840 19656 47904
rect 19720 47840 19736 47904
rect 19800 47840 19816 47904
rect 19880 47840 19888 47904
rect 19568 46816 19888 47840
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 45728 19888 46752
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 44640 19888 45664
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 43552 19888 44576
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 42464 19888 43488
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 41376 19888 42400
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 40288 19888 41312
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 39200 19888 40224
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 38112 19888 39136
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 37024 19888 38048
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 16803 11524 16869 11525
rect 16803 11460 16804 11524
rect 16868 11460 16869 11524
rect 16803 11459 16869 11460
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 6867 8396 6933 8397
rect 6867 8332 6868 8396
rect 6932 8332 6933 8396
rect 6867 8331 6933 8332
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 6870 4045 6930 8331
rect 12755 6220 12821 6221
rect 12755 6156 12756 6220
rect 12820 6156 12821 6220
rect 12755 6155 12821 6156
rect 6867 4044 6933 4045
rect 6867 3980 6868 4044
rect 6932 3980 6933 4044
rect 6867 3979 6933 3980
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 12758 3365 12818 6155
rect 13123 5676 13189 5677
rect 13123 5612 13124 5676
rect 13188 5612 13189 5676
rect 13123 5611 13189 5612
rect 12755 3364 12821 3365
rect 12755 3300 12756 3364
rect 12820 3300 12821 3364
rect 12755 3299 12821 3300
rect 13126 3093 13186 5611
rect 16806 4861 16866 11459
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 17907 5676 17973 5677
rect 17907 5612 17908 5676
rect 17972 5612 17973 5676
rect 17907 5611 17973 5612
rect 16803 4860 16869 4861
rect 16803 4796 16804 4860
rect 16868 4796 16869 4860
rect 16803 4795 16869 4796
rect 17910 4045 17970 5611
rect 19568 5472 19888 6496
rect 34928 57152 35248 57712
rect 34928 57088 34936 57152
rect 35000 57088 35016 57152
rect 35080 57088 35096 57152
rect 35160 57088 35176 57152
rect 35240 57088 35248 57152
rect 34928 56064 35248 57088
rect 34928 56000 34936 56064
rect 35000 56000 35016 56064
rect 35080 56000 35096 56064
rect 35160 56000 35176 56064
rect 35240 56000 35248 56064
rect 34928 54976 35248 56000
rect 34928 54912 34936 54976
rect 35000 54912 35016 54976
rect 35080 54912 35096 54976
rect 35160 54912 35176 54976
rect 35240 54912 35248 54976
rect 34928 53888 35248 54912
rect 34928 53824 34936 53888
rect 35000 53824 35016 53888
rect 35080 53824 35096 53888
rect 35160 53824 35176 53888
rect 35240 53824 35248 53888
rect 34928 52800 35248 53824
rect 34928 52736 34936 52800
rect 35000 52736 35016 52800
rect 35080 52736 35096 52800
rect 35160 52736 35176 52800
rect 35240 52736 35248 52800
rect 34928 51712 35248 52736
rect 34928 51648 34936 51712
rect 35000 51648 35016 51712
rect 35080 51648 35096 51712
rect 35160 51648 35176 51712
rect 35240 51648 35248 51712
rect 34928 50624 35248 51648
rect 34928 50560 34936 50624
rect 35000 50560 35016 50624
rect 35080 50560 35096 50624
rect 35160 50560 35176 50624
rect 35240 50560 35248 50624
rect 34928 49536 35248 50560
rect 34928 49472 34936 49536
rect 35000 49472 35016 49536
rect 35080 49472 35096 49536
rect 35160 49472 35176 49536
rect 35240 49472 35248 49536
rect 34928 48448 35248 49472
rect 34928 48384 34936 48448
rect 35000 48384 35016 48448
rect 35080 48384 35096 48448
rect 35160 48384 35176 48448
rect 35240 48384 35248 48448
rect 34928 47360 35248 48384
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 46272 35248 47296
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 45184 35248 46208
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 44096 35248 45120
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 43008 35248 44032
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 41920 35248 42944
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 40832 35248 41856
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 39744 35248 40768
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 38656 35248 39680
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 20667 6356 20733 6357
rect 20667 6292 20668 6356
rect 20732 6292 20733 6356
rect 20667 6291 20733 6292
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19379 4996 19445 4997
rect 19379 4932 19380 4996
rect 19444 4932 19445 4996
rect 19379 4931 19445 4932
rect 17907 4044 17973 4045
rect 17907 3980 17908 4044
rect 17972 3980 17973 4044
rect 17907 3979 17973 3980
rect 19382 3501 19442 4931
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19379 3500 19445 3501
rect 19379 3436 19380 3500
rect 19444 3436 19445 3500
rect 19379 3435 19445 3436
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 13123 3092 13189 3093
rect 13123 3028 13124 3092
rect 13188 3028 13189 3092
rect 13123 3027 13189 3028
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 2208 19888 3232
rect 20670 3093 20730 6291
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 20667 3092 20733 3093
rect 20667 3028 20668 3092
rect 20732 3028 20733 3092
rect 20667 3027 20733 3028
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
rect 50288 57696 50608 57712
rect 50288 57632 50296 57696
rect 50360 57632 50376 57696
rect 50440 57632 50456 57696
rect 50520 57632 50536 57696
rect 50600 57632 50608 57696
rect 50288 56608 50608 57632
rect 50288 56544 50296 56608
rect 50360 56544 50376 56608
rect 50440 56544 50456 56608
rect 50520 56544 50536 56608
rect 50600 56544 50608 56608
rect 50288 55520 50608 56544
rect 50288 55456 50296 55520
rect 50360 55456 50376 55520
rect 50440 55456 50456 55520
rect 50520 55456 50536 55520
rect 50600 55456 50608 55520
rect 50288 54432 50608 55456
rect 50288 54368 50296 54432
rect 50360 54368 50376 54432
rect 50440 54368 50456 54432
rect 50520 54368 50536 54432
rect 50600 54368 50608 54432
rect 50288 53344 50608 54368
rect 50288 53280 50296 53344
rect 50360 53280 50376 53344
rect 50440 53280 50456 53344
rect 50520 53280 50536 53344
rect 50600 53280 50608 53344
rect 50288 52256 50608 53280
rect 50288 52192 50296 52256
rect 50360 52192 50376 52256
rect 50440 52192 50456 52256
rect 50520 52192 50536 52256
rect 50600 52192 50608 52256
rect 50288 51168 50608 52192
rect 50288 51104 50296 51168
rect 50360 51104 50376 51168
rect 50440 51104 50456 51168
rect 50520 51104 50536 51168
rect 50600 51104 50608 51168
rect 50288 50080 50608 51104
rect 50288 50016 50296 50080
rect 50360 50016 50376 50080
rect 50440 50016 50456 50080
rect 50520 50016 50536 50080
rect 50600 50016 50608 50080
rect 50288 48992 50608 50016
rect 50288 48928 50296 48992
rect 50360 48928 50376 48992
rect 50440 48928 50456 48992
rect 50520 48928 50536 48992
rect 50600 48928 50608 48992
rect 50288 47904 50608 48928
rect 50288 47840 50296 47904
rect 50360 47840 50376 47904
rect 50440 47840 50456 47904
rect 50520 47840 50536 47904
rect 50600 47840 50608 47904
rect 50288 46816 50608 47840
rect 50288 46752 50296 46816
rect 50360 46752 50376 46816
rect 50440 46752 50456 46816
rect 50520 46752 50536 46816
rect 50600 46752 50608 46816
rect 50288 45728 50608 46752
rect 50288 45664 50296 45728
rect 50360 45664 50376 45728
rect 50440 45664 50456 45728
rect 50520 45664 50536 45728
rect 50600 45664 50608 45728
rect 50288 44640 50608 45664
rect 50288 44576 50296 44640
rect 50360 44576 50376 44640
rect 50440 44576 50456 44640
rect 50520 44576 50536 44640
rect 50600 44576 50608 44640
rect 50288 43552 50608 44576
rect 50288 43488 50296 43552
rect 50360 43488 50376 43552
rect 50440 43488 50456 43552
rect 50520 43488 50536 43552
rect 50600 43488 50608 43552
rect 50288 42464 50608 43488
rect 50288 42400 50296 42464
rect 50360 42400 50376 42464
rect 50440 42400 50456 42464
rect 50520 42400 50536 42464
rect 50600 42400 50608 42464
rect 50288 41376 50608 42400
rect 50288 41312 50296 41376
rect 50360 41312 50376 41376
rect 50440 41312 50456 41376
rect 50520 41312 50536 41376
rect 50600 41312 50608 41376
rect 50288 40288 50608 41312
rect 50288 40224 50296 40288
rect 50360 40224 50376 40288
rect 50440 40224 50456 40288
rect 50520 40224 50536 40288
rect 50600 40224 50608 40288
rect 50288 39200 50608 40224
rect 50288 39136 50296 39200
rect 50360 39136 50376 39200
rect 50440 39136 50456 39200
rect 50520 39136 50536 39200
rect 50600 39136 50608 39200
rect 50288 38112 50608 39136
rect 50288 38048 50296 38112
rect 50360 38048 50376 38112
rect 50440 38048 50456 38112
rect 50520 38048 50536 38112
rect 50600 38048 50608 38112
rect 50288 37024 50608 38048
rect 50288 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50608 37024
rect 50288 35936 50608 36960
rect 50288 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50608 35936
rect 50288 34848 50608 35872
rect 50288 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50608 34848
rect 50288 33760 50608 34784
rect 50288 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50608 33760
rect 50288 32672 50608 33696
rect 50288 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50608 32672
rect 50288 31584 50608 32608
rect 50288 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50608 31584
rect 50288 30496 50608 31520
rect 50288 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50608 30496
rect 50288 29408 50608 30432
rect 50288 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50608 29408
rect 50288 28320 50608 29344
rect 50288 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50608 28320
rect 50288 27232 50608 28256
rect 50288 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50608 27232
rect 50288 26144 50608 27168
rect 50288 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50608 26144
rect 50288 25056 50608 26080
rect 50288 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50608 25056
rect 50288 23968 50608 24992
rect 50288 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50608 23968
rect 50288 22880 50608 23904
rect 50288 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50608 22880
rect 50288 21792 50608 22816
rect 50288 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50608 21792
rect 50288 20704 50608 21728
rect 50288 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50608 20704
rect 50288 19616 50608 20640
rect 50288 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50608 19616
rect 50288 18528 50608 19552
rect 50288 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50608 18528
rect 50288 17440 50608 18464
rect 50288 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50608 17440
rect 50288 16352 50608 17376
rect 50288 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50608 16352
rect 50288 15264 50608 16288
rect 50288 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50608 15264
rect 50288 14176 50608 15200
rect 50288 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50608 14176
rect 50288 13088 50608 14112
rect 50288 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50608 13088
rect 50288 12000 50608 13024
rect 50288 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50608 12000
rect 50288 10912 50608 11936
rect 50288 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50608 10912
rect 50288 9824 50608 10848
rect 50288 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50608 9824
rect 50288 8736 50608 9760
rect 50288 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50608 8736
rect 50288 7648 50608 8672
rect 50288 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50608 7648
rect 50288 6560 50608 7584
rect 50288 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50608 6560
rect 50288 5472 50608 6496
rect 50288 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50608 5472
rect 50288 4384 50608 5408
rect 50288 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50608 4384
rect 50288 3296 50608 4320
rect 50288 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50608 3296
rect 50288 2208 50608 3232
rect 50288 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50608 2208
rect 50288 2128 50608 2144
rect 65648 57152 65968 57712
rect 65648 57088 65656 57152
rect 65720 57088 65736 57152
rect 65800 57088 65816 57152
rect 65880 57088 65896 57152
rect 65960 57088 65968 57152
rect 65648 56064 65968 57088
rect 65648 56000 65656 56064
rect 65720 56000 65736 56064
rect 65800 56000 65816 56064
rect 65880 56000 65896 56064
rect 65960 56000 65968 56064
rect 65648 54976 65968 56000
rect 65648 54912 65656 54976
rect 65720 54912 65736 54976
rect 65800 54912 65816 54976
rect 65880 54912 65896 54976
rect 65960 54912 65968 54976
rect 65648 53888 65968 54912
rect 65648 53824 65656 53888
rect 65720 53824 65736 53888
rect 65800 53824 65816 53888
rect 65880 53824 65896 53888
rect 65960 53824 65968 53888
rect 65648 52800 65968 53824
rect 65648 52736 65656 52800
rect 65720 52736 65736 52800
rect 65800 52736 65816 52800
rect 65880 52736 65896 52800
rect 65960 52736 65968 52800
rect 65648 51712 65968 52736
rect 65648 51648 65656 51712
rect 65720 51648 65736 51712
rect 65800 51648 65816 51712
rect 65880 51648 65896 51712
rect 65960 51648 65968 51712
rect 65648 50624 65968 51648
rect 65648 50560 65656 50624
rect 65720 50560 65736 50624
rect 65800 50560 65816 50624
rect 65880 50560 65896 50624
rect 65960 50560 65968 50624
rect 65648 49536 65968 50560
rect 65648 49472 65656 49536
rect 65720 49472 65736 49536
rect 65800 49472 65816 49536
rect 65880 49472 65896 49536
rect 65960 49472 65968 49536
rect 65648 48448 65968 49472
rect 65648 48384 65656 48448
rect 65720 48384 65736 48448
rect 65800 48384 65816 48448
rect 65880 48384 65896 48448
rect 65960 48384 65968 48448
rect 65648 47360 65968 48384
rect 65648 47296 65656 47360
rect 65720 47296 65736 47360
rect 65800 47296 65816 47360
rect 65880 47296 65896 47360
rect 65960 47296 65968 47360
rect 65648 46272 65968 47296
rect 65648 46208 65656 46272
rect 65720 46208 65736 46272
rect 65800 46208 65816 46272
rect 65880 46208 65896 46272
rect 65960 46208 65968 46272
rect 65648 45184 65968 46208
rect 65648 45120 65656 45184
rect 65720 45120 65736 45184
rect 65800 45120 65816 45184
rect 65880 45120 65896 45184
rect 65960 45120 65968 45184
rect 65648 44096 65968 45120
rect 65648 44032 65656 44096
rect 65720 44032 65736 44096
rect 65800 44032 65816 44096
rect 65880 44032 65896 44096
rect 65960 44032 65968 44096
rect 65648 43008 65968 44032
rect 65648 42944 65656 43008
rect 65720 42944 65736 43008
rect 65800 42944 65816 43008
rect 65880 42944 65896 43008
rect 65960 42944 65968 43008
rect 65648 41920 65968 42944
rect 65648 41856 65656 41920
rect 65720 41856 65736 41920
rect 65800 41856 65816 41920
rect 65880 41856 65896 41920
rect 65960 41856 65968 41920
rect 65648 40832 65968 41856
rect 65648 40768 65656 40832
rect 65720 40768 65736 40832
rect 65800 40768 65816 40832
rect 65880 40768 65896 40832
rect 65960 40768 65968 40832
rect 65648 39744 65968 40768
rect 65648 39680 65656 39744
rect 65720 39680 65736 39744
rect 65800 39680 65816 39744
rect 65880 39680 65896 39744
rect 65960 39680 65968 39744
rect 65648 38656 65968 39680
rect 65648 38592 65656 38656
rect 65720 38592 65736 38656
rect 65800 38592 65816 38656
rect 65880 38592 65896 38656
rect 65960 38592 65968 38656
rect 65648 37568 65968 38592
rect 65648 37504 65656 37568
rect 65720 37504 65736 37568
rect 65800 37504 65816 37568
rect 65880 37504 65896 37568
rect 65960 37504 65968 37568
rect 65648 36480 65968 37504
rect 65648 36416 65656 36480
rect 65720 36416 65736 36480
rect 65800 36416 65816 36480
rect 65880 36416 65896 36480
rect 65960 36416 65968 36480
rect 65648 35392 65968 36416
rect 65648 35328 65656 35392
rect 65720 35328 65736 35392
rect 65800 35328 65816 35392
rect 65880 35328 65896 35392
rect 65960 35328 65968 35392
rect 65648 34304 65968 35328
rect 65648 34240 65656 34304
rect 65720 34240 65736 34304
rect 65800 34240 65816 34304
rect 65880 34240 65896 34304
rect 65960 34240 65968 34304
rect 65648 33216 65968 34240
rect 65648 33152 65656 33216
rect 65720 33152 65736 33216
rect 65800 33152 65816 33216
rect 65880 33152 65896 33216
rect 65960 33152 65968 33216
rect 65648 32128 65968 33152
rect 65648 32064 65656 32128
rect 65720 32064 65736 32128
rect 65800 32064 65816 32128
rect 65880 32064 65896 32128
rect 65960 32064 65968 32128
rect 65648 31040 65968 32064
rect 65648 30976 65656 31040
rect 65720 30976 65736 31040
rect 65800 30976 65816 31040
rect 65880 30976 65896 31040
rect 65960 30976 65968 31040
rect 65648 29952 65968 30976
rect 65648 29888 65656 29952
rect 65720 29888 65736 29952
rect 65800 29888 65816 29952
rect 65880 29888 65896 29952
rect 65960 29888 65968 29952
rect 65648 28864 65968 29888
rect 65648 28800 65656 28864
rect 65720 28800 65736 28864
rect 65800 28800 65816 28864
rect 65880 28800 65896 28864
rect 65960 28800 65968 28864
rect 65648 27776 65968 28800
rect 65648 27712 65656 27776
rect 65720 27712 65736 27776
rect 65800 27712 65816 27776
rect 65880 27712 65896 27776
rect 65960 27712 65968 27776
rect 65648 26688 65968 27712
rect 65648 26624 65656 26688
rect 65720 26624 65736 26688
rect 65800 26624 65816 26688
rect 65880 26624 65896 26688
rect 65960 26624 65968 26688
rect 65648 25600 65968 26624
rect 65648 25536 65656 25600
rect 65720 25536 65736 25600
rect 65800 25536 65816 25600
rect 65880 25536 65896 25600
rect 65960 25536 65968 25600
rect 65648 24512 65968 25536
rect 65648 24448 65656 24512
rect 65720 24448 65736 24512
rect 65800 24448 65816 24512
rect 65880 24448 65896 24512
rect 65960 24448 65968 24512
rect 65648 23424 65968 24448
rect 65648 23360 65656 23424
rect 65720 23360 65736 23424
rect 65800 23360 65816 23424
rect 65880 23360 65896 23424
rect 65960 23360 65968 23424
rect 65648 22336 65968 23360
rect 65648 22272 65656 22336
rect 65720 22272 65736 22336
rect 65800 22272 65816 22336
rect 65880 22272 65896 22336
rect 65960 22272 65968 22336
rect 65648 21248 65968 22272
rect 65648 21184 65656 21248
rect 65720 21184 65736 21248
rect 65800 21184 65816 21248
rect 65880 21184 65896 21248
rect 65960 21184 65968 21248
rect 65648 20160 65968 21184
rect 65648 20096 65656 20160
rect 65720 20096 65736 20160
rect 65800 20096 65816 20160
rect 65880 20096 65896 20160
rect 65960 20096 65968 20160
rect 65648 19072 65968 20096
rect 65648 19008 65656 19072
rect 65720 19008 65736 19072
rect 65800 19008 65816 19072
rect 65880 19008 65896 19072
rect 65960 19008 65968 19072
rect 65648 17984 65968 19008
rect 65648 17920 65656 17984
rect 65720 17920 65736 17984
rect 65800 17920 65816 17984
rect 65880 17920 65896 17984
rect 65960 17920 65968 17984
rect 65648 16896 65968 17920
rect 65648 16832 65656 16896
rect 65720 16832 65736 16896
rect 65800 16832 65816 16896
rect 65880 16832 65896 16896
rect 65960 16832 65968 16896
rect 65648 15808 65968 16832
rect 65648 15744 65656 15808
rect 65720 15744 65736 15808
rect 65800 15744 65816 15808
rect 65880 15744 65896 15808
rect 65960 15744 65968 15808
rect 65648 14720 65968 15744
rect 65648 14656 65656 14720
rect 65720 14656 65736 14720
rect 65800 14656 65816 14720
rect 65880 14656 65896 14720
rect 65960 14656 65968 14720
rect 65648 13632 65968 14656
rect 65648 13568 65656 13632
rect 65720 13568 65736 13632
rect 65800 13568 65816 13632
rect 65880 13568 65896 13632
rect 65960 13568 65968 13632
rect 65648 12544 65968 13568
rect 65648 12480 65656 12544
rect 65720 12480 65736 12544
rect 65800 12480 65816 12544
rect 65880 12480 65896 12544
rect 65960 12480 65968 12544
rect 65648 11456 65968 12480
rect 65648 11392 65656 11456
rect 65720 11392 65736 11456
rect 65800 11392 65816 11456
rect 65880 11392 65896 11456
rect 65960 11392 65968 11456
rect 65648 10368 65968 11392
rect 65648 10304 65656 10368
rect 65720 10304 65736 10368
rect 65800 10304 65816 10368
rect 65880 10304 65896 10368
rect 65960 10304 65968 10368
rect 65648 9280 65968 10304
rect 65648 9216 65656 9280
rect 65720 9216 65736 9280
rect 65800 9216 65816 9280
rect 65880 9216 65896 9280
rect 65960 9216 65968 9280
rect 65648 8192 65968 9216
rect 65648 8128 65656 8192
rect 65720 8128 65736 8192
rect 65800 8128 65816 8192
rect 65880 8128 65896 8192
rect 65960 8128 65968 8192
rect 65648 7104 65968 8128
rect 65648 7040 65656 7104
rect 65720 7040 65736 7104
rect 65800 7040 65816 7104
rect 65880 7040 65896 7104
rect 65960 7040 65968 7104
rect 65648 6016 65968 7040
rect 65648 5952 65656 6016
rect 65720 5952 65736 6016
rect 65800 5952 65816 6016
rect 65880 5952 65896 6016
rect 65960 5952 65968 6016
rect 65648 4928 65968 5952
rect 65648 4864 65656 4928
rect 65720 4864 65736 4928
rect 65800 4864 65816 4928
rect 65880 4864 65896 4928
rect 65960 4864 65968 4928
rect 65648 3840 65968 4864
rect 65648 3776 65656 3840
rect 65720 3776 65736 3840
rect 65800 3776 65816 3840
rect 65880 3776 65896 3840
rect 65960 3776 65968 3840
rect 65648 2752 65968 3776
rect 65648 2688 65656 2752
rect 65720 2688 65736 2752
rect 65800 2688 65816 2752
rect 65880 2688 65896 2752
rect 65960 2688 65968 2752
rect 65648 2128 65968 2688
use sky130_fd_sc_hd__diode_2  ANTENNA__169__A dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 8004 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__174__B
timestamp 1649977179
transform 1 0 3772 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__176__A
timestamp 1649977179
transform -1 0 8740 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__177__A
timestamp 1649977179
transform -1 0 3312 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__179__A
timestamp 1649977179
transform 1 0 7268 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__195__A
timestamp 1649977179
transform 1 0 4876 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__196__A
timestamp 1649977179
transform -1 0 5520 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__210__A
timestamp 1649977179
transform 1 0 9200 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__211__A
timestamp 1649977179
transform 1 0 8924 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__225__A
timestamp 1649977179
transform 1 0 7636 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__240__A
timestamp 1649977179
transform 1 0 20056 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__254__B
timestamp 1649977179
transform 1 0 4876 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__255__A
timestamp 1649977179
transform 1 0 14168 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__257__A
timestamp 1649977179
transform 1 0 7544 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__260__A
timestamp 1649977179
transform 1 0 11408 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__270__A
timestamp 1649977179
transform -1 0 2944 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__272__A
timestamp 1649977179
transform 1 0 4784 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__274__A
timestamp 1649977179
transform 1 0 4416 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__284__A
timestamp 1649977179
transform 1 0 8924 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__286__A
timestamp 1649977179
transform 1 0 8924 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__288__A
timestamp 1649977179
transform -1 0 11684 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__298__A
timestamp 1649977179
transform 1 0 23736 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__299__A
timestamp 1649977179
transform -1 0 25208 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__300__A
timestamp 1649977179
transform -1 0 22264 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__302__A
timestamp 1649977179
transform -1 0 23368 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__312__A
timestamp 1649977179
transform -1 0 24472 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__313__A
timestamp 1649977179
transform -1 0 21804 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__314__A
timestamp 1649977179
transform 1 0 20516 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__316__A
timestamp 1649977179
transform 1 0 21160 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_wb_clk_i_A
timestamp 1649977179
transform -1 0 12328 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1649977179
transform -1 0 3128 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1649977179
transform -1 0 24564 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1649977179
transform -1 0 24840 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1649977179
transform -1 0 24564 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1649977179
transform -1 0 21988 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1649977179
transform -1 0 7268 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1649977179
transform -1 0 7452 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1649977179
transform -1 0 14628 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1649977179
transform -1 0 4876 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1649977179
transform -1 0 12788 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1649977179
transform -1 0 14260 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1649977179
transform -1 0 8372 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1649977179
transform -1 0 14260 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1649977179
transform -1 0 17940 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1649977179
transform -1 0 6716 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1649977179
transform -1 0 18676 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1649977179
transform -1 0 18492 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1649977179
transform -1 0 11040 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1649977179
transform -1 0 18768 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1649977179
transform -1 0 18124 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1649977179
transform -1 0 18124 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1649977179
transform -1 0 19412 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1649977179
transform -1 0 16836 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1649977179
transform -1 0 11224 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1649977179
transform -1 0 2760 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1649977179
transform -1 0 3680 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1649977179
transform -1 0 13156 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1649977179
transform -1 0 8924 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1649977179
transform -1 0 9108 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1649977179
transform -1 0 14812 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1649977179
transform -1 0 4324 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1649977179
transform -1 0 13616 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1649977179
transform -1 0 12052 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1649977179
transform -1 0 3312 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output35_A
timestamp 1649977179
transform -1 0 27140 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2484 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2760 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24
timestamp 1649977179
transform 1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29
timestamp 1649977179
transform 1 0 3772 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33
timestamp 1649977179
transform 1 0 4140 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40
timestamp 1649977179
transform 1 0 4784 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52
timestamp 1649977179
transform 1 0 5888 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_60
timestamp 1649977179
transform 1 0 6624 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_80
timestamp 1649977179
transform 1 0 8464 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_85 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 8924 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_92
timestamp 1649977179
transform 1 0 9568 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_100
timestamp 1649977179
transform 1 0 10304 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_108
timestamp 1649977179
transform 1 0 11040 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_113
timestamp 1649977179
transform 1 0 11500 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_120
timestamp 1649977179
transform 1 0 12144 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_128
timestamp 1649977179
transform 1 0 12880 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_136
timestamp 1649977179
transform 1 0 13616 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_141
timestamp 1649977179
transform 1 0 14076 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_148
timestamp 1649977179
transform 1 0 14720 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_156
timestamp 1649977179
transform 1 0 15456 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_164
timestamp 1649977179
transform 1 0 16192 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_169
timestamp 1649977179
transform 1 0 16652 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_189 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 18492 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_195
timestamp 1649977179
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_203
timestamp 1649977179
transform 1 0 19780 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_211
timestamp 1649977179
transform 1 0 20516 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_219
timestamp 1649977179
transform 1 0 21252 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_223
timestamp 1649977179
transform 1 0 21620 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_229 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 22172 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_237
timestamp 1649977179
transform 1 0 22908 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_241
timestamp 1649977179
transform 1 0 23276 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_248
timestamp 1649977179
transform 1 0 23920 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_253
timestamp 1649977179
transform 1 0 24380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_257
timestamp 1649977179
transform 1 0 24748 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_261
timestamp 1649977179
transform 1 0 25116 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_268
timestamp 1649977179
transform 1 0 25760 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_276
timestamp 1649977179
transform 1 0 26496 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_285
timestamp 1649977179
transform 1 0 27324 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_293
timestamp 1649977179
transform 1 0 28060 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_297
timestamp 1649977179
transform 1 0 28428 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_304
timestamp 1649977179
transform 1 0 29072 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_309
timestamp 1649977179
transform 1 0 29532 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_318
timestamp 1649977179
transform 1 0 30360 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_325
timestamp 1649977179
transform 1 0 31004 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_332
timestamp 1649977179
transform 1 0 31648 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_337
timestamp 1649977179
transform 1 0 32108 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_346
timestamp 1649977179
transform 1 0 32936 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_353
timestamp 1649977179
transform 1 0 33580 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_360
timestamp 1649977179
transform 1 0 34224 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_365
timestamp 1649977179
transform 1 0 34684 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_369
timestamp 1649977179
transform 1 0 35052 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_376
timestamp 1649977179
transform 1 0 35696 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_383
timestamp 1649977179
transform 1 0 36340 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_391
timestamp 1649977179
transform 1 0 37076 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_396
timestamp 1649977179
transform 1 0 37536 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_403
timestamp 1649977179
transform 1 0 38180 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_410
timestamp 1649977179
transform 1 0 38824 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_418
timestamp 1649977179
transform 1 0 39560 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_424
timestamp 1649977179
transform 1 0 40112 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_431
timestamp 1649977179
transform 1 0 40756 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_438
timestamp 1649977179
transform 1 0 41400 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_446
timestamp 1649977179
transform 1 0 42136 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_452
timestamp 1649977179
transform 1 0 42688 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_459
timestamp 1649977179
transform 1 0 43332 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_466
timestamp 1649977179
transform 1 0 43976 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_474
timestamp 1649977179
transform 1 0 44712 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_480
timestamp 1649977179
transform 1 0 45264 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_487
timestamp 1649977179
transform 1 0 45908 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_494
timestamp 1649977179
transform 1 0 46552 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_502
timestamp 1649977179
transform 1 0 47288 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_508
timestamp 1649977179
transform 1 0 47840 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_515
timestamp 1649977179
transform 1 0 48484 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_522
timestamp 1649977179
transform 1 0 49128 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_530
timestamp 1649977179
transform 1 0 49864 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_536
timestamp 1649977179
transform 1 0 50416 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_543
timestamp 1649977179
transform 1 0 51060 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_550
timestamp 1649977179
transform 1 0 51704 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_558
timestamp 1649977179
transform 1 0 52440 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_564
timestamp 1649977179
transform 1 0 52992 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_571
timestamp 1649977179
transform 1 0 53636 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_578
timestamp 1649977179
transform 1 0 54280 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_586
timestamp 1649977179
transform 1 0 55016 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_592
timestamp 1649977179
transform 1 0 55568 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_599
timestamp 1649977179
transform 1 0 56212 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_606
timestamp 1649977179
transform 1 0 56856 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_614
timestamp 1649977179
transform 1 0 57592 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_620
timestamp 1649977179
transform 1 0 58144 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_627
timestamp 1649977179
transform 1 0 58788 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_634
timestamp 1649977179
transform 1 0 59432 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_642
timestamp 1649977179
transform 1 0 60168 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_645
timestamp 1649977179
transform 1 0 60444 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_657
timestamp 1649977179
transform 1 0 61548 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_669
timestamp 1649977179
transform 1 0 62652 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_673
timestamp 1649977179
transform 1 0 63020 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_685
timestamp 1649977179
transform 1 0 64124 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_697
timestamp 1649977179
transform 1 0 65228 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_701
timestamp 1649977179
transform 1 0 65596 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_713
timestamp 1649977179
transform 1 0 66700 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_725
timestamp 1649977179
transform 1 0 67804 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_729
timestamp 1649977179
transform 1 0 68172 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1649977179
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_15
timestamp 1649977179
transform 1 0 2484 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_19
timestamp 1649977179
transform 1 0 2852 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_22
timestamp 1649977179
transform 1 0 3128 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_28
timestamp 1649977179
transform 1 0 3680 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_40
timestamp 1649977179
transform 1 0 4784 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_52
timestamp 1649977179
transform 1 0 5888 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_57
timestamp 1649977179
transform 1 0 6348 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_62
timestamp 1649977179
transform 1 0 6808 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_82
timestamp 1649977179
transform 1 0 8648 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_88
timestamp 1649977179
transform 1 0 9200 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1649977179
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1649977179
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_113
timestamp 1649977179
transform 1 0 11500 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_117
timestamp 1649977179
transform 1 0 11868 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_122
timestamp 1649977179
transform 1 0 12328 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_131
timestamp 1649977179
transform 1 0 13156 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_143
timestamp 1649977179
transform 1 0 14260 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_163
timestamp 1649977179
transform 1 0 16100 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1649977179
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_177
timestamp 1649977179
transform 1 0 17388 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_184
timestamp 1649977179
transform 1 0 18032 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_204
timestamp 1649977179
transform 1 0 19872 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_212
timestamp 1649977179
transform 1 0 20608 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_216
timestamp 1649977179
transform 1 0 20976 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_220
timestamp 1649977179
transform 1 0 21344 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_227
timestamp 1649977179
transform 1 0 21988 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_234
timestamp 1649977179
transform 1 0 22632 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_241
timestamp 1649977179
transform 1 0 23276 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_248
timestamp 1649977179
transform 1 0 23920 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_255
timestamp 1649977179
transform 1 0 24564 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_262
timestamp 1649977179
transform 1 0 25208 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_269
timestamp 1649977179
transform 1 0 25852 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_276
timestamp 1649977179
transform 1 0 26496 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_283
timestamp 1649977179
transform 1 0 27140 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_290
timestamp 1649977179
transform 1 0 27784 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_297
timestamp 1649977179
transform 1 0 28428 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_304
timestamp 1649977179
transform 1 0 29072 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_311
timestamp 1649977179
transform 1 0 29716 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_318
timestamp 1649977179
transform 1 0 30360 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_325
timestamp 1649977179
transform 1 0 31004 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_332
timestamp 1649977179
transform 1 0 31648 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_337
timestamp 1649977179
transform 1 0 32108 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_342
timestamp 1649977179
transform 1 0 32568 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_349
timestamp 1649977179
transform 1 0 33212 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_356
timestamp 1649977179
transform 1 0 33856 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_363
timestamp 1649977179
transform 1 0 34500 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_370
timestamp 1649977179
transform 1 0 35144 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_377
timestamp 1649977179
transform 1 0 35788 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_1_386
timestamp 1649977179
transform 1 0 36616 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_396
timestamp 1649977179
transform 1 0 37536 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_403
timestamp 1649977179
transform 1 0 38180 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_410
timestamp 1649977179
transform 1 0 38824 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_417
timestamp 1649977179
transform 1 0 39468 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_424
timestamp 1649977179
transform 1 0 40112 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_431
timestamp 1649977179
transform 1 0 40756 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_438
timestamp 1649977179
transform 1 0 41400 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_446
timestamp 1649977179
transform 1 0 42136 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_452
timestamp 1649977179
transform 1 0 42688 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_459
timestamp 1649977179
transform 1 0 43332 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_466
timestamp 1649977179
transform 1 0 43976 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_473
timestamp 1649977179
transform 1 0 44620 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_480
timestamp 1649977179
transform 1 0 45264 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_487
timestamp 1649977179
transform 1 0 45908 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_494
timestamp 1649977179
transform 1 0 46552 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_502
timestamp 1649977179
transform 1 0 47288 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_508
timestamp 1649977179
transform 1 0 47840 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_515
timestamp 1649977179
transform 1 0 48484 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_522
timestamp 1649977179
transform 1 0 49128 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_529
timestamp 1649977179
transform 1 0 49772 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_536
timestamp 1649977179
transform 1 0 50416 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_543
timestamp 1649977179
transform 1 0 51060 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_550
timestamp 1649977179
transform 1 0 51704 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_558
timestamp 1649977179
transform 1 0 52440 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_564
timestamp 1649977179
transform 1 0 52992 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_571
timestamp 1649977179
transform 1 0 53636 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_578
timestamp 1649977179
transform 1 0 54280 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_585
timestamp 1649977179
transform 1 0 54924 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_592
timestamp 1649977179
transform 1 0 55568 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_599
timestamp 1649977179
transform 1 0 56212 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_606
timestamp 1649977179
transform 1 0 56856 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_614
timestamp 1649977179
transform 1 0 57592 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_620
timestamp 1649977179
transform 1 0 58144 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_627
timestamp 1649977179
transform 1 0 58788 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_639
timestamp 1649977179
transform 1 0 59892 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_651
timestamp 1649977179
transform 1 0 60996 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_663
timestamp 1649977179
transform 1 0 62100 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_671
timestamp 1649977179
transform 1 0 62836 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_673
timestamp 1649977179
transform 1 0 63020 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_685
timestamp 1649977179
transform 1 0 64124 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_697
timestamp 1649977179
transform 1 0 65228 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_709
timestamp 1649977179
transform 1 0 66332 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_721
timestamp 1649977179
transform 1 0 67436 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_727
timestamp 1649977179
transform 1 0 67988 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_729
timestamp 1649977179
transform 1 0 68172 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1649977179
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1649977179
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1649977179
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_29
timestamp 1649977179
transform 1 0 3772 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_35
timestamp 1649977179
transform 1 0 4324 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_41
timestamp 1649977179
transform 1 0 4876 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_53
timestamp 1649977179
transform 1 0 5980 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_65
timestamp 1649977179
transform 1 0 7084 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_69
timestamp 1649977179
transform 1 0 7452 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_73
timestamp 1649977179
transform 1 0 7820 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_80
timestamp 1649977179
transform 1 0 8464 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_87
timestamp 1649977179
transform 1 0 9108 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_94
timestamp 1649977179
transform 1 0 9752 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_2_116
timestamp 1649977179
transform 1 0 11776 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_122
timestamp 1649977179
transform 1 0 12328 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1649977179
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1649977179
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_141
timestamp 1649977179
transform 1 0 14076 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_147
timestamp 1649977179
transform 1 0 14628 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_155
timestamp 1649977179
transform 1 0 15364 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_167
timestamp 1649977179
transform 1 0 16468 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_191
timestamp 1649977179
transform 1 0 18676 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1649977179
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_201
timestamp 1649977179
transform 1 0 19596 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_209
timestamp 1649977179
transform 1 0 20332 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_217
timestamp 1649977179
transform 1 0 21068 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_227
timestamp 1649977179
transform 1 0 21988 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_235
timestamp 1649977179
transform 1 0 22724 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_239
timestamp 1649977179
transform 1 0 23092 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_248
timestamp 1649977179
transform 1 0 23920 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_256
timestamp 1649977179
transform 1 0 24656 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_263
timestamp 1649977179
transform 1 0 25300 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_271
timestamp 1649977179
transform 1 0 26036 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_275
timestamp 1649977179
transform 1 0 26404 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_281
timestamp 1649977179
transform 1 0 26956 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_285
timestamp 1649977179
transform 1 0 27324 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_292
timestamp 1649977179
transform 1 0 27968 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_299
timestamp 1649977179
transform 1 0 28612 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1649977179
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_312
timestamp 1649977179
transform 1 0 29808 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_316
timestamp 1649977179
transform 1 0 30176 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_320
timestamp 1649977179
transform 1 0 30544 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_328
timestamp 1649977179
transform 1 0 31280 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_332
timestamp 1649977179
transform 1 0 31648 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_2_341
timestamp 1649977179
transform 1 0 32476 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_2_350
timestamp 1649977179
transform 1 0 33304 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_362
timestamp 1649977179
transform 1 0 34408 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1649977179
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_377
timestamp 1649977179
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_389
timestamp 1649977179
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_401
timestamp 1649977179
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_413
timestamp 1649977179
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp 1649977179
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_421
timestamp 1649977179
transform 1 0 39836 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_425
timestamp 1649977179
transform 1 0 40204 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_432
timestamp 1649977179
transform 1 0 40848 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_439
timestamp 1649977179
transform 1 0 41492 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_446
timestamp 1649977179
transform 1 0 42136 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_2_455
timestamp 1649977179
transform 1 0 42964 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_463
timestamp 1649977179
transform 1 0 43700 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_467
timestamp 1649977179
transform 1 0 44068 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_475
timestamp 1649977179
transform 1 0 44804 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_477
timestamp 1649977179
transform 1 0 44988 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_482
timestamp 1649977179
transform 1 0 45448 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_489
timestamp 1649977179
transform 1 0 46092 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_496
timestamp 1649977179
transform 1 0 46736 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_504
timestamp 1649977179
transform 1 0 47472 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_509
timestamp 1649977179
transform 1 0 47932 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_516
timestamp 1649977179
transform 1 0 48576 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_528
timestamp 1649977179
transform 1 0 49680 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_536
timestamp 1649977179
transform 1 0 50416 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_543
timestamp 1649977179
transform 1 0 51060 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_550
timestamp 1649977179
transform 1 0 51704 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_557
timestamp 1649977179
transform 1 0 52348 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_566
timestamp 1649977179
transform 1 0 53176 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_573
timestamp 1649977179
transform 1 0 53820 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_585
timestamp 1649977179
transform 1 0 54924 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_589
timestamp 1649977179
transform 1 0 55292 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_593
timestamp 1649977179
transform 1 0 55660 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_600
timestamp 1649977179
transform 1 0 56304 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_607
timestamp 1649977179
transform 1 0 56948 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_614
timestamp 1649977179
transform 1 0 57592 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_621
timestamp 1649977179
transform 1 0 58236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_633
timestamp 1649977179
transform 1 0 59340 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_641
timestamp 1649977179
transform 1 0 60076 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_645
timestamp 1649977179
transform 1 0 60444 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_657
timestamp 1649977179
transform 1 0 61548 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_669
timestamp 1649977179
transform 1 0 62652 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_681
timestamp 1649977179
transform 1 0 63756 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_693
timestamp 1649977179
transform 1 0 64860 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_699
timestamp 1649977179
transform 1 0 65412 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_701
timestamp 1649977179
transform 1 0 65596 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_713
timestamp 1649977179
transform 1 0 66700 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_725
timestamp 1649977179
transform 1 0 67804 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1649977179
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_15
timestamp 1649977179
transform 1 0 2484 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_20
timestamp 1649977179
transform 1 0 2944 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_29
timestamp 1649977179
transform 1 0 3772 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_43
timestamp 1649977179
transform 1 0 5060 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_52
timestamp 1649977179
transform 1 0 5888 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_57
timestamp 1649977179
transform 1 0 6348 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_75
timestamp 1649977179
transform 1 0 8004 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_95
timestamp 1649977179
transform 1 0 9844 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_103
timestamp 1649977179
transform 1 0 10580 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_108
timestamp 1649977179
transform 1 0 11040 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_115
timestamp 1649977179
transform 1 0 11684 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_127
timestamp 1649977179
transform 1 0 12788 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_147
timestamp 1649977179
transform 1 0 14628 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_151
timestamp 1649977179
transform 1 0 14996 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_156
timestamp 1649977179
transform 1 0 15456 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_164
timestamp 1649977179
transform 1 0 16192 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_171
timestamp 1649977179
transform 1 0 16836 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_179
timestamp 1649977179
transform 1 0 17572 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_199
timestamp 1649977179
transform 1 0 19412 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_206
timestamp 1649977179
transform 1 0 20056 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_213
timestamp 1649977179
transform 1 0 20700 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_220
timestamp 1649977179
transform 1 0 21344 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_231
timestamp 1649977179
transform 1 0 22356 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_238
timestamp 1649977179
transform 1 0 23000 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_245
timestamp 1649977179
transform 1 0 23644 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_252
timestamp 1649977179
transform 1 0 24288 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_258
timestamp 1649977179
transform 1 0 24840 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_270
timestamp 1649977179
transform 1 0 25944 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_278
timestamp 1649977179
transform 1 0 26680 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1649977179
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1649977179
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1649977179
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_317
timestamp 1649977179
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1649977179
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1649977179
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1649977179
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1649977179
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1649977179
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1649977179
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1649977179
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1649977179
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1649977179
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_405
timestamp 1649977179
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_417
timestamp 1649977179
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_429
timestamp 1649977179
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_441
timestamp 1649977179
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 1649977179
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_449
timestamp 1649977179
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_461
timestamp 1649977179
transform 1 0 43516 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_473
timestamp 1649977179
transform 1 0 44620 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_485
timestamp 1649977179
transform 1 0 45724 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_497
timestamp 1649977179
transform 1 0 46828 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_503
timestamp 1649977179
transform 1 0 47380 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_505
timestamp 1649977179
transform 1 0 47564 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_517
timestamp 1649977179
transform 1 0 48668 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_529
timestamp 1649977179
transform 1 0 49772 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_541
timestamp 1649977179
transform 1 0 50876 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_553
timestamp 1649977179
transform 1 0 51980 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_559
timestamp 1649977179
transform 1 0 52532 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_561
timestamp 1649977179
transform 1 0 52716 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_573
timestamp 1649977179
transform 1 0 53820 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_585
timestamp 1649977179
transform 1 0 54924 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_597
timestamp 1649977179
transform 1 0 56028 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_609
timestamp 1649977179
transform 1 0 57132 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_615
timestamp 1649977179
transform 1 0 57684 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_617
timestamp 1649977179
transform 1 0 57868 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_629
timestamp 1649977179
transform 1 0 58972 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_641
timestamp 1649977179
transform 1 0 60076 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_653
timestamp 1649977179
transform 1 0 61180 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_665
timestamp 1649977179
transform 1 0 62284 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_671
timestamp 1649977179
transform 1 0 62836 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_673
timestamp 1649977179
transform 1 0 63020 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_685
timestamp 1649977179
transform 1 0 64124 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_697
timestamp 1649977179
transform 1 0 65228 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_709
timestamp 1649977179
transform 1 0 66332 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_721
timestamp 1649977179
transform 1 0 67436 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_727
timestamp 1649977179
transform 1 0 67988 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_729
timestamp 1649977179
transform 1 0 68172 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1649977179
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1649977179
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1649977179
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_34
timestamp 1649977179
transform 1 0 4232 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_43
timestamp 1649977179
transform 1 0 5060 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_53
timestamp 1649977179
transform 1 0 5980 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_60
timestamp 1649977179
transform 1 0 6624 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_80
timestamp 1649977179
transform 1 0 8464 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_87
timestamp 1649977179
transform 1 0 9108 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_94
timestamp 1649977179
transform 1 0 9752 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_114
timestamp 1649977179
transform 1 0 11592 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_127
timestamp 1649977179
transform 1 0 12788 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_131
timestamp 1649977179
transform 1 0 13156 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_136
timestamp 1649977179
transform 1 0 13616 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_141
timestamp 1649977179
transform 1 0 14076 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_145
timestamp 1649977179
transform 1 0 14444 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_152
timestamp 1649977179
transform 1 0 15088 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_162
timestamp 1649977179
transform 1 0 16008 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_172
timestamp 1649977179
transform 1 0 16928 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_182
timestamp 1649977179
transform 1 0 17848 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_190
timestamp 1649977179
transform 1 0 18584 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_197
timestamp 1649977179
transform 1 0 19228 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_204
timestamp 1649977179
transform 1 0 19872 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_211
timestamp 1649977179
transform 1 0 20516 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_221
timestamp 1649977179
transform 1 0 21436 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_231
timestamp 1649977179
transform 1 0 22356 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_237
timestamp 1649977179
transform 1 0 22908 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_246
timestamp 1649977179
transform 1 0 23736 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_4_255
timestamp 1649977179
transform 1 0 24564 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_267
timestamp 1649977179
transform 1 0 25668 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_279
timestamp 1649977179
transform 1 0 26772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_291
timestamp 1649977179
transform 1 0 27876 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_303
timestamp 1649977179
transform 1 0 28980 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1649977179
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1649977179
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1649977179
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1649977179
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1649977179
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1649977179
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1649977179
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1649977179
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1649977179
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_389
timestamp 1649977179
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_401
timestamp 1649977179
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp 1649977179
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1649977179
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_421
timestamp 1649977179
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_433
timestamp 1649977179
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_445
timestamp 1649977179
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_457
timestamp 1649977179
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_469
timestamp 1649977179
transform 1 0 44252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 1649977179
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_477
timestamp 1649977179
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_489
timestamp 1649977179
transform 1 0 46092 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_501
timestamp 1649977179
transform 1 0 47196 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_513
timestamp 1649977179
transform 1 0 48300 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_525
timestamp 1649977179
transform 1 0 49404 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_531
timestamp 1649977179
transform 1 0 49956 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_533
timestamp 1649977179
transform 1 0 50140 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_545
timestamp 1649977179
transform 1 0 51244 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_557
timestamp 1649977179
transform 1 0 52348 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_569
timestamp 1649977179
transform 1 0 53452 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_581
timestamp 1649977179
transform 1 0 54556 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_587
timestamp 1649977179
transform 1 0 55108 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_589
timestamp 1649977179
transform 1 0 55292 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_601
timestamp 1649977179
transform 1 0 56396 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_613
timestamp 1649977179
transform 1 0 57500 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_625
timestamp 1649977179
transform 1 0 58604 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_637
timestamp 1649977179
transform 1 0 59708 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_643
timestamp 1649977179
transform 1 0 60260 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_645
timestamp 1649977179
transform 1 0 60444 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_657
timestamp 1649977179
transform 1 0 61548 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_669
timestamp 1649977179
transform 1 0 62652 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_681
timestamp 1649977179
transform 1 0 63756 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_693
timestamp 1649977179
transform 1 0 64860 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_699
timestamp 1649977179
transform 1 0 65412 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_701
timestamp 1649977179
transform 1 0 65596 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_713
timestamp 1649977179
transform 1 0 66700 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_725
timestamp 1649977179
transform 1 0 67804 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1649977179
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_15
timestamp 1649977179
transform 1 0 2484 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_23
timestamp 1649977179
transform 1 0 3220 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_31
timestamp 1649977179
transform 1 0 3956 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_35
timestamp 1649977179
transform 1 0 4324 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_38
timestamp 1649977179
transform 1 0 4600 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_52
timestamp 1649977179
transform 1 0 5888 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_65
timestamp 1649977179
transform 1 0 7084 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_93
timestamp 1649977179
transform 1 0 9660 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_103
timestamp 1649977179
transform 1 0 10580 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1649977179
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_113
timestamp 1649977179
transform 1 0 11500 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_120
timestamp 1649977179
transform 1 0 12144 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_132
timestamp 1649977179
transform 1 0 13248 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_146
timestamp 1649977179
transform 1 0 14536 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_5_160
timestamp 1649977179
transform 1 0 15824 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_5_185
timestamp 1649977179
transform 1 0 18124 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_193
timestamp 1649977179
transform 1 0 18860 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_197
timestamp 1649977179
transform 1 0 19228 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_207
timestamp 1649977179
transform 1 0 20148 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1649977179
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1649977179
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_228
timestamp 1649977179
transform 1 0 22080 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_235
timestamp 1649977179
transform 1 0 22724 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_249
timestamp 1649977179
transform 1 0 24012 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_255
timestamp 1649977179
transform 1 0 24564 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_267
timestamp 1649977179
transform 1 0 25668 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1649977179
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1649977179
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_293
timestamp 1649977179
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_305
timestamp 1649977179
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_317
timestamp 1649977179
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1649977179
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1649977179
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1649977179
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1649977179
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1649977179
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1649977179
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1649977179
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1649977179
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_393
timestamp 1649977179
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_405
timestamp 1649977179
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_417
timestamp 1649977179
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_429
timestamp 1649977179
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_441
timestamp 1649977179
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1649977179
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_449
timestamp 1649977179
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_461
timestamp 1649977179
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_473
timestamp 1649977179
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_485
timestamp 1649977179
transform 1 0 45724 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_497
timestamp 1649977179
transform 1 0 46828 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_503
timestamp 1649977179
transform 1 0 47380 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_505
timestamp 1649977179
transform 1 0 47564 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_517
timestamp 1649977179
transform 1 0 48668 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_529
timestamp 1649977179
transform 1 0 49772 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_541
timestamp 1649977179
transform 1 0 50876 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_553
timestamp 1649977179
transform 1 0 51980 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_559
timestamp 1649977179
transform 1 0 52532 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_561
timestamp 1649977179
transform 1 0 52716 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_573
timestamp 1649977179
transform 1 0 53820 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_585
timestamp 1649977179
transform 1 0 54924 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_597
timestamp 1649977179
transform 1 0 56028 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_609
timestamp 1649977179
transform 1 0 57132 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_615
timestamp 1649977179
transform 1 0 57684 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_617
timestamp 1649977179
transform 1 0 57868 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_629
timestamp 1649977179
transform 1 0 58972 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_641
timestamp 1649977179
transform 1 0 60076 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_653
timestamp 1649977179
transform 1 0 61180 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_665
timestamp 1649977179
transform 1 0 62284 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_671
timestamp 1649977179
transform 1 0 62836 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_673
timestamp 1649977179
transform 1 0 63020 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_685
timestamp 1649977179
transform 1 0 64124 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_697
timestamp 1649977179
transform 1 0 65228 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_709
timestamp 1649977179
transform 1 0 66332 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_721
timestamp 1649977179
transform 1 0 67436 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_727
timestamp 1649977179
transform 1 0 67988 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_729
timestamp 1649977179
transform 1 0 68172 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1649977179
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1649977179
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1649977179
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_34
timestamp 1649977179
transform 1 0 4232 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_42
timestamp 1649977179
transform 1 0 4968 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_51
timestamp 1649977179
transform 1 0 5796 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_63
timestamp 1649977179
transform 1 0 6900 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_71
timestamp 1649977179
transform 1 0 7636 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_75
timestamp 1649977179
transform 1 0 8004 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1649977179
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_87
timestamp 1649977179
transform 1 0 9108 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_94
timestamp 1649977179
transform 1 0 9752 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_101
timestamp 1649977179
transform 1 0 10396 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_121
timestamp 1649977179
transform 1 0 12236 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_127
timestamp 1649977179
transform 1 0 12788 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_135
timestamp 1649977179
transform 1 0 13524 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1649977179
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_141
timestamp 1649977179
transform 1 0 14076 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_145
timestamp 1649977179
transform 1 0 14444 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_154
timestamp 1649977179
transform 1 0 15272 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_178
timestamp 1649977179
transform 1 0 17480 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_185
timestamp 1649977179
transform 1 0 18124 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_192
timestamp 1649977179
transform 1 0 18768 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_213
timestamp 1649977179
transform 1 0 20700 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_222
timestamp 1649977179
transform 1 0 21528 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_236
timestamp 1649977179
transform 1 0 22816 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_242
timestamp 1649977179
transform 1 0 23368 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_248
timestamp 1649977179
transform 1 0 23920 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1649977179
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1649977179
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_277
timestamp 1649977179
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_289
timestamp 1649977179
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1649977179
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1649977179
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1649977179
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1649977179
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1649977179
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1649977179
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1649977179
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1649977179
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1649977179
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1649977179
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_389
timestamp 1649977179
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_401
timestamp 1649977179
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 1649977179
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1649977179
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_421
timestamp 1649977179
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_433
timestamp 1649977179
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_445
timestamp 1649977179
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_457
timestamp 1649977179
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_469
timestamp 1649977179
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 1649977179
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_477
timestamp 1649977179
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_489
timestamp 1649977179
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_501
timestamp 1649977179
transform 1 0 47196 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_513
timestamp 1649977179
transform 1 0 48300 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_525
timestamp 1649977179
transform 1 0 49404 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_531
timestamp 1649977179
transform 1 0 49956 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_533
timestamp 1649977179
transform 1 0 50140 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_545
timestamp 1649977179
transform 1 0 51244 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_557
timestamp 1649977179
transform 1 0 52348 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_569
timestamp 1649977179
transform 1 0 53452 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_581
timestamp 1649977179
transform 1 0 54556 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_587
timestamp 1649977179
transform 1 0 55108 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_589
timestamp 1649977179
transform 1 0 55292 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_601
timestamp 1649977179
transform 1 0 56396 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_613
timestamp 1649977179
transform 1 0 57500 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_625
timestamp 1649977179
transform 1 0 58604 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_637
timestamp 1649977179
transform 1 0 59708 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_643
timestamp 1649977179
transform 1 0 60260 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_645
timestamp 1649977179
transform 1 0 60444 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_657
timestamp 1649977179
transform 1 0 61548 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_669
timestamp 1649977179
transform 1 0 62652 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_681
timestamp 1649977179
transform 1 0 63756 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_693
timestamp 1649977179
transform 1 0 64860 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_699
timestamp 1649977179
transform 1 0 65412 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_701
timestamp 1649977179
transform 1 0 65596 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_713
timestamp 1649977179
transform 1 0 66700 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_725
timestamp 1649977179
transform 1 0 67804 0 1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1649977179
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_15
timestamp 1649977179
transform 1 0 2484 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_20
timestamp 1649977179
transform 1 0 2944 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_27
timestamp 1649977179
transform 1 0 3588 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_36
timestamp 1649977179
transform 1 0 4416 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_42
timestamp 1649977179
transform 1 0 4968 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_52
timestamp 1649977179
transform 1 0 5888 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_57
timestamp 1649977179
transform 1 0 6348 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_61
timestamp 1649977179
transform 1 0 6716 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_67
timestamp 1649977179
transform 1 0 7268 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_73
timestamp 1649977179
transform 1 0 7820 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_79
timestamp 1649977179
transform 1 0 8372 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_85
timestamp 1649977179
transform 1 0 8924 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_92
timestamp 1649977179
transform 1 0 9568 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_106
timestamp 1649977179
transform 1 0 10856 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_113
timestamp 1649977179
transform 1 0 11500 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_117
timestamp 1649977179
transform 1 0 11868 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_124
timestamp 1649977179
transform 1 0 12512 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_144
timestamp 1649977179
transform 1 0 14352 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_150
timestamp 1649977179
transform 1 0 14904 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_156
timestamp 1649977179
transform 1 0 15456 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_160
timestamp 1649977179
transform 1 0 15824 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_164
timestamp 1649977179
transform 1 0 16192 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_169
timestamp 1649977179
transform 1 0 16652 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_174
timestamp 1649977179
transform 1 0 17112 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_181
timestamp 1649977179
transform 1 0 17756 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_201
timestamp 1649977179
transform 1 0 19596 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_213
timestamp 1649977179
transform 1 0 20700 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_220
timestamp 1649977179
transform 1 0 21344 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_233
timestamp 1649977179
transform 1 0 22540 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_247
timestamp 1649977179
transform 1 0 23828 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_259
timestamp 1649977179
transform 1 0 24932 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_271
timestamp 1649977179
transform 1 0 26036 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1649977179
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1649977179
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1649977179
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1649977179
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_317
timestamp 1649977179
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1649977179
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1649977179
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1649977179
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1649977179
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1649977179
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1649977179
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1649977179
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1649977179
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_393
timestamp 1649977179
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_405
timestamp 1649977179
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_417
timestamp 1649977179
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_429
timestamp 1649977179
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_441
timestamp 1649977179
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1649977179
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_449
timestamp 1649977179
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_461
timestamp 1649977179
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_473
timestamp 1649977179
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_485
timestamp 1649977179
transform 1 0 45724 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_497
timestamp 1649977179
transform 1 0 46828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_503
timestamp 1649977179
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_505
timestamp 1649977179
transform 1 0 47564 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_517
timestamp 1649977179
transform 1 0 48668 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_529
timestamp 1649977179
transform 1 0 49772 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_541
timestamp 1649977179
transform 1 0 50876 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_553
timestamp 1649977179
transform 1 0 51980 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_559
timestamp 1649977179
transform 1 0 52532 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_561
timestamp 1649977179
transform 1 0 52716 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_573
timestamp 1649977179
transform 1 0 53820 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_585
timestamp 1649977179
transform 1 0 54924 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_597
timestamp 1649977179
transform 1 0 56028 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_609
timestamp 1649977179
transform 1 0 57132 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_615
timestamp 1649977179
transform 1 0 57684 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_617
timestamp 1649977179
transform 1 0 57868 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_629
timestamp 1649977179
transform 1 0 58972 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_641
timestamp 1649977179
transform 1 0 60076 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_653
timestamp 1649977179
transform 1 0 61180 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_665
timestamp 1649977179
transform 1 0 62284 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_671
timestamp 1649977179
transform 1 0 62836 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_673
timestamp 1649977179
transform 1 0 63020 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_685
timestamp 1649977179
transform 1 0 64124 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_697
timestamp 1649977179
transform 1 0 65228 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_709
timestamp 1649977179
transform 1 0 66332 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_721
timestamp 1649977179
transform 1 0 67436 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_727
timestamp 1649977179
transform 1 0 67988 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_729
timestamp 1649977179
transform 1 0 68172 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1649977179
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1649977179
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1649977179
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_39
timestamp 1649977179
transform 1 0 4692 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_45
timestamp 1649977179
transform 1 0 5244 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_48
timestamp 1649977179
transform 1 0 5520 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_60
timestamp 1649977179
transform 1 0 6624 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_80
timestamp 1649977179
transform 1 0 8464 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_8_85
timestamp 1649977179
transform 1 0 8924 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_94
timestamp 1649977179
transform 1 0 9752 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_101
timestamp 1649977179
transform 1 0 10396 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_108
timestamp 1649977179
transform 1 0 11040 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_115
timestamp 1649977179
transform 1 0 11684 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_122
timestamp 1649977179
transform 1 0 12328 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_129
timestamp 1649977179
transform 1 0 12972 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_136
timestamp 1649977179
transform 1 0 13616 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_143
timestamp 1649977179
transform 1 0 14260 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_152
timestamp 1649977179
transform 1 0 15088 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_159
timestamp 1649977179
transform 1 0 15732 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_179
timestamp 1649977179
transform 1 0 17572 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_185
timestamp 1649977179
transform 1 0 18124 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_192
timestamp 1649977179
transform 1 0 18768 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_200
timestamp 1649977179
transform 1 0 19504 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_212
timestamp 1649977179
transform 1 0 20608 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_224
timestamp 1649977179
transform 1 0 21712 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_230
timestamp 1649977179
transform 1 0 22264 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_238
timestamp 1649977179
transform 1 0 23000 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_247
timestamp 1649977179
transform 1 0 23828 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1649977179
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_258
timestamp 1649977179
transform 1 0 24840 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_270
timestamp 1649977179
transform 1 0 25944 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_282
timestamp 1649977179
transform 1 0 27048 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_294
timestamp 1649977179
transform 1 0 28152 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_306
timestamp 1649977179
transform 1 0 29256 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1649977179
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1649977179
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1649977179
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_345
timestamp 1649977179
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1649977179
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1649977179
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1649977179
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1649977179
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_389
timestamp 1649977179
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_401
timestamp 1649977179
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 1649977179
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1649977179
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_421
timestamp 1649977179
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_433
timestamp 1649977179
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_445
timestamp 1649977179
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_457
timestamp 1649977179
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 1649977179
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1649977179
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_477
timestamp 1649977179
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_489
timestamp 1649977179
transform 1 0 46092 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_501
timestamp 1649977179
transform 1 0 47196 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_513
timestamp 1649977179
transform 1 0 48300 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_525
timestamp 1649977179
transform 1 0 49404 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_531
timestamp 1649977179
transform 1 0 49956 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_533
timestamp 1649977179
transform 1 0 50140 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_545
timestamp 1649977179
transform 1 0 51244 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_557
timestamp 1649977179
transform 1 0 52348 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_569
timestamp 1649977179
transform 1 0 53452 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_581
timestamp 1649977179
transform 1 0 54556 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_587
timestamp 1649977179
transform 1 0 55108 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_589
timestamp 1649977179
transform 1 0 55292 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_601
timestamp 1649977179
transform 1 0 56396 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_613
timestamp 1649977179
transform 1 0 57500 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_625
timestamp 1649977179
transform 1 0 58604 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_637
timestamp 1649977179
transform 1 0 59708 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_643
timestamp 1649977179
transform 1 0 60260 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_645
timestamp 1649977179
transform 1 0 60444 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_657
timestamp 1649977179
transform 1 0 61548 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_669
timestamp 1649977179
transform 1 0 62652 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_681
timestamp 1649977179
transform 1 0 63756 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_693
timestamp 1649977179
transform 1 0 64860 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_699
timestamp 1649977179
transform 1 0 65412 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_701
timestamp 1649977179
transform 1 0 65596 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_713
timestamp 1649977179
transform 1 0 66700 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_725
timestamp 1649977179
transform 1 0 67804 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1649977179
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1649977179
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_27
timestamp 1649977179
transform 1 0 3588 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_31
timestamp 1649977179
transform 1 0 3956 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_35
timestamp 1649977179
transform 1 0 4324 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_45
timestamp 1649977179
transform 1 0 5244 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_52
timestamp 1649977179
transform 1 0 5888 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_63
timestamp 1649977179
transform 1 0 6900 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_69
timestamp 1649977179
transform 1 0 7452 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_93
timestamp 1649977179
transform 1 0 9660 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1649977179
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1649977179
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_113
timestamp 1649977179
transform 1 0 11500 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_117
timestamp 1649977179
transform 1 0 11868 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_129
timestamp 1649977179
transform 1 0 12972 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_153
timestamp 1649977179
transform 1 0 15180 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_164
timestamp 1649977179
transform 1 0 16192 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_177
timestamp 1649977179
transform 1 0 17388 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_201
timestamp 1649977179
transform 1 0 19596 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_205
timestamp 1649977179
transform 1 0 19964 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_208
timestamp 1649977179
transform 1 0 20240 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1649977179
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1649977179
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_228
timestamp 1649977179
transform 1 0 22080 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_237
timestamp 1649977179
transform 1 0 22908 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_246
timestamp 1649977179
transform 1 0 23736 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_258
timestamp 1649977179
transform 1 0 24840 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_270
timestamp 1649977179
transform 1 0 25944 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_278
timestamp 1649977179
transform 1 0 26680 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1649977179
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1649977179
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_305
timestamp 1649977179
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_317
timestamp 1649977179
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1649977179
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1649977179
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1649977179
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_349
timestamp 1649977179
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_361
timestamp 1649977179
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_373
timestamp 1649977179
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1649977179
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1649977179
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_393
timestamp 1649977179
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_405
timestamp 1649977179
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_417
timestamp 1649977179
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_429
timestamp 1649977179
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_441
timestamp 1649977179
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 1649977179
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_449
timestamp 1649977179
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_461
timestamp 1649977179
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_473
timestamp 1649977179
transform 1 0 44620 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_485
timestamp 1649977179
transform 1 0 45724 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_497
timestamp 1649977179
transform 1 0 46828 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_503
timestamp 1649977179
transform 1 0 47380 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_505
timestamp 1649977179
transform 1 0 47564 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_517
timestamp 1649977179
transform 1 0 48668 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_529
timestamp 1649977179
transform 1 0 49772 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_541
timestamp 1649977179
transform 1 0 50876 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_553
timestamp 1649977179
transform 1 0 51980 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_559
timestamp 1649977179
transform 1 0 52532 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_561
timestamp 1649977179
transform 1 0 52716 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_573
timestamp 1649977179
transform 1 0 53820 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_585
timestamp 1649977179
transform 1 0 54924 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_597
timestamp 1649977179
transform 1 0 56028 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_609
timestamp 1649977179
transform 1 0 57132 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_615
timestamp 1649977179
transform 1 0 57684 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_617
timestamp 1649977179
transform 1 0 57868 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_629
timestamp 1649977179
transform 1 0 58972 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_641
timestamp 1649977179
transform 1 0 60076 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_653
timestamp 1649977179
transform 1 0 61180 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_665
timestamp 1649977179
transform 1 0 62284 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_671
timestamp 1649977179
transform 1 0 62836 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_673
timestamp 1649977179
transform 1 0 63020 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_685
timestamp 1649977179
transform 1 0 64124 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_697
timestamp 1649977179
transform 1 0 65228 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_709
timestamp 1649977179
transform 1 0 66332 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_721
timestamp 1649977179
transform 1 0 67436 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_727
timestamp 1649977179
transform 1 0 67988 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_729
timestamp 1649977179
transform 1 0 68172 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1649977179
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1649977179
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1649977179
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_29
timestamp 1649977179
transform 1 0 3772 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_37
timestamp 1649977179
transform 1 0 4508 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_43
timestamp 1649977179
transform 1 0 5060 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_55
timestamp 1649977179
transform 1 0 6164 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_63
timestamp 1649977179
transform 1 0 6900 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_80
timestamp 1649977179
transform 1 0 8464 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_10_85
timestamp 1649977179
transform 1 0 8924 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_94
timestamp 1649977179
transform 1 0 9752 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_104
timestamp 1649977179
transform 1 0 10672 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_114
timestamp 1649977179
transform 1 0 11592 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_124
timestamp 1649977179
transform 1 0 12512 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_136
timestamp 1649977179
transform 1 0 13616 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_10_141
timestamp 1649977179
transform 1 0 14076 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_147
timestamp 1649977179
transform 1 0 14628 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_154
timestamp 1649977179
transform 1 0 15272 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_178
timestamp 1649977179
transform 1 0 17480 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_185
timestamp 1649977179
transform 1 0 18124 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_189
timestamp 1649977179
transform 1 0 18492 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_192
timestamp 1649977179
transform 1 0 18768 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_213
timestamp 1649977179
transform 1 0 20700 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_226
timestamp 1649977179
transform 1 0 21896 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_242
timestamp 1649977179
transform 1 0 23368 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_250
timestamp 1649977179
transform 1 0 24104 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_256
timestamp 1649977179
transform 1 0 24656 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_262
timestamp 1649977179
transform 1 0 25208 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_274
timestamp 1649977179
transform 1 0 26312 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_286
timestamp 1649977179
transform 1 0 27416 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_298
timestamp 1649977179
transform 1 0 28520 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_306
timestamp 1649977179
transform 1 0 29256 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_309
timestamp 1649977179
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_321
timestamp 1649977179
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_333
timestamp 1649977179
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_345
timestamp 1649977179
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1649977179
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1649977179
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_365
timestamp 1649977179
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_377
timestamp 1649977179
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_389
timestamp 1649977179
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_401
timestamp 1649977179
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_413
timestamp 1649977179
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_419
timestamp 1649977179
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_421
timestamp 1649977179
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_433
timestamp 1649977179
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_445
timestamp 1649977179
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_457
timestamp 1649977179
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_469
timestamp 1649977179
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp 1649977179
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_477
timestamp 1649977179
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_489
timestamp 1649977179
transform 1 0 46092 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_501
timestamp 1649977179
transform 1 0 47196 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_513
timestamp 1649977179
transform 1 0 48300 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_525
timestamp 1649977179
transform 1 0 49404 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_531
timestamp 1649977179
transform 1 0 49956 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_533
timestamp 1649977179
transform 1 0 50140 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_545
timestamp 1649977179
transform 1 0 51244 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_557
timestamp 1649977179
transform 1 0 52348 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_569
timestamp 1649977179
transform 1 0 53452 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_581
timestamp 1649977179
transform 1 0 54556 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_587
timestamp 1649977179
transform 1 0 55108 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_589
timestamp 1649977179
transform 1 0 55292 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_601
timestamp 1649977179
transform 1 0 56396 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_613
timestamp 1649977179
transform 1 0 57500 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_625
timestamp 1649977179
transform 1 0 58604 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_637
timestamp 1649977179
transform 1 0 59708 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_643
timestamp 1649977179
transform 1 0 60260 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_645
timestamp 1649977179
transform 1 0 60444 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_657
timestamp 1649977179
transform 1 0 61548 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_669
timestamp 1649977179
transform 1 0 62652 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_681
timestamp 1649977179
transform 1 0 63756 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_693
timestamp 1649977179
transform 1 0 64860 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_699
timestamp 1649977179
transform 1 0 65412 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_701
timestamp 1649977179
transform 1 0 65596 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_713
timestamp 1649977179
transform 1 0 66700 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_725
timestamp 1649977179
transform 1 0 67804 0 1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1649977179
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1649977179
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_27
timestamp 1649977179
transform 1 0 3588 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_33
timestamp 1649977179
transform 1 0 4140 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_44
timestamp 1649977179
transform 1 0 5152 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1649977179
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1649977179
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_65
timestamp 1649977179
transform 1 0 7084 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_73
timestamp 1649977179
transform 1 0 7820 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_81
timestamp 1649977179
transform 1 0 8556 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_87
timestamp 1649977179
transform 1 0 9108 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_94
timestamp 1649977179
transform 1 0 9752 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_106
timestamp 1649977179
transform 1 0 10856 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_113
timestamp 1649977179
transform 1 0 11500 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_120
timestamp 1649977179
transform 1 0 12144 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_132
timestamp 1649977179
transform 1 0 13248 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_139
timestamp 1649977179
transform 1 0 13892 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_159
timestamp 1649977179
transform 1 0 15732 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1649977179
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_179
timestamp 1649977179
transform 1 0 17572 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_201
timestamp 1649977179
transform 1 0 19596 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_211
timestamp 1649977179
transform 1 0 20516 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_217
timestamp 1649977179
transform 1 0 21068 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_220
timestamp 1649977179
transform 1 0 21344 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_235
timestamp 1649977179
transform 1 0 22724 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_239
timestamp 1649977179
transform 1 0 23092 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_248
timestamp 1649977179
transform 1 0 23920 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_254
timestamp 1649977179
transform 1 0 24472 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_266
timestamp 1649977179
transform 1 0 25576 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_278
timestamp 1649977179
transform 1 0 26680 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1649977179
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_293
timestamp 1649977179
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_305
timestamp 1649977179
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_317
timestamp 1649977179
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1649977179
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1649977179
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_337
timestamp 1649977179
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_349
timestamp 1649977179
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_361
timestamp 1649977179
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_373
timestamp 1649977179
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1649977179
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1649977179
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_393
timestamp 1649977179
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_405
timestamp 1649977179
transform 1 0 38364 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_417
timestamp 1649977179
transform 1 0 39468 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_429
timestamp 1649977179
transform 1 0 40572 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_441
timestamp 1649977179
transform 1 0 41676 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 1649977179
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_449
timestamp 1649977179
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_461
timestamp 1649977179
transform 1 0 43516 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_473
timestamp 1649977179
transform 1 0 44620 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_485
timestamp 1649977179
transform 1 0 45724 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_497
timestamp 1649977179
transform 1 0 46828 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_503
timestamp 1649977179
transform 1 0 47380 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_505
timestamp 1649977179
transform 1 0 47564 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_517
timestamp 1649977179
transform 1 0 48668 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_529
timestamp 1649977179
transform 1 0 49772 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_541
timestamp 1649977179
transform 1 0 50876 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_553
timestamp 1649977179
transform 1 0 51980 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_559
timestamp 1649977179
transform 1 0 52532 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_561
timestamp 1649977179
transform 1 0 52716 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_573
timestamp 1649977179
transform 1 0 53820 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_585
timestamp 1649977179
transform 1 0 54924 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_597
timestamp 1649977179
transform 1 0 56028 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_609
timestamp 1649977179
transform 1 0 57132 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_615
timestamp 1649977179
transform 1 0 57684 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_617
timestamp 1649977179
transform 1 0 57868 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_629
timestamp 1649977179
transform 1 0 58972 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_641
timestamp 1649977179
transform 1 0 60076 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_653
timestamp 1649977179
transform 1 0 61180 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_665
timestamp 1649977179
transform 1 0 62284 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_671
timestamp 1649977179
transform 1 0 62836 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_673
timestamp 1649977179
transform 1 0 63020 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_685
timestamp 1649977179
transform 1 0 64124 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_697
timestamp 1649977179
transform 1 0 65228 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_709
timestamp 1649977179
transform 1 0 66332 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_721
timestamp 1649977179
transform 1 0 67436 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_727
timestamp 1649977179
transform 1 0 67988 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_729
timestamp 1649977179
transform 1 0 68172 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1649977179
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_15
timestamp 1649977179
transform 1 0 2484 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_24
timestamp 1649977179
transform 1 0 3312 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_31
timestamp 1649977179
transform 1 0 3956 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_35
timestamp 1649977179
transform 1 0 4324 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_46
timestamp 1649977179
transform 1 0 5336 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_60
timestamp 1649977179
transform 1 0 6624 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_80
timestamp 1649977179
transform 1 0 8464 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_85
timestamp 1649977179
transform 1 0 8924 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_89
timestamp 1649977179
transform 1 0 9292 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_93
timestamp 1649977179
transform 1 0 9660 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_99
timestamp 1649977179
transform 1 0 10212 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_116
timestamp 1649977179
transform 1 0 11776 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_122
timestamp 1649977179
transform 1 0 12328 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_136
timestamp 1649977179
transform 1 0 13616 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_157
timestamp 1649977179
transform 1 0 15548 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_177
timestamp 1649977179
transform 1 0 17388 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_183
timestamp 1649977179
transform 1 0 17940 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1649977179
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1649977179
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_199
timestamp 1649977179
transform 1 0 19412 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_207
timestamp 1649977179
transform 1 0 20148 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_216
timestamp 1649977179
transform 1 0 20976 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_230
timestamp 1649977179
transform 1 0 22264 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_234
timestamp 1649977179
transform 1 0 22632 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_243
timestamp 1649977179
transform 1 0 23460 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1649977179
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_253
timestamp 1649977179
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_265
timestamp 1649977179
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_277
timestamp 1649977179
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_289
timestamp 1649977179
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1649977179
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1649977179
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_309
timestamp 1649977179
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_321
timestamp 1649977179
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_333
timestamp 1649977179
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_345
timestamp 1649977179
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1649977179
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1649977179
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_365
timestamp 1649977179
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_377
timestamp 1649977179
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_389
timestamp 1649977179
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_401
timestamp 1649977179
transform 1 0 37996 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_413
timestamp 1649977179
transform 1 0 39100 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_419
timestamp 1649977179
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_421
timestamp 1649977179
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_433
timestamp 1649977179
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_445
timestamp 1649977179
transform 1 0 42044 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_457
timestamp 1649977179
transform 1 0 43148 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_469
timestamp 1649977179
transform 1 0 44252 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 1649977179
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_477
timestamp 1649977179
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_489
timestamp 1649977179
transform 1 0 46092 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_501
timestamp 1649977179
transform 1 0 47196 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_513
timestamp 1649977179
transform 1 0 48300 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_525
timestamp 1649977179
transform 1 0 49404 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_531
timestamp 1649977179
transform 1 0 49956 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_533
timestamp 1649977179
transform 1 0 50140 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_545
timestamp 1649977179
transform 1 0 51244 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_557
timestamp 1649977179
transform 1 0 52348 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_569
timestamp 1649977179
transform 1 0 53452 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_581
timestamp 1649977179
transform 1 0 54556 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_587
timestamp 1649977179
transform 1 0 55108 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_589
timestamp 1649977179
transform 1 0 55292 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_601
timestamp 1649977179
transform 1 0 56396 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_613
timestamp 1649977179
transform 1 0 57500 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_625
timestamp 1649977179
transform 1 0 58604 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_637
timestamp 1649977179
transform 1 0 59708 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_643
timestamp 1649977179
transform 1 0 60260 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_645
timestamp 1649977179
transform 1 0 60444 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_657
timestamp 1649977179
transform 1 0 61548 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_669
timestamp 1649977179
transform 1 0 62652 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_681
timestamp 1649977179
transform 1 0 63756 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_693
timestamp 1649977179
transform 1 0 64860 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_699
timestamp 1649977179
transform 1 0 65412 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_701
timestamp 1649977179
transform 1 0 65596 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_713
timestamp 1649977179
transform 1 0 66700 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_725
timestamp 1649977179
transform 1 0 67804 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1649977179
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_15
timestamp 1649977179
transform 1 0 2484 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_23
timestamp 1649977179
transform 1 0 3220 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_27
timestamp 1649977179
transform 1 0 3588 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_41
timestamp 1649977179
transform 1 0 4876 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_48
timestamp 1649977179
transform 1 0 5520 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_63
timestamp 1649977179
transform 1 0 6900 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_69
timestamp 1649977179
transform 1 0 7452 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_75
timestamp 1649977179
transform 1 0 8004 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_83
timestamp 1649977179
transform 1 0 8740 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_87
timestamp 1649977179
transform 1 0 9108 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_90
timestamp 1649977179
transform 1 0 9384 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_102
timestamp 1649977179
transform 1 0 10488 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_108
timestamp 1649977179
transform 1 0 11040 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_113
timestamp 1649977179
transform 1 0 11500 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_117
timestamp 1649977179
transform 1 0 11868 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_128
timestamp 1649977179
transform 1 0 12880 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_13_136
timestamp 1649977179
transform 1 0 13616 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_144
timestamp 1649977179
transform 1 0 14352 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_147
timestamp 1649977179
transform 1 0 14628 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1649977179
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1649977179
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_179
timestamp 1649977179
transform 1 0 17572 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_185
timestamp 1649977179
transform 1 0 18124 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_191
timestamp 1649977179
transform 1 0 18676 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_203
timestamp 1649977179
transform 1 0 19780 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_213
timestamp 1649977179
transform 1 0 20700 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_220
timestamp 1649977179
transform 1 0 21344 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_228
timestamp 1649977179
transform 1 0 22080 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_234
timestamp 1649977179
transform 1 0 22632 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_243
timestamp 1649977179
transform 1 0 23460 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_255
timestamp 1649977179
transform 1 0 24564 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_267
timestamp 1649977179
transform 1 0 25668 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1649977179
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_281
timestamp 1649977179
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_293
timestamp 1649977179
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_305
timestamp 1649977179
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_317
timestamp 1649977179
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1649977179
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1649977179
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_337
timestamp 1649977179
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_349
timestamp 1649977179
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_361
timestamp 1649977179
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_373
timestamp 1649977179
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1649977179
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1649977179
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_393
timestamp 1649977179
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_405
timestamp 1649977179
transform 1 0 38364 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_417
timestamp 1649977179
transform 1 0 39468 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_429
timestamp 1649977179
transform 1 0 40572 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_441
timestamp 1649977179
transform 1 0 41676 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_447
timestamp 1649977179
transform 1 0 42228 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_449
timestamp 1649977179
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_461
timestamp 1649977179
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_473
timestamp 1649977179
transform 1 0 44620 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_485
timestamp 1649977179
transform 1 0 45724 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_497
timestamp 1649977179
transform 1 0 46828 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_503
timestamp 1649977179
transform 1 0 47380 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_505
timestamp 1649977179
transform 1 0 47564 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_517
timestamp 1649977179
transform 1 0 48668 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_529
timestamp 1649977179
transform 1 0 49772 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_541
timestamp 1649977179
transform 1 0 50876 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_553
timestamp 1649977179
transform 1 0 51980 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_559
timestamp 1649977179
transform 1 0 52532 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_561
timestamp 1649977179
transform 1 0 52716 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_573
timestamp 1649977179
transform 1 0 53820 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_585
timestamp 1649977179
transform 1 0 54924 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_597
timestamp 1649977179
transform 1 0 56028 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_609
timestamp 1649977179
transform 1 0 57132 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_615
timestamp 1649977179
transform 1 0 57684 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_617
timestamp 1649977179
transform 1 0 57868 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_629
timestamp 1649977179
transform 1 0 58972 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_641
timestamp 1649977179
transform 1 0 60076 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_653
timestamp 1649977179
transform 1 0 61180 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_665
timestamp 1649977179
transform 1 0 62284 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_671
timestamp 1649977179
transform 1 0 62836 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_673
timestamp 1649977179
transform 1 0 63020 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_685
timestamp 1649977179
transform 1 0 64124 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_697
timestamp 1649977179
transform 1 0 65228 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_709
timestamp 1649977179
transform 1 0 66332 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_721
timestamp 1649977179
transform 1 0 67436 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_727
timestamp 1649977179
transform 1 0 67988 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_729
timestamp 1649977179
transform 1 0 68172 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1649977179
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_15
timestamp 1649977179
transform 1 0 2484 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_21
timestamp 1649977179
transform 1 0 3036 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_24
timestamp 1649977179
transform 1 0 3312 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_29
timestamp 1649977179
transform 1 0 3772 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_36
timestamp 1649977179
transform 1 0 4416 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_48
timestamp 1649977179
transform 1 0 5520 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_60
timestamp 1649977179
transform 1 0 6624 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_80
timestamp 1649977179
transform 1 0 8464 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1649977179
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_97
timestamp 1649977179
transform 1 0 10028 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_105
timestamp 1649977179
transform 1 0 10764 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_14_110
timestamp 1649977179
transform 1 0 11224 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_116
timestamp 1649977179
transform 1 0 11776 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_119
timestamp 1649977179
transform 1 0 12052 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_127
timestamp 1649977179
transform 1 0 12788 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_131
timestamp 1649977179
transform 1 0 13156 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1649977179
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_143
timestamp 1649977179
transform 1 0 14260 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_149
timestamp 1649977179
transform 1 0 14812 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_171
timestamp 1649977179
transform 1 0 16836 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_175
timestamp 1649977179
transform 1 0 17204 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_192
timestamp 1649977179
transform 1 0 18768 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_197
timestamp 1649977179
transform 1 0 19228 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_205
timestamp 1649977179
transform 1 0 19964 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_215
timestamp 1649977179
transform 1 0 20884 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_225
timestamp 1649977179
transform 1 0 21804 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_233
timestamp 1649977179
transform 1 0 22540 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_239
timestamp 1649977179
transform 1 0 23092 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_248
timestamp 1649977179
transform 1 0 23920 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_253
timestamp 1649977179
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_265
timestamp 1649977179
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_277
timestamp 1649977179
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_289
timestamp 1649977179
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_301
timestamp 1649977179
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1649977179
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_309
timestamp 1649977179
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_321
timestamp 1649977179
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_333
timestamp 1649977179
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_345
timestamp 1649977179
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1649977179
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1649977179
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_365
timestamp 1649977179
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_377
timestamp 1649977179
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_389
timestamp 1649977179
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_401
timestamp 1649977179
transform 1 0 37996 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_413
timestamp 1649977179
transform 1 0 39100 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_419
timestamp 1649977179
transform 1 0 39652 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_421
timestamp 1649977179
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_433
timestamp 1649977179
transform 1 0 40940 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_445
timestamp 1649977179
transform 1 0 42044 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_457
timestamp 1649977179
transform 1 0 43148 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_469
timestamp 1649977179
transform 1 0 44252 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_475
timestamp 1649977179
transform 1 0 44804 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_477
timestamp 1649977179
transform 1 0 44988 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_489
timestamp 1649977179
transform 1 0 46092 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_501
timestamp 1649977179
transform 1 0 47196 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_513
timestamp 1649977179
transform 1 0 48300 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_525
timestamp 1649977179
transform 1 0 49404 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_531
timestamp 1649977179
transform 1 0 49956 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_533
timestamp 1649977179
transform 1 0 50140 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_545
timestamp 1649977179
transform 1 0 51244 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_557
timestamp 1649977179
transform 1 0 52348 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_569
timestamp 1649977179
transform 1 0 53452 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_581
timestamp 1649977179
transform 1 0 54556 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_587
timestamp 1649977179
transform 1 0 55108 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_589
timestamp 1649977179
transform 1 0 55292 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_601
timestamp 1649977179
transform 1 0 56396 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_613
timestamp 1649977179
transform 1 0 57500 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_625
timestamp 1649977179
transform 1 0 58604 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_637
timestamp 1649977179
transform 1 0 59708 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_643
timestamp 1649977179
transform 1 0 60260 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_645
timestamp 1649977179
transform 1 0 60444 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_657
timestamp 1649977179
transform 1 0 61548 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_669
timestamp 1649977179
transform 1 0 62652 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_681
timestamp 1649977179
transform 1 0 63756 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_693
timestamp 1649977179
transform 1 0 64860 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_699
timestamp 1649977179
transform 1 0 65412 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_701
timestamp 1649977179
transform 1 0 65596 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_713
timestamp 1649977179
transform 1 0 66700 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_725
timestamp 1649977179
transform 1 0 67804 0 1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1649977179
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1649977179
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_27
timestamp 1649977179
transform 1 0 3588 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_15_39
timestamp 1649977179
transform 1 0 4692 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_45
timestamp 1649977179
transform 1 0 5244 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_52
timestamp 1649977179
transform 1 0 5888 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_65
timestamp 1649977179
transform 1 0 7084 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_71
timestamp 1649977179
transform 1 0 7636 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_88
timestamp 1649977179
transform 1 0 9200 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_108
timestamp 1649977179
transform 1 0 11040 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1649977179
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_125
timestamp 1649977179
transform 1 0 12604 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_145
timestamp 1649977179
transform 1 0 14444 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_157
timestamp 1649977179
transform 1 0 15548 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_165
timestamp 1649977179
transform 1 0 16284 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_177
timestamp 1649977179
transform 1 0 17388 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_15_201
timestamp 1649977179
transform 1 0 19596 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_209
timestamp 1649977179
transform 1 0 20332 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_218
timestamp 1649977179
transform 1 0 21160 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_15_230
timestamp 1649977179
transform 1 0 22264 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_243
timestamp 1649977179
transform 1 0 23460 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_252
timestamp 1649977179
transform 1 0 24288 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_264
timestamp 1649977179
transform 1 0 25392 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_276
timestamp 1649977179
transform 1 0 26496 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_281
timestamp 1649977179
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_293
timestamp 1649977179
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_305
timestamp 1649977179
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_317
timestamp 1649977179
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_329
timestamp 1649977179
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1649977179
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_337
timestamp 1649977179
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_349
timestamp 1649977179
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_361
timestamp 1649977179
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_373
timestamp 1649977179
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1649977179
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1649977179
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_393
timestamp 1649977179
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_405
timestamp 1649977179
transform 1 0 38364 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_417
timestamp 1649977179
transform 1 0 39468 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_429
timestamp 1649977179
transform 1 0 40572 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_441
timestamp 1649977179
transform 1 0 41676 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_447
timestamp 1649977179
transform 1 0 42228 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_449
timestamp 1649977179
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_461
timestamp 1649977179
transform 1 0 43516 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_473
timestamp 1649977179
transform 1 0 44620 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_485
timestamp 1649977179
transform 1 0 45724 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_497
timestamp 1649977179
transform 1 0 46828 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_503
timestamp 1649977179
transform 1 0 47380 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_505
timestamp 1649977179
transform 1 0 47564 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_517
timestamp 1649977179
transform 1 0 48668 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_529
timestamp 1649977179
transform 1 0 49772 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_541
timestamp 1649977179
transform 1 0 50876 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_553
timestamp 1649977179
transform 1 0 51980 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_559
timestamp 1649977179
transform 1 0 52532 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_561
timestamp 1649977179
transform 1 0 52716 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_573
timestamp 1649977179
transform 1 0 53820 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_585
timestamp 1649977179
transform 1 0 54924 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_597
timestamp 1649977179
transform 1 0 56028 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_609
timestamp 1649977179
transform 1 0 57132 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_615
timestamp 1649977179
transform 1 0 57684 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_617
timestamp 1649977179
transform 1 0 57868 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_629
timestamp 1649977179
transform 1 0 58972 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_641
timestamp 1649977179
transform 1 0 60076 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_653
timestamp 1649977179
transform 1 0 61180 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_665
timestamp 1649977179
transform 1 0 62284 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_671
timestamp 1649977179
transform 1 0 62836 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_673
timestamp 1649977179
transform 1 0 63020 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_685
timestamp 1649977179
transform 1 0 64124 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_697
timestamp 1649977179
transform 1 0 65228 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_709
timestamp 1649977179
transform 1 0 66332 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_721
timestamp 1649977179
transform 1 0 67436 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_727
timestamp 1649977179
transform 1 0 67988 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_729
timestamp 1649977179
transform 1 0 68172 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1649977179
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1649977179
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1649977179
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_29
timestamp 1649977179
transform 1 0 3772 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_39
timestamp 1649977179
transform 1 0 4692 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_47
timestamp 1649977179
transform 1 0 5428 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_58
timestamp 1649977179
transform 1 0 6440 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_70
timestamp 1649977179
transform 1 0 7544 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_82
timestamp 1649977179
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1649977179
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_97
timestamp 1649977179
transform 1 0 10028 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_116
timestamp 1649977179
transform 1 0 11776 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_136
timestamp 1649977179
transform 1 0 13616 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1649977179
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_153
timestamp 1649977179
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_165
timestamp 1649977179
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_177
timestamp 1649977179
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1649977179
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1649977179
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_197
timestamp 1649977179
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_209
timestamp 1649977179
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_221
timestamp 1649977179
transform 1 0 21436 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_229
timestamp 1649977179
transform 1 0 22172 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_236
timestamp 1649977179
transform 1 0 22816 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_246
timestamp 1649977179
transform 1 0 23736 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_16_253
timestamp 1649977179
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_265
timestamp 1649977179
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_277
timestamp 1649977179
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_289
timestamp 1649977179
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 1649977179
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1649977179
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_309
timestamp 1649977179
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_321
timestamp 1649977179
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_333
timestamp 1649977179
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_345
timestamp 1649977179
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_357
timestamp 1649977179
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1649977179
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_365
timestamp 1649977179
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_377
timestamp 1649977179
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_389
timestamp 1649977179
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_401
timestamp 1649977179
transform 1 0 37996 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_413
timestamp 1649977179
transform 1 0 39100 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_419
timestamp 1649977179
transform 1 0 39652 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_421
timestamp 1649977179
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_433
timestamp 1649977179
transform 1 0 40940 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_445
timestamp 1649977179
transform 1 0 42044 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_457
timestamp 1649977179
transform 1 0 43148 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_469
timestamp 1649977179
transform 1 0 44252 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_475
timestamp 1649977179
transform 1 0 44804 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_477
timestamp 1649977179
transform 1 0 44988 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_489
timestamp 1649977179
transform 1 0 46092 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_501
timestamp 1649977179
transform 1 0 47196 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_513
timestamp 1649977179
transform 1 0 48300 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_525
timestamp 1649977179
transform 1 0 49404 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_531
timestamp 1649977179
transform 1 0 49956 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_533
timestamp 1649977179
transform 1 0 50140 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_545
timestamp 1649977179
transform 1 0 51244 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_557
timestamp 1649977179
transform 1 0 52348 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_569
timestamp 1649977179
transform 1 0 53452 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_581
timestamp 1649977179
transform 1 0 54556 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_587
timestamp 1649977179
transform 1 0 55108 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_589
timestamp 1649977179
transform 1 0 55292 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_601
timestamp 1649977179
transform 1 0 56396 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_613
timestamp 1649977179
transform 1 0 57500 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_625
timestamp 1649977179
transform 1 0 58604 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_637
timestamp 1649977179
transform 1 0 59708 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_643
timestamp 1649977179
transform 1 0 60260 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_645
timestamp 1649977179
transform 1 0 60444 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_657
timestamp 1649977179
transform 1 0 61548 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_669
timestamp 1649977179
transform 1 0 62652 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_681
timestamp 1649977179
transform 1 0 63756 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_693
timestamp 1649977179
transform 1 0 64860 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_699
timestamp 1649977179
transform 1 0 65412 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_701
timestamp 1649977179
transform 1 0 65596 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_713
timestamp 1649977179
transform 1 0 66700 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_725
timestamp 1649977179
transform 1 0 67804 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1649977179
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1649977179
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1649977179
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_47
timestamp 1649977179
transform 1 0 5428 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1649977179
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_57
timestamp 1649977179
transform 1 0 6348 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_65
timestamp 1649977179
transform 1 0 7084 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_82
timestamp 1649977179
transform 1 0 8648 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_102
timestamp 1649977179
transform 1 0 10488 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_110
timestamp 1649977179
transform 1 0 11224 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1649977179
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_125
timestamp 1649977179
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_137
timestamp 1649977179
transform 1 0 13708 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_145
timestamp 1649977179
transform 1 0 14444 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_163
timestamp 1649977179
transform 1 0 16100 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1649977179
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1649977179
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_181
timestamp 1649977179
transform 1 0 17756 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_187
timestamp 1649977179
transform 1 0 18308 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_204
timestamp 1649977179
transform 1 0 19872 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_220
timestamp 1649977179
transform 1 0 21344 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_225
timestamp 1649977179
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_237
timestamp 1649977179
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_249
timestamp 1649977179
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_261
timestamp 1649977179
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1649977179
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1649977179
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_281
timestamp 1649977179
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_293
timestamp 1649977179
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_305
timestamp 1649977179
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_317
timestamp 1649977179
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_329
timestamp 1649977179
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1649977179
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_337
timestamp 1649977179
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_349
timestamp 1649977179
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_361
timestamp 1649977179
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_373
timestamp 1649977179
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1649977179
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1649977179
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_393
timestamp 1649977179
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_405
timestamp 1649977179
transform 1 0 38364 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_417
timestamp 1649977179
transform 1 0 39468 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_429
timestamp 1649977179
transform 1 0 40572 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_441
timestamp 1649977179
transform 1 0 41676 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_447
timestamp 1649977179
transform 1 0 42228 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_449
timestamp 1649977179
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_461
timestamp 1649977179
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_473
timestamp 1649977179
transform 1 0 44620 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_485
timestamp 1649977179
transform 1 0 45724 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_497
timestamp 1649977179
transform 1 0 46828 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_503
timestamp 1649977179
transform 1 0 47380 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_505
timestamp 1649977179
transform 1 0 47564 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_517
timestamp 1649977179
transform 1 0 48668 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_529
timestamp 1649977179
transform 1 0 49772 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_541
timestamp 1649977179
transform 1 0 50876 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_553
timestamp 1649977179
transform 1 0 51980 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_559
timestamp 1649977179
transform 1 0 52532 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_561
timestamp 1649977179
transform 1 0 52716 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_573
timestamp 1649977179
transform 1 0 53820 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_585
timestamp 1649977179
transform 1 0 54924 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_597
timestamp 1649977179
transform 1 0 56028 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_609
timestamp 1649977179
transform 1 0 57132 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_615
timestamp 1649977179
transform 1 0 57684 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_617
timestamp 1649977179
transform 1 0 57868 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_629
timestamp 1649977179
transform 1 0 58972 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_641
timestamp 1649977179
transform 1 0 60076 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_653
timestamp 1649977179
transform 1 0 61180 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_665
timestamp 1649977179
transform 1 0 62284 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_671
timestamp 1649977179
transform 1 0 62836 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_673
timestamp 1649977179
transform 1 0 63020 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_685
timestamp 1649977179
transform 1 0 64124 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_697
timestamp 1649977179
transform 1 0 65228 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_709
timestamp 1649977179
transform 1 0 66332 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_721
timestamp 1649977179
transform 1 0 67436 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_727
timestamp 1649977179
transform 1 0 67988 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_729
timestamp 1649977179
transform 1 0 68172 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1649977179
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1649977179
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1649977179
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_29
timestamp 1649977179
transform 1 0 3772 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_37
timestamp 1649977179
transform 1 0 4508 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_49
timestamp 1649977179
transform 1 0 5612 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_61
timestamp 1649977179
transform 1 0 6716 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_80
timestamp 1649977179
transform 1 0 8464 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1649977179
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_97
timestamp 1649977179
transform 1 0 10028 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_114
timestamp 1649977179
transform 1 0 11592 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_134
timestamp 1649977179
transform 1 0 13432 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1649977179
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_153
timestamp 1649977179
transform 1 0 15180 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_172
timestamp 1649977179
transform 1 0 16928 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_192
timestamp 1649977179
transform 1 0 18768 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_213
timestamp 1649977179
transform 1 0 20700 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_225
timestamp 1649977179
transform 1 0 21804 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_237
timestamp 1649977179
transform 1 0 22908 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_249
timestamp 1649977179
transform 1 0 24012 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_253
timestamp 1649977179
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_265
timestamp 1649977179
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_277
timestamp 1649977179
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_289
timestamp 1649977179
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_301
timestamp 1649977179
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1649977179
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_309
timestamp 1649977179
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_321
timestamp 1649977179
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_333
timestamp 1649977179
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_345
timestamp 1649977179
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1649977179
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1649977179
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_365
timestamp 1649977179
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_377
timestamp 1649977179
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_389
timestamp 1649977179
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_401
timestamp 1649977179
transform 1 0 37996 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_413
timestamp 1649977179
transform 1 0 39100 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_419
timestamp 1649977179
transform 1 0 39652 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_421
timestamp 1649977179
transform 1 0 39836 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_433
timestamp 1649977179
transform 1 0 40940 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_445
timestamp 1649977179
transform 1 0 42044 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_457
timestamp 1649977179
transform 1 0 43148 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_469
timestamp 1649977179
transform 1 0 44252 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_475
timestamp 1649977179
transform 1 0 44804 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_477
timestamp 1649977179
transform 1 0 44988 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_489
timestamp 1649977179
transform 1 0 46092 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_501
timestamp 1649977179
transform 1 0 47196 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_513
timestamp 1649977179
transform 1 0 48300 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_525
timestamp 1649977179
transform 1 0 49404 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_531
timestamp 1649977179
transform 1 0 49956 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_533
timestamp 1649977179
transform 1 0 50140 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_545
timestamp 1649977179
transform 1 0 51244 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_557
timestamp 1649977179
transform 1 0 52348 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_569
timestamp 1649977179
transform 1 0 53452 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_581
timestamp 1649977179
transform 1 0 54556 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_587
timestamp 1649977179
transform 1 0 55108 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_589
timestamp 1649977179
transform 1 0 55292 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_601
timestamp 1649977179
transform 1 0 56396 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_613
timestamp 1649977179
transform 1 0 57500 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_625
timestamp 1649977179
transform 1 0 58604 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_637
timestamp 1649977179
transform 1 0 59708 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_643
timestamp 1649977179
transform 1 0 60260 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_645
timestamp 1649977179
transform 1 0 60444 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_657
timestamp 1649977179
transform 1 0 61548 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_669
timestamp 1649977179
transform 1 0 62652 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_681
timestamp 1649977179
transform 1 0 63756 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_693
timestamp 1649977179
transform 1 0 64860 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_699
timestamp 1649977179
transform 1 0 65412 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_701
timestamp 1649977179
transform 1 0 65596 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_713
timestamp 1649977179
transform 1 0 66700 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_725
timestamp 1649977179
transform 1 0 67804 0 1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1649977179
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1649977179
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1649977179
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_47
timestamp 1649977179
transform 1 0 5428 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1649977179
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1649977179
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_69
timestamp 1649977179
transform 1 0 7452 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_72
timestamp 1649977179
transform 1 0 7728 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_84
timestamp 1649977179
transform 1 0 8832 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_91
timestamp 1649977179
transform 1 0 9476 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_103
timestamp 1649977179
transform 1 0 10580 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1649977179
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1649977179
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_125
timestamp 1649977179
transform 1 0 12604 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_133
timestamp 1649977179
transform 1 0 13340 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_150
timestamp 1649977179
transform 1 0 14904 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_164
timestamp 1649977179
transform 1 0 16192 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_169
timestamp 1649977179
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_181
timestamp 1649977179
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_193
timestamp 1649977179
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_205
timestamp 1649977179
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_217
timestamp 1649977179
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1649977179
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_225
timestamp 1649977179
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_237
timestamp 1649977179
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_249
timestamp 1649977179
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_261
timestamp 1649977179
transform 1 0 25116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_273
timestamp 1649977179
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1649977179
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_281
timestamp 1649977179
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_293
timestamp 1649977179
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_305
timestamp 1649977179
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_317
timestamp 1649977179
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 1649977179
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1649977179
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_337
timestamp 1649977179
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_349
timestamp 1649977179
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_361
timestamp 1649977179
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_373
timestamp 1649977179
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_385
timestamp 1649977179
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1649977179
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_393
timestamp 1649977179
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_405
timestamp 1649977179
transform 1 0 38364 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_417
timestamp 1649977179
transform 1 0 39468 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_429
timestamp 1649977179
transform 1 0 40572 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_441
timestamp 1649977179
transform 1 0 41676 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_447
timestamp 1649977179
transform 1 0 42228 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_449
timestamp 1649977179
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_461
timestamp 1649977179
transform 1 0 43516 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_473
timestamp 1649977179
transform 1 0 44620 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_485
timestamp 1649977179
transform 1 0 45724 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_497
timestamp 1649977179
transform 1 0 46828 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_503
timestamp 1649977179
transform 1 0 47380 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_505
timestamp 1649977179
transform 1 0 47564 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_517
timestamp 1649977179
transform 1 0 48668 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_529
timestamp 1649977179
transform 1 0 49772 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_541
timestamp 1649977179
transform 1 0 50876 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_553
timestamp 1649977179
transform 1 0 51980 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_559
timestamp 1649977179
transform 1 0 52532 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_561
timestamp 1649977179
transform 1 0 52716 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_573
timestamp 1649977179
transform 1 0 53820 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_585
timestamp 1649977179
transform 1 0 54924 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_597
timestamp 1649977179
transform 1 0 56028 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_609
timestamp 1649977179
transform 1 0 57132 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_615
timestamp 1649977179
transform 1 0 57684 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_617
timestamp 1649977179
transform 1 0 57868 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_629
timestamp 1649977179
transform 1 0 58972 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_641
timestamp 1649977179
transform 1 0 60076 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_653
timestamp 1649977179
transform 1 0 61180 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_665
timestamp 1649977179
transform 1 0 62284 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_671
timestamp 1649977179
transform 1 0 62836 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_673
timestamp 1649977179
transform 1 0 63020 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_685
timestamp 1649977179
transform 1 0 64124 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_697
timestamp 1649977179
transform 1 0 65228 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_709
timestamp 1649977179
transform 1 0 66332 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_721
timestamp 1649977179
transform 1 0 67436 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_727
timestamp 1649977179
transform 1 0 67988 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_729
timestamp 1649977179
transform 1 0 68172 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1649977179
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1649977179
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1649977179
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1649977179
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1649977179
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1649977179
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_65
timestamp 1649977179
transform 1 0 7084 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_70
timestamp 1649977179
transform 1 0 7544 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_79
timestamp 1649977179
transform 1 0 8372 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1649977179
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_90
timestamp 1649977179
transform 1 0 9384 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_98
timestamp 1649977179
transform 1 0 10120 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_108
timestamp 1649977179
transform 1 0 11040 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_114
timestamp 1649977179
transform 1 0 11592 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_122
timestamp 1649977179
transform 1 0 12328 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_132
timestamp 1649977179
transform 1 0 13248 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_141
timestamp 1649977179
transform 1 0 14076 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_149
timestamp 1649977179
transform 1 0 14812 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_160
timestamp 1649977179
transform 1 0 15824 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_172
timestamp 1649977179
transform 1 0 16928 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_184
timestamp 1649977179
transform 1 0 18032 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_197
timestamp 1649977179
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_209
timestamp 1649977179
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_221
timestamp 1649977179
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_233
timestamp 1649977179
transform 1 0 22540 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_245
timestamp 1649977179
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1649977179
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_253
timestamp 1649977179
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_265
timestamp 1649977179
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_277
timestamp 1649977179
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_289
timestamp 1649977179
transform 1 0 27692 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_301
timestamp 1649977179
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1649977179
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_309
timestamp 1649977179
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_321
timestamp 1649977179
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_333
timestamp 1649977179
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_345
timestamp 1649977179
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_357
timestamp 1649977179
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1649977179
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_365
timestamp 1649977179
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_377
timestamp 1649977179
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_389
timestamp 1649977179
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_401
timestamp 1649977179
transform 1 0 37996 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_413
timestamp 1649977179
transform 1 0 39100 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_419
timestamp 1649977179
transform 1 0 39652 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_421
timestamp 1649977179
transform 1 0 39836 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_433
timestamp 1649977179
transform 1 0 40940 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_445
timestamp 1649977179
transform 1 0 42044 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_457
timestamp 1649977179
transform 1 0 43148 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_469
timestamp 1649977179
transform 1 0 44252 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_475
timestamp 1649977179
transform 1 0 44804 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_477
timestamp 1649977179
transform 1 0 44988 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_489
timestamp 1649977179
transform 1 0 46092 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_501
timestamp 1649977179
transform 1 0 47196 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_513
timestamp 1649977179
transform 1 0 48300 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_525
timestamp 1649977179
transform 1 0 49404 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_531
timestamp 1649977179
transform 1 0 49956 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_533
timestamp 1649977179
transform 1 0 50140 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_545
timestamp 1649977179
transform 1 0 51244 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_557
timestamp 1649977179
transform 1 0 52348 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_569
timestamp 1649977179
transform 1 0 53452 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_581
timestamp 1649977179
transform 1 0 54556 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_587
timestamp 1649977179
transform 1 0 55108 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_589
timestamp 1649977179
transform 1 0 55292 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_601
timestamp 1649977179
transform 1 0 56396 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_613
timestamp 1649977179
transform 1 0 57500 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_625
timestamp 1649977179
transform 1 0 58604 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_637
timestamp 1649977179
transform 1 0 59708 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_643
timestamp 1649977179
transform 1 0 60260 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_645
timestamp 1649977179
transform 1 0 60444 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_657
timestamp 1649977179
transform 1 0 61548 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_669
timestamp 1649977179
transform 1 0 62652 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_681
timestamp 1649977179
transform 1 0 63756 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_693
timestamp 1649977179
transform 1 0 64860 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_699
timestamp 1649977179
transform 1 0 65412 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_701
timestamp 1649977179
transform 1 0 65596 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_713
timestamp 1649977179
transform 1 0 66700 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_725
timestamp 1649977179
transform 1 0 67804 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1649977179
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1649977179
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_27
timestamp 1649977179
transform 1 0 3588 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_31
timestamp 1649977179
transform 1 0 3956 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_37
timestamp 1649977179
transform 1 0 4508 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_43
timestamp 1649977179
transform 1 0 5060 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1649977179
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_57
timestamp 1649977179
transform 1 0 6348 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_65
timestamp 1649977179
transform 1 0 7084 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_70
timestamp 1649977179
transform 1 0 7544 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_74
timestamp 1649977179
transform 1 0 7912 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_80
timestamp 1649977179
transform 1 0 8464 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_89
timestamp 1649977179
transform 1 0 9292 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_97
timestamp 1649977179
transform 1 0 10028 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_108
timestamp 1649977179
transform 1 0 11040 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_123
timestamp 1649977179
transform 1 0 12420 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_129
timestamp 1649977179
transform 1 0 12972 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_138
timestamp 1649977179
transform 1 0 13800 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_144
timestamp 1649977179
transform 1 0 14352 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_158
timestamp 1649977179
transform 1 0 15640 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp 1649977179
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_169
timestamp 1649977179
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_181
timestamp 1649977179
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_193
timestamp 1649977179
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_205
timestamp 1649977179
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_217
timestamp 1649977179
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1649977179
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_225
timestamp 1649977179
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_237
timestamp 1649977179
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_249
timestamp 1649977179
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_261
timestamp 1649977179
transform 1 0 25116 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_273
timestamp 1649977179
transform 1 0 26220 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1649977179
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_281
timestamp 1649977179
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_293
timestamp 1649977179
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_305
timestamp 1649977179
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_317
timestamp 1649977179
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_329
timestamp 1649977179
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1649977179
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_337
timestamp 1649977179
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_349
timestamp 1649977179
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_361
timestamp 1649977179
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_373
timestamp 1649977179
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1649977179
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1649977179
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_393
timestamp 1649977179
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_405
timestamp 1649977179
transform 1 0 38364 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_417
timestamp 1649977179
transform 1 0 39468 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_429
timestamp 1649977179
transform 1 0 40572 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_441
timestamp 1649977179
transform 1 0 41676 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_447
timestamp 1649977179
transform 1 0 42228 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_449
timestamp 1649977179
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_461
timestamp 1649977179
transform 1 0 43516 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_473
timestamp 1649977179
transform 1 0 44620 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_485
timestamp 1649977179
transform 1 0 45724 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_497
timestamp 1649977179
transform 1 0 46828 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_503
timestamp 1649977179
transform 1 0 47380 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_505
timestamp 1649977179
transform 1 0 47564 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_517
timestamp 1649977179
transform 1 0 48668 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_529
timestamp 1649977179
transform 1 0 49772 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_541
timestamp 1649977179
transform 1 0 50876 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_553
timestamp 1649977179
transform 1 0 51980 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_559
timestamp 1649977179
transform 1 0 52532 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_561
timestamp 1649977179
transform 1 0 52716 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_573
timestamp 1649977179
transform 1 0 53820 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_585
timestamp 1649977179
transform 1 0 54924 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_597
timestamp 1649977179
transform 1 0 56028 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_609
timestamp 1649977179
transform 1 0 57132 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_615
timestamp 1649977179
transform 1 0 57684 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_617
timestamp 1649977179
transform 1 0 57868 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_629
timestamp 1649977179
transform 1 0 58972 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_641
timestamp 1649977179
transform 1 0 60076 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_653
timestamp 1649977179
transform 1 0 61180 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_665
timestamp 1649977179
transform 1 0 62284 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_671
timestamp 1649977179
transform 1 0 62836 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_673
timestamp 1649977179
transform 1 0 63020 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_685
timestamp 1649977179
transform 1 0 64124 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_697
timestamp 1649977179
transform 1 0 65228 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_709
timestamp 1649977179
transform 1 0 66332 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_721
timestamp 1649977179
transform 1 0 67436 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_727
timestamp 1649977179
transform 1 0 67988 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_729
timestamp 1649977179
transform 1 0 68172 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1649977179
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1649977179
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1649977179
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1649977179
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1649977179
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1649977179
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1649977179
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1649977179
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1649977179
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1649977179
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_97
timestamp 1649977179
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_109
timestamp 1649977179
transform 1 0 11132 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_113
timestamp 1649977179
transform 1 0 11500 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_122
timestamp 1649977179
transform 1 0 12328 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_134
timestamp 1649977179
transform 1 0 13432 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_22_141
timestamp 1649977179
transform 1 0 14076 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_149
timestamp 1649977179
transform 1 0 14812 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_159
timestamp 1649977179
transform 1 0 15732 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_171
timestamp 1649977179
transform 1 0 16836 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_183
timestamp 1649977179
transform 1 0 17940 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1649977179
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_197
timestamp 1649977179
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_209
timestamp 1649977179
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_221
timestamp 1649977179
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_233
timestamp 1649977179
transform 1 0 22540 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_245
timestamp 1649977179
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1649977179
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_253
timestamp 1649977179
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_265
timestamp 1649977179
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_277
timestamp 1649977179
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_289
timestamp 1649977179
transform 1 0 27692 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_301
timestamp 1649977179
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1649977179
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_309
timestamp 1649977179
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_321
timestamp 1649977179
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_333
timestamp 1649977179
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_345
timestamp 1649977179
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 1649977179
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1649977179
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_365
timestamp 1649977179
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_377
timestamp 1649977179
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_389
timestamp 1649977179
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_401
timestamp 1649977179
transform 1 0 37996 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_413
timestamp 1649977179
transform 1 0 39100 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_419
timestamp 1649977179
transform 1 0 39652 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_421
timestamp 1649977179
transform 1 0 39836 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_433
timestamp 1649977179
transform 1 0 40940 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_445
timestamp 1649977179
transform 1 0 42044 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_457
timestamp 1649977179
transform 1 0 43148 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_469
timestamp 1649977179
transform 1 0 44252 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_475
timestamp 1649977179
transform 1 0 44804 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_477
timestamp 1649977179
transform 1 0 44988 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_489
timestamp 1649977179
transform 1 0 46092 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_501
timestamp 1649977179
transform 1 0 47196 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_513
timestamp 1649977179
transform 1 0 48300 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_525
timestamp 1649977179
transform 1 0 49404 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_531
timestamp 1649977179
transform 1 0 49956 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_533
timestamp 1649977179
transform 1 0 50140 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_545
timestamp 1649977179
transform 1 0 51244 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_557
timestamp 1649977179
transform 1 0 52348 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_569
timestamp 1649977179
transform 1 0 53452 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_581
timestamp 1649977179
transform 1 0 54556 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_587
timestamp 1649977179
transform 1 0 55108 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_589
timestamp 1649977179
transform 1 0 55292 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_601
timestamp 1649977179
transform 1 0 56396 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_613
timestamp 1649977179
transform 1 0 57500 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_625
timestamp 1649977179
transform 1 0 58604 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_637
timestamp 1649977179
transform 1 0 59708 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_643
timestamp 1649977179
transform 1 0 60260 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_645
timestamp 1649977179
transform 1 0 60444 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_657
timestamp 1649977179
transform 1 0 61548 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_669
timestamp 1649977179
transform 1 0 62652 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_681
timestamp 1649977179
transform 1 0 63756 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_693
timestamp 1649977179
transform 1 0 64860 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_699
timestamp 1649977179
transform 1 0 65412 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_701
timestamp 1649977179
transform 1 0 65596 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_713
timestamp 1649977179
transform 1 0 66700 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_725
timestamp 1649977179
transform 1 0 67804 0 1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1649977179
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1649977179
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1649977179
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1649977179
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1649977179
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1649977179
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1649977179
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1649977179
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 1649977179
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_93
timestamp 1649977179
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1649977179
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1649977179
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1649977179
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1649977179
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_137
timestamp 1649977179
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_149
timestamp 1649977179
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1649977179
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1649977179
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_169
timestamp 1649977179
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_181
timestamp 1649977179
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_193
timestamp 1649977179
transform 1 0 18860 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_205
timestamp 1649977179
transform 1 0 19964 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_217
timestamp 1649977179
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1649977179
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_225
timestamp 1649977179
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_237
timestamp 1649977179
transform 1 0 22908 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_249
timestamp 1649977179
transform 1 0 24012 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_261
timestamp 1649977179
transform 1 0 25116 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_273
timestamp 1649977179
transform 1 0 26220 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 1649977179
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_281
timestamp 1649977179
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_293
timestamp 1649977179
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_305
timestamp 1649977179
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_317
timestamp 1649977179
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_329
timestamp 1649977179
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1649977179
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_337
timestamp 1649977179
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_349
timestamp 1649977179
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_361
timestamp 1649977179
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_373
timestamp 1649977179
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1649977179
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1649977179
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_393
timestamp 1649977179
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_405
timestamp 1649977179
transform 1 0 38364 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_417
timestamp 1649977179
transform 1 0 39468 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_429
timestamp 1649977179
transform 1 0 40572 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_441
timestamp 1649977179
transform 1 0 41676 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_447
timestamp 1649977179
transform 1 0 42228 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_449
timestamp 1649977179
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_461
timestamp 1649977179
transform 1 0 43516 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_473
timestamp 1649977179
transform 1 0 44620 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_485
timestamp 1649977179
transform 1 0 45724 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_497
timestamp 1649977179
transform 1 0 46828 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_503
timestamp 1649977179
transform 1 0 47380 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_505
timestamp 1649977179
transform 1 0 47564 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_517
timestamp 1649977179
transform 1 0 48668 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_529
timestamp 1649977179
transform 1 0 49772 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_541
timestamp 1649977179
transform 1 0 50876 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_553
timestamp 1649977179
transform 1 0 51980 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_559
timestamp 1649977179
transform 1 0 52532 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_561
timestamp 1649977179
transform 1 0 52716 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_573
timestamp 1649977179
transform 1 0 53820 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_585
timestamp 1649977179
transform 1 0 54924 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_597
timestamp 1649977179
transform 1 0 56028 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_609
timestamp 1649977179
transform 1 0 57132 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_615
timestamp 1649977179
transform 1 0 57684 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_617
timestamp 1649977179
transform 1 0 57868 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_629
timestamp 1649977179
transform 1 0 58972 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_641
timestamp 1649977179
transform 1 0 60076 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_653
timestamp 1649977179
transform 1 0 61180 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_665
timestamp 1649977179
transform 1 0 62284 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_671
timestamp 1649977179
transform 1 0 62836 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_673
timestamp 1649977179
transform 1 0 63020 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_685
timestamp 1649977179
transform 1 0 64124 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_697
timestamp 1649977179
transform 1 0 65228 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_709
timestamp 1649977179
transform 1 0 66332 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_721
timestamp 1649977179
transform 1 0 67436 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_727
timestamp 1649977179
transform 1 0 67988 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_729
timestamp 1649977179
transform 1 0 68172 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1649977179
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1649977179
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1649977179
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1649977179
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1649977179
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1649977179
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1649977179
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1649977179
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1649977179
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1649977179
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_97
timestamp 1649977179
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_109
timestamp 1649977179
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_121
timestamp 1649977179
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1649977179
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1649977179
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1649977179
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_153
timestamp 1649977179
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_165
timestamp 1649977179
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_177
timestamp 1649977179
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_189
timestamp 1649977179
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1649977179
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_197
timestamp 1649977179
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_209
timestamp 1649977179
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_221
timestamp 1649977179
transform 1 0 21436 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_233
timestamp 1649977179
transform 1 0 22540 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_245
timestamp 1649977179
transform 1 0 23644 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1649977179
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_253
timestamp 1649977179
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_265
timestamp 1649977179
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_277
timestamp 1649977179
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_289
timestamp 1649977179
transform 1 0 27692 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_301
timestamp 1649977179
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1649977179
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_309
timestamp 1649977179
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_321
timestamp 1649977179
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_333
timestamp 1649977179
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_345
timestamp 1649977179
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_357
timestamp 1649977179
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1649977179
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_365
timestamp 1649977179
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_377
timestamp 1649977179
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_389
timestamp 1649977179
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_401
timestamp 1649977179
transform 1 0 37996 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_413
timestamp 1649977179
transform 1 0 39100 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_419
timestamp 1649977179
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_421
timestamp 1649977179
transform 1 0 39836 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_433
timestamp 1649977179
transform 1 0 40940 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_445
timestamp 1649977179
transform 1 0 42044 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_457
timestamp 1649977179
transform 1 0 43148 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_469
timestamp 1649977179
transform 1 0 44252 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_475
timestamp 1649977179
transform 1 0 44804 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_477
timestamp 1649977179
transform 1 0 44988 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_489
timestamp 1649977179
transform 1 0 46092 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_501
timestamp 1649977179
transform 1 0 47196 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_513
timestamp 1649977179
transform 1 0 48300 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_525
timestamp 1649977179
transform 1 0 49404 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_531
timestamp 1649977179
transform 1 0 49956 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_533
timestamp 1649977179
transform 1 0 50140 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_545
timestamp 1649977179
transform 1 0 51244 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_557
timestamp 1649977179
transform 1 0 52348 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_569
timestamp 1649977179
transform 1 0 53452 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_581
timestamp 1649977179
transform 1 0 54556 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_587
timestamp 1649977179
transform 1 0 55108 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_589
timestamp 1649977179
transform 1 0 55292 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_601
timestamp 1649977179
transform 1 0 56396 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_613
timestamp 1649977179
transform 1 0 57500 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_625
timestamp 1649977179
transform 1 0 58604 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_637
timestamp 1649977179
transform 1 0 59708 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_643
timestamp 1649977179
transform 1 0 60260 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_645
timestamp 1649977179
transform 1 0 60444 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_657
timestamp 1649977179
transform 1 0 61548 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_669
timestamp 1649977179
transform 1 0 62652 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_681
timestamp 1649977179
transform 1 0 63756 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_693
timestamp 1649977179
transform 1 0 64860 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_699
timestamp 1649977179
transform 1 0 65412 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_701
timestamp 1649977179
transform 1 0 65596 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_713
timestamp 1649977179
transform 1 0 66700 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_725
timestamp 1649977179
transform 1 0 67804 0 1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1649977179
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1649977179
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_27
timestamp 1649977179
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_39
timestamp 1649977179
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1649977179
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1649977179
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1649977179
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1649977179
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 1649977179
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_93
timestamp 1649977179
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1649977179
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1649977179
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1649977179
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 1649977179
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_137
timestamp 1649977179
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_149
timestamp 1649977179
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1649977179
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1649977179
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1649977179
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_181
timestamp 1649977179
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_193
timestamp 1649977179
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_205
timestamp 1649977179
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp 1649977179
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1649977179
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_225
timestamp 1649977179
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_237
timestamp 1649977179
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_249
timestamp 1649977179
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_261
timestamp 1649977179
transform 1 0 25116 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_273
timestamp 1649977179
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1649977179
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_281
timestamp 1649977179
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_293
timestamp 1649977179
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_305
timestamp 1649977179
transform 1 0 29164 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_317
timestamp 1649977179
transform 1 0 30268 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_329
timestamp 1649977179
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1649977179
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_337
timestamp 1649977179
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_349
timestamp 1649977179
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_361
timestamp 1649977179
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_373
timestamp 1649977179
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_385
timestamp 1649977179
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1649977179
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_393
timestamp 1649977179
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_405
timestamp 1649977179
transform 1 0 38364 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_417
timestamp 1649977179
transform 1 0 39468 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_429
timestamp 1649977179
transform 1 0 40572 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_441
timestamp 1649977179
transform 1 0 41676 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_447
timestamp 1649977179
transform 1 0 42228 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_449
timestamp 1649977179
transform 1 0 42412 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_461
timestamp 1649977179
transform 1 0 43516 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_473
timestamp 1649977179
transform 1 0 44620 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_485
timestamp 1649977179
transform 1 0 45724 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_497
timestamp 1649977179
transform 1 0 46828 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_503
timestamp 1649977179
transform 1 0 47380 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_505
timestamp 1649977179
transform 1 0 47564 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_517
timestamp 1649977179
transform 1 0 48668 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_529
timestamp 1649977179
transform 1 0 49772 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_541
timestamp 1649977179
transform 1 0 50876 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_553
timestamp 1649977179
transform 1 0 51980 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_559
timestamp 1649977179
transform 1 0 52532 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_561
timestamp 1649977179
transform 1 0 52716 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_573
timestamp 1649977179
transform 1 0 53820 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_585
timestamp 1649977179
transform 1 0 54924 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_597
timestamp 1649977179
transform 1 0 56028 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_609
timestamp 1649977179
transform 1 0 57132 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_615
timestamp 1649977179
transform 1 0 57684 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_617
timestamp 1649977179
transform 1 0 57868 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_629
timestamp 1649977179
transform 1 0 58972 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_641
timestamp 1649977179
transform 1 0 60076 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_653
timestamp 1649977179
transform 1 0 61180 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_665
timestamp 1649977179
transform 1 0 62284 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_671
timestamp 1649977179
transform 1 0 62836 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_673
timestamp 1649977179
transform 1 0 63020 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_685
timestamp 1649977179
transform 1 0 64124 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_697
timestamp 1649977179
transform 1 0 65228 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_709
timestamp 1649977179
transform 1 0 66332 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_721
timestamp 1649977179
transform 1 0 67436 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_727
timestamp 1649977179
transform 1 0 67988 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_729
timestamp 1649977179
transform 1 0 68172 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1649977179
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1649977179
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1649977179
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1649977179
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1649977179
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1649977179
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1649977179
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1649977179
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1649977179
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1649977179
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1649977179
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_109
timestamp 1649977179
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_121
timestamp 1649977179
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1649977179
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1649977179
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1649977179
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_153
timestamp 1649977179
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_165
timestamp 1649977179
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_177
timestamp 1649977179
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_189
timestamp 1649977179
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1649977179
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_197
timestamp 1649977179
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_209
timestamp 1649977179
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_221
timestamp 1649977179
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_233
timestamp 1649977179
transform 1 0 22540 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_245
timestamp 1649977179
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1649977179
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_253
timestamp 1649977179
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_265
timestamp 1649977179
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_277
timestamp 1649977179
transform 1 0 26588 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_289
timestamp 1649977179
transform 1 0 27692 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_301
timestamp 1649977179
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1649977179
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_309
timestamp 1649977179
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_321
timestamp 1649977179
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_333
timestamp 1649977179
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_345
timestamp 1649977179
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_357
timestamp 1649977179
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1649977179
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_365
timestamp 1649977179
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_377
timestamp 1649977179
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_389
timestamp 1649977179
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_401
timestamp 1649977179
transform 1 0 37996 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_413
timestamp 1649977179
transform 1 0 39100 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_419
timestamp 1649977179
transform 1 0 39652 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_421
timestamp 1649977179
transform 1 0 39836 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_433
timestamp 1649977179
transform 1 0 40940 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_445
timestamp 1649977179
transform 1 0 42044 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_457
timestamp 1649977179
transform 1 0 43148 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_469
timestamp 1649977179
transform 1 0 44252 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_475
timestamp 1649977179
transform 1 0 44804 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_477
timestamp 1649977179
transform 1 0 44988 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_489
timestamp 1649977179
transform 1 0 46092 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_501
timestamp 1649977179
transform 1 0 47196 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_513
timestamp 1649977179
transform 1 0 48300 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_525
timestamp 1649977179
transform 1 0 49404 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_531
timestamp 1649977179
transform 1 0 49956 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_533
timestamp 1649977179
transform 1 0 50140 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_545
timestamp 1649977179
transform 1 0 51244 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_557
timestamp 1649977179
transform 1 0 52348 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_569
timestamp 1649977179
transform 1 0 53452 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_581
timestamp 1649977179
transform 1 0 54556 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_587
timestamp 1649977179
transform 1 0 55108 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_589
timestamp 1649977179
transform 1 0 55292 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_601
timestamp 1649977179
transform 1 0 56396 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_613
timestamp 1649977179
transform 1 0 57500 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_625
timestamp 1649977179
transform 1 0 58604 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_637
timestamp 1649977179
transform 1 0 59708 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_643
timestamp 1649977179
transform 1 0 60260 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_645
timestamp 1649977179
transform 1 0 60444 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_657
timestamp 1649977179
transform 1 0 61548 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_669
timestamp 1649977179
transform 1 0 62652 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_681
timestamp 1649977179
transform 1 0 63756 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_693
timestamp 1649977179
transform 1 0 64860 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_699
timestamp 1649977179
transform 1 0 65412 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_701
timestamp 1649977179
transform 1 0 65596 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_713
timestamp 1649977179
transform 1 0 66700 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_725
timestamp 1649977179
transform 1 0 67804 0 1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1649977179
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1649977179
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 1649977179
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_39
timestamp 1649977179
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1649977179
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1649977179
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1649977179
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1649977179
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_81
timestamp 1649977179
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_93
timestamp 1649977179
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1649977179
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1649977179
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1649977179
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1649977179
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_137
timestamp 1649977179
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_149
timestamp 1649977179
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1649977179
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1649977179
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_169
timestamp 1649977179
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_181
timestamp 1649977179
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_193
timestamp 1649977179
transform 1 0 18860 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_205
timestamp 1649977179
transform 1 0 19964 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_217
timestamp 1649977179
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1649977179
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_225
timestamp 1649977179
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_237
timestamp 1649977179
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_249
timestamp 1649977179
transform 1 0 24012 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_261
timestamp 1649977179
transform 1 0 25116 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_273
timestamp 1649977179
transform 1 0 26220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1649977179
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_281
timestamp 1649977179
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_293
timestamp 1649977179
transform 1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_305
timestamp 1649977179
transform 1 0 29164 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_317
timestamp 1649977179
transform 1 0 30268 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_329
timestamp 1649977179
transform 1 0 31372 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1649977179
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_337
timestamp 1649977179
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_349
timestamp 1649977179
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_361
timestamp 1649977179
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_373
timestamp 1649977179
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_385
timestamp 1649977179
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1649977179
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_393
timestamp 1649977179
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_405
timestamp 1649977179
transform 1 0 38364 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_417
timestamp 1649977179
transform 1 0 39468 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_429
timestamp 1649977179
transform 1 0 40572 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_441
timestamp 1649977179
transform 1 0 41676 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_447
timestamp 1649977179
transform 1 0 42228 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_449
timestamp 1649977179
transform 1 0 42412 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_461
timestamp 1649977179
transform 1 0 43516 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_473
timestamp 1649977179
transform 1 0 44620 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_485
timestamp 1649977179
transform 1 0 45724 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_497
timestamp 1649977179
transform 1 0 46828 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_503
timestamp 1649977179
transform 1 0 47380 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_505
timestamp 1649977179
transform 1 0 47564 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_517
timestamp 1649977179
transform 1 0 48668 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_529
timestamp 1649977179
transform 1 0 49772 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_541
timestamp 1649977179
transform 1 0 50876 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_553
timestamp 1649977179
transform 1 0 51980 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_559
timestamp 1649977179
transform 1 0 52532 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_561
timestamp 1649977179
transform 1 0 52716 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_573
timestamp 1649977179
transform 1 0 53820 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_585
timestamp 1649977179
transform 1 0 54924 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_597
timestamp 1649977179
transform 1 0 56028 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_609
timestamp 1649977179
transform 1 0 57132 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_615
timestamp 1649977179
transform 1 0 57684 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_617
timestamp 1649977179
transform 1 0 57868 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_629
timestamp 1649977179
transform 1 0 58972 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_641
timestamp 1649977179
transform 1 0 60076 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_653
timestamp 1649977179
transform 1 0 61180 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_665
timestamp 1649977179
transform 1 0 62284 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_671
timestamp 1649977179
transform 1 0 62836 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_673
timestamp 1649977179
transform 1 0 63020 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_685
timestamp 1649977179
transform 1 0 64124 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_697
timestamp 1649977179
transform 1 0 65228 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_709
timestamp 1649977179
transform 1 0 66332 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_721
timestamp 1649977179
transform 1 0 67436 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_727
timestamp 1649977179
transform 1 0 67988 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_729
timestamp 1649977179
transform 1 0 68172 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1649977179
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1649977179
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1649977179
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1649977179
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1649977179
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1649977179
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1649977179
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1649977179
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1649977179
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1649977179
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1649977179
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_109
timestamp 1649977179
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_121
timestamp 1649977179
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1649977179
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1649977179
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1649977179
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_153
timestamp 1649977179
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_165
timestamp 1649977179
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_177
timestamp 1649977179
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp 1649977179
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1649977179
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_197
timestamp 1649977179
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_209
timestamp 1649977179
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_221
timestamp 1649977179
transform 1 0 21436 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_233
timestamp 1649977179
transform 1 0 22540 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_245
timestamp 1649977179
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1649977179
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_253
timestamp 1649977179
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_265
timestamp 1649977179
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_277
timestamp 1649977179
transform 1 0 26588 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_289
timestamp 1649977179
transform 1 0 27692 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_301
timestamp 1649977179
transform 1 0 28796 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 1649977179
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_309
timestamp 1649977179
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_321
timestamp 1649977179
transform 1 0 30636 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_333
timestamp 1649977179
transform 1 0 31740 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_345
timestamp 1649977179
transform 1 0 32844 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_357
timestamp 1649977179
transform 1 0 33948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1649977179
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_365
timestamp 1649977179
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_377
timestamp 1649977179
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_389
timestamp 1649977179
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_401
timestamp 1649977179
transform 1 0 37996 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_413
timestamp 1649977179
transform 1 0 39100 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_419
timestamp 1649977179
transform 1 0 39652 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_421
timestamp 1649977179
transform 1 0 39836 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_433
timestamp 1649977179
transform 1 0 40940 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_445
timestamp 1649977179
transform 1 0 42044 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_457
timestamp 1649977179
transform 1 0 43148 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_469
timestamp 1649977179
transform 1 0 44252 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_475
timestamp 1649977179
transform 1 0 44804 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_477
timestamp 1649977179
transform 1 0 44988 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_489
timestamp 1649977179
transform 1 0 46092 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_501
timestamp 1649977179
transform 1 0 47196 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_513
timestamp 1649977179
transform 1 0 48300 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_525
timestamp 1649977179
transform 1 0 49404 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_531
timestamp 1649977179
transform 1 0 49956 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_533
timestamp 1649977179
transform 1 0 50140 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_545
timestamp 1649977179
transform 1 0 51244 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_557
timestamp 1649977179
transform 1 0 52348 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_569
timestamp 1649977179
transform 1 0 53452 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_581
timestamp 1649977179
transform 1 0 54556 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_587
timestamp 1649977179
transform 1 0 55108 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_589
timestamp 1649977179
transform 1 0 55292 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_601
timestamp 1649977179
transform 1 0 56396 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_613
timestamp 1649977179
transform 1 0 57500 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_625
timestamp 1649977179
transform 1 0 58604 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_637
timestamp 1649977179
transform 1 0 59708 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_643
timestamp 1649977179
transform 1 0 60260 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_645
timestamp 1649977179
transform 1 0 60444 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_657
timestamp 1649977179
transform 1 0 61548 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_669
timestamp 1649977179
transform 1 0 62652 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_681
timestamp 1649977179
transform 1 0 63756 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_693
timestamp 1649977179
transform 1 0 64860 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_699
timestamp 1649977179
transform 1 0 65412 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_701
timestamp 1649977179
transform 1 0 65596 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_713
timestamp 1649977179
transform 1 0 66700 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_725
timestamp 1649977179
transform 1 0 67804 0 1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1649977179
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_15
timestamp 1649977179
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_27
timestamp 1649977179
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_39
timestamp 1649977179
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1649977179
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1649977179
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1649977179
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_69
timestamp 1649977179
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_81
timestamp 1649977179
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_93
timestamp 1649977179
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1649977179
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1649977179
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1649977179
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_125
timestamp 1649977179
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_137
timestamp 1649977179
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_149
timestamp 1649977179
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1649977179
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1649977179
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 1649977179
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_181
timestamp 1649977179
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_193
timestamp 1649977179
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_205
timestamp 1649977179
transform 1 0 19964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_217
timestamp 1649977179
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1649977179
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_225
timestamp 1649977179
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_237
timestamp 1649977179
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_249
timestamp 1649977179
transform 1 0 24012 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_261
timestamp 1649977179
transform 1 0 25116 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_273
timestamp 1649977179
transform 1 0 26220 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 1649977179
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_281
timestamp 1649977179
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_293
timestamp 1649977179
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_305
timestamp 1649977179
transform 1 0 29164 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_317
timestamp 1649977179
transform 1 0 30268 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_329
timestamp 1649977179
transform 1 0 31372 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 1649977179
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_337
timestamp 1649977179
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_349
timestamp 1649977179
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_361
timestamp 1649977179
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_373
timestamp 1649977179
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_385
timestamp 1649977179
transform 1 0 36524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1649977179
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_393
timestamp 1649977179
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_405
timestamp 1649977179
transform 1 0 38364 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_417
timestamp 1649977179
transform 1 0 39468 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_429
timestamp 1649977179
transform 1 0 40572 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_441
timestamp 1649977179
transform 1 0 41676 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_447
timestamp 1649977179
transform 1 0 42228 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_449
timestamp 1649977179
transform 1 0 42412 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_461
timestamp 1649977179
transform 1 0 43516 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_473
timestamp 1649977179
transform 1 0 44620 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_485
timestamp 1649977179
transform 1 0 45724 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_497
timestamp 1649977179
transform 1 0 46828 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_503
timestamp 1649977179
transform 1 0 47380 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_505
timestamp 1649977179
transform 1 0 47564 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_517
timestamp 1649977179
transform 1 0 48668 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_529
timestamp 1649977179
transform 1 0 49772 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_541
timestamp 1649977179
transform 1 0 50876 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_553
timestamp 1649977179
transform 1 0 51980 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_559
timestamp 1649977179
transform 1 0 52532 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_561
timestamp 1649977179
transform 1 0 52716 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_573
timestamp 1649977179
transform 1 0 53820 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_585
timestamp 1649977179
transform 1 0 54924 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_597
timestamp 1649977179
transform 1 0 56028 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_609
timestamp 1649977179
transform 1 0 57132 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_615
timestamp 1649977179
transform 1 0 57684 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_617
timestamp 1649977179
transform 1 0 57868 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_629
timestamp 1649977179
transform 1 0 58972 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_641
timestamp 1649977179
transform 1 0 60076 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_653
timestamp 1649977179
transform 1 0 61180 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_665
timestamp 1649977179
transform 1 0 62284 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_671
timestamp 1649977179
transform 1 0 62836 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_673
timestamp 1649977179
transform 1 0 63020 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_685
timestamp 1649977179
transform 1 0 64124 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_697
timestamp 1649977179
transform 1 0 65228 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_709
timestamp 1649977179
transform 1 0 66332 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_721
timestamp 1649977179
transform 1 0 67436 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_727
timestamp 1649977179
transform 1 0 67988 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_729
timestamp 1649977179
transform 1 0 68172 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1649977179
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1649977179
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1649977179
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1649977179
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1649977179
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1649977179
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_65
timestamp 1649977179
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1649977179
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1649977179
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1649977179
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_97
timestamp 1649977179
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_109
timestamp 1649977179
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_121
timestamp 1649977179
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1649977179
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1649977179
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1649977179
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_153
timestamp 1649977179
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_165
timestamp 1649977179
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_177
timestamp 1649977179
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1649977179
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1649977179
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_197
timestamp 1649977179
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_209
timestamp 1649977179
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_221
timestamp 1649977179
transform 1 0 21436 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_233
timestamp 1649977179
transform 1 0 22540 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_245
timestamp 1649977179
transform 1 0 23644 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 1649977179
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_253
timestamp 1649977179
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_265
timestamp 1649977179
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_277
timestamp 1649977179
transform 1 0 26588 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_289
timestamp 1649977179
transform 1 0 27692 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_301
timestamp 1649977179
transform 1 0 28796 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_307
timestamp 1649977179
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_309
timestamp 1649977179
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_321
timestamp 1649977179
transform 1 0 30636 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_333
timestamp 1649977179
transform 1 0 31740 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_345
timestamp 1649977179
transform 1 0 32844 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_357
timestamp 1649977179
transform 1 0 33948 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 1649977179
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_365
timestamp 1649977179
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_377
timestamp 1649977179
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_389
timestamp 1649977179
transform 1 0 36892 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_401
timestamp 1649977179
transform 1 0 37996 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_413
timestamp 1649977179
transform 1 0 39100 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_419
timestamp 1649977179
transform 1 0 39652 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_421
timestamp 1649977179
transform 1 0 39836 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_433
timestamp 1649977179
transform 1 0 40940 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_445
timestamp 1649977179
transform 1 0 42044 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_457
timestamp 1649977179
transform 1 0 43148 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_469
timestamp 1649977179
transform 1 0 44252 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_475
timestamp 1649977179
transform 1 0 44804 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_477
timestamp 1649977179
transform 1 0 44988 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_489
timestamp 1649977179
transform 1 0 46092 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_501
timestamp 1649977179
transform 1 0 47196 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_513
timestamp 1649977179
transform 1 0 48300 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_525
timestamp 1649977179
transform 1 0 49404 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_531
timestamp 1649977179
transform 1 0 49956 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_533
timestamp 1649977179
transform 1 0 50140 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_545
timestamp 1649977179
transform 1 0 51244 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_557
timestamp 1649977179
transform 1 0 52348 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_569
timestamp 1649977179
transform 1 0 53452 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_581
timestamp 1649977179
transform 1 0 54556 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_587
timestamp 1649977179
transform 1 0 55108 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_589
timestamp 1649977179
transform 1 0 55292 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_601
timestamp 1649977179
transform 1 0 56396 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_613
timestamp 1649977179
transform 1 0 57500 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_625
timestamp 1649977179
transform 1 0 58604 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_637
timestamp 1649977179
transform 1 0 59708 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_643
timestamp 1649977179
transform 1 0 60260 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_645
timestamp 1649977179
transform 1 0 60444 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_657
timestamp 1649977179
transform 1 0 61548 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_669
timestamp 1649977179
transform 1 0 62652 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_681
timestamp 1649977179
transform 1 0 63756 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_693
timestamp 1649977179
transform 1 0 64860 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_699
timestamp 1649977179
transform 1 0 65412 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_701
timestamp 1649977179
transform 1 0 65596 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_713
timestamp 1649977179
transform 1 0 66700 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_725
timestamp 1649977179
transform 1 0 67804 0 1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1649977179
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1649977179
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_27
timestamp 1649977179
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_39
timestamp 1649977179
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1649977179
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1649977179
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1649977179
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1649977179
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 1649977179
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_93
timestamp 1649977179
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1649977179
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1649977179
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1649977179
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_125
timestamp 1649977179
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_137
timestamp 1649977179
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_149
timestamp 1649977179
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 1649977179
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1649977179
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_169
timestamp 1649977179
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_181
timestamp 1649977179
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_193
timestamp 1649977179
transform 1 0 18860 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_205
timestamp 1649977179
transform 1 0 19964 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_217
timestamp 1649977179
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1649977179
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_225
timestamp 1649977179
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_237
timestamp 1649977179
transform 1 0 22908 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_249
timestamp 1649977179
transform 1 0 24012 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_261
timestamp 1649977179
transform 1 0 25116 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_273
timestamp 1649977179
transform 1 0 26220 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 1649977179
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_281
timestamp 1649977179
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_293
timestamp 1649977179
transform 1 0 28060 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_305
timestamp 1649977179
transform 1 0 29164 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_317
timestamp 1649977179
transform 1 0 30268 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_329
timestamp 1649977179
transform 1 0 31372 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_335
timestamp 1649977179
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_337
timestamp 1649977179
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_349
timestamp 1649977179
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_361
timestamp 1649977179
transform 1 0 34316 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_373
timestamp 1649977179
transform 1 0 35420 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_385
timestamp 1649977179
transform 1 0 36524 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1649977179
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_393
timestamp 1649977179
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_405
timestamp 1649977179
transform 1 0 38364 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_417
timestamp 1649977179
transform 1 0 39468 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_429
timestamp 1649977179
transform 1 0 40572 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_441
timestamp 1649977179
transform 1 0 41676 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_447
timestamp 1649977179
transform 1 0 42228 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_449
timestamp 1649977179
transform 1 0 42412 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_461
timestamp 1649977179
transform 1 0 43516 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_473
timestamp 1649977179
transform 1 0 44620 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_485
timestamp 1649977179
transform 1 0 45724 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_497
timestamp 1649977179
transform 1 0 46828 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_503
timestamp 1649977179
transform 1 0 47380 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_505
timestamp 1649977179
transform 1 0 47564 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_517
timestamp 1649977179
transform 1 0 48668 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_529
timestamp 1649977179
transform 1 0 49772 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_541
timestamp 1649977179
transform 1 0 50876 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_553
timestamp 1649977179
transform 1 0 51980 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_559
timestamp 1649977179
transform 1 0 52532 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_561
timestamp 1649977179
transform 1 0 52716 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_573
timestamp 1649977179
transform 1 0 53820 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_585
timestamp 1649977179
transform 1 0 54924 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_597
timestamp 1649977179
transform 1 0 56028 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_609
timestamp 1649977179
transform 1 0 57132 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_615
timestamp 1649977179
transform 1 0 57684 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_617
timestamp 1649977179
transform 1 0 57868 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_629
timestamp 1649977179
transform 1 0 58972 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_641
timestamp 1649977179
transform 1 0 60076 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_653
timestamp 1649977179
transform 1 0 61180 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_665
timestamp 1649977179
transform 1 0 62284 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_671
timestamp 1649977179
transform 1 0 62836 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_673
timestamp 1649977179
transform 1 0 63020 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_685
timestamp 1649977179
transform 1 0 64124 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_697
timestamp 1649977179
transform 1 0 65228 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_709
timestamp 1649977179
transform 1 0 66332 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_721
timestamp 1649977179
transform 1 0 67436 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_727
timestamp 1649977179
transform 1 0 67988 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_729
timestamp 1649977179
transform 1 0 68172 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1649977179
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1649977179
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1649977179
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1649977179
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1649977179
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1649977179
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_65
timestamp 1649977179
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1649977179
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1649977179
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1649977179
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_97
timestamp 1649977179
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_109
timestamp 1649977179
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_121
timestamp 1649977179
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 1649977179
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1649977179
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_141
timestamp 1649977179
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_153
timestamp 1649977179
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_165
timestamp 1649977179
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_177
timestamp 1649977179
transform 1 0 17388 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_189
timestamp 1649977179
transform 1 0 18492 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1649977179
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_197
timestamp 1649977179
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_209
timestamp 1649977179
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_221
timestamp 1649977179
transform 1 0 21436 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_233
timestamp 1649977179
transform 1 0 22540 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_245
timestamp 1649977179
transform 1 0 23644 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1649977179
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_253
timestamp 1649977179
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_265
timestamp 1649977179
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_277
timestamp 1649977179
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_289
timestamp 1649977179
transform 1 0 27692 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_301
timestamp 1649977179
transform 1 0 28796 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 1649977179
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_309
timestamp 1649977179
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_321
timestamp 1649977179
transform 1 0 30636 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_333
timestamp 1649977179
transform 1 0 31740 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_345
timestamp 1649977179
transform 1 0 32844 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_357
timestamp 1649977179
transform 1 0 33948 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1649977179
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_365
timestamp 1649977179
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_377
timestamp 1649977179
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_389
timestamp 1649977179
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_401
timestamp 1649977179
transform 1 0 37996 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_413
timestamp 1649977179
transform 1 0 39100 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_419
timestamp 1649977179
transform 1 0 39652 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_421
timestamp 1649977179
transform 1 0 39836 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_433
timestamp 1649977179
transform 1 0 40940 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_445
timestamp 1649977179
transform 1 0 42044 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_457
timestamp 1649977179
transform 1 0 43148 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_469
timestamp 1649977179
transform 1 0 44252 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_475
timestamp 1649977179
transform 1 0 44804 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_477
timestamp 1649977179
transform 1 0 44988 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_489
timestamp 1649977179
transform 1 0 46092 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_501
timestamp 1649977179
transform 1 0 47196 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_513
timestamp 1649977179
transform 1 0 48300 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_525
timestamp 1649977179
transform 1 0 49404 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_531
timestamp 1649977179
transform 1 0 49956 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_533
timestamp 1649977179
transform 1 0 50140 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_545
timestamp 1649977179
transform 1 0 51244 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_557
timestamp 1649977179
transform 1 0 52348 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_569
timestamp 1649977179
transform 1 0 53452 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_581
timestamp 1649977179
transform 1 0 54556 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_587
timestamp 1649977179
transform 1 0 55108 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_589
timestamp 1649977179
transform 1 0 55292 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_601
timestamp 1649977179
transform 1 0 56396 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_613
timestamp 1649977179
transform 1 0 57500 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_625
timestamp 1649977179
transform 1 0 58604 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_637
timestamp 1649977179
transform 1 0 59708 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_643
timestamp 1649977179
transform 1 0 60260 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_645
timestamp 1649977179
transform 1 0 60444 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_657
timestamp 1649977179
transform 1 0 61548 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_669
timestamp 1649977179
transform 1 0 62652 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_681
timestamp 1649977179
transform 1 0 63756 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_693
timestamp 1649977179
transform 1 0 64860 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_699
timestamp 1649977179
transform 1 0 65412 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_701
timestamp 1649977179
transform 1 0 65596 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_713
timestamp 1649977179
transform 1 0 66700 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_725
timestamp 1649977179
transform 1 0 67804 0 1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1649977179
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1649977179
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_27
timestamp 1649977179
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_39
timestamp 1649977179
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1649977179
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1649977179
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1649977179
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_69
timestamp 1649977179
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_81
timestamp 1649977179
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_93
timestamp 1649977179
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1649977179
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1649977179
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1649977179
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_125
timestamp 1649977179
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_137
timestamp 1649977179
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_149
timestamp 1649977179
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_161
timestamp 1649977179
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1649977179
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_169
timestamp 1649977179
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_181
timestamp 1649977179
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_193
timestamp 1649977179
transform 1 0 18860 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_205
timestamp 1649977179
transform 1 0 19964 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_217
timestamp 1649977179
transform 1 0 21068 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1649977179
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_225
timestamp 1649977179
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_237
timestamp 1649977179
transform 1 0 22908 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_249
timestamp 1649977179
transform 1 0 24012 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_261
timestamp 1649977179
transform 1 0 25116 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_273
timestamp 1649977179
transform 1 0 26220 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1649977179
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_281
timestamp 1649977179
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_293
timestamp 1649977179
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_305
timestamp 1649977179
transform 1 0 29164 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_317
timestamp 1649977179
transform 1 0 30268 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_329
timestamp 1649977179
transform 1 0 31372 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 1649977179
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_337
timestamp 1649977179
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_349
timestamp 1649977179
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_361
timestamp 1649977179
transform 1 0 34316 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_373
timestamp 1649977179
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_385
timestamp 1649977179
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 1649977179
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_393
timestamp 1649977179
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_405
timestamp 1649977179
transform 1 0 38364 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_417
timestamp 1649977179
transform 1 0 39468 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_429
timestamp 1649977179
transform 1 0 40572 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_441
timestamp 1649977179
transform 1 0 41676 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_447
timestamp 1649977179
transform 1 0 42228 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_449
timestamp 1649977179
transform 1 0 42412 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_461
timestamp 1649977179
transform 1 0 43516 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_473
timestamp 1649977179
transform 1 0 44620 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_485
timestamp 1649977179
transform 1 0 45724 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_497
timestamp 1649977179
transform 1 0 46828 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_503
timestamp 1649977179
transform 1 0 47380 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_505
timestamp 1649977179
transform 1 0 47564 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_517
timestamp 1649977179
transform 1 0 48668 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_529
timestamp 1649977179
transform 1 0 49772 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_541
timestamp 1649977179
transform 1 0 50876 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_553
timestamp 1649977179
transform 1 0 51980 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_559
timestamp 1649977179
transform 1 0 52532 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_561
timestamp 1649977179
transform 1 0 52716 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_573
timestamp 1649977179
transform 1 0 53820 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_585
timestamp 1649977179
transform 1 0 54924 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_597
timestamp 1649977179
transform 1 0 56028 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_609
timestamp 1649977179
transform 1 0 57132 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_615
timestamp 1649977179
transform 1 0 57684 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_617
timestamp 1649977179
transform 1 0 57868 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_629
timestamp 1649977179
transform 1 0 58972 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_641
timestamp 1649977179
transform 1 0 60076 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_653
timestamp 1649977179
transform 1 0 61180 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_665
timestamp 1649977179
transform 1 0 62284 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_671
timestamp 1649977179
transform 1 0 62836 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_673
timestamp 1649977179
transform 1 0 63020 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_685
timestamp 1649977179
transform 1 0 64124 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_697
timestamp 1649977179
transform 1 0 65228 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_709
timestamp 1649977179
transform 1 0 66332 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_721
timestamp 1649977179
transform 1 0 67436 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_727
timestamp 1649977179
transform 1 0 67988 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_729
timestamp 1649977179
transform 1 0 68172 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1649977179
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_15
timestamp 1649977179
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1649977179
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1649977179
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1649977179
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_53
timestamp 1649977179
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_65
timestamp 1649977179
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1649977179
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1649977179
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1649977179
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_97
timestamp 1649977179
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_109
timestamp 1649977179
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_121
timestamp 1649977179
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1649977179
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1649977179
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_141
timestamp 1649977179
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_153
timestamp 1649977179
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_165
timestamp 1649977179
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_177
timestamp 1649977179
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_189
timestamp 1649977179
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1649977179
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_197
timestamp 1649977179
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_209
timestamp 1649977179
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_221
timestamp 1649977179
transform 1 0 21436 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_233
timestamp 1649977179
transform 1 0 22540 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_245
timestamp 1649977179
transform 1 0 23644 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1649977179
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_253
timestamp 1649977179
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_265
timestamp 1649977179
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_277
timestamp 1649977179
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_289
timestamp 1649977179
transform 1 0 27692 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_301
timestamp 1649977179
transform 1 0 28796 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 1649977179
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_309
timestamp 1649977179
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_321
timestamp 1649977179
transform 1 0 30636 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_333
timestamp 1649977179
transform 1 0 31740 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_345
timestamp 1649977179
transform 1 0 32844 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_357
timestamp 1649977179
transform 1 0 33948 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1649977179
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_365
timestamp 1649977179
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_377
timestamp 1649977179
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_389
timestamp 1649977179
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_401
timestamp 1649977179
transform 1 0 37996 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_413
timestamp 1649977179
transform 1 0 39100 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_419
timestamp 1649977179
transform 1 0 39652 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_421
timestamp 1649977179
transform 1 0 39836 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_433
timestamp 1649977179
transform 1 0 40940 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_445
timestamp 1649977179
transform 1 0 42044 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_457
timestamp 1649977179
transform 1 0 43148 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_469
timestamp 1649977179
transform 1 0 44252 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_475
timestamp 1649977179
transform 1 0 44804 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_477
timestamp 1649977179
transform 1 0 44988 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_489
timestamp 1649977179
transform 1 0 46092 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_501
timestamp 1649977179
transform 1 0 47196 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_513
timestamp 1649977179
transform 1 0 48300 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_525
timestamp 1649977179
transform 1 0 49404 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_531
timestamp 1649977179
transform 1 0 49956 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_533
timestamp 1649977179
transform 1 0 50140 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_545
timestamp 1649977179
transform 1 0 51244 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_557
timestamp 1649977179
transform 1 0 52348 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_569
timestamp 1649977179
transform 1 0 53452 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_581
timestamp 1649977179
transform 1 0 54556 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_587
timestamp 1649977179
transform 1 0 55108 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_589
timestamp 1649977179
transform 1 0 55292 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_601
timestamp 1649977179
transform 1 0 56396 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_613
timestamp 1649977179
transform 1 0 57500 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_625
timestamp 1649977179
transform 1 0 58604 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_637
timestamp 1649977179
transform 1 0 59708 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_643
timestamp 1649977179
transform 1 0 60260 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_645
timestamp 1649977179
transform 1 0 60444 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_657
timestamp 1649977179
transform 1 0 61548 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_669
timestamp 1649977179
transform 1 0 62652 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_681
timestamp 1649977179
transform 1 0 63756 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_693
timestamp 1649977179
transform 1 0 64860 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_699
timestamp 1649977179
transform 1 0 65412 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_701
timestamp 1649977179
transform 1 0 65596 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_713
timestamp 1649977179
transform 1 0 66700 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_725
timestamp 1649977179
transform 1 0 67804 0 1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 1649977179
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_15
timestamp 1649977179
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_27
timestamp 1649977179
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_39
timestamp 1649977179
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1649977179
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1649977179
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1649977179
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_69
timestamp 1649977179
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_81
timestamp 1649977179
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_93
timestamp 1649977179
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1649977179
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1649977179
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 1649977179
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_125
timestamp 1649977179
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_137
timestamp 1649977179
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_149
timestamp 1649977179
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 1649977179
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1649977179
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_169
timestamp 1649977179
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_181
timestamp 1649977179
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_193
timestamp 1649977179
transform 1 0 18860 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_205
timestamp 1649977179
transform 1 0 19964 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_217
timestamp 1649977179
transform 1 0 21068 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1649977179
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_225
timestamp 1649977179
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_237
timestamp 1649977179
transform 1 0 22908 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_249
timestamp 1649977179
transform 1 0 24012 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_261
timestamp 1649977179
transform 1 0 25116 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_273
timestamp 1649977179
transform 1 0 26220 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1649977179
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_281
timestamp 1649977179
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_293
timestamp 1649977179
transform 1 0 28060 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_305
timestamp 1649977179
transform 1 0 29164 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_317
timestamp 1649977179
transform 1 0 30268 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_329
timestamp 1649977179
transform 1 0 31372 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1649977179
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_337
timestamp 1649977179
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_349
timestamp 1649977179
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_361
timestamp 1649977179
transform 1 0 34316 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_373
timestamp 1649977179
transform 1 0 35420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_385
timestamp 1649977179
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1649977179
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_393
timestamp 1649977179
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_405
timestamp 1649977179
transform 1 0 38364 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_417
timestamp 1649977179
transform 1 0 39468 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_429
timestamp 1649977179
transform 1 0 40572 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_441
timestamp 1649977179
transform 1 0 41676 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_447
timestamp 1649977179
transform 1 0 42228 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_449
timestamp 1649977179
transform 1 0 42412 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_461
timestamp 1649977179
transform 1 0 43516 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_473
timestamp 1649977179
transform 1 0 44620 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_485
timestamp 1649977179
transform 1 0 45724 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_497
timestamp 1649977179
transform 1 0 46828 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_503
timestamp 1649977179
transform 1 0 47380 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_505
timestamp 1649977179
transform 1 0 47564 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_517
timestamp 1649977179
transform 1 0 48668 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_529
timestamp 1649977179
transform 1 0 49772 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_541
timestamp 1649977179
transform 1 0 50876 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_553
timestamp 1649977179
transform 1 0 51980 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_559
timestamp 1649977179
transform 1 0 52532 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_561
timestamp 1649977179
transform 1 0 52716 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_573
timestamp 1649977179
transform 1 0 53820 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_585
timestamp 1649977179
transform 1 0 54924 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_597
timestamp 1649977179
transform 1 0 56028 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_609
timestamp 1649977179
transform 1 0 57132 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_615
timestamp 1649977179
transform 1 0 57684 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_617
timestamp 1649977179
transform 1 0 57868 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_629
timestamp 1649977179
transform 1 0 58972 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_641
timestamp 1649977179
transform 1 0 60076 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_653
timestamp 1649977179
transform 1 0 61180 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_665
timestamp 1649977179
transform 1 0 62284 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_671
timestamp 1649977179
transform 1 0 62836 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_673
timestamp 1649977179
transform 1 0 63020 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_685
timestamp 1649977179
transform 1 0 64124 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_697
timestamp 1649977179
transform 1 0 65228 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_709
timestamp 1649977179
transform 1 0 66332 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_721
timestamp 1649977179
transform 1 0 67436 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_727
timestamp 1649977179
transform 1 0 67988 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_729
timestamp 1649977179
transform 1 0 68172 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1649977179
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1649977179
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1649977179
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1649977179
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1649977179
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_53
timestamp 1649977179
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_65
timestamp 1649977179
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1649977179
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1649977179
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1649977179
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_97
timestamp 1649977179
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_109
timestamp 1649977179
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_121
timestamp 1649977179
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1649977179
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1649977179
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_141
timestamp 1649977179
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_153
timestamp 1649977179
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_165
timestamp 1649977179
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_177
timestamp 1649977179
transform 1 0 17388 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_189
timestamp 1649977179
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1649977179
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_197
timestamp 1649977179
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_209
timestamp 1649977179
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_221
timestamp 1649977179
transform 1 0 21436 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_233
timestamp 1649977179
transform 1 0 22540 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_245
timestamp 1649977179
transform 1 0 23644 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1649977179
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_253
timestamp 1649977179
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_265
timestamp 1649977179
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_277
timestamp 1649977179
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_289
timestamp 1649977179
transform 1 0 27692 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_301
timestamp 1649977179
transform 1 0 28796 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1649977179
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_309
timestamp 1649977179
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_321
timestamp 1649977179
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_333
timestamp 1649977179
transform 1 0 31740 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_345
timestamp 1649977179
transform 1 0 32844 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_357
timestamp 1649977179
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1649977179
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_365
timestamp 1649977179
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_377
timestamp 1649977179
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_389
timestamp 1649977179
transform 1 0 36892 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_401
timestamp 1649977179
transform 1 0 37996 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_413
timestamp 1649977179
transform 1 0 39100 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_419
timestamp 1649977179
transform 1 0 39652 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_421
timestamp 1649977179
transform 1 0 39836 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_433
timestamp 1649977179
transform 1 0 40940 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_445
timestamp 1649977179
transform 1 0 42044 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_457
timestamp 1649977179
transform 1 0 43148 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_469
timestamp 1649977179
transform 1 0 44252 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_475
timestamp 1649977179
transform 1 0 44804 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_477
timestamp 1649977179
transform 1 0 44988 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_489
timestamp 1649977179
transform 1 0 46092 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_501
timestamp 1649977179
transform 1 0 47196 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_513
timestamp 1649977179
transform 1 0 48300 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_525
timestamp 1649977179
transform 1 0 49404 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_531
timestamp 1649977179
transform 1 0 49956 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_533
timestamp 1649977179
transform 1 0 50140 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_545
timestamp 1649977179
transform 1 0 51244 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_557
timestamp 1649977179
transform 1 0 52348 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_569
timestamp 1649977179
transform 1 0 53452 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_581
timestamp 1649977179
transform 1 0 54556 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_587
timestamp 1649977179
transform 1 0 55108 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_589
timestamp 1649977179
transform 1 0 55292 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_601
timestamp 1649977179
transform 1 0 56396 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_613
timestamp 1649977179
transform 1 0 57500 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_625
timestamp 1649977179
transform 1 0 58604 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_637
timestamp 1649977179
transform 1 0 59708 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_643
timestamp 1649977179
transform 1 0 60260 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_645
timestamp 1649977179
transform 1 0 60444 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_657
timestamp 1649977179
transform 1 0 61548 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_669
timestamp 1649977179
transform 1 0 62652 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_681
timestamp 1649977179
transform 1 0 63756 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_693
timestamp 1649977179
transform 1 0 64860 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_699
timestamp 1649977179
transform 1 0 65412 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_701
timestamp 1649977179
transform 1 0 65596 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_713
timestamp 1649977179
transform 1 0 66700 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_725
timestamp 1649977179
transform 1 0 67804 0 1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_37_3
timestamp 1649977179
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_15
timestamp 1649977179
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_27
timestamp 1649977179
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_39
timestamp 1649977179
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1649977179
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1649977179
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1649977179
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_69
timestamp 1649977179
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_81
timestamp 1649977179
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_93
timestamp 1649977179
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1649977179
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1649977179
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_113
timestamp 1649977179
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_125
timestamp 1649977179
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_137
timestamp 1649977179
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_149
timestamp 1649977179
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1649977179
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1649977179
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_169
timestamp 1649977179
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_181
timestamp 1649977179
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_193
timestamp 1649977179
transform 1 0 18860 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_205
timestamp 1649977179
transform 1 0 19964 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_217
timestamp 1649977179
transform 1 0 21068 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1649977179
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_225
timestamp 1649977179
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_237
timestamp 1649977179
transform 1 0 22908 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_249
timestamp 1649977179
transform 1 0 24012 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_261
timestamp 1649977179
transform 1 0 25116 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_273
timestamp 1649977179
transform 1 0 26220 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1649977179
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_281
timestamp 1649977179
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_293
timestamp 1649977179
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_305
timestamp 1649977179
transform 1 0 29164 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_317
timestamp 1649977179
transform 1 0 30268 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_329
timestamp 1649977179
transform 1 0 31372 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1649977179
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_337
timestamp 1649977179
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_349
timestamp 1649977179
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_361
timestamp 1649977179
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_373
timestamp 1649977179
transform 1 0 35420 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_385
timestamp 1649977179
transform 1 0 36524 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 1649977179
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_393
timestamp 1649977179
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_405
timestamp 1649977179
transform 1 0 38364 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_417
timestamp 1649977179
transform 1 0 39468 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_429
timestamp 1649977179
transform 1 0 40572 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_441
timestamp 1649977179
transform 1 0 41676 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_447
timestamp 1649977179
transform 1 0 42228 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_449
timestamp 1649977179
transform 1 0 42412 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_461
timestamp 1649977179
transform 1 0 43516 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_473
timestamp 1649977179
transform 1 0 44620 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_485
timestamp 1649977179
transform 1 0 45724 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_497
timestamp 1649977179
transform 1 0 46828 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_503
timestamp 1649977179
transform 1 0 47380 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_505
timestamp 1649977179
transform 1 0 47564 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_517
timestamp 1649977179
transform 1 0 48668 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_529
timestamp 1649977179
transform 1 0 49772 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_541
timestamp 1649977179
transform 1 0 50876 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_553
timestamp 1649977179
transform 1 0 51980 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_559
timestamp 1649977179
transform 1 0 52532 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_561
timestamp 1649977179
transform 1 0 52716 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_573
timestamp 1649977179
transform 1 0 53820 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_585
timestamp 1649977179
transform 1 0 54924 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_597
timestamp 1649977179
transform 1 0 56028 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_609
timestamp 1649977179
transform 1 0 57132 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_615
timestamp 1649977179
transform 1 0 57684 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_617
timestamp 1649977179
transform 1 0 57868 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_629
timestamp 1649977179
transform 1 0 58972 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_641
timestamp 1649977179
transform 1 0 60076 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_653
timestamp 1649977179
transform 1 0 61180 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_665
timestamp 1649977179
transform 1 0 62284 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_671
timestamp 1649977179
transform 1 0 62836 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_673
timestamp 1649977179
transform 1 0 63020 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_685
timestamp 1649977179
transform 1 0 64124 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_697
timestamp 1649977179
transform 1 0 65228 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_709
timestamp 1649977179
transform 1 0 66332 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_721
timestamp 1649977179
transform 1 0 67436 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_727
timestamp 1649977179
transform 1 0 67988 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_729
timestamp 1649977179
transform 1 0 68172 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1649977179
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1649977179
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1649977179
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1649977179
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1649977179
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1649977179
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_65
timestamp 1649977179
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1649977179
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1649977179
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1649977179
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_97
timestamp 1649977179
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_109
timestamp 1649977179
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_121
timestamp 1649977179
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 1649977179
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1649977179
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_141
timestamp 1649977179
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_153
timestamp 1649977179
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_165
timestamp 1649977179
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_177
timestamp 1649977179
transform 1 0 17388 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_189
timestamp 1649977179
transform 1 0 18492 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1649977179
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_197
timestamp 1649977179
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_209
timestamp 1649977179
transform 1 0 20332 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_221
timestamp 1649977179
transform 1 0 21436 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_233
timestamp 1649977179
transform 1 0 22540 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_245
timestamp 1649977179
transform 1 0 23644 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 1649977179
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_253
timestamp 1649977179
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_265
timestamp 1649977179
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_277
timestamp 1649977179
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_289
timestamp 1649977179
transform 1 0 27692 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_301
timestamp 1649977179
transform 1 0 28796 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1649977179
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_309
timestamp 1649977179
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_321
timestamp 1649977179
transform 1 0 30636 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_333
timestamp 1649977179
transform 1 0 31740 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_345
timestamp 1649977179
transform 1 0 32844 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_357
timestamp 1649977179
transform 1 0 33948 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1649977179
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_365
timestamp 1649977179
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_377
timestamp 1649977179
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_389
timestamp 1649977179
transform 1 0 36892 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_401
timestamp 1649977179
transform 1 0 37996 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_413
timestamp 1649977179
transform 1 0 39100 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_419
timestamp 1649977179
transform 1 0 39652 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_421
timestamp 1649977179
transform 1 0 39836 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_433
timestamp 1649977179
transform 1 0 40940 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_445
timestamp 1649977179
transform 1 0 42044 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_457
timestamp 1649977179
transform 1 0 43148 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_469
timestamp 1649977179
transform 1 0 44252 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_475
timestamp 1649977179
transform 1 0 44804 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_477
timestamp 1649977179
transform 1 0 44988 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_489
timestamp 1649977179
transform 1 0 46092 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_501
timestamp 1649977179
transform 1 0 47196 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_513
timestamp 1649977179
transform 1 0 48300 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_525
timestamp 1649977179
transform 1 0 49404 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_531
timestamp 1649977179
transform 1 0 49956 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_533
timestamp 1649977179
transform 1 0 50140 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_545
timestamp 1649977179
transform 1 0 51244 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_557
timestamp 1649977179
transform 1 0 52348 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_569
timestamp 1649977179
transform 1 0 53452 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_581
timestamp 1649977179
transform 1 0 54556 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_587
timestamp 1649977179
transform 1 0 55108 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_589
timestamp 1649977179
transform 1 0 55292 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_601
timestamp 1649977179
transform 1 0 56396 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_613
timestamp 1649977179
transform 1 0 57500 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_625
timestamp 1649977179
transform 1 0 58604 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_637
timestamp 1649977179
transform 1 0 59708 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_643
timestamp 1649977179
transform 1 0 60260 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_645
timestamp 1649977179
transform 1 0 60444 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_657
timestamp 1649977179
transform 1 0 61548 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_669
timestamp 1649977179
transform 1 0 62652 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_681
timestamp 1649977179
transform 1 0 63756 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_693
timestamp 1649977179
transform 1 0 64860 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_699
timestamp 1649977179
transform 1 0 65412 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_701
timestamp 1649977179
transform 1 0 65596 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_713
timestamp 1649977179
transform 1 0 66700 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_725
timestamp 1649977179
transform 1 0 67804 0 1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1649977179
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_15
timestamp 1649977179
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_27
timestamp 1649977179
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_39
timestamp 1649977179
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1649977179
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1649977179
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1649977179
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_69
timestamp 1649977179
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_81
timestamp 1649977179
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_93
timestamp 1649977179
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1649977179
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1649977179
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_113
timestamp 1649977179
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_125
timestamp 1649977179
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_137
timestamp 1649977179
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_149
timestamp 1649977179
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1649977179
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1649977179
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_169
timestamp 1649977179
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_181
timestamp 1649977179
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_193
timestamp 1649977179
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_205
timestamp 1649977179
transform 1 0 19964 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_217
timestamp 1649977179
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1649977179
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_225
timestamp 1649977179
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_237
timestamp 1649977179
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_249
timestamp 1649977179
transform 1 0 24012 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_261
timestamp 1649977179
transform 1 0 25116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_273
timestamp 1649977179
transform 1 0 26220 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1649977179
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_281
timestamp 1649977179
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_293
timestamp 1649977179
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_305
timestamp 1649977179
transform 1 0 29164 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_317
timestamp 1649977179
transform 1 0 30268 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_329
timestamp 1649977179
transform 1 0 31372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 1649977179
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_337
timestamp 1649977179
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_349
timestamp 1649977179
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_361
timestamp 1649977179
transform 1 0 34316 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_373
timestamp 1649977179
transform 1 0 35420 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_385
timestamp 1649977179
transform 1 0 36524 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1649977179
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_393
timestamp 1649977179
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_405
timestamp 1649977179
transform 1 0 38364 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_417
timestamp 1649977179
transform 1 0 39468 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_429
timestamp 1649977179
transform 1 0 40572 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_441
timestamp 1649977179
transform 1 0 41676 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_447
timestamp 1649977179
transform 1 0 42228 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_449
timestamp 1649977179
transform 1 0 42412 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_461
timestamp 1649977179
transform 1 0 43516 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_473
timestamp 1649977179
transform 1 0 44620 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_485
timestamp 1649977179
transform 1 0 45724 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_497
timestamp 1649977179
transform 1 0 46828 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_503
timestamp 1649977179
transform 1 0 47380 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_505
timestamp 1649977179
transform 1 0 47564 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_517
timestamp 1649977179
transform 1 0 48668 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_529
timestamp 1649977179
transform 1 0 49772 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_541
timestamp 1649977179
transform 1 0 50876 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_553
timestamp 1649977179
transform 1 0 51980 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_559
timestamp 1649977179
transform 1 0 52532 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_561
timestamp 1649977179
transform 1 0 52716 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_573
timestamp 1649977179
transform 1 0 53820 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_585
timestamp 1649977179
transform 1 0 54924 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_597
timestamp 1649977179
transform 1 0 56028 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_609
timestamp 1649977179
transform 1 0 57132 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_615
timestamp 1649977179
transform 1 0 57684 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_617
timestamp 1649977179
transform 1 0 57868 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_629
timestamp 1649977179
transform 1 0 58972 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_641
timestamp 1649977179
transform 1 0 60076 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_653
timestamp 1649977179
transform 1 0 61180 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_665
timestamp 1649977179
transform 1 0 62284 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_671
timestamp 1649977179
transform 1 0 62836 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_673
timestamp 1649977179
transform 1 0 63020 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_685
timestamp 1649977179
transform 1 0 64124 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_697
timestamp 1649977179
transform 1 0 65228 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_709
timestamp 1649977179
transform 1 0 66332 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_721
timestamp 1649977179
transform 1 0 67436 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_727
timestamp 1649977179
transform 1 0 67988 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_729
timestamp 1649977179
transform 1 0 68172 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_3
timestamp 1649977179
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_15
timestamp 1649977179
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1649977179
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1649977179
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1649977179
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1649977179
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_65
timestamp 1649977179
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1649977179
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1649977179
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 1649977179
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_97
timestamp 1649977179
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_109
timestamp 1649977179
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_121
timestamp 1649977179
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1649977179
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1649977179
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_141
timestamp 1649977179
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_153
timestamp 1649977179
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_165
timestamp 1649977179
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_177
timestamp 1649977179
transform 1 0 17388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_189
timestamp 1649977179
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1649977179
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_197
timestamp 1649977179
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_209
timestamp 1649977179
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_221
timestamp 1649977179
transform 1 0 21436 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_233
timestamp 1649977179
transform 1 0 22540 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_245
timestamp 1649977179
transform 1 0 23644 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1649977179
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_253
timestamp 1649977179
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_265
timestamp 1649977179
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_277
timestamp 1649977179
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_289
timestamp 1649977179
transform 1 0 27692 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_301
timestamp 1649977179
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 1649977179
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_309
timestamp 1649977179
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_321
timestamp 1649977179
transform 1 0 30636 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_333
timestamp 1649977179
transform 1 0 31740 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_345
timestamp 1649977179
transform 1 0 32844 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_357
timestamp 1649977179
transform 1 0 33948 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 1649977179
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_365
timestamp 1649977179
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_377
timestamp 1649977179
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_389
timestamp 1649977179
transform 1 0 36892 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_401
timestamp 1649977179
transform 1 0 37996 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_413
timestamp 1649977179
transform 1 0 39100 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_419
timestamp 1649977179
transform 1 0 39652 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_421
timestamp 1649977179
transform 1 0 39836 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_433
timestamp 1649977179
transform 1 0 40940 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_445
timestamp 1649977179
transform 1 0 42044 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_457
timestamp 1649977179
transform 1 0 43148 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_469
timestamp 1649977179
transform 1 0 44252 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_475
timestamp 1649977179
transform 1 0 44804 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_477
timestamp 1649977179
transform 1 0 44988 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_489
timestamp 1649977179
transform 1 0 46092 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_501
timestamp 1649977179
transform 1 0 47196 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_513
timestamp 1649977179
transform 1 0 48300 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_525
timestamp 1649977179
transform 1 0 49404 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_531
timestamp 1649977179
transform 1 0 49956 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_533
timestamp 1649977179
transform 1 0 50140 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_545
timestamp 1649977179
transform 1 0 51244 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_557
timestamp 1649977179
transform 1 0 52348 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_569
timestamp 1649977179
transform 1 0 53452 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_581
timestamp 1649977179
transform 1 0 54556 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_587
timestamp 1649977179
transform 1 0 55108 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_589
timestamp 1649977179
transform 1 0 55292 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_601
timestamp 1649977179
transform 1 0 56396 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_613
timestamp 1649977179
transform 1 0 57500 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_625
timestamp 1649977179
transform 1 0 58604 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_637
timestamp 1649977179
transform 1 0 59708 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_643
timestamp 1649977179
transform 1 0 60260 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_645
timestamp 1649977179
transform 1 0 60444 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_657
timestamp 1649977179
transform 1 0 61548 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_669
timestamp 1649977179
transform 1 0 62652 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_681
timestamp 1649977179
transform 1 0 63756 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_693
timestamp 1649977179
transform 1 0 64860 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_699
timestamp 1649977179
transform 1 0 65412 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_701
timestamp 1649977179
transform 1 0 65596 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_713
timestamp 1649977179
transform 1 0 66700 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_725
timestamp 1649977179
transform 1 0 67804 0 1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_41_3
timestamp 1649977179
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_15
timestamp 1649977179
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_27
timestamp 1649977179
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_39
timestamp 1649977179
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1649977179
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1649977179
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1649977179
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_69
timestamp 1649977179
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_81
timestamp 1649977179
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_93
timestamp 1649977179
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1649977179
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1649977179
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_113
timestamp 1649977179
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_125
timestamp 1649977179
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_137
timestamp 1649977179
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_149
timestamp 1649977179
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 1649977179
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1649977179
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_169
timestamp 1649977179
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_181
timestamp 1649977179
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_193
timestamp 1649977179
transform 1 0 18860 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_205
timestamp 1649977179
transform 1 0 19964 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_217
timestamp 1649977179
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1649977179
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_225
timestamp 1649977179
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_237
timestamp 1649977179
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_249
timestamp 1649977179
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_261
timestamp 1649977179
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_273
timestamp 1649977179
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1649977179
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_281
timestamp 1649977179
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_293
timestamp 1649977179
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_305
timestamp 1649977179
transform 1 0 29164 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_317
timestamp 1649977179
transform 1 0 30268 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_329
timestamp 1649977179
transform 1 0 31372 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1649977179
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_337
timestamp 1649977179
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_349
timestamp 1649977179
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_361
timestamp 1649977179
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_373
timestamp 1649977179
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_385
timestamp 1649977179
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 1649977179
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_393
timestamp 1649977179
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_405
timestamp 1649977179
transform 1 0 38364 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_417
timestamp 1649977179
transform 1 0 39468 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_429
timestamp 1649977179
transform 1 0 40572 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_441
timestamp 1649977179
transform 1 0 41676 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_447
timestamp 1649977179
transform 1 0 42228 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_449
timestamp 1649977179
transform 1 0 42412 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_461
timestamp 1649977179
transform 1 0 43516 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_473
timestamp 1649977179
transform 1 0 44620 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_485
timestamp 1649977179
transform 1 0 45724 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_497
timestamp 1649977179
transform 1 0 46828 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_503
timestamp 1649977179
transform 1 0 47380 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_505
timestamp 1649977179
transform 1 0 47564 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_517
timestamp 1649977179
transform 1 0 48668 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_529
timestamp 1649977179
transform 1 0 49772 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_541
timestamp 1649977179
transform 1 0 50876 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_553
timestamp 1649977179
transform 1 0 51980 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_559
timestamp 1649977179
transform 1 0 52532 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_561
timestamp 1649977179
transform 1 0 52716 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_573
timestamp 1649977179
transform 1 0 53820 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_585
timestamp 1649977179
transform 1 0 54924 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_597
timestamp 1649977179
transform 1 0 56028 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_609
timestamp 1649977179
transform 1 0 57132 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_615
timestamp 1649977179
transform 1 0 57684 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_617
timestamp 1649977179
transform 1 0 57868 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_629
timestamp 1649977179
transform 1 0 58972 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_641
timestamp 1649977179
transform 1 0 60076 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_653
timestamp 1649977179
transform 1 0 61180 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_665
timestamp 1649977179
transform 1 0 62284 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_671
timestamp 1649977179
transform 1 0 62836 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_673
timestamp 1649977179
transform 1 0 63020 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_685
timestamp 1649977179
transform 1 0 64124 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_697
timestamp 1649977179
transform 1 0 65228 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_709
timestamp 1649977179
transform 1 0 66332 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_721
timestamp 1649977179
transform 1 0 67436 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_727
timestamp 1649977179
transform 1 0 67988 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_729
timestamp 1649977179
transform 1 0 68172 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1649977179
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1649977179
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1649977179
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1649977179
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1649977179
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_53
timestamp 1649977179
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_65
timestamp 1649977179
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1649977179
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1649977179
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_85
timestamp 1649977179
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_97
timestamp 1649977179
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_109
timestamp 1649977179
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_121
timestamp 1649977179
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp 1649977179
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1649977179
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_141
timestamp 1649977179
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_153
timestamp 1649977179
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_165
timestamp 1649977179
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_177
timestamp 1649977179
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_189
timestamp 1649977179
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1649977179
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_197
timestamp 1649977179
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_209
timestamp 1649977179
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_221
timestamp 1649977179
transform 1 0 21436 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_233
timestamp 1649977179
transform 1 0 22540 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_245
timestamp 1649977179
transform 1 0 23644 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1649977179
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_253
timestamp 1649977179
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_265
timestamp 1649977179
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_277
timestamp 1649977179
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_289
timestamp 1649977179
transform 1 0 27692 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_301
timestamp 1649977179
transform 1 0 28796 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1649977179
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_309
timestamp 1649977179
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_321
timestamp 1649977179
transform 1 0 30636 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_333
timestamp 1649977179
transform 1 0 31740 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_345
timestamp 1649977179
transform 1 0 32844 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_357
timestamp 1649977179
transform 1 0 33948 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_363
timestamp 1649977179
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_365
timestamp 1649977179
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_377
timestamp 1649977179
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_389
timestamp 1649977179
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_401
timestamp 1649977179
transform 1 0 37996 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_413
timestamp 1649977179
transform 1 0 39100 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_419
timestamp 1649977179
transform 1 0 39652 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_421
timestamp 1649977179
transform 1 0 39836 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_433
timestamp 1649977179
transform 1 0 40940 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_445
timestamp 1649977179
transform 1 0 42044 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_457
timestamp 1649977179
transform 1 0 43148 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_469
timestamp 1649977179
transform 1 0 44252 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_475
timestamp 1649977179
transform 1 0 44804 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_477
timestamp 1649977179
transform 1 0 44988 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_489
timestamp 1649977179
transform 1 0 46092 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_501
timestamp 1649977179
transform 1 0 47196 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_513
timestamp 1649977179
transform 1 0 48300 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_525
timestamp 1649977179
transform 1 0 49404 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_531
timestamp 1649977179
transform 1 0 49956 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_533
timestamp 1649977179
transform 1 0 50140 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_545
timestamp 1649977179
transform 1 0 51244 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_557
timestamp 1649977179
transform 1 0 52348 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_569
timestamp 1649977179
transform 1 0 53452 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_581
timestamp 1649977179
transform 1 0 54556 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_587
timestamp 1649977179
transform 1 0 55108 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_589
timestamp 1649977179
transform 1 0 55292 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_601
timestamp 1649977179
transform 1 0 56396 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_613
timestamp 1649977179
transform 1 0 57500 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_625
timestamp 1649977179
transform 1 0 58604 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_637
timestamp 1649977179
transform 1 0 59708 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_643
timestamp 1649977179
transform 1 0 60260 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_645
timestamp 1649977179
transform 1 0 60444 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_657
timestamp 1649977179
transform 1 0 61548 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_669
timestamp 1649977179
transform 1 0 62652 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_681
timestamp 1649977179
transform 1 0 63756 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_693
timestamp 1649977179
transform 1 0 64860 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_699
timestamp 1649977179
transform 1 0 65412 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_701
timestamp 1649977179
transform 1 0 65596 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_713
timestamp 1649977179
transform 1 0 66700 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_725
timestamp 1649977179
transform 1 0 67804 0 1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1649977179
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1649977179
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_27
timestamp 1649977179
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_39
timestamp 1649977179
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1649977179
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1649977179
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1649977179
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_69
timestamp 1649977179
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_81
timestamp 1649977179
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_93
timestamp 1649977179
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1649977179
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1649977179
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_113
timestamp 1649977179
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_125
timestamp 1649977179
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_137
timestamp 1649977179
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_149
timestamp 1649977179
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_161
timestamp 1649977179
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1649977179
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_169
timestamp 1649977179
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_181
timestamp 1649977179
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_193
timestamp 1649977179
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_205
timestamp 1649977179
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_217
timestamp 1649977179
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1649977179
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_225
timestamp 1649977179
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_237
timestamp 1649977179
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_249
timestamp 1649977179
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_261
timestamp 1649977179
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_273
timestamp 1649977179
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1649977179
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_281
timestamp 1649977179
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_293
timestamp 1649977179
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_305
timestamp 1649977179
transform 1 0 29164 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_317
timestamp 1649977179
transform 1 0 30268 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_329
timestamp 1649977179
transform 1 0 31372 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1649977179
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_337
timestamp 1649977179
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_349
timestamp 1649977179
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_361
timestamp 1649977179
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_373
timestamp 1649977179
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_385
timestamp 1649977179
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1649977179
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_393
timestamp 1649977179
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_405
timestamp 1649977179
transform 1 0 38364 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_417
timestamp 1649977179
transform 1 0 39468 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_429
timestamp 1649977179
transform 1 0 40572 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_441
timestamp 1649977179
transform 1 0 41676 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_447
timestamp 1649977179
transform 1 0 42228 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_449
timestamp 1649977179
transform 1 0 42412 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_461
timestamp 1649977179
transform 1 0 43516 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_473
timestamp 1649977179
transform 1 0 44620 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_485
timestamp 1649977179
transform 1 0 45724 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_497
timestamp 1649977179
transform 1 0 46828 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_503
timestamp 1649977179
transform 1 0 47380 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_505
timestamp 1649977179
transform 1 0 47564 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_517
timestamp 1649977179
transform 1 0 48668 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_529
timestamp 1649977179
transform 1 0 49772 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_541
timestamp 1649977179
transform 1 0 50876 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_553
timestamp 1649977179
transform 1 0 51980 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_559
timestamp 1649977179
transform 1 0 52532 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_561
timestamp 1649977179
transform 1 0 52716 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_573
timestamp 1649977179
transform 1 0 53820 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_585
timestamp 1649977179
transform 1 0 54924 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_597
timestamp 1649977179
transform 1 0 56028 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_609
timestamp 1649977179
transform 1 0 57132 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_615
timestamp 1649977179
transform 1 0 57684 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_617
timestamp 1649977179
transform 1 0 57868 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_629
timestamp 1649977179
transform 1 0 58972 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_641
timestamp 1649977179
transform 1 0 60076 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_653
timestamp 1649977179
transform 1 0 61180 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_665
timestamp 1649977179
transform 1 0 62284 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_671
timestamp 1649977179
transform 1 0 62836 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_673
timestamp 1649977179
transform 1 0 63020 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_685
timestamp 1649977179
transform 1 0 64124 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_697
timestamp 1649977179
transform 1 0 65228 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_709
timestamp 1649977179
transform 1 0 66332 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_721
timestamp 1649977179
transform 1 0 67436 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_727
timestamp 1649977179
transform 1 0 67988 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_729
timestamp 1649977179
transform 1 0 68172 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1649977179
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_15
timestamp 1649977179
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1649977179
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1649977179
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1649977179
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1649977179
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_65
timestamp 1649977179
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1649977179
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1649977179
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_85
timestamp 1649977179
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_97
timestamp 1649977179
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_109
timestamp 1649977179
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_121
timestamp 1649977179
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1649977179
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1649977179
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_141
timestamp 1649977179
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_153
timestamp 1649977179
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_165
timestamp 1649977179
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_177
timestamp 1649977179
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_189
timestamp 1649977179
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1649977179
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_197
timestamp 1649977179
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_209
timestamp 1649977179
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_221
timestamp 1649977179
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_233
timestamp 1649977179
transform 1 0 22540 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_245
timestamp 1649977179
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1649977179
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_253
timestamp 1649977179
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_265
timestamp 1649977179
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_277
timestamp 1649977179
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_289
timestamp 1649977179
transform 1 0 27692 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_301
timestamp 1649977179
transform 1 0 28796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1649977179
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_309
timestamp 1649977179
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_321
timestamp 1649977179
transform 1 0 30636 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_333
timestamp 1649977179
transform 1 0 31740 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_345
timestamp 1649977179
transform 1 0 32844 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_357
timestamp 1649977179
transform 1 0 33948 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1649977179
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_365
timestamp 1649977179
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_377
timestamp 1649977179
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_389
timestamp 1649977179
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_401
timestamp 1649977179
transform 1 0 37996 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_413
timestamp 1649977179
transform 1 0 39100 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_419
timestamp 1649977179
transform 1 0 39652 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_421
timestamp 1649977179
transform 1 0 39836 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_433
timestamp 1649977179
transform 1 0 40940 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_445
timestamp 1649977179
transform 1 0 42044 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_457
timestamp 1649977179
transform 1 0 43148 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_469
timestamp 1649977179
transform 1 0 44252 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_475
timestamp 1649977179
transform 1 0 44804 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_477
timestamp 1649977179
transform 1 0 44988 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_489
timestamp 1649977179
transform 1 0 46092 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_501
timestamp 1649977179
transform 1 0 47196 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_513
timestamp 1649977179
transform 1 0 48300 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_525
timestamp 1649977179
transform 1 0 49404 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_531
timestamp 1649977179
transform 1 0 49956 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_533
timestamp 1649977179
transform 1 0 50140 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_545
timestamp 1649977179
transform 1 0 51244 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_557
timestamp 1649977179
transform 1 0 52348 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_569
timestamp 1649977179
transform 1 0 53452 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_581
timestamp 1649977179
transform 1 0 54556 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_587
timestamp 1649977179
transform 1 0 55108 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_589
timestamp 1649977179
transform 1 0 55292 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_601
timestamp 1649977179
transform 1 0 56396 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_613
timestamp 1649977179
transform 1 0 57500 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_625
timestamp 1649977179
transform 1 0 58604 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_637
timestamp 1649977179
transform 1 0 59708 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_643
timestamp 1649977179
transform 1 0 60260 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_645
timestamp 1649977179
transform 1 0 60444 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_657
timestamp 1649977179
transform 1 0 61548 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_669
timestamp 1649977179
transform 1 0 62652 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_681
timestamp 1649977179
transform 1 0 63756 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_693
timestamp 1649977179
transform 1 0 64860 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_699
timestamp 1649977179
transform 1 0 65412 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_701
timestamp 1649977179
transform 1 0 65596 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_713
timestamp 1649977179
transform 1 0 66700 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_725
timestamp 1649977179
transform 1 0 67804 0 1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1649977179
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_15
timestamp 1649977179
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_27
timestamp 1649977179
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_39
timestamp 1649977179
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1649977179
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1649977179
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1649977179
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_69
timestamp 1649977179
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_81
timestamp 1649977179
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_93
timestamp 1649977179
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1649977179
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1649977179
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_113
timestamp 1649977179
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_125
timestamp 1649977179
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_137
timestamp 1649977179
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_149
timestamp 1649977179
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp 1649977179
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1649977179
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_169
timestamp 1649977179
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_181
timestamp 1649977179
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_193
timestamp 1649977179
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_205
timestamp 1649977179
transform 1 0 19964 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_217
timestamp 1649977179
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1649977179
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_225
timestamp 1649977179
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_237
timestamp 1649977179
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_249
timestamp 1649977179
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_261
timestamp 1649977179
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_273
timestamp 1649977179
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1649977179
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_281
timestamp 1649977179
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_293
timestamp 1649977179
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_305
timestamp 1649977179
transform 1 0 29164 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_317
timestamp 1649977179
transform 1 0 30268 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_329
timestamp 1649977179
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1649977179
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_337
timestamp 1649977179
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_349
timestamp 1649977179
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_361
timestamp 1649977179
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_373
timestamp 1649977179
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_385
timestamp 1649977179
transform 1 0 36524 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1649977179
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_393
timestamp 1649977179
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_405
timestamp 1649977179
transform 1 0 38364 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_417
timestamp 1649977179
transform 1 0 39468 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_429
timestamp 1649977179
transform 1 0 40572 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_441
timestamp 1649977179
transform 1 0 41676 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_447
timestamp 1649977179
transform 1 0 42228 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_449
timestamp 1649977179
transform 1 0 42412 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_461
timestamp 1649977179
transform 1 0 43516 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_473
timestamp 1649977179
transform 1 0 44620 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_485
timestamp 1649977179
transform 1 0 45724 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_497
timestamp 1649977179
transform 1 0 46828 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_503
timestamp 1649977179
transform 1 0 47380 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_505
timestamp 1649977179
transform 1 0 47564 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_517
timestamp 1649977179
transform 1 0 48668 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_529
timestamp 1649977179
transform 1 0 49772 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_541
timestamp 1649977179
transform 1 0 50876 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_553
timestamp 1649977179
transform 1 0 51980 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_559
timestamp 1649977179
transform 1 0 52532 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_561
timestamp 1649977179
transform 1 0 52716 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_573
timestamp 1649977179
transform 1 0 53820 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_585
timestamp 1649977179
transform 1 0 54924 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_597
timestamp 1649977179
transform 1 0 56028 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_609
timestamp 1649977179
transform 1 0 57132 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_615
timestamp 1649977179
transform 1 0 57684 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_617
timestamp 1649977179
transform 1 0 57868 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_629
timestamp 1649977179
transform 1 0 58972 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_641
timestamp 1649977179
transform 1 0 60076 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_653
timestamp 1649977179
transform 1 0 61180 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_665
timestamp 1649977179
transform 1 0 62284 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_671
timestamp 1649977179
transform 1 0 62836 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_673
timestamp 1649977179
transform 1 0 63020 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_685
timestamp 1649977179
transform 1 0 64124 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_697
timestamp 1649977179
transform 1 0 65228 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_709
timestamp 1649977179
transform 1 0 66332 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_721
timestamp 1649977179
transform 1 0 67436 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_727
timestamp 1649977179
transform 1 0 67988 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_729
timestamp 1649977179
transform 1 0 68172 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1649977179
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1649977179
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1649977179
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1649977179
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1649977179
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_53
timestamp 1649977179
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_65
timestamp 1649977179
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1649977179
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1649977179
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_85
timestamp 1649977179
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_97
timestamp 1649977179
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_109
timestamp 1649977179
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_121
timestamp 1649977179
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1649977179
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1649977179
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_141
timestamp 1649977179
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_153
timestamp 1649977179
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_165
timestamp 1649977179
transform 1 0 16284 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_177
timestamp 1649977179
transform 1 0 17388 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_189
timestamp 1649977179
transform 1 0 18492 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1649977179
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_197
timestamp 1649977179
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_209
timestamp 1649977179
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_221
timestamp 1649977179
transform 1 0 21436 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_233
timestamp 1649977179
transform 1 0 22540 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_245
timestamp 1649977179
transform 1 0 23644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1649977179
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_253
timestamp 1649977179
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_265
timestamp 1649977179
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_277
timestamp 1649977179
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_289
timestamp 1649977179
transform 1 0 27692 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_301
timestamp 1649977179
transform 1 0 28796 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 1649977179
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_309
timestamp 1649977179
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_321
timestamp 1649977179
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_333
timestamp 1649977179
transform 1 0 31740 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_345
timestamp 1649977179
transform 1 0 32844 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_357
timestamp 1649977179
transform 1 0 33948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1649977179
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_365
timestamp 1649977179
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_377
timestamp 1649977179
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_389
timestamp 1649977179
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_401
timestamp 1649977179
transform 1 0 37996 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_413
timestamp 1649977179
transform 1 0 39100 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_419
timestamp 1649977179
transform 1 0 39652 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_421
timestamp 1649977179
transform 1 0 39836 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_433
timestamp 1649977179
transform 1 0 40940 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_445
timestamp 1649977179
transform 1 0 42044 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_457
timestamp 1649977179
transform 1 0 43148 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_469
timestamp 1649977179
transform 1 0 44252 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_475
timestamp 1649977179
transform 1 0 44804 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_477
timestamp 1649977179
transform 1 0 44988 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_489
timestamp 1649977179
transform 1 0 46092 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_501
timestamp 1649977179
transform 1 0 47196 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_513
timestamp 1649977179
transform 1 0 48300 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_525
timestamp 1649977179
transform 1 0 49404 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_531
timestamp 1649977179
transform 1 0 49956 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_533
timestamp 1649977179
transform 1 0 50140 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_545
timestamp 1649977179
transform 1 0 51244 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_557
timestamp 1649977179
transform 1 0 52348 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_569
timestamp 1649977179
transform 1 0 53452 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_581
timestamp 1649977179
transform 1 0 54556 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_587
timestamp 1649977179
transform 1 0 55108 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_589
timestamp 1649977179
transform 1 0 55292 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_601
timestamp 1649977179
transform 1 0 56396 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_613
timestamp 1649977179
transform 1 0 57500 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_625
timestamp 1649977179
transform 1 0 58604 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_637
timestamp 1649977179
transform 1 0 59708 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_643
timestamp 1649977179
transform 1 0 60260 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_645
timestamp 1649977179
transform 1 0 60444 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_657
timestamp 1649977179
transform 1 0 61548 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_669
timestamp 1649977179
transform 1 0 62652 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_681
timestamp 1649977179
transform 1 0 63756 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_693
timestamp 1649977179
transform 1 0 64860 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_699
timestamp 1649977179
transform 1 0 65412 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_701
timestamp 1649977179
transform 1 0 65596 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_713
timestamp 1649977179
transform 1 0 66700 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_725
timestamp 1649977179
transform 1 0 67804 0 1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_47_3
timestamp 1649977179
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_15
timestamp 1649977179
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_27
timestamp 1649977179
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_39
timestamp 1649977179
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1649977179
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1649977179
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1649977179
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_69
timestamp 1649977179
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_81
timestamp 1649977179
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_93
timestamp 1649977179
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 1649977179
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1649977179
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_113
timestamp 1649977179
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_125
timestamp 1649977179
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_137
timestamp 1649977179
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_149
timestamp 1649977179
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_161
timestamp 1649977179
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1649977179
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_169
timestamp 1649977179
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_181
timestamp 1649977179
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_193
timestamp 1649977179
transform 1 0 18860 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_205
timestamp 1649977179
transform 1 0 19964 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_217
timestamp 1649977179
transform 1 0 21068 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1649977179
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_225
timestamp 1649977179
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_237
timestamp 1649977179
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_249
timestamp 1649977179
transform 1 0 24012 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_261
timestamp 1649977179
transform 1 0 25116 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_273
timestamp 1649977179
transform 1 0 26220 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 1649977179
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_281
timestamp 1649977179
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_293
timestamp 1649977179
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_305
timestamp 1649977179
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_317
timestamp 1649977179
transform 1 0 30268 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_329
timestamp 1649977179
transform 1 0 31372 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 1649977179
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_337
timestamp 1649977179
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_349
timestamp 1649977179
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_361
timestamp 1649977179
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_373
timestamp 1649977179
transform 1 0 35420 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_385
timestamp 1649977179
transform 1 0 36524 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_391
timestamp 1649977179
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_393
timestamp 1649977179
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_405
timestamp 1649977179
transform 1 0 38364 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_417
timestamp 1649977179
transform 1 0 39468 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_429
timestamp 1649977179
transform 1 0 40572 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_441
timestamp 1649977179
transform 1 0 41676 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_447
timestamp 1649977179
transform 1 0 42228 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_449
timestamp 1649977179
transform 1 0 42412 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_461
timestamp 1649977179
transform 1 0 43516 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_473
timestamp 1649977179
transform 1 0 44620 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_485
timestamp 1649977179
transform 1 0 45724 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_497
timestamp 1649977179
transform 1 0 46828 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_503
timestamp 1649977179
transform 1 0 47380 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_505
timestamp 1649977179
transform 1 0 47564 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_517
timestamp 1649977179
transform 1 0 48668 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_529
timestamp 1649977179
transform 1 0 49772 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_541
timestamp 1649977179
transform 1 0 50876 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_553
timestamp 1649977179
transform 1 0 51980 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_559
timestamp 1649977179
transform 1 0 52532 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_561
timestamp 1649977179
transform 1 0 52716 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_573
timestamp 1649977179
transform 1 0 53820 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_585
timestamp 1649977179
transform 1 0 54924 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_597
timestamp 1649977179
transform 1 0 56028 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_609
timestamp 1649977179
transform 1 0 57132 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_615
timestamp 1649977179
transform 1 0 57684 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_617
timestamp 1649977179
transform 1 0 57868 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_629
timestamp 1649977179
transform 1 0 58972 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_641
timestamp 1649977179
transform 1 0 60076 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_653
timestamp 1649977179
transform 1 0 61180 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_665
timestamp 1649977179
transform 1 0 62284 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_671
timestamp 1649977179
transform 1 0 62836 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_673
timestamp 1649977179
transform 1 0 63020 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_685
timestamp 1649977179
transform 1 0 64124 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_697
timestamp 1649977179
transform 1 0 65228 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_709
timestamp 1649977179
transform 1 0 66332 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_721
timestamp 1649977179
transform 1 0 67436 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_727
timestamp 1649977179
transform 1 0 67988 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_729
timestamp 1649977179
transform 1 0 68172 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1649977179
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1649977179
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1649977179
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1649977179
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_41
timestamp 1649977179
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_53
timestamp 1649977179
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_65
timestamp 1649977179
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1649977179
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1649977179
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_85
timestamp 1649977179
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_97
timestamp 1649977179
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_109
timestamp 1649977179
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_121
timestamp 1649977179
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1649977179
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1649977179
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_141
timestamp 1649977179
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_153
timestamp 1649977179
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_165
timestamp 1649977179
transform 1 0 16284 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_177
timestamp 1649977179
transform 1 0 17388 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_189
timestamp 1649977179
transform 1 0 18492 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1649977179
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_197
timestamp 1649977179
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_209
timestamp 1649977179
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_221
timestamp 1649977179
transform 1 0 21436 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_233
timestamp 1649977179
transform 1 0 22540 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_245
timestamp 1649977179
transform 1 0 23644 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1649977179
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_253
timestamp 1649977179
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_265
timestamp 1649977179
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_277
timestamp 1649977179
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_289
timestamp 1649977179
transform 1 0 27692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_301
timestamp 1649977179
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 1649977179
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_309
timestamp 1649977179
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_321
timestamp 1649977179
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_333
timestamp 1649977179
transform 1 0 31740 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_345
timestamp 1649977179
transform 1 0 32844 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_357
timestamp 1649977179
transform 1 0 33948 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 1649977179
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_365
timestamp 1649977179
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_377
timestamp 1649977179
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_389
timestamp 1649977179
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_401
timestamp 1649977179
transform 1 0 37996 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_413
timestamp 1649977179
transform 1 0 39100 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_419
timestamp 1649977179
transform 1 0 39652 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_421
timestamp 1649977179
transform 1 0 39836 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_433
timestamp 1649977179
transform 1 0 40940 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_445
timestamp 1649977179
transform 1 0 42044 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_457
timestamp 1649977179
transform 1 0 43148 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_469
timestamp 1649977179
transform 1 0 44252 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_475
timestamp 1649977179
transform 1 0 44804 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_477
timestamp 1649977179
transform 1 0 44988 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_489
timestamp 1649977179
transform 1 0 46092 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_501
timestamp 1649977179
transform 1 0 47196 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_513
timestamp 1649977179
transform 1 0 48300 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_525
timestamp 1649977179
transform 1 0 49404 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_531
timestamp 1649977179
transform 1 0 49956 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_533
timestamp 1649977179
transform 1 0 50140 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_545
timestamp 1649977179
transform 1 0 51244 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_557
timestamp 1649977179
transform 1 0 52348 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_569
timestamp 1649977179
transform 1 0 53452 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_581
timestamp 1649977179
transform 1 0 54556 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_587
timestamp 1649977179
transform 1 0 55108 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_589
timestamp 1649977179
transform 1 0 55292 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_601
timestamp 1649977179
transform 1 0 56396 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_613
timestamp 1649977179
transform 1 0 57500 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_625
timestamp 1649977179
transform 1 0 58604 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_637
timestamp 1649977179
transform 1 0 59708 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_643
timestamp 1649977179
transform 1 0 60260 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_645
timestamp 1649977179
transform 1 0 60444 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_657
timestamp 1649977179
transform 1 0 61548 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_669
timestamp 1649977179
transform 1 0 62652 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_681
timestamp 1649977179
transform 1 0 63756 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_693
timestamp 1649977179
transform 1 0 64860 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_699
timestamp 1649977179
transform 1 0 65412 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_701
timestamp 1649977179
transform 1 0 65596 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_713
timestamp 1649977179
transform 1 0 66700 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_725
timestamp 1649977179
transform 1 0 67804 0 1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1649977179
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 1649977179
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_27
timestamp 1649977179
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_39
timestamp 1649977179
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1649977179
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1649977179
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1649977179
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_69
timestamp 1649977179
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_81
timestamp 1649977179
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_93
timestamp 1649977179
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1649977179
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1649977179
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_113
timestamp 1649977179
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_125
timestamp 1649977179
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_137
timestamp 1649977179
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_149
timestamp 1649977179
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_161
timestamp 1649977179
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1649977179
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_169
timestamp 1649977179
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_181
timestamp 1649977179
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_193
timestamp 1649977179
transform 1 0 18860 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_205
timestamp 1649977179
transform 1 0 19964 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_217
timestamp 1649977179
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1649977179
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_225
timestamp 1649977179
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_237
timestamp 1649977179
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_249
timestamp 1649977179
transform 1 0 24012 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_261
timestamp 1649977179
transform 1 0 25116 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_273
timestamp 1649977179
transform 1 0 26220 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1649977179
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_281
timestamp 1649977179
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_293
timestamp 1649977179
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_305
timestamp 1649977179
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_317
timestamp 1649977179
transform 1 0 30268 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_329
timestamp 1649977179
transform 1 0 31372 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1649977179
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_337
timestamp 1649977179
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_349
timestamp 1649977179
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_361
timestamp 1649977179
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_373
timestamp 1649977179
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_385
timestamp 1649977179
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 1649977179
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_393
timestamp 1649977179
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_405
timestamp 1649977179
transform 1 0 38364 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_417
timestamp 1649977179
transform 1 0 39468 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_429
timestamp 1649977179
transform 1 0 40572 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_441
timestamp 1649977179
transform 1 0 41676 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_447
timestamp 1649977179
transform 1 0 42228 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_449
timestamp 1649977179
transform 1 0 42412 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_461
timestamp 1649977179
transform 1 0 43516 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_473
timestamp 1649977179
transform 1 0 44620 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_485
timestamp 1649977179
transform 1 0 45724 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_497
timestamp 1649977179
transform 1 0 46828 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_503
timestamp 1649977179
transform 1 0 47380 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_505
timestamp 1649977179
transform 1 0 47564 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_517
timestamp 1649977179
transform 1 0 48668 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_529
timestamp 1649977179
transform 1 0 49772 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_541
timestamp 1649977179
transform 1 0 50876 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_553
timestamp 1649977179
transform 1 0 51980 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_559
timestamp 1649977179
transform 1 0 52532 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_561
timestamp 1649977179
transform 1 0 52716 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_573
timestamp 1649977179
transform 1 0 53820 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_585
timestamp 1649977179
transform 1 0 54924 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_597
timestamp 1649977179
transform 1 0 56028 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_609
timestamp 1649977179
transform 1 0 57132 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_615
timestamp 1649977179
transform 1 0 57684 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_617
timestamp 1649977179
transform 1 0 57868 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_629
timestamp 1649977179
transform 1 0 58972 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_641
timestamp 1649977179
transform 1 0 60076 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_653
timestamp 1649977179
transform 1 0 61180 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_665
timestamp 1649977179
transform 1 0 62284 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_671
timestamp 1649977179
transform 1 0 62836 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_673
timestamp 1649977179
transform 1 0 63020 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_685
timestamp 1649977179
transform 1 0 64124 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_697
timestamp 1649977179
transform 1 0 65228 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_709
timestamp 1649977179
transform 1 0 66332 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_721
timestamp 1649977179
transform 1 0 67436 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_727
timestamp 1649977179
transform 1 0 67988 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_729
timestamp 1649977179
transform 1 0 68172 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_3
timestamp 1649977179
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_15
timestamp 1649977179
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1649977179
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1649977179
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_41
timestamp 1649977179
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_53
timestamp 1649977179
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_65
timestamp 1649977179
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1649977179
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1649977179
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_85
timestamp 1649977179
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_97
timestamp 1649977179
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_109
timestamp 1649977179
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_121
timestamp 1649977179
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1649977179
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1649977179
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_141
timestamp 1649977179
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_153
timestamp 1649977179
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_165
timestamp 1649977179
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_177
timestamp 1649977179
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_189
timestamp 1649977179
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1649977179
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_197
timestamp 1649977179
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_209
timestamp 1649977179
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_221
timestamp 1649977179
transform 1 0 21436 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_233
timestamp 1649977179
transform 1 0 22540 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_245
timestamp 1649977179
transform 1 0 23644 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1649977179
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_253
timestamp 1649977179
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_265
timestamp 1649977179
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_277
timestamp 1649977179
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_289
timestamp 1649977179
transform 1 0 27692 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_301
timestamp 1649977179
transform 1 0 28796 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 1649977179
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_309
timestamp 1649977179
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_321
timestamp 1649977179
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_333
timestamp 1649977179
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_345
timestamp 1649977179
transform 1 0 32844 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_357
timestamp 1649977179
transform 1 0 33948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1649977179
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_365
timestamp 1649977179
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_377
timestamp 1649977179
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_389
timestamp 1649977179
transform 1 0 36892 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_401
timestamp 1649977179
transform 1 0 37996 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_413
timestamp 1649977179
transform 1 0 39100 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_419
timestamp 1649977179
transform 1 0 39652 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_421
timestamp 1649977179
transform 1 0 39836 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_433
timestamp 1649977179
transform 1 0 40940 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_445
timestamp 1649977179
transform 1 0 42044 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_457
timestamp 1649977179
transform 1 0 43148 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_469
timestamp 1649977179
transform 1 0 44252 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_475
timestamp 1649977179
transform 1 0 44804 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_477
timestamp 1649977179
transform 1 0 44988 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_489
timestamp 1649977179
transform 1 0 46092 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_501
timestamp 1649977179
transform 1 0 47196 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_513
timestamp 1649977179
transform 1 0 48300 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_525
timestamp 1649977179
transform 1 0 49404 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_531
timestamp 1649977179
transform 1 0 49956 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_533
timestamp 1649977179
transform 1 0 50140 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_545
timestamp 1649977179
transform 1 0 51244 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_557
timestamp 1649977179
transform 1 0 52348 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_569
timestamp 1649977179
transform 1 0 53452 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_581
timestamp 1649977179
transform 1 0 54556 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_587
timestamp 1649977179
transform 1 0 55108 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_589
timestamp 1649977179
transform 1 0 55292 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_601
timestamp 1649977179
transform 1 0 56396 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_613
timestamp 1649977179
transform 1 0 57500 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_625
timestamp 1649977179
transform 1 0 58604 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_637
timestamp 1649977179
transform 1 0 59708 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_643
timestamp 1649977179
transform 1 0 60260 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_645
timestamp 1649977179
transform 1 0 60444 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_657
timestamp 1649977179
transform 1 0 61548 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_669
timestamp 1649977179
transform 1 0 62652 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_681
timestamp 1649977179
transform 1 0 63756 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_693
timestamp 1649977179
transform 1 0 64860 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_699
timestamp 1649977179
transform 1 0 65412 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_701
timestamp 1649977179
transform 1 0 65596 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_713
timestamp 1649977179
transform 1 0 66700 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_725
timestamp 1649977179
transform 1 0 67804 0 1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1649977179
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1649977179
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_27
timestamp 1649977179
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_39
timestamp 1649977179
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1649977179
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1649977179
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1649977179
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_69
timestamp 1649977179
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_81
timestamp 1649977179
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_93
timestamp 1649977179
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1649977179
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1649977179
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_113
timestamp 1649977179
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_125
timestamp 1649977179
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_137
timestamp 1649977179
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_149
timestamp 1649977179
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_161
timestamp 1649977179
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1649977179
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_169
timestamp 1649977179
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_181
timestamp 1649977179
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_193
timestamp 1649977179
transform 1 0 18860 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_205
timestamp 1649977179
transform 1 0 19964 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_217
timestamp 1649977179
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1649977179
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_225
timestamp 1649977179
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_237
timestamp 1649977179
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_249
timestamp 1649977179
transform 1 0 24012 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_261
timestamp 1649977179
transform 1 0 25116 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_273
timestamp 1649977179
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1649977179
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_281
timestamp 1649977179
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_293
timestamp 1649977179
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_305
timestamp 1649977179
transform 1 0 29164 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_317
timestamp 1649977179
transform 1 0 30268 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_329
timestamp 1649977179
transform 1 0 31372 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_335
timestamp 1649977179
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_337
timestamp 1649977179
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_349
timestamp 1649977179
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_361
timestamp 1649977179
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_373
timestamp 1649977179
transform 1 0 35420 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_385
timestamp 1649977179
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1649977179
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_393
timestamp 1649977179
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_405
timestamp 1649977179
transform 1 0 38364 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_417
timestamp 1649977179
transform 1 0 39468 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_429
timestamp 1649977179
transform 1 0 40572 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_441
timestamp 1649977179
transform 1 0 41676 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_447
timestamp 1649977179
transform 1 0 42228 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_449
timestamp 1649977179
transform 1 0 42412 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_461
timestamp 1649977179
transform 1 0 43516 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_473
timestamp 1649977179
transform 1 0 44620 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_485
timestamp 1649977179
transform 1 0 45724 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_497
timestamp 1649977179
transform 1 0 46828 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_503
timestamp 1649977179
transform 1 0 47380 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_505
timestamp 1649977179
transform 1 0 47564 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_517
timestamp 1649977179
transform 1 0 48668 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_529
timestamp 1649977179
transform 1 0 49772 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_541
timestamp 1649977179
transform 1 0 50876 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_553
timestamp 1649977179
transform 1 0 51980 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_559
timestamp 1649977179
transform 1 0 52532 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_561
timestamp 1649977179
transform 1 0 52716 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_573
timestamp 1649977179
transform 1 0 53820 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_585
timestamp 1649977179
transform 1 0 54924 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_597
timestamp 1649977179
transform 1 0 56028 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_609
timestamp 1649977179
transform 1 0 57132 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_615
timestamp 1649977179
transform 1 0 57684 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_617
timestamp 1649977179
transform 1 0 57868 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_629
timestamp 1649977179
transform 1 0 58972 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_641
timestamp 1649977179
transform 1 0 60076 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_653
timestamp 1649977179
transform 1 0 61180 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_665
timestamp 1649977179
transform 1 0 62284 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_671
timestamp 1649977179
transform 1 0 62836 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_673
timestamp 1649977179
transform 1 0 63020 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_685
timestamp 1649977179
transform 1 0 64124 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_697
timestamp 1649977179
transform 1 0 65228 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_709
timestamp 1649977179
transform 1 0 66332 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_721
timestamp 1649977179
transform 1 0 67436 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_727
timestamp 1649977179
transform 1 0 67988 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_729
timestamp 1649977179
transform 1 0 68172 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_3
timestamp 1649977179
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_15
timestamp 1649977179
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1649977179
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1649977179
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1649977179
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_53
timestamp 1649977179
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_65
timestamp 1649977179
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1649977179
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1649977179
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_85
timestamp 1649977179
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_97
timestamp 1649977179
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_109
timestamp 1649977179
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_121
timestamp 1649977179
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1649977179
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1649977179
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_141
timestamp 1649977179
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_153
timestamp 1649977179
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_165
timestamp 1649977179
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_177
timestamp 1649977179
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_189
timestamp 1649977179
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1649977179
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_197
timestamp 1649977179
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_209
timestamp 1649977179
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_221
timestamp 1649977179
transform 1 0 21436 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_233
timestamp 1649977179
transform 1 0 22540 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_245
timestamp 1649977179
transform 1 0 23644 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1649977179
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_253
timestamp 1649977179
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_265
timestamp 1649977179
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_277
timestamp 1649977179
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_289
timestamp 1649977179
transform 1 0 27692 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_301
timestamp 1649977179
transform 1 0 28796 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1649977179
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_309
timestamp 1649977179
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_321
timestamp 1649977179
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_333
timestamp 1649977179
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_345
timestamp 1649977179
transform 1 0 32844 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_357
timestamp 1649977179
transform 1 0 33948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_363
timestamp 1649977179
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_365
timestamp 1649977179
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_377
timestamp 1649977179
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_389
timestamp 1649977179
transform 1 0 36892 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_401
timestamp 1649977179
transform 1 0 37996 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_413
timestamp 1649977179
transform 1 0 39100 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_419
timestamp 1649977179
transform 1 0 39652 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_421
timestamp 1649977179
transform 1 0 39836 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_433
timestamp 1649977179
transform 1 0 40940 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_445
timestamp 1649977179
transform 1 0 42044 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_457
timestamp 1649977179
transform 1 0 43148 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_469
timestamp 1649977179
transform 1 0 44252 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_475
timestamp 1649977179
transform 1 0 44804 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_477
timestamp 1649977179
transform 1 0 44988 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_489
timestamp 1649977179
transform 1 0 46092 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_501
timestamp 1649977179
transform 1 0 47196 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_513
timestamp 1649977179
transform 1 0 48300 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_525
timestamp 1649977179
transform 1 0 49404 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_531
timestamp 1649977179
transform 1 0 49956 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_533
timestamp 1649977179
transform 1 0 50140 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_545
timestamp 1649977179
transform 1 0 51244 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_557
timestamp 1649977179
transform 1 0 52348 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_569
timestamp 1649977179
transform 1 0 53452 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_581
timestamp 1649977179
transform 1 0 54556 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_587
timestamp 1649977179
transform 1 0 55108 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_589
timestamp 1649977179
transform 1 0 55292 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_601
timestamp 1649977179
transform 1 0 56396 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_613
timestamp 1649977179
transform 1 0 57500 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_625
timestamp 1649977179
transform 1 0 58604 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_637
timestamp 1649977179
transform 1 0 59708 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_643
timestamp 1649977179
transform 1 0 60260 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_645
timestamp 1649977179
transform 1 0 60444 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_657
timestamp 1649977179
transform 1 0 61548 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_669
timestamp 1649977179
transform 1 0 62652 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_681
timestamp 1649977179
transform 1 0 63756 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_693
timestamp 1649977179
transform 1 0 64860 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_699
timestamp 1649977179
transform 1 0 65412 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_701
timestamp 1649977179
transform 1 0 65596 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_713
timestamp 1649977179
transform 1 0 66700 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_725
timestamp 1649977179
transform 1 0 67804 0 1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1649977179
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 1649977179
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_27
timestamp 1649977179
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_39
timestamp 1649977179
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1649977179
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1649977179
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1649977179
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_69
timestamp 1649977179
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_81
timestamp 1649977179
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_93
timestamp 1649977179
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1649977179
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1649977179
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_113
timestamp 1649977179
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_125
timestamp 1649977179
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_137
timestamp 1649977179
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_149
timestamp 1649977179
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 1649977179
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1649977179
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_169
timestamp 1649977179
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_181
timestamp 1649977179
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_193
timestamp 1649977179
transform 1 0 18860 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_205
timestamp 1649977179
transform 1 0 19964 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_217
timestamp 1649977179
transform 1 0 21068 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1649977179
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_225
timestamp 1649977179
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_237
timestamp 1649977179
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_249
timestamp 1649977179
transform 1 0 24012 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_261
timestamp 1649977179
transform 1 0 25116 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_273
timestamp 1649977179
transform 1 0 26220 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1649977179
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_281
timestamp 1649977179
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_293
timestamp 1649977179
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_305
timestamp 1649977179
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_317
timestamp 1649977179
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_329
timestamp 1649977179
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1649977179
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_337
timestamp 1649977179
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_349
timestamp 1649977179
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_361
timestamp 1649977179
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_373
timestamp 1649977179
transform 1 0 35420 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_385
timestamp 1649977179
transform 1 0 36524 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 1649977179
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_393
timestamp 1649977179
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_405
timestamp 1649977179
transform 1 0 38364 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_417
timestamp 1649977179
transform 1 0 39468 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_429
timestamp 1649977179
transform 1 0 40572 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_441
timestamp 1649977179
transform 1 0 41676 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_447
timestamp 1649977179
transform 1 0 42228 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_449
timestamp 1649977179
transform 1 0 42412 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_461
timestamp 1649977179
transform 1 0 43516 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_473
timestamp 1649977179
transform 1 0 44620 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_485
timestamp 1649977179
transform 1 0 45724 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_497
timestamp 1649977179
transform 1 0 46828 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_503
timestamp 1649977179
transform 1 0 47380 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_505
timestamp 1649977179
transform 1 0 47564 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_517
timestamp 1649977179
transform 1 0 48668 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_529
timestamp 1649977179
transform 1 0 49772 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_541
timestamp 1649977179
transform 1 0 50876 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_553
timestamp 1649977179
transform 1 0 51980 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_559
timestamp 1649977179
transform 1 0 52532 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_561
timestamp 1649977179
transform 1 0 52716 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_573
timestamp 1649977179
transform 1 0 53820 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_585
timestamp 1649977179
transform 1 0 54924 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_597
timestamp 1649977179
transform 1 0 56028 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_609
timestamp 1649977179
transform 1 0 57132 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_615
timestamp 1649977179
transform 1 0 57684 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_617
timestamp 1649977179
transform 1 0 57868 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_629
timestamp 1649977179
transform 1 0 58972 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_641
timestamp 1649977179
transform 1 0 60076 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_653
timestamp 1649977179
transform 1 0 61180 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_665
timestamp 1649977179
transform 1 0 62284 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_671
timestamp 1649977179
transform 1 0 62836 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_673
timestamp 1649977179
transform 1 0 63020 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_685
timestamp 1649977179
transform 1 0 64124 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_697
timestamp 1649977179
transform 1 0 65228 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_709
timestamp 1649977179
transform 1 0 66332 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_721
timestamp 1649977179
transform 1 0 67436 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_727
timestamp 1649977179
transform 1 0 67988 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_729
timestamp 1649977179
transform 1 0 68172 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1649977179
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1649977179
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1649977179
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1649977179
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1649977179
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_53
timestamp 1649977179
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_65
timestamp 1649977179
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1649977179
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1649977179
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_85
timestamp 1649977179
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_97
timestamp 1649977179
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_109
timestamp 1649977179
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_121
timestamp 1649977179
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1649977179
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1649977179
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_141
timestamp 1649977179
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_153
timestamp 1649977179
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_165
timestamp 1649977179
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_177
timestamp 1649977179
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_189
timestamp 1649977179
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1649977179
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_197
timestamp 1649977179
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_209
timestamp 1649977179
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_221
timestamp 1649977179
transform 1 0 21436 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_233
timestamp 1649977179
transform 1 0 22540 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_245
timestamp 1649977179
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1649977179
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_253
timestamp 1649977179
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_265
timestamp 1649977179
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_277
timestamp 1649977179
transform 1 0 26588 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_289
timestamp 1649977179
transform 1 0 27692 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_301
timestamp 1649977179
transform 1 0 28796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1649977179
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_309
timestamp 1649977179
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_321
timestamp 1649977179
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_333
timestamp 1649977179
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_345
timestamp 1649977179
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_357
timestamp 1649977179
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1649977179
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_365
timestamp 1649977179
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_377
timestamp 1649977179
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_389
timestamp 1649977179
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_401
timestamp 1649977179
transform 1 0 37996 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_413
timestamp 1649977179
transform 1 0 39100 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_419
timestamp 1649977179
transform 1 0 39652 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_421
timestamp 1649977179
transform 1 0 39836 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_433
timestamp 1649977179
transform 1 0 40940 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_445
timestamp 1649977179
transform 1 0 42044 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_457
timestamp 1649977179
transform 1 0 43148 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_469
timestamp 1649977179
transform 1 0 44252 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_475
timestamp 1649977179
transform 1 0 44804 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_477
timestamp 1649977179
transform 1 0 44988 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_489
timestamp 1649977179
transform 1 0 46092 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_501
timestamp 1649977179
transform 1 0 47196 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_513
timestamp 1649977179
transform 1 0 48300 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_525
timestamp 1649977179
transform 1 0 49404 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_531
timestamp 1649977179
transform 1 0 49956 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_533
timestamp 1649977179
transform 1 0 50140 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_545
timestamp 1649977179
transform 1 0 51244 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_557
timestamp 1649977179
transform 1 0 52348 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_569
timestamp 1649977179
transform 1 0 53452 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_581
timestamp 1649977179
transform 1 0 54556 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_587
timestamp 1649977179
transform 1 0 55108 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_589
timestamp 1649977179
transform 1 0 55292 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_601
timestamp 1649977179
transform 1 0 56396 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_613
timestamp 1649977179
transform 1 0 57500 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_625
timestamp 1649977179
transform 1 0 58604 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_637
timestamp 1649977179
transform 1 0 59708 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_643
timestamp 1649977179
transform 1 0 60260 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_645
timestamp 1649977179
transform 1 0 60444 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_657
timestamp 1649977179
transform 1 0 61548 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_669
timestamp 1649977179
transform 1 0 62652 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_681
timestamp 1649977179
transform 1 0 63756 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_693
timestamp 1649977179
transform 1 0 64860 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_699
timestamp 1649977179
transform 1 0 65412 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_701
timestamp 1649977179
transform 1 0 65596 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_713
timestamp 1649977179
transform 1 0 66700 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_725
timestamp 1649977179
transform 1 0 67804 0 1 31552
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_55_3
timestamp 1649977179
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_15
timestamp 1649977179
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_27
timestamp 1649977179
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_39
timestamp 1649977179
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 1649977179
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1649977179
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 1649977179
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_69
timestamp 1649977179
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_81
timestamp 1649977179
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_93
timestamp 1649977179
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1649977179
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1649977179
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_113
timestamp 1649977179
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_125
timestamp 1649977179
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_137
timestamp 1649977179
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_149
timestamp 1649977179
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1649977179
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1649977179
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_169
timestamp 1649977179
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_181
timestamp 1649977179
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_193
timestamp 1649977179
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_205
timestamp 1649977179
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_217
timestamp 1649977179
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1649977179
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_225
timestamp 1649977179
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_237
timestamp 1649977179
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_249
timestamp 1649977179
transform 1 0 24012 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_261
timestamp 1649977179
transform 1 0 25116 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_273
timestamp 1649977179
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1649977179
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_281
timestamp 1649977179
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_293
timestamp 1649977179
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_305
timestamp 1649977179
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_317
timestamp 1649977179
transform 1 0 30268 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_329
timestamp 1649977179
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 1649977179
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_337
timestamp 1649977179
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_349
timestamp 1649977179
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_361
timestamp 1649977179
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_373
timestamp 1649977179
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_385
timestamp 1649977179
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1649977179
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_393
timestamp 1649977179
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_405
timestamp 1649977179
transform 1 0 38364 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_417
timestamp 1649977179
transform 1 0 39468 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_429
timestamp 1649977179
transform 1 0 40572 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_441
timestamp 1649977179
transform 1 0 41676 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_447
timestamp 1649977179
transform 1 0 42228 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_449
timestamp 1649977179
transform 1 0 42412 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_461
timestamp 1649977179
transform 1 0 43516 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_473
timestamp 1649977179
transform 1 0 44620 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_485
timestamp 1649977179
transform 1 0 45724 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_497
timestamp 1649977179
transform 1 0 46828 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_503
timestamp 1649977179
transform 1 0 47380 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_505
timestamp 1649977179
transform 1 0 47564 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_517
timestamp 1649977179
transform 1 0 48668 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_529
timestamp 1649977179
transform 1 0 49772 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_541
timestamp 1649977179
transform 1 0 50876 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_553
timestamp 1649977179
transform 1 0 51980 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_559
timestamp 1649977179
transform 1 0 52532 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_561
timestamp 1649977179
transform 1 0 52716 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_573
timestamp 1649977179
transform 1 0 53820 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_585
timestamp 1649977179
transform 1 0 54924 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_597
timestamp 1649977179
transform 1 0 56028 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_609
timestamp 1649977179
transform 1 0 57132 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_615
timestamp 1649977179
transform 1 0 57684 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_617
timestamp 1649977179
transform 1 0 57868 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_629
timestamp 1649977179
transform 1 0 58972 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_641
timestamp 1649977179
transform 1 0 60076 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_653
timestamp 1649977179
transform 1 0 61180 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_665
timestamp 1649977179
transform 1 0 62284 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_671
timestamp 1649977179
transform 1 0 62836 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_673
timestamp 1649977179
transform 1 0 63020 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_685
timestamp 1649977179
transform 1 0 64124 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_697
timestamp 1649977179
transform 1 0 65228 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_709
timestamp 1649977179
transform 1 0 66332 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_721
timestamp 1649977179
transform 1 0 67436 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_727
timestamp 1649977179
transform 1 0 67988 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_729
timestamp 1649977179
transform 1 0 68172 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1649977179
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1649977179
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1649977179
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1649977179
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1649977179
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_53
timestamp 1649977179
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_65
timestamp 1649977179
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1649977179
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1649977179
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_85
timestamp 1649977179
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_97
timestamp 1649977179
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_109
timestamp 1649977179
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_121
timestamp 1649977179
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1649977179
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1649977179
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_141
timestamp 1649977179
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_153
timestamp 1649977179
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_165
timestamp 1649977179
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_177
timestamp 1649977179
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_189
timestamp 1649977179
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1649977179
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_197
timestamp 1649977179
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_209
timestamp 1649977179
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_221
timestamp 1649977179
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_233
timestamp 1649977179
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_245
timestamp 1649977179
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1649977179
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_253
timestamp 1649977179
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_265
timestamp 1649977179
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_277
timestamp 1649977179
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_289
timestamp 1649977179
transform 1 0 27692 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_301
timestamp 1649977179
transform 1 0 28796 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_307
timestamp 1649977179
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_309
timestamp 1649977179
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_321
timestamp 1649977179
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_333
timestamp 1649977179
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_345
timestamp 1649977179
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_357
timestamp 1649977179
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1649977179
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_365
timestamp 1649977179
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_377
timestamp 1649977179
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_389
timestamp 1649977179
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_401
timestamp 1649977179
transform 1 0 37996 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_413
timestamp 1649977179
transform 1 0 39100 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_419
timestamp 1649977179
transform 1 0 39652 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_421
timestamp 1649977179
transform 1 0 39836 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_433
timestamp 1649977179
transform 1 0 40940 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_445
timestamp 1649977179
transform 1 0 42044 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_457
timestamp 1649977179
transform 1 0 43148 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_469
timestamp 1649977179
transform 1 0 44252 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_475
timestamp 1649977179
transform 1 0 44804 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_477
timestamp 1649977179
transform 1 0 44988 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_489
timestamp 1649977179
transform 1 0 46092 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_501
timestamp 1649977179
transform 1 0 47196 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_513
timestamp 1649977179
transform 1 0 48300 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_525
timestamp 1649977179
transform 1 0 49404 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_531
timestamp 1649977179
transform 1 0 49956 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_533
timestamp 1649977179
transform 1 0 50140 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_545
timestamp 1649977179
transform 1 0 51244 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_557
timestamp 1649977179
transform 1 0 52348 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_569
timestamp 1649977179
transform 1 0 53452 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_581
timestamp 1649977179
transform 1 0 54556 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_587
timestamp 1649977179
transform 1 0 55108 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_589
timestamp 1649977179
transform 1 0 55292 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_601
timestamp 1649977179
transform 1 0 56396 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_613
timestamp 1649977179
transform 1 0 57500 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_625
timestamp 1649977179
transform 1 0 58604 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_637
timestamp 1649977179
transform 1 0 59708 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_643
timestamp 1649977179
transform 1 0 60260 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_645
timestamp 1649977179
transform 1 0 60444 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_657
timestamp 1649977179
transform 1 0 61548 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_669
timestamp 1649977179
transform 1 0 62652 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_681
timestamp 1649977179
transform 1 0 63756 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_693
timestamp 1649977179
transform 1 0 64860 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_699
timestamp 1649977179
transform 1 0 65412 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_701
timestamp 1649977179
transform 1 0 65596 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_713
timestamp 1649977179
transform 1 0 66700 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_725
timestamp 1649977179
transform 1 0 67804 0 1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1649977179
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_15
timestamp 1649977179
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_27
timestamp 1649977179
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_39
timestamp 1649977179
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1649977179
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1649977179
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1649977179
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_69
timestamp 1649977179
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_81
timestamp 1649977179
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_93
timestamp 1649977179
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1649977179
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1649977179
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_113
timestamp 1649977179
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_125
timestamp 1649977179
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_137
timestamp 1649977179
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_149
timestamp 1649977179
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1649977179
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1649977179
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_169
timestamp 1649977179
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_181
timestamp 1649977179
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_193
timestamp 1649977179
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_205
timestamp 1649977179
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_217
timestamp 1649977179
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1649977179
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_225
timestamp 1649977179
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_237
timestamp 1649977179
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_249
timestamp 1649977179
transform 1 0 24012 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_261
timestamp 1649977179
transform 1 0 25116 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_273
timestamp 1649977179
transform 1 0 26220 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1649977179
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_281
timestamp 1649977179
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_293
timestamp 1649977179
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_305
timestamp 1649977179
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_317
timestamp 1649977179
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_329
timestamp 1649977179
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1649977179
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_337
timestamp 1649977179
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_349
timestamp 1649977179
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_361
timestamp 1649977179
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_373
timestamp 1649977179
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_385
timestamp 1649977179
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1649977179
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_393
timestamp 1649977179
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_405
timestamp 1649977179
transform 1 0 38364 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_417
timestamp 1649977179
transform 1 0 39468 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_429
timestamp 1649977179
transform 1 0 40572 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_441
timestamp 1649977179
transform 1 0 41676 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_447
timestamp 1649977179
transform 1 0 42228 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_449
timestamp 1649977179
transform 1 0 42412 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_461
timestamp 1649977179
transform 1 0 43516 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_473
timestamp 1649977179
transform 1 0 44620 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_485
timestamp 1649977179
transform 1 0 45724 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_497
timestamp 1649977179
transform 1 0 46828 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_503
timestamp 1649977179
transform 1 0 47380 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_505
timestamp 1649977179
transform 1 0 47564 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_517
timestamp 1649977179
transform 1 0 48668 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_529
timestamp 1649977179
transform 1 0 49772 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_541
timestamp 1649977179
transform 1 0 50876 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_553
timestamp 1649977179
transform 1 0 51980 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_559
timestamp 1649977179
transform 1 0 52532 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_561
timestamp 1649977179
transform 1 0 52716 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_573
timestamp 1649977179
transform 1 0 53820 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_585
timestamp 1649977179
transform 1 0 54924 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_597
timestamp 1649977179
transform 1 0 56028 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_609
timestamp 1649977179
transform 1 0 57132 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_615
timestamp 1649977179
transform 1 0 57684 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_617
timestamp 1649977179
transform 1 0 57868 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_629
timestamp 1649977179
transform 1 0 58972 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_641
timestamp 1649977179
transform 1 0 60076 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_653
timestamp 1649977179
transform 1 0 61180 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_665
timestamp 1649977179
transform 1 0 62284 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_671
timestamp 1649977179
transform 1 0 62836 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_673
timestamp 1649977179
transform 1 0 63020 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_685
timestamp 1649977179
transform 1 0 64124 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_697
timestamp 1649977179
transform 1 0 65228 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_709
timestamp 1649977179
transform 1 0 66332 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_721
timestamp 1649977179
transform 1 0 67436 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_727
timestamp 1649977179
transform 1 0 67988 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_729
timestamp 1649977179
transform 1 0 68172 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1649977179
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1649977179
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1649977179
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1649977179
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1649977179
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_53
timestamp 1649977179
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_65
timestamp 1649977179
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1649977179
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1649977179
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_85
timestamp 1649977179
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_97
timestamp 1649977179
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_109
timestamp 1649977179
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_121
timestamp 1649977179
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1649977179
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1649977179
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_141
timestamp 1649977179
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_153
timestamp 1649977179
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_165
timestamp 1649977179
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_177
timestamp 1649977179
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1649977179
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1649977179
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_197
timestamp 1649977179
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_209
timestamp 1649977179
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_221
timestamp 1649977179
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_233
timestamp 1649977179
transform 1 0 22540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_245
timestamp 1649977179
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1649977179
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_253
timestamp 1649977179
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_265
timestamp 1649977179
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_277
timestamp 1649977179
transform 1 0 26588 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_289
timestamp 1649977179
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_301
timestamp 1649977179
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1649977179
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_309
timestamp 1649977179
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_321
timestamp 1649977179
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_333
timestamp 1649977179
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_345
timestamp 1649977179
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_357
timestamp 1649977179
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1649977179
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_365
timestamp 1649977179
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_377
timestamp 1649977179
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_389
timestamp 1649977179
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_401
timestamp 1649977179
transform 1 0 37996 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_413
timestamp 1649977179
transform 1 0 39100 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_419
timestamp 1649977179
transform 1 0 39652 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_421
timestamp 1649977179
transform 1 0 39836 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_433
timestamp 1649977179
transform 1 0 40940 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_445
timestamp 1649977179
transform 1 0 42044 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_457
timestamp 1649977179
transform 1 0 43148 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_469
timestamp 1649977179
transform 1 0 44252 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_475
timestamp 1649977179
transform 1 0 44804 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_477
timestamp 1649977179
transform 1 0 44988 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_489
timestamp 1649977179
transform 1 0 46092 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_501
timestamp 1649977179
transform 1 0 47196 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_513
timestamp 1649977179
transform 1 0 48300 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_525
timestamp 1649977179
transform 1 0 49404 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_531
timestamp 1649977179
transform 1 0 49956 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_533
timestamp 1649977179
transform 1 0 50140 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_545
timestamp 1649977179
transform 1 0 51244 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_557
timestamp 1649977179
transform 1 0 52348 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_569
timestamp 1649977179
transform 1 0 53452 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_581
timestamp 1649977179
transform 1 0 54556 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_587
timestamp 1649977179
transform 1 0 55108 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_589
timestamp 1649977179
transform 1 0 55292 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_601
timestamp 1649977179
transform 1 0 56396 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_613
timestamp 1649977179
transform 1 0 57500 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_625
timestamp 1649977179
transform 1 0 58604 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_637
timestamp 1649977179
transform 1 0 59708 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_643
timestamp 1649977179
transform 1 0 60260 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_645
timestamp 1649977179
transform 1 0 60444 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_657
timestamp 1649977179
transform 1 0 61548 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_669
timestamp 1649977179
transform 1 0 62652 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_681
timestamp 1649977179
transform 1 0 63756 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_693
timestamp 1649977179
transform 1 0 64860 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_699
timestamp 1649977179
transform 1 0 65412 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_701
timestamp 1649977179
transform 1 0 65596 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_713
timestamp 1649977179
transform 1 0 66700 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_725
timestamp 1649977179
transform 1 0 67804 0 1 33728
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_59_3
timestamp 1649977179
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_15
timestamp 1649977179
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_27
timestamp 1649977179
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_39
timestamp 1649977179
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1649977179
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1649977179
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1649977179
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_69
timestamp 1649977179
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_81
timestamp 1649977179
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_93
timestamp 1649977179
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1649977179
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1649977179
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_113
timestamp 1649977179
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_125
timestamp 1649977179
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_137
timestamp 1649977179
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_149
timestamp 1649977179
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1649977179
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1649977179
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_169
timestamp 1649977179
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_181
timestamp 1649977179
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_193
timestamp 1649977179
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_205
timestamp 1649977179
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 1649977179
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1649977179
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_225
timestamp 1649977179
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_237
timestamp 1649977179
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_249
timestamp 1649977179
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_261
timestamp 1649977179
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_273
timestamp 1649977179
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1649977179
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_281
timestamp 1649977179
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_293
timestamp 1649977179
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_305
timestamp 1649977179
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_317
timestamp 1649977179
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_329
timestamp 1649977179
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1649977179
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_337
timestamp 1649977179
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_349
timestamp 1649977179
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_361
timestamp 1649977179
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_373
timestamp 1649977179
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_385
timestamp 1649977179
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 1649977179
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_393
timestamp 1649977179
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_405
timestamp 1649977179
transform 1 0 38364 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_417
timestamp 1649977179
transform 1 0 39468 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_429
timestamp 1649977179
transform 1 0 40572 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_441
timestamp 1649977179
transform 1 0 41676 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_447
timestamp 1649977179
transform 1 0 42228 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_449
timestamp 1649977179
transform 1 0 42412 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_461
timestamp 1649977179
transform 1 0 43516 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_473
timestamp 1649977179
transform 1 0 44620 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_485
timestamp 1649977179
transform 1 0 45724 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_497
timestamp 1649977179
transform 1 0 46828 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_503
timestamp 1649977179
transform 1 0 47380 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_505
timestamp 1649977179
transform 1 0 47564 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_517
timestamp 1649977179
transform 1 0 48668 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_529
timestamp 1649977179
transform 1 0 49772 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_541
timestamp 1649977179
transform 1 0 50876 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_553
timestamp 1649977179
transform 1 0 51980 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_559
timestamp 1649977179
transform 1 0 52532 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_561
timestamp 1649977179
transform 1 0 52716 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_573
timestamp 1649977179
transform 1 0 53820 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_585
timestamp 1649977179
transform 1 0 54924 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_597
timestamp 1649977179
transform 1 0 56028 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_609
timestamp 1649977179
transform 1 0 57132 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_615
timestamp 1649977179
transform 1 0 57684 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_617
timestamp 1649977179
transform 1 0 57868 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_629
timestamp 1649977179
transform 1 0 58972 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_641
timestamp 1649977179
transform 1 0 60076 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_653
timestamp 1649977179
transform 1 0 61180 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_665
timestamp 1649977179
transform 1 0 62284 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_671
timestamp 1649977179
transform 1 0 62836 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_673
timestamp 1649977179
transform 1 0 63020 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_685
timestamp 1649977179
transform 1 0 64124 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_697
timestamp 1649977179
transform 1 0 65228 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_709
timestamp 1649977179
transform 1 0 66332 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_721
timestamp 1649977179
transform 1 0 67436 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_727
timestamp 1649977179
transform 1 0 67988 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_729
timestamp 1649977179
transform 1 0 68172 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 1649977179
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_15
timestamp 1649977179
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1649977179
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1649977179
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1649977179
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_53
timestamp 1649977179
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_65
timestamp 1649977179
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1649977179
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1649977179
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_85
timestamp 1649977179
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_97
timestamp 1649977179
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_109
timestamp 1649977179
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_121
timestamp 1649977179
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1649977179
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1649977179
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_141
timestamp 1649977179
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_153
timestamp 1649977179
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_165
timestamp 1649977179
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_177
timestamp 1649977179
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_189
timestamp 1649977179
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1649977179
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_197
timestamp 1649977179
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_209
timestamp 1649977179
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_221
timestamp 1649977179
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_233
timestamp 1649977179
transform 1 0 22540 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_245
timestamp 1649977179
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1649977179
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_253
timestamp 1649977179
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_265
timestamp 1649977179
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_277
timestamp 1649977179
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_289
timestamp 1649977179
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_301
timestamp 1649977179
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1649977179
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_309
timestamp 1649977179
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_321
timestamp 1649977179
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_333
timestamp 1649977179
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_345
timestamp 1649977179
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_357
timestamp 1649977179
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 1649977179
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_365
timestamp 1649977179
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_377
timestamp 1649977179
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_389
timestamp 1649977179
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_401
timestamp 1649977179
transform 1 0 37996 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_413
timestamp 1649977179
transform 1 0 39100 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_419
timestamp 1649977179
transform 1 0 39652 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_421
timestamp 1649977179
transform 1 0 39836 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_433
timestamp 1649977179
transform 1 0 40940 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_445
timestamp 1649977179
transform 1 0 42044 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_457
timestamp 1649977179
transform 1 0 43148 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_469
timestamp 1649977179
transform 1 0 44252 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_475
timestamp 1649977179
transform 1 0 44804 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_477
timestamp 1649977179
transform 1 0 44988 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_489
timestamp 1649977179
transform 1 0 46092 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_501
timestamp 1649977179
transform 1 0 47196 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_513
timestamp 1649977179
transform 1 0 48300 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_525
timestamp 1649977179
transform 1 0 49404 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_531
timestamp 1649977179
transform 1 0 49956 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_533
timestamp 1649977179
transform 1 0 50140 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_545
timestamp 1649977179
transform 1 0 51244 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_557
timestamp 1649977179
transform 1 0 52348 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_569
timestamp 1649977179
transform 1 0 53452 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_581
timestamp 1649977179
transform 1 0 54556 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_587
timestamp 1649977179
transform 1 0 55108 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_589
timestamp 1649977179
transform 1 0 55292 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_601
timestamp 1649977179
transform 1 0 56396 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_613
timestamp 1649977179
transform 1 0 57500 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_625
timestamp 1649977179
transform 1 0 58604 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_637
timestamp 1649977179
transform 1 0 59708 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_643
timestamp 1649977179
transform 1 0 60260 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_645
timestamp 1649977179
transform 1 0 60444 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_657
timestamp 1649977179
transform 1 0 61548 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_669
timestamp 1649977179
transform 1 0 62652 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_681
timestamp 1649977179
transform 1 0 63756 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_693
timestamp 1649977179
transform 1 0 64860 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_699
timestamp 1649977179
transform 1 0 65412 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_701
timestamp 1649977179
transform 1 0 65596 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_713
timestamp 1649977179
transform 1 0 66700 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_725
timestamp 1649977179
transform 1 0 67804 0 1 34816
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_61_3
timestamp 1649977179
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_15
timestamp 1649977179
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_27
timestamp 1649977179
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_39
timestamp 1649977179
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 1649977179
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1649977179
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1649977179
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_69
timestamp 1649977179
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_81
timestamp 1649977179
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_93
timestamp 1649977179
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1649977179
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1649977179
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_113
timestamp 1649977179
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_125
timestamp 1649977179
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_137
timestamp 1649977179
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_149
timestamp 1649977179
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1649977179
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1649977179
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_169
timestamp 1649977179
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_181
timestamp 1649977179
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_193
timestamp 1649977179
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_205
timestamp 1649977179
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_217
timestamp 1649977179
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1649977179
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_225
timestamp 1649977179
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_237
timestamp 1649977179
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_249
timestamp 1649977179
transform 1 0 24012 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_261
timestamp 1649977179
transform 1 0 25116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_273
timestamp 1649977179
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1649977179
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_281
timestamp 1649977179
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_293
timestamp 1649977179
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_305
timestamp 1649977179
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_317
timestamp 1649977179
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_329
timestamp 1649977179
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1649977179
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_337
timestamp 1649977179
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_349
timestamp 1649977179
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_361
timestamp 1649977179
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_373
timestamp 1649977179
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_385
timestamp 1649977179
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_391
timestamp 1649977179
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_393
timestamp 1649977179
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_405
timestamp 1649977179
transform 1 0 38364 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_417
timestamp 1649977179
transform 1 0 39468 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_429
timestamp 1649977179
transform 1 0 40572 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_441
timestamp 1649977179
transform 1 0 41676 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_447
timestamp 1649977179
transform 1 0 42228 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_449
timestamp 1649977179
transform 1 0 42412 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_461
timestamp 1649977179
transform 1 0 43516 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_473
timestamp 1649977179
transform 1 0 44620 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_485
timestamp 1649977179
transform 1 0 45724 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_497
timestamp 1649977179
transform 1 0 46828 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_503
timestamp 1649977179
transform 1 0 47380 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_505
timestamp 1649977179
transform 1 0 47564 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_517
timestamp 1649977179
transform 1 0 48668 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_529
timestamp 1649977179
transform 1 0 49772 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_541
timestamp 1649977179
transform 1 0 50876 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_553
timestamp 1649977179
transform 1 0 51980 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_559
timestamp 1649977179
transform 1 0 52532 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_561
timestamp 1649977179
transform 1 0 52716 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_573
timestamp 1649977179
transform 1 0 53820 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_585
timestamp 1649977179
transform 1 0 54924 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_597
timestamp 1649977179
transform 1 0 56028 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_609
timestamp 1649977179
transform 1 0 57132 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_615
timestamp 1649977179
transform 1 0 57684 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_617
timestamp 1649977179
transform 1 0 57868 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_629
timestamp 1649977179
transform 1 0 58972 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_641
timestamp 1649977179
transform 1 0 60076 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_653
timestamp 1649977179
transform 1 0 61180 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_665
timestamp 1649977179
transform 1 0 62284 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_671
timestamp 1649977179
transform 1 0 62836 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_673
timestamp 1649977179
transform 1 0 63020 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_685
timestamp 1649977179
transform 1 0 64124 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_697
timestamp 1649977179
transform 1 0 65228 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_709
timestamp 1649977179
transform 1 0 66332 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_721
timestamp 1649977179
transform 1 0 67436 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_727
timestamp 1649977179
transform 1 0 67988 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_729
timestamp 1649977179
transform 1 0 68172 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_3
timestamp 1649977179
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_15
timestamp 1649977179
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1649977179
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1649977179
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_41
timestamp 1649977179
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_53
timestamp 1649977179
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_65
timestamp 1649977179
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1649977179
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1649977179
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_85
timestamp 1649977179
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_97
timestamp 1649977179
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_109
timestamp 1649977179
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_121
timestamp 1649977179
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1649977179
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1649977179
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_141
timestamp 1649977179
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_153
timestamp 1649977179
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_165
timestamp 1649977179
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_177
timestamp 1649977179
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1649977179
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1649977179
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_197
timestamp 1649977179
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_209
timestamp 1649977179
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_221
timestamp 1649977179
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_233
timestamp 1649977179
transform 1 0 22540 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_245
timestamp 1649977179
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1649977179
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_253
timestamp 1649977179
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_265
timestamp 1649977179
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_277
timestamp 1649977179
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_289
timestamp 1649977179
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_301
timestamp 1649977179
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 1649977179
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_309
timestamp 1649977179
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_321
timestamp 1649977179
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_333
timestamp 1649977179
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_345
timestamp 1649977179
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 1649977179
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1649977179
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_365
timestamp 1649977179
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_377
timestamp 1649977179
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_389
timestamp 1649977179
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_401
timestamp 1649977179
transform 1 0 37996 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_413
timestamp 1649977179
transform 1 0 39100 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_419
timestamp 1649977179
transform 1 0 39652 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_421
timestamp 1649977179
transform 1 0 39836 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_433
timestamp 1649977179
transform 1 0 40940 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_445
timestamp 1649977179
transform 1 0 42044 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_457
timestamp 1649977179
transform 1 0 43148 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_469
timestamp 1649977179
transform 1 0 44252 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_475
timestamp 1649977179
transform 1 0 44804 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_477
timestamp 1649977179
transform 1 0 44988 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_489
timestamp 1649977179
transform 1 0 46092 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_501
timestamp 1649977179
transform 1 0 47196 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_513
timestamp 1649977179
transform 1 0 48300 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_525
timestamp 1649977179
transform 1 0 49404 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_531
timestamp 1649977179
transform 1 0 49956 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_533
timestamp 1649977179
transform 1 0 50140 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_545
timestamp 1649977179
transform 1 0 51244 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_557
timestamp 1649977179
transform 1 0 52348 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_569
timestamp 1649977179
transform 1 0 53452 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_581
timestamp 1649977179
transform 1 0 54556 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_587
timestamp 1649977179
transform 1 0 55108 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_589
timestamp 1649977179
transform 1 0 55292 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_601
timestamp 1649977179
transform 1 0 56396 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_613
timestamp 1649977179
transform 1 0 57500 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_625
timestamp 1649977179
transform 1 0 58604 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_637
timestamp 1649977179
transform 1 0 59708 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_643
timestamp 1649977179
transform 1 0 60260 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_645
timestamp 1649977179
transform 1 0 60444 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_657
timestamp 1649977179
transform 1 0 61548 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_669
timestamp 1649977179
transform 1 0 62652 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_681
timestamp 1649977179
transform 1 0 63756 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_693
timestamp 1649977179
transform 1 0 64860 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_699
timestamp 1649977179
transform 1 0 65412 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_701
timestamp 1649977179
transform 1 0 65596 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_713
timestamp 1649977179
transform 1 0 66700 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_725
timestamp 1649977179
transform 1 0 67804 0 1 35904
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_63_3
timestamp 1649977179
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_15
timestamp 1649977179
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_27
timestamp 1649977179
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_39
timestamp 1649977179
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_51
timestamp 1649977179
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1649977179
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_57
timestamp 1649977179
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_69
timestamp 1649977179
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_81
timestamp 1649977179
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_93
timestamp 1649977179
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1649977179
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1649977179
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_113
timestamp 1649977179
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_125
timestamp 1649977179
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_137
timestamp 1649977179
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_149
timestamp 1649977179
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1649977179
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1649977179
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_169
timestamp 1649977179
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_181
timestamp 1649977179
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_193
timestamp 1649977179
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_205
timestamp 1649977179
transform 1 0 19964 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_217
timestamp 1649977179
transform 1 0 21068 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1649977179
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_225
timestamp 1649977179
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_237
timestamp 1649977179
transform 1 0 22908 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_249
timestamp 1649977179
transform 1 0 24012 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_261
timestamp 1649977179
transform 1 0 25116 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_273
timestamp 1649977179
transform 1 0 26220 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_279
timestamp 1649977179
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_281
timestamp 1649977179
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_293
timestamp 1649977179
transform 1 0 28060 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_305
timestamp 1649977179
transform 1 0 29164 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_317
timestamp 1649977179
transform 1 0 30268 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_329
timestamp 1649977179
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_335
timestamp 1649977179
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_337
timestamp 1649977179
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_349
timestamp 1649977179
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_361
timestamp 1649977179
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_373
timestamp 1649977179
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_385
timestamp 1649977179
transform 1 0 36524 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_391
timestamp 1649977179
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_393
timestamp 1649977179
transform 1 0 37260 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_405
timestamp 1649977179
transform 1 0 38364 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_417
timestamp 1649977179
transform 1 0 39468 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_429
timestamp 1649977179
transform 1 0 40572 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_441
timestamp 1649977179
transform 1 0 41676 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_447
timestamp 1649977179
transform 1 0 42228 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_449
timestamp 1649977179
transform 1 0 42412 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_461
timestamp 1649977179
transform 1 0 43516 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_473
timestamp 1649977179
transform 1 0 44620 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_485
timestamp 1649977179
transform 1 0 45724 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_497
timestamp 1649977179
transform 1 0 46828 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_503
timestamp 1649977179
transform 1 0 47380 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_505
timestamp 1649977179
transform 1 0 47564 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_517
timestamp 1649977179
transform 1 0 48668 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_529
timestamp 1649977179
transform 1 0 49772 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_541
timestamp 1649977179
transform 1 0 50876 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_553
timestamp 1649977179
transform 1 0 51980 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_559
timestamp 1649977179
transform 1 0 52532 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_561
timestamp 1649977179
transform 1 0 52716 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_573
timestamp 1649977179
transform 1 0 53820 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_585
timestamp 1649977179
transform 1 0 54924 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_597
timestamp 1649977179
transform 1 0 56028 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_609
timestamp 1649977179
transform 1 0 57132 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_615
timestamp 1649977179
transform 1 0 57684 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_617
timestamp 1649977179
transform 1 0 57868 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_629
timestamp 1649977179
transform 1 0 58972 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_641
timestamp 1649977179
transform 1 0 60076 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_653
timestamp 1649977179
transform 1 0 61180 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_665
timestamp 1649977179
transform 1 0 62284 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_671
timestamp 1649977179
transform 1 0 62836 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_673
timestamp 1649977179
transform 1 0 63020 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_685
timestamp 1649977179
transform 1 0 64124 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_697
timestamp 1649977179
transform 1 0 65228 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_709
timestamp 1649977179
transform 1 0 66332 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_721
timestamp 1649977179
transform 1 0 67436 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_727
timestamp 1649977179
transform 1 0 67988 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_729
timestamp 1649977179
transform 1 0 68172 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_3
timestamp 1649977179
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_15
timestamp 1649977179
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1649977179
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_29
timestamp 1649977179
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_41
timestamp 1649977179
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_53
timestamp 1649977179
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_65
timestamp 1649977179
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1649977179
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1649977179
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_85
timestamp 1649977179
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_97
timestamp 1649977179
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_109
timestamp 1649977179
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_121
timestamp 1649977179
transform 1 0 12236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_133
timestamp 1649977179
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1649977179
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_141
timestamp 1649977179
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_153
timestamp 1649977179
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_165
timestamp 1649977179
transform 1 0 16284 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_177
timestamp 1649977179
transform 1 0 17388 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_189
timestamp 1649977179
transform 1 0 18492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 1649977179
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_197
timestamp 1649977179
transform 1 0 19228 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_209
timestamp 1649977179
transform 1 0 20332 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_221
timestamp 1649977179
transform 1 0 21436 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_233
timestamp 1649977179
transform 1 0 22540 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_245
timestamp 1649977179
transform 1 0 23644 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_251
timestamp 1649977179
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_253
timestamp 1649977179
transform 1 0 24380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_265
timestamp 1649977179
transform 1 0 25484 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_277
timestamp 1649977179
transform 1 0 26588 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_289
timestamp 1649977179
transform 1 0 27692 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_301
timestamp 1649977179
transform 1 0 28796 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_307
timestamp 1649977179
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_309
timestamp 1649977179
transform 1 0 29532 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_321
timestamp 1649977179
transform 1 0 30636 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_333
timestamp 1649977179
transform 1 0 31740 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_345
timestamp 1649977179
transform 1 0 32844 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_357
timestamp 1649977179
transform 1 0 33948 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_363
timestamp 1649977179
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_365
timestamp 1649977179
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_377
timestamp 1649977179
transform 1 0 35788 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_389
timestamp 1649977179
transform 1 0 36892 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_401
timestamp 1649977179
transform 1 0 37996 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_413
timestamp 1649977179
transform 1 0 39100 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_419
timestamp 1649977179
transform 1 0 39652 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_421
timestamp 1649977179
transform 1 0 39836 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_433
timestamp 1649977179
transform 1 0 40940 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_445
timestamp 1649977179
transform 1 0 42044 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_457
timestamp 1649977179
transform 1 0 43148 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_469
timestamp 1649977179
transform 1 0 44252 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_475
timestamp 1649977179
transform 1 0 44804 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_477
timestamp 1649977179
transform 1 0 44988 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_489
timestamp 1649977179
transform 1 0 46092 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_501
timestamp 1649977179
transform 1 0 47196 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_513
timestamp 1649977179
transform 1 0 48300 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_525
timestamp 1649977179
transform 1 0 49404 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_531
timestamp 1649977179
transform 1 0 49956 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_533
timestamp 1649977179
transform 1 0 50140 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_545
timestamp 1649977179
transform 1 0 51244 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_557
timestamp 1649977179
transform 1 0 52348 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_569
timestamp 1649977179
transform 1 0 53452 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_581
timestamp 1649977179
transform 1 0 54556 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_587
timestamp 1649977179
transform 1 0 55108 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_589
timestamp 1649977179
transform 1 0 55292 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_601
timestamp 1649977179
transform 1 0 56396 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_613
timestamp 1649977179
transform 1 0 57500 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_625
timestamp 1649977179
transform 1 0 58604 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_637
timestamp 1649977179
transform 1 0 59708 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_643
timestamp 1649977179
transform 1 0 60260 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_645
timestamp 1649977179
transform 1 0 60444 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_657
timestamp 1649977179
transform 1 0 61548 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_669
timestamp 1649977179
transform 1 0 62652 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_681
timestamp 1649977179
transform 1 0 63756 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_693
timestamp 1649977179
transform 1 0 64860 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_699
timestamp 1649977179
transform 1 0 65412 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_701
timestamp 1649977179
transform 1 0 65596 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_713
timestamp 1649977179
transform 1 0 66700 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_725
timestamp 1649977179
transform 1 0 67804 0 1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_65_3
timestamp 1649977179
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_15
timestamp 1649977179
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_27
timestamp 1649977179
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_39
timestamp 1649977179
transform 1 0 4692 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_51
timestamp 1649977179
transform 1 0 5796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1649977179
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_57
timestamp 1649977179
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_69
timestamp 1649977179
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_81
timestamp 1649977179
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_93
timestamp 1649977179
transform 1 0 9660 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_105
timestamp 1649977179
transform 1 0 10764 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_111
timestamp 1649977179
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_113
timestamp 1649977179
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_125
timestamp 1649977179
transform 1 0 12604 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_137
timestamp 1649977179
transform 1 0 13708 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_149
timestamp 1649977179
transform 1 0 14812 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_161
timestamp 1649977179
transform 1 0 15916 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_167
timestamp 1649977179
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_169
timestamp 1649977179
transform 1 0 16652 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_181
timestamp 1649977179
transform 1 0 17756 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_193
timestamp 1649977179
transform 1 0 18860 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_205
timestamp 1649977179
transform 1 0 19964 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_217
timestamp 1649977179
transform 1 0 21068 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_223
timestamp 1649977179
transform 1 0 21620 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_225
timestamp 1649977179
transform 1 0 21804 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_237
timestamp 1649977179
transform 1 0 22908 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_249
timestamp 1649977179
transform 1 0 24012 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_261
timestamp 1649977179
transform 1 0 25116 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_273
timestamp 1649977179
transform 1 0 26220 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_279
timestamp 1649977179
transform 1 0 26772 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_281
timestamp 1649977179
transform 1 0 26956 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_293
timestamp 1649977179
transform 1 0 28060 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_305
timestamp 1649977179
transform 1 0 29164 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_317
timestamp 1649977179
transform 1 0 30268 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_329
timestamp 1649977179
transform 1 0 31372 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_335
timestamp 1649977179
transform 1 0 31924 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_337
timestamp 1649977179
transform 1 0 32108 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_349
timestamp 1649977179
transform 1 0 33212 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_361
timestamp 1649977179
transform 1 0 34316 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_373
timestamp 1649977179
transform 1 0 35420 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_385
timestamp 1649977179
transform 1 0 36524 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_391
timestamp 1649977179
transform 1 0 37076 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_393
timestamp 1649977179
transform 1 0 37260 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_405
timestamp 1649977179
transform 1 0 38364 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_417
timestamp 1649977179
transform 1 0 39468 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_429
timestamp 1649977179
transform 1 0 40572 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_441
timestamp 1649977179
transform 1 0 41676 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_447
timestamp 1649977179
transform 1 0 42228 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_449
timestamp 1649977179
transform 1 0 42412 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_461
timestamp 1649977179
transform 1 0 43516 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_473
timestamp 1649977179
transform 1 0 44620 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_485
timestamp 1649977179
transform 1 0 45724 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_497
timestamp 1649977179
transform 1 0 46828 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_503
timestamp 1649977179
transform 1 0 47380 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_505
timestamp 1649977179
transform 1 0 47564 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_517
timestamp 1649977179
transform 1 0 48668 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_529
timestamp 1649977179
transform 1 0 49772 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_541
timestamp 1649977179
transform 1 0 50876 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_553
timestamp 1649977179
transform 1 0 51980 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_559
timestamp 1649977179
transform 1 0 52532 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_561
timestamp 1649977179
transform 1 0 52716 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_573
timestamp 1649977179
transform 1 0 53820 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_585
timestamp 1649977179
transform 1 0 54924 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_597
timestamp 1649977179
transform 1 0 56028 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_609
timestamp 1649977179
transform 1 0 57132 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_615
timestamp 1649977179
transform 1 0 57684 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_617
timestamp 1649977179
transform 1 0 57868 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_629
timestamp 1649977179
transform 1 0 58972 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_641
timestamp 1649977179
transform 1 0 60076 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_653
timestamp 1649977179
transform 1 0 61180 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_665
timestamp 1649977179
transform 1 0 62284 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_671
timestamp 1649977179
transform 1 0 62836 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_673
timestamp 1649977179
transform 1 0 63020 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_685
timestamp 1649977179
transform 1 0 64124 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_697
timestamp 1649977179
transform 1 0 65228 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_709
timestamp 1649977179
transform 1 0 66332 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_721
timestamp 1649977179
transform 1 0 67436 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_727
timestamp 1649977179
transform 1 0 67988 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_729
timestamp 1649977179
transform 1 0 68172 0 -1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_66_3
timestamp 1649977179
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_15
timestamp 1649977179
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1649977179
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_29
timestamp 1649977179
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_41
timestamp 1649977179
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_53
timestamp 1649977179
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_65
timestamp 1649977179
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_77
timestamp 1649977179
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1649977179
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_85
timestamp 1649977179
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_97
timestamp 1649977179
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_109
timestamp 1649977179
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_121
timestamp 1649977179
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_133
timestamp 1649977179
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 1649977179
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_141
timestamp 1649977179
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_153
timestamp 1649977179
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_165
timestamp 1649977179
transform 1 0 16284 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_177
timestamp 1649977179
transform 1 0 17388 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_189
timestamp 1649977179
transform 1 0 18492 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_195
timestamp 1649977179
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_197
timestamp 1649977179
transform 1 0 19228 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_209
timestamp 1649977179
transform 1 0 20332 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_221
timestamp 1649977179
transform 1 0 21436 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_233
timestamp 1649977179
transform 1 0 22540 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_245
timestamp 1649977179
transform 1 0 23644 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_251
timestamp 1649977179
transform 1 0 24196 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_253
timestamp 1649977179
transform 1 0 24380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_265
timestamp 1649977179
transform 1 0 25484 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_277
timestamp 1649977179
transform 1 0 26588 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_289
timestamp 1649977179
transform 1 0 27692 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_301
timestamp 1649977179
transform 1 0 28796 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_307
timestamp 1649977179
transform 1 0 29348 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_309
timestamp 1649977179
transform 1 0 29532 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_321
timestamp 1649977179
transform 1 0 30636 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_333
timestamp 1649977179
transform 1 0 31740 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_345
timestamp 1649977179
transform 1 0 32844 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_357
timestamp 1649977179
transform 1 0 33948 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_363
timestamp 1649977179
transform 1 0 34500 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_365
timestamp 1649977179
transform 1 0 34684 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_377
timestamp 1649977179
transform 1 0 35788 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_389
timestamp 1649977179
transform 1 0 36892 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_401
timestamp 1649977179
transform 1 0 37996 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_413
timestamp 1649977179
transform 1 0 39100 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_419
timestamp 1649977179
transform 1 0 39652 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_421
timestamp 1649977179
transform 1 0 39836 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_433
timestamp 1649977179
transform 1 0 40940 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_445
timestamp 1649977179
transform 1 0 42044 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_457
timestamp 1649977179
transform 1 0 43148 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_469
timestamp 1649977179
transform 1 0 44252 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_475
timestamp 1649977179
transform 1 0 44804 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_477
timestamp 1649977179
transform 1 0 44988 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_489
timestamp 1649977179
transform 1 0 46092 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_501
timestamp 1649977179
transform 1 0 47196 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_513
timestamp 1649977179
transform 1 0 48300 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_525
timestamp 1649977179
transform 1 0 49404 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_531
timestamp 1649977179
transform 1 0 49956 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_533
timestamp 1649977179
transform 1 0 50140 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_545
timestamp 1649977179
transform 1 0 51244 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_557
timestamp 1649977179
transform 1 0 52348 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_569
timestamp 1649977179
transform 1 0 53452 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_581
timestamp 1649977179
transform 1 0 54556 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_587
timestamp 1649977179
transform 1 0 55108 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_589
timestamp 1649977179
transform 1 0 55292 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_601
timestamp 1649977179
transform 1 0 56396 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_613
timestamp 1649977179
transform 1 0 57500 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_625
timestamp 1649977179
transform 1 0 58604 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_637
timestamp 1649977179
transform 1 0 59708 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_643
timestamp 1649977179
transform 1 0 60260 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_645
timestamp 1649977179
transform 1 0 60444 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_657
timestamp 1649977179
transform 1 0 61548 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_669
timestamp 1649977179
transform 1 0 62652 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_681
timestamp 1649977179
transform 1 0 63756 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_693
timestamp 1649977179
transform 1 0 64860 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_699
timestamp 1649977179
transform 1 0 65412 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_701
timestamp 1649977179
transform 1 0 65596 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_713
timestamp 1649977179
transform 1 0 66700 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_725
timestamp 1649977179
transform 1 0 67804 0 1 38080
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_67_3
timestamp 1649977179
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_15
timestamp 1649977179
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_27
timestamp 1649977179
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_39
timestamp 1649977179
transform 1 0 4692 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_51
timestamp 1649977179
transform 1 0 5796 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_55
timestamp 1649977179
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_57
timestamp 1649977179
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_69
timestamp 1649977179
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_81
timestamp 1649977179
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_93
timestamp 1649977179
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_105
timestamp 1649977179
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 1649977179
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_113
timestamp 1649977179
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_125
timestamp 1649977179
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_137
timestamp 1649977179
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_149
timestamp 1649977179
transform 1 0 14812 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_161
timestamp 1649977179
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_167
timestamp 1649977179
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_169
timestamp 1649977179
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_181
timestamp 1649977179
transform 1 0 17756 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_193
timestamp 1649977179
transform 1 0 18860 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_205
timestamp 1649977179
transform 1 0 19964 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_217
timestamp 1649977179
transform 1 0 21068 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_223
timestamp 1649977179
transform 1 0 21620 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_225
timestamp 1649977179
transform 1 0 21804 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_237
timestamp 1649977179
transform 1 0 22908 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_249
timestamp 1649977179
transform 1 0 24012 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_261
timestamp 1649977179
transform 1 0 25116 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_273
timestamp 1649977179
transform 1 0 26220 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_279
timestamp 1649977179
transform 1 0 26772 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_281
timestamp 1649977179
transform 1 0 26956 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_293
timestamp 1649977179
transform 1 0 28060 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_305
timestamp 1649977179
transform 1 0 29164 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_317
timestamp 1649977179
transform 1 0 30268 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_329
timestamp 1649977179
transform 1 0 31372 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_335
timestamp 1649977179
transform 1 0 31924 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_337
timestamp 1649977179
transform 1 0 32108 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_349
timestamp 1649977179
transform 1 0 33212 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_361
timestamp 1649977179
transform 1 0 34316 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_373
timestamp 1649977179
transform 1 0 35420 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_385
timestamp 1649977179
transform 1 0 36524 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_391
timestamp 1649977179
transform 1 0 37076 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_393
timestamp 1649977179
transform 1 0 37260 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_405
timestamp 1649977179
transform 1 0 38364 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_417
timestamp 1649977179
transform 1 0 39468 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_429
timestamp 1649977179
transform 1 0 40572 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_441
timestamp 1649977179
transform 1 0 41676 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_447
timestamp 1649977179
transform 1 0 42228 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_449
timestamp 1649977179
transform 1 0 42412 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_461
timestamp 1649977179
transform 1 0 43516 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_473
timestamp 1649977179
transform 1 0 44620 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_485
timestamp 1649977179
transform 1 0 45724 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_497
timestamp 1649977179
transform 1 0 46828 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_503
timestamp 1649977179
transform 1 0 47380 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_505
timestamp 1649977179
transform 1 0 47564 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_517
timestamp 1649977179
transform 1 0 48668 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_529
timestamp 1649977179
transform 1 0 49772 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_541
timestamp 1649977179
transform 1 0 50876 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_553
timestamp 1649977179
transform 1 0 51980 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_559
timestamp 1649977179
transform 1 0 52532 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_561
timestamp 1649977179
transform 1 0 52716 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_573
timestamp 1649977179
transform 1 0 53820 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_585
timestamp 1649977179
transform 1 0 54924 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_597
timestamp 1649977179
transform 1 0 56028 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_609
timestamp 1649977179
transform 1 0 57132 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_615
timestamp 1649977179
transform 1 0 57684 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_617
timestamp 1649977179
transform 1 0 57868 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_629
timestamp 1649977179
transform 1 0 58972 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_641
timestamp 1649977179
transform 1 0 60076 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_653
timestamp 1649977179
transform 1 0 61180 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_665
timestamp 1649977179
transform 1 0 62284 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_671
timestamp 1649977179
transform 1 0 62836 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_673
timestamp 1649977179
transform 1 0 63020 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_685
timestamp 1649977179
transform 1 0 64124 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_697
timestamp 1649977179
transform 1 0 65228 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_709
timestamp 1649977179
transform 1 0 66332 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_721
timestamp 1649977179
transform 1 0 67436 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_727
timestamp 1649977179
transform 1 0 67988 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_729
timestamp 1649977179
transform 1 0 68172 0 -1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_68_3
timestamp 1649977179
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_15
timestamp 1649977179
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1649977179
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_29
timestamp 1649977179
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_41
timestamp 1649977179
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_53
timestamp 1649977179
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_65
timestamp 1649977179
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_77
timestamp 1649977179
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 1649977179
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_85
timestamp 1649977179
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_97
timestamp 1649977179
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_109
timestamp 1649977179
transform 1 0 11132 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_121
timestamp 1649977179
transform 1 0 12236 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_133
timestamp 1649977179
transform 1 0 13340 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_139
timestamp 1649977179
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_141
timestamp 1649977179
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_153
timestamp 1649977179
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_165
timestamp 1649977179
transform 1 0 16284 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_177
timestamp 1649977179
transform 1 0 17388 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_189
timestamp 1649977179
transform 1 0 18492 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_195
timestamp 1649977179
transform 1 0 19044 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_197
timestamp 1649977179
transform 1 0 19228 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_209
timestamp 1649977179
transform 1 0 20332 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_221
timestamp 1649977179
transform 1 0 21436 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_233
timestamp 1649977179
transform 1 0 22540 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_245
timestamp 1649977179
transform 1 0 23644 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_251
timestamp 1649977179
transform 1 0 24196 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_253
timestamp 1649977179
transform 1 0 24380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_265
timestamp 1649977179
transform 1 0 25484 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_277
timestamp 1649977179
transform 1 0 26588 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_289
timestamp 1649977179
transform 1 0 27692 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_301
timestamp 1649977179
transform 1 0 28796 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_307
timestamp 1649977179
transform 1 0 29348 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_309
timestamp 1649977179
transform 1 0 29532 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_321
timestamp 1649977179
transform 1 0 30636 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_333
timestamp 1649977179
transform 1 0 31740 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_345
timestamp 1649977179
transform 1 0 32844 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_357
timestamp 1649977179
transform 1 0 33948 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_363
timestamp 1649977179
transform 1 0 34500 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_365
timestamp 1649977179
transform 1 0 34684 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_377
timestamp 1649977179
transform 1 0 35788 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_389
timestamp 1649977179
transform 1 0 36892 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_401
timestamp 1649977179
transform 1 0 37996 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_413
timestamp 1649977179
transform 1 0 39100 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_419
timestamp 1649977179
transform 1 0 39652 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_421
timestamp 1649977179
transform 1 0 39836 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_433
timestamp 1649977179
transform 1 0 40940 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_445
timestamp 1649977179
transform 1 0 42044 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_457
timestamp 1649977179
transform 1 0 43148 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_469
timestamp 1649977179
transform 1 0 44252 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_475
timestamp 1649977179
transform 1 0 44804 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_477
timestamp 1649977179
transform 1 0 44988 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_489
timestamp 1649977179
transform 1 0 46092 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_501
timestamp 1649977179
transform 1 0 47196 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_513
timestamp 1649977179
transform 1 0 48300 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_525
timestamp 1649977179
transform 1 0 49404 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_531
timestamp 1649977179
transform 1 0 49956 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_533
timestamp 1649977179
transform 1 0 50140 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_545
timestamp 1649977179
transform 1 0 51244 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_557
timestamp 1649977179
transform 1 0 52348 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_569
timestamp 1649977179
transform 1 0 53452 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_581
timestamp 1649977179
transform 1 0 54556 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_587
timestamp 1649977179
transform 1 0 55108 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_589
timestamp 1649977179
transform 1 0 55292 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_601
timestamp 1649977179
transform 1 0 56396 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_613
timestamp 1649977179
transform 1 0 57500 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_625
timestamp 1649977179
transform 1 0 58604 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_637
timestamp 1649977179
transform 1 0 59708 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_643
timestamp 1649977179
transform 1 0 60260 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_645
timestamp 1649977179
transform 1 0 60444 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_657
timestamp 1649977179
transform 1 0 61548 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_669
timestamp 1649977179
transform 1 0 62652 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_681
timestamp 1649977179
transform 1 0 63756 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_693
timestamp 1649977179
transform 1 0 64860 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_699
timestamp 1649977179
transform 1 0 65412 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_701
timestamp 1649977179
transform 1 0 65596 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_713
timestamp 1649977179
transform 1 0 66700 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_725
timestamp 1649977179
transform 1 0 67804 0 1 39168
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_69_3
timestamp 1649977179
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_15
timestamp 1649977179
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_27
timestamp 1649977179
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_39
timestamp 1649977179
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_51
timestamp 1649977179
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1649977179
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_57
timestamp 1649977179
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_69
timestamp 1649977179
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_81
timestamp 1649977179
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_93
timestamp 1649977179
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_105
timestamp 1649977179
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_111
timestamp 1649977179
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_113
timestamp 1649977179
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_125
timestamp 1649977179
transform 1 0 12604 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_137
timestamp 1649977179
transform 1 0 13708 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_149
timestamp 1649977179
transform 1 0 14812 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_161
timestamp 1649977179
transform 1 0 15916 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_167
timestamp 1649977179
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_169
timestamp 1649977179
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_181
timestamp 1649977179
transform 1 0 17756 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_193
timestamp 1649977179
transform 1 0 18860 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_205
timestamp 1649977179
transform 1 0 19964 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_217
timestamp 1649977179
transform 1 0 21068 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_223
timestamp 1649977179
transform 1 0 21620 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_225
timestamp 1649977179
transform 1 0 21804 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_237
timestamp 1649977179
transform 1 0 22908 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_249
timestamp 1649977179
transform 1 0 24012 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_261
timestamp 1649977179
transform 1 0 25116 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_273
timestamp 1649977179
transform 1 0 26220 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_279
timestamp 1649977179
transform 1 0 26772 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_281
timestamp 1649977179
transform 1 0 26956 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_293
timestamp 1649977179
transform 1 0 28060 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_305
timestamp 1649977179
transform 1 0 29164 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_317
timestamp 1649977179
transform 1 0 30268 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_329
timestamp 1649977179
transform 1 0 31372 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_335
timestamp 1649977179
transform 1 0 31924 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_337
timestamp 1649977179
transform 1 0 32108 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_349
timestamp 1649977179
transform 1 0 33212 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_361
timestamp 1649977179
transform 1 0 34316 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_373
timestamp 1649977179
transform 1 0 35420 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_385
timestamp 1649977179
transform 1 0 36524 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_391
timestamp 1649977179
transform 1 0 37076 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_393
timestamp 1649977179
transform 1 0 37260 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_405
timestamp 1649977179
transform 1 0 38364 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_417
timestamp 1649977179
transform 1 0 39468 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_429
timestamp 1649977179
transform 1 0 40572 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_441
timestamp 1649977179
transform 1 0 41676 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_447
timestamp 1649977179
transform 1 0 42228 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_449
timestamp 1649977179
transform 1 0 42412 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_461
timestamp 1649977179
transform 1 0 43516 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_473
timestamp 1649977179
transform 1 0 44620 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_485
timestamp 1649977179
transform 1 0 45724 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_497
timestamp 1649977179
transform 1 0 46828 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_503
timestamp 1649977179
transform 1 0 47380 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_505
timestamp 1649977179
transform 1 0 47564 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_517
timestamp 1649977179
transform 1 0 48668 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_529
timestamp 1649977179
transform 1 0 49772 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_541
timestamp 1649977179
transform 1 0 50876 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_553
timestamp 1649977179
transform 1 0 51980 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_559
timestamp 1649977179
transform 1 0 52532 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_561
timestamp 1649977179
transform 1 0 52716 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_573
timestamp 1649977179
transform 1 0 53820 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_585
timestamp 1649977179
transform 1 0 54924 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_597
timestamp 1649977179
transform 1 0 56028 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_609
timestamp 1649977179
transform 1 0 57132 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_615
timestamp 1649977179
transform 1 0 57684 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_617
timestamp 1649977179
transform 1 0 57868 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_629
timestamp 1649977179
transform 1 0 58972 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_641
timestamp 1649977179
transform 1 0 60076 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_653
timestamp 1649977179
transform 1 0 61180 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_665
timestamp 1649977179
transform 1 0 62284 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_671
timestamp 1649977179
transform 1 0 62836 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_673
timestamp 1649977179
transform 1 0 63020 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_685
timestamp 1649977179
transform 1 0 64124 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_697
timestamp 1649977179
transform 1 0 65228 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_709
timestamp 1649977179
transform 1 0 66332 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_721
timestamp 1649977179
transform 1 0 67436 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_727
timestamp 1649977179
transform 1 0 67988 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_729
timestamp 1649977179
transform 1 0 68172 0 -1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_70_3
timestamp 1649977179
transform 1 0 1380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_15
timestamp 1649977179
transform 1 0 2484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1649977179
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_29
timestamp 1649977179
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_41
timestamp 1649977179
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_53
timestamp 1649977179
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_65
timestamp 1649977179
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_77
timestamp 1649977179
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1649977179
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_85
timestamp 1649977179
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_97
timestamp 1649977179
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_109
timestamp 1649977179
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_121
timestamp 1649977179
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_133
timestamp 1649977179
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_139
timestamp 1649977179
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_141
timestamp 1649977179
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_153
timestamp 1649977179
transform 1 0 15180 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_165
timestamp 1649977179
transform 1 0 16284 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_177
timestamp 1649977179
transform 1 0 17388 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_189
timestamp 1649977179
transform 1 0 18492 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_195
timestamp 1649977179
transform 1 0 19044 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_197
timestamp 1649977179
transform 1 0 19228 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_209
timestamp 1649977179
transform 1 0 20332 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_221
timestamp 1649977179
transform 1 0 21436 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_233
timestamp 1649977179
transform 1 0 22540 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_245
timestamp 1649977179
transform 1 0 23644 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_251
timestamp 1649977179
transform 1 0 24196 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_253
timestamp 1649977179
transform 1 0 24380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_265
timestamp 1649977179
transform 1 0 25484 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_277
timestamp 1649977179
transform 1 0 26588 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_289
timestamp 1649977179
transform 1 0 27692 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_301
timestamp 1649977179
transform 1 0 28796 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_307
timestamp 1649977179
transform 1 0 29348 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_309
timestamp 1649977179
transform 1 0 29532 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_321
timestamp 1649977179
transform 1 0 30636 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_333
timestamp 1649977179
transform 1 0 31740 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_345
timestamp 1649977179
transform 1 0 32844 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_357
timestamp 1649977179
transform 1 0 33948 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_363
timestamp 1649977179
transform 1 0 34500 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_365
timestamp 1649977179
transform 1 0 34684 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_377
timestamp 1649977179
transform 1 0 35788 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_389
timestamp 1649977179
transform 1 0 36892 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_401
timestamp 1649977179
transform 1 0 37996 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_413
timestamp 1649977179
transform 1 0 39100 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_419
timestamp 1649977179
transform 1 0 39652 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_421
timestamp 1649977179
transform 1 0 39836 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_433
timestamp 1649977179
transform 1 0 40940 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_445
timestamp 1649977179
transform 1 0 42044 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_457
timestamp 1649977179
transform 1 0 43148 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_469
timestamp 1649977179
transform 1 0 44252 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_475
timestamp 1649977179
transform 1 0 44804 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_477
timestamp 1649977179
transform 1 0 44988 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_489
timestamp 1649977179
transform 1 0 46092 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_501
timestamp 1649977179
transform 1 0 47196 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_513
timestamp 1649977179
transform 1 0 48300 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_525
timestamp 1649977179
transform 1 0 49404 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_531
timestamp 1649977179
transform 1 0 49956 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_533
timestamp 1649977179
transform 1 0 50140 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_545
timestamp 1649977179
transform 1 0 51244 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_557
timestamp 1649977179
transform 1 0 52348 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_569
timestamp 1649977179
transform 1 0 53452 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_581
timestamp 1649977179
transform 1 0 54556 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_587
timestamp 1649977179
transform 1 0 55108 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_589
timestamp 1649977179
transform 1 0 55292 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_601
timestamp 1649977179
transform 1 0 56396 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_613
timestamp 1649977179
transform 1 0 57500 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_625
timestamp 1649977179
transform 1 0 58604 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_637
timestamp 1649977179
transform 1 0 59708 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_643
timestamp 1649977179
transform 1 0 60260 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_645
timestamp 1649977179
transform 1 0 60444 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_657
timestamp 1649977179
transform 1 0 61548 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_669
timestamp 1649977179
transform 1 0 62652 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_681
timestamp 1649977179
transform 1 0 63756 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_693
timestamp 1649977179
transform 1 0 64860 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_699
timestamp 1649977179
transform 1 0 65412 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_701
timestamp 1649977179
transform 1 0 65596 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_713
timestamp 1649977179
transform 1 0 66700 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_725
timestamp 1649977179
transform 1 0 67804 0 1 40256
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_71_3
timestamp 1649977179
transform 1 0 1380 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_15
timestamp 1649977179
transform 1 0 2484 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_27
timestamp 1649977179
transform 1 0 3588 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_39
timestamp 1649977179
transform 1 0 4692 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_51
timestamp 1649977179
transform 1 0 5796 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_55
timestamp 1649977179
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_57
timestamp 1649977179
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_69
timestamp 1649977179
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_81
timestamp 1649977179
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_93
timestamp 1649977179
transform 1 0 9660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_105
timestamp 1649977179
transform 1 0 10764 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_111
timestamp 1649977179
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_113
timestamp 1649977179
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_125
timestamp 1649977179
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_137
timestamp 1649977179
transform 1 0 13708 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_149
timestamp 1649977179
transform 1 0 14812 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_161
timestamp 1649977179
transform 1 0 15916 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_167
timestamp 1649977179
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_169
timestamp 1649977179
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_181
timestamp 1649977179
transform 1 0 17756 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_193
timestamp 1649977179
transform 1 0 18860 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_205
timestamp 1649977179
transform 1 0 19964 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_217
timestamp 1649977179
transform 1 0 21068 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_223
timestamp 1649977179
transform 1 0 21620 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_225
timestamp 1649977179
transform 1 0 21804 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_237
timestamp 1649977179
transform 1 0 22908 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_249
timestamp 1649977179
transform 1 0 24012 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_261
timestamp 1649977179
transform 1 0 25116 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_273
timestamp 1649977179
transform 1 0 26220 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_279
timestamp 1649977179
transform 1 0 26772 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_281
timestamp 1649977179
transform 1 0 26956 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_293
timestamp 1649977179
transform 1 0 28060 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_305
timestamp 1649977179
transform 1 0 29164 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_317
timestamp 1649977179
transform 1 0 30268 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_329
timestamp 1649977179
transform 1 0 31372 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_335
timestamp 1649977179
transform 1 0 31924 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_337
timestamp 1649977179
transform 1 0 32108 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_349
timestamp 1649977179
transform 1 0 33212 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_361
timestamp 1649977179
transform 1 0 34316 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_373
timestamp 1649977179
transform 1 0 35420 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_385
timestamp 1649977179
transform 1 0 36524 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_391
timestamp 1649977179
transform 1 0 37076 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_393
timestamp 1649977179
transform 1 0 37260 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_405
timestamp 1649977179
transform 1 0 38364 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_417
timestamp 1649977179
transform 1 0 39468 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_429
timestamp 1649977179
transform 1 0 40572 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_441
timestamp 1649977179
transform 1 0 41676 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_447
timestamp 1649977179
transform 1 0 42228 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_449
timestamp 1649977179
transform 1 0 42412 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_461
timestamp 1649977179
transform 1 0 43516 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_473
timestamp 1649977179
transform 1 0 44620 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_485
timestamp 1649977179
transform 1 0 45724 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_497
timestamp 1649977179
transform 1 0 46828 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_503
timestamp 1649977179
transform 1 0 47380 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_505
timestamp 1649977179
transform 1 0 47564 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_517
timestamp 1649977179
transform 1 0 48668 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_529
timestamp 1649977179
transform 1 0 49772 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_541
timestamp 1649977179
transform 1 0 50876 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_553
timestamp 1649977179
transform 1 0 51980 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_559
timestamp 1649977179
transform 1 0 52532 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_561
timestamp 1649977179
transform 1 0 52716 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_573
timestamp 1649977179
transform 1 0 53820 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_585
timestamp 1649977179
transform 1 0 54924 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_597
timestamp 1649977179
transform 1 0 56028 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_609
timestamp 1649977179
transform 1 0 57132 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_615
timestamp 1649977179
transform 1 0 57684 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_617
timestamp 1649977179
transform 1 0 57868 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_629
timestamp 1649977179
transform 1 0 58972 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_641
timestamp 1649977179
transform 1 0 60076 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_653
timestamp 1649977179
transform 1 0 61180 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_665
timestamp 1649977179
transform 1 0 62284 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_671
timestamp 1649977179
transform 1 0 62836 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_673
timestamp 1649977179
transform 1 0 63020 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_685
timestamp 1649977179
transform 1 0 64124 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_697
timestamp 1649977179
transform 1 0 65228 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_709
timestamp 1649977179
transform 1 0 66332 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_721
timestamp 1649977179
transform 1 0 67436 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_727
timestamp 1649977179
transform 1 0 67988 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_729
timestamp 1649977179
transform 1 0 68172 0 -1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_72_3
timestamp 1649977179
transform 1 0 1380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_15
timestamp 1649977179
transform 1 0 2484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_27
timestamp 1649977179
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_29
timestamp 1649977179
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_41
timestamp 1649977179
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_53
timestamp 1649977179
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_65
timestamp 1649977179
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_77
timestamp 1649977179
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1649977179
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_85
timestamp 1649977179
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_97
timestamp 1649977179
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_109
timestamp 1649977179
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_121
timestamp 1649977179
transform 1 0 12236 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_133
timestamp 1649977179
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 1649977179
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_141
timestamp 1649977179
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_153
timestamp 1649977179
transform 1 0 15180 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_165
timestamp 1649977179
transform 1 0 16284 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_177
timestamp 1649977179
transform 1 0 17388 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_189
timestamp 1649977179
transform 1 0 18492 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_195
timestamp 1649977179
transform 1 0 19044 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_197
timestamp 1649977179
transform 1 0 19228 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_209
timestamp 1649977179
transform 1 0 20332 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_221
timestamp 1649977179
transform 1 0 21436 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_233
timestamp 1649977179
transform 1 0 22540 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_245
timestamp 1649977179
transform 1 0 23644 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_251
timestamp 1649977179
transform 1 0 24196 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_253
timestamp 1649977179
transform 1 0 24380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_265
timestamp 1649977179
transform 1 0 25484 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_277
timestamp 1649977179
transform 1 0 26588 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_289
timestamp 1649977179
transform 1 0 27692 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_301
timestamp 1649977179
transform 1 0 28796 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_307
timestamp 1649977179
transform 1 0 29348 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_309
timestamp 1649977179
transform 1 0 29532 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_321
timestamp 1649977179
transform 1 0 30636 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_333
timestamp 1649977179
transform 1 0 31740 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_345
timestamp 1649977179
transform 1 0 32844 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_357
timestamp 1649977179
transform 1 0 33948 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_363
timestamp 1649977179
transform 1 0 34500 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_365
timestamp 1649977179
transform 1 0 34684 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_377
timestamp 1649977179
transform 1 0 35788 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_389
timestamp 1649977179
transform 1 0 36892 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_401
timestamp 1649977179
transform 1 0 37996 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_413
timestamp 1649977179
transform 1 0 39100 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_419
timestamp 1649977179
transform 1 0 39652 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_421
timestamp 1649977179
transform 1 0 39836 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_433
timestamp 1649977179
transform 1 0 40940 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_445
timestamp 1649977179
transform 1 0 42044 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_457
timestamp 1649977179
transform 1 0 43148 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_469
timestamp 1649977179
transform 1 0 44252 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_475
timestamp 1649977179
transform 1 0 44804 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_477
timestamp 1649977179
transform 1 0 44988 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_489
timestamp 1649977179
transform 1 0 46092 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_501
timestamp 1649977179
transform 1 0 47196 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_513
timestamp 1649977179
transform 1 0 48300 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_525
timestamp 1649977179
transform 1 0 49404 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_531
timestamp 1649977179
transform 1 0 49956 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_533
timestamp 1649977179
transform 1 0 50140 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_545
timestamp 1649977179
transform 1 0 51244 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_557
timestamp 1649977179
transform 1 0 52348 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_569
timestamp 1649977179
transform 1 0 53452 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_581
timestamp 1649977179
transform 1 0 54556 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_587
timestamp 1649977179
transform 1 0 55108 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_589
timestamp 1649977179
transform 1 0 55292 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_601
timestamp 1649977179
transform 1 0 56396 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_613
timestamp 1649977179
transform 1 0 57500 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_625
timestamp 1649977179
transform 1 0 58604 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_637
timestamp 1649977179
transform 1 0 59708 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_643
timestamp 1649977179
transform 1 0 60260 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_645
timestamp 1649977179
transform 1 0 60444 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_657
timestamp 1649977179
transform 1 0 61548 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_669
timestamp 1649977179
transform 1 0 62652 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_681
timestamp 1649977179
transform 1 0 63756 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_693
timestamp 1649977179
transform 1 0 64860 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_699
timestamp 1649977179
transform 1 0 65412 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_701
timestamp 1649977179
transform 1 0 65596 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_713
timestamp 1649977179
transform 1 0 66700 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_725
timestamp 1649977179
transform 1 0 67804 0 1 41344
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_73_3
timestamp 1649977179
transform 1 0 1380 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_15
timestamp 1649977179
transform 1 0 2484 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_27
timestamp 1649977179
transform 1 0 3588 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_39
timestamp 1649977179
transform 1 0 4692 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_51
timestamp 1649977179
transform 1 0 5796 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 1649977179
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_57
timestamp 1649977179
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_69
timestamp 1649977179
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_81
timestamp 1649977179
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_93
timestamp 1649977179
transform 1 0 9660 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_105
timestamp 1649977179
transform 1 0 10764 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_111
timestamp 1649977179
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_113
timestamp 1649977179
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_125
timestamp 1649977179
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_137
timestamp 1649977179
transform 1 0 13708 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_149
timestamp 1649977179
transform 1 0 14812 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_161
timestamp 1649977179
transform 1 0 15916 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_167
timestamp 1649977179
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_169
timestamp 1649977179
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_181
timestamp 1649977179
transform 1 0 17756 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_193
timestamp 1649977179
transform 1 0 18860 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_205
timestamp 1649977179
transform 1 0 19964 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_217
timestamp 1649977179
transform 1 0 21068 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_223
timestamp 1649977179
transform 1 0 21620 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_225
timestamp 1649977179
transform 1 0 21804 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_237
timestamp 1649977179
transform 1 0 22908 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_249
timestamp 1649977179
transform 1 0 24012 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_261
timestamp 1649977179
transform 1 0 25116 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_273
timestamp 1649977179
transform 1 0 26220 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_279
timestamp 1649977179
transform 1 0 26772 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_281
timestamp 1649977179
transform 1 0 26956 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_293
timestamp 1649977179
transform 1 0 28060 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_305
timestamp 1649977179
transform 1 0 29164 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_317
timestamp 1649977179
transform 1 0 30268 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_329
timestamp 1649977179
transform 1 0 31372 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_335
timestamp 1649977179
transform 1 0 31924 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_337
timestamp 1649977179
transform 1 0 32108 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_349
timestamp 1649977179
transform 1 0 33212 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_361
timestamp 1649977179
transform 1 0 34316 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_373
timestamp 1649977179
transform 1 0 35420 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_385
timestamp 1649977179
transform 1 0 36524 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_391
timestamp 1649977179
transform 1 0 37076 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_393
timestamp 1649977179
transform 1 0 37260 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_405
timestamp 1649977179
transform 1 0 38364 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_417
timestamp 1649977179
transform 1 0 39468 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_429
timestamp 1649977179
transform 1 0 40572 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_441
timestamp 1649977179
transform 1 0 41676 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_447
timestamp 1649977179
transform 1 0 42228 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_449
timestamp 1649977179
transform 1 0 42412 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_461
timestamp 1649977179
transform 1 0 43516 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_473
timestamp 1649977179
transform 1 0 44620 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_485
timestamp 1649977179
transform 1 0 45724 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_497
timestamp 1649977179
transform 1 0 46828 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_503
timestamp 1649977179
transform 1 0 47380 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_505
timestamp 1649977179
transform 1 0 47564 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_517
timestamp 1649977179
transform 1 0 48668 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_529
timestamp 1649977179
transform 1 0 49772 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_541
timestamp 1649977179
transform 1 0 50876 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_553
timestamp 1649977179
transform 1 0 51980 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_559
timestamp 1649977179
transform 1 0 52532 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_561
timestamp 1649977179
transform 1 0 52716 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_573
timestamp 1649977179
transform 1 0 53820 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_585
timestamp 1649977179
transform 1 0 54924 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_597
timestamp 1649977179
transform 1 0 56028 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_609
timestamp 1649977179
transform 1 0 57132 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_615
timestamp 1649977179
transform 1 0 57684 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_617
timestamp 1649977179
transform 1 0 57868 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_629
timestamp 1649977179
transform 1 0 58972 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_641
timestamp 1649977179
transform 1 0 60076 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_653
timestamp 1649977179
transform 1 0 61180 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_665
timestamp 1649977179
transform 1 0 62284 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_671
timestamp 1649977179
transform 1 0 62836 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_673
timestamp 1649977179
transform 1 0 63020 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_685
timestamp 1649977179
transform 1 0 64124 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_697
timestamp 1649977179
transform 1 0 65228 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_709
timestamp 1649977179
transform 1 0 66332 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_721
timestamp 1649977179
transform 1 0 67436 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_727
timestamp 1649977179
transform 1 0 67988 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_729
timestamp 1649977179
transform 1 0 68172 0 -1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_74_3
timestamp 1649977179
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_15
timestamp 1649977179
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1649977179
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_29
timestamp 1649977179
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_41
timestamp 1649977179
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_53
timestamp 1649977179
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_65
timestamp 1649977179
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_77
timestamp 1649977179
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 1649977179
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_85
timestamp 1649977179
transform 1 0 8924 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_97
timestamp 1649977179
transform 1 0 10028 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_109
timestamp 1649977179
transform 1 0 11132 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_121
timestamp 1649977179
transform 1 0 12236 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_133
timestamp 1649977179
transform 1 0 13340 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_139
timestamp 1649977179
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_141
timestamp 1649977179
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_153
timestamp 1649977179
transform 1 0 15180 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_165
timestamp 1649977179
transform 1 0 16284 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_177
timestamp 1649977179
transform 1 0 17388 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_189
timestamp 1649977179
transform 1 0 18492 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_195
timestamp 1649977179
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_197
timestamp 1649977179
transform 1 0 19228 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_209
timestamp 1649977179
transform 1 0 20332 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_221
timestamp 1649977179
transform 1 0 21436 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_233
timestamp 1649977179
transform 1 0 22540 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_245
timestamp 1649977179
transform 1 0 23644 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_251
timestamp 1649977179
transform 1 0 24196 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_253
timestamp 1649977179
transform 1 0 24380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_265
timestamp 1649977179
transform 1 0 25484 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_277
timestamp 1649977179
transform 1 0 26588 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_289
timestamp 1649977179
transform 1 0 27692 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_301
timestamp 1649977179
transform 1 0 28796 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_307
timestamp 1649977179
transform 1 0 29348 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_309
timestamp 1649977179
transform 1 0 29532 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_321
timestamp 1649977179
transform 1 0 30636 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_333
timestamp 1649977179
transform 1 0 31740 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_345
timestamp 1649977179
transform 1 0 32844 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_357
timestamp 1649977179
transform 1 0 33948 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_363
timestamp 1649977179
transform 1 0 34500 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_365
timestamp 1649977179
transform 1 0 34684 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_377
timestamp 1649977179
transform 1 0 35788 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_389
timestamp 1649977179
transform 1 0 36892 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_401
timestamp 1649977179
transform 1 0 37996 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_413
timestamp 1649977179
transform 1 0 39100 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_419
timestamp 1649977179
transform 1 0 39652 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_421
timestamp 1649977179
transform 1 0 39836 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_433
timestamp 1649977179
transform 1 0 40940 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_445
timestamp 1649977179
transform 1 0 42044 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_457
timestamp 1649977179
transform 1 0 43148 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_469
timestamp 1649977179
transform 1 0 44252 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_475
timestamp 1649977179
transform 1 0 44804 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_477
timestamp 1649977179
transform 1 0 44988 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_489
timestamp 1649977179
transform 1 0 46092 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_501
timestamp 1649977179
transform 1 0 47196 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_513
timestamp 1649977179
transform 1 0 48300 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_525
timestamp 1649977179
transform 1 0 49404 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_531
timestamp 1649977179
transform 1 0 49956 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_533
timestamp 1649977179
transform 1 0 50140 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_545
timestamp 1649977179
transform 1 0 51244 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_557
timestamp 1649977179
transform 1 0 52348 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_569
timestamp 1649977179
transform 1 0 53452 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_581
timestamp 1649977179
transform 1 0 54556 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_587
timestamp 1649977179
transform 1 0 55108 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_589
timestamp 1649977179
transform 1 0 55292 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_601
timestamp 1649977179
transform 1 0 56396 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_613
timestamp 1649977179
transform 1 0 57500 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_625
timestamp 1649977179
transform 1 0 58604 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_637
timestamp 1649977179
transform 1 0 59708 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_643
timestamp 1649977179
transform 1 0 60260 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_645
timestamp 1649977179
transform 1 0 60444 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_657
timestamp 1649977179
transform 1 0 61548 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_669
timestamp 1649977179
transform 1 0 62652 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_681
timestamp 1649977179
transform 1 0 63756 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_693
timestamp 1649977179
transform 1 0 64860 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_699
timestamp 1649977179
transform 1 0 65412 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_701
timestamp 1649977179
transform 1 0 65596 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_713
timestamp 1649977179
transform 1 0 66700 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_725
timestamp 1649977179
transform 1 0 67804 0 1 42432
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_75_3
timestamp 1649977179
transform 1 0 1380 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_15
timestamp 1649977179
transform 1 0 2484 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_27
timestamp 1649977179
transform 1 0 3588 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_39
timestamp 1649977179
transform 1 0 4692 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_51
timestamp 1649977179
transform 1 0 5796 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_55
timestamp 1649977179
transform 1 0 6164 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_57
timestamp 1649977179
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_69
timestamp 1649977179
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_81
timestamp 1649977179
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_93
timestamp 1649977179
transform 1 0 9660 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_105
timestamp 1649977179
transform 1 0 10764 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_111
timestamp 1649977179
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_113
timestamp 1649977179
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_125
timestamp 1649977179
transform 1 0 12604 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_137
timestamp 1649977179
transform 1 0 13708 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_149
timestamp 1649977179
transform 1 0 14812 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_161
timestamp 1649977179
transform 1 0 15916 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_167
timestamp 1649977179
transform 1 0 16468 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_169
timestamp 1649977179
transform 1 0 16652 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_181
timestamp 1649977179
transform 1 0 17756 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_193
timestamp 1649977179
transform 1 0 18860 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_205
timestamp 1649977179
transform 1 0 19964 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_217
timestamp 1649977179
transform 1 0 21068 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_223
timestamp 1649977179
transform 1 0 21620 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_225
timestamp 1649977179
transform 1 0 21804 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_237
timestamp 1649977179
transform 1 0 22908 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_249
timestamp 1649977179
transform 1 0 24012 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_261
timestamp 1649977179
transform 1 0 25116 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_273
timestamp 1649977179
transform 1 0 26220 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_279
timestamp 1649977179
transform 1 0 26772 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_281
timestamp 1649977179
transform 1 0 26956 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_293
timestamp 1649977179
transform 1 0 28060 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_305
timestamp 1649977179
transform 1 0 29164 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_317
timestamp 1649977179
transform 1 0 30268 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_329
timestamp 1649977179
transform 1 0 31372 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_335
timestamp 1649977179
transform 1 0 31924 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_337
timestamp 1649977179
transform 1 0 32108 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_349
timestamp 1649977179
transform 1 0 33212 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_361
timestamp 1649977179
transform 1 0 34316 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_373
timestamp 1649977179
transform 1 0 35420 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_385
timestamp 1649977179
transform 1 0 36524 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_391
timestamp 1649977179
transform 1 0 37076 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_393
timestamp 1649977179
transform 1 0 37260 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_405
timestamp 1649977179
transform 1 0 38364 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_417
timestamp 1649977179
transform 1 0 39468 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_429
timestamp 1649977179
transform 1 0 40572 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_441
timestamp 1649977179
transform 1 0 41676 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_447
timestamp 1649977179
transform 1 0 42228 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_449
timestamp 1649977179
transform 1 0 42412 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_461
timestamp 1649977179
transform 1 0 43516 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_473
timestamp 1649977179
transform 1 0 44620 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_485
timestamp 1649977179
transform 1 0 45724 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_497
timestamp 1649977179
transform 1 0 46828 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_503
timestamp 1649977179
transform 1 0 47380 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_505
timestamp 1649977179
transform 1 0 47564 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_517
timestamp 1649977179
transform 1 0 48668 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_529
timestamp 1649977179
transform 1 0 49772 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_541
timestamp 1649977179
transform 1 0 50876 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_553
timestamp 1649977179
transform 1 0 51980 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_559
timestamp 1649977179
transform 1 0 52532 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_561
timestamp 1649977179
transform 1 0 52716 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_573
timestamp 1649977179
transform 1 0 53820 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_585
timestamp 1649977179
transform 1 0 54924 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_597
timestamp 1649977179
transform 1 0 56028 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_609
timestamp 1649977179
transform 1 0 57132 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_615
timestamp 1649977179
transform 1 0 57684 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_617
timestamp 1649977179
transform 1 0 57868 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_629
timestamp 1649977179
transform 1 0 58972 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_641
timestamp 1649977179
transform 1 0 60076 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_653
timestamp 1649977179
transform 1 0 61180 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_665
timestamp 1649977179
transform 1 0 62284 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_671
timestamp 1649977179
transform 1 0 62836 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_673
timestamp 1649977179
transform 1 0 63020 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_685
timestamp 1649977179
transform 1 0 64124 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_697
timestamp 1649977179
transform 1 0 65228 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_709
timestamp 1649977179
transform 1 0 66332 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_721
timestamp 1649977179
transform 1 0 67436 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_727
timestamp 1649977179
transform 1 0 67988 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_729
timestamp 1649977179
transform 1 0 68172 0 -1 43520
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_76_3
timestamp 1649977179
transform 1 0 1380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_15
timestamp 1649977179
transform 1 0 2484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 1649977179
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_29
timestamp 1649977179
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_41
timestamp 1649977179
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_53
timestamp 1649977179
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_65
timestamp 1649977179
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_77
timestamp 1649977179
transform 1 0 8188 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_83
timestamp 1649977179
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_85
timestamp 1649977179
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_97
timestamp 1649977179
transform 1 0 10028 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_109
timestamp 1649977179
transform 1 0 11132 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_121
timestamp 1649977179
transform 1 0 12236 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_133
timestamp 1649977179
transform 1 0 13340 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_139
timestamp 1649977179
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_141
timestamp 1649977179
transform 1 0 14076 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_153
timestamp 1649977179
transform 1 0 15180 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_165
timestamp 1649977179
transform 1 0 16284 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_177
timestamp 1649977179
transform 1 0 17388 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_189
timestamp 1649977179
transform 1 0 18492 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_195
timestamp 1649977179
transform 1 0 19044 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_197
timestamp 1649977179
transform 1 0 19228 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_209
timestamp 1649977179
transform 1 0 20332 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_221
timestamp 1649977179
transform 1 0 21436 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_233
timestamp 1649977179
transform 1 0 22540 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_245
timestamp 1649977179
transform 1 0 23644 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_251
timestamp 1649977179
transform 1 0 24196 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_253
timestamp 1649977179
transform 1 0 24380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_265
timestamp 1649977179
transform 1 0 25484 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_277
timestamp 1649977179
transform 1 0 26588 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_289
timestamp 1649977179
transform 1 0 27692 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_301
timestamp 1649977179
transform 1 0 28796 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_307
timestamp 1649977179
transform 1 0 29348 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_309
timestamp 1649977179
transform 1 0 29532 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_321
timestamp 1649977179
transform 1 0 30636 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_333
timestamp 1649977179
transform 1 0 31740 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_345
timestamp 1649977179
transform 1 0 32844 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_357
timestamp 1649977179
transform 1 0 33948 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_363
timestamp 1649977179
transform 1 0 34500 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_365
timestamp 1649977179
transform 1 0 34684 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_377
timestamp 1649977179
transform 1 0 35788 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_389
timestamp 1649977179
transform 1 0 36892 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_401
timestamp 1649977179
transform 1 0 37996 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_413
timestamp 1649977179
transform 1 0 39100 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_419
timestamp 1649977179
transform 1 0 39652 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_421
timestamp 1649977179
transform 1 0 39836 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_433
timestamp 1649977179
transform 1 0 40940 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_445
timestamp 1649977179
transform 1 0 42044 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_457
timestamp 1649977179
transform 1 0 43148 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_469
timestamp 1649977179
transform 1 0 44252 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_475
timestamp 1649977179
transform 1 0 44804 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_477
timestamp 1649977179
transform 1 0 44988 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_489
timestamp 1649977179
transform 1 0 46092 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_501
timestamp 1649977179
transform 1 0 47196 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_513
timestamp 1649977179
transform 1 0 48300 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_525
timestamp 1649977179
transform 1 0 49404 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_531
timestamp 1649977179
transform 1 0 49956 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_533
timestamp 1649977179
transform 1 0 50140 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_545
timestamp 1649977179
transform 1 0 51244 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_557
timestamp 1649977179
transform 1 0 52348 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_569
timestamp 1649977179
transform 1 0 53452 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_581
timestamp 1649977179
transform 1 0 54556 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_587
timestamp 1649977179
transform 1 0 55108 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_589
timestamp 1649977179
transform 1 0 55292 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_601
timestamp 1649977179
transform 1 0 56396 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_613
timestamp 1649977179
transform 1 0 57500 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_625
timestamp 1649977179
transform 1 0 58604 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_637
timestamp 1649977179
transform 1 0 59708 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_643
timestamp 1649977179
transform 1 0 60260 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_645
timestamp 1649977179
transform 1 0 60444 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_657
timestamp 1649977179
transform 1 0 61548 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_669
timestamp 1649977179
transform 1 0 62652 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_681
timestamp 1649977179
transform 1 0 63756 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_693
timestamp 1649977179
transform 1 0 64860 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_699
timestamp 1649977179
transform 1 0 65412 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_701
timestamp 1649977179
transform 1 0 65596 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_713
timestamp 1649977179
transform 1 0 66700 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_725
timestamp 1649977179
transform 1 0 67804 0 1 43520
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_77_3
timestamp 1649977179
transform 1 0 1380 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_15
timestamp 1649977179
transform 1 0 2484 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_27
timestamp 1649977179
transform 1 0 3588 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_39
timestamp 1649977179
transform 1 0 4692 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_51
timestamp 1649977179
transform 1 0 5796 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_55
timestamp 1649977179
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_57
timestamp 1649977179
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_69
timestamp 1649977179
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_81
timestamp 1649977179
transform 1 0 8556 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_93
timestamp 1649977179
transform 1 0 9660 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_105
timestamp 1649977179
transform 1 0 10764 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_111
timestamp 1649977179
transform 1 0 11316 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_113
timestamp 1649977179
transform 1 0 11500 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_125
timestamp 1649977179
transform 1 0 12604 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_137
timestamp 1649977179
transform 1 0 13708 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_149
timestamp 1649977179
transform 1 0 14812 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_161
timestamp 1649977179
transform 1 0 15916 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_167
timestamp 1649977179
transform 1 0 16468 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_169
timestamp 1649977179
transform 1 0 16652 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_181
timestamp 1649977179
transform 1 0 17756 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_193
timestamp 1649977179
transform 1 0 18860 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_205
timestamp 1649977179
transform 1 0 19964 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_217
timestamp 1649977179
transform 1 0 21068 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_223
timestamp 1649977179
transform 1 0 21620 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_225
timestamp 1649977179
transform 1 0 21804 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_237
timestamp 1649977179
transform 1 0 22908 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_249
timestamp 1649977179
transform 1 0 24012 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_261
timestamp 1649977179
transform 1 0 25116 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_273
timestamp 1649977179
transform 1 0 26220 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_279
timestamp 1649977179
transform 1 0 26772 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_281
timestamp 1649977179
transform 1 0 26956 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_293
timestamp 1649977179
transform 1 0 28060 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_305
timestamp 1649977179
transform 1 0 29164 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_317
timestamp 1649977179
transform 1 0 30268 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_329
timestamp 1649977179
transform 1 0 31372 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_335
timestamp 1649977179
transform 1 0 31924 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_337
timestamp 1649977179
transform 1 0 32108 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_349
timestamp 1649977179
transform 1 0 33212 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_361
timestamp 1649977179
transform 1 0 34316 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_373
timestamp 1649977179
transform 1 0 35420 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_385
timestamp 1649977179
transform 1 0 36524 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_391
timestamp 1649977179
transform 1 0 37076 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_393
timestamp 1649977179
transform 1 0 37260 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_405
timestamp 1649977179
transform 1 0 38364 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_417
timestamp 1649977179
transform 1 0 39468 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_429
timestamp 1649977179
transform 1 0 40572 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_441
timestamp 1649977179
transform 1 0 41676 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_447
timestamp 1649977179
transform 1 0 42228 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_449
timestamp 1649977179
transform 1 0 42412 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_461
timestamp 1649977179
transform 1 0 43516 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_473
timestamp 1649977179
transform 1 0 44620 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_485
timestamp 1649977179
transform 1 0 45724 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_497
timestamp 1649977179
transform 1 0 46828 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_503
timestamp 1649977179
transform 1 0 47380 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_505
timestamp 1649977179
transform 1 0 47564 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_517
timestamp 1649977179
transform 1 0 48668 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_529
timestamp 1649977179
transform 1 0 49772 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_541
timestamp 1649977179
transform 1 0 50876 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_553
timestamp 1649977179
transform 1 0 51980 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_559
timestamp 1649977179
transform 1 0 52532 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_561
timestamp 1649977179
transform 1 0 52716 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_573
timestamp 1649977179
transform 1 0 53820 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_585
timestamp 1649977179
transform 1 0 54924 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_597
timestamp 1649977179
transform 1 0 56028 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_609
timestamp 1649977179
transform 1 0 57132 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_615
timestamp 1649977179
transform 1 0 57684 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_617
timestamp 1649977179
transform 1 0 57868 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_629
timestamp 1649977179
transform 1 0 58972 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_641
timestamp 1649977179
transform 1 0 60076 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_653
timestamp 1649977179
transform 1 0 61180 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_665
timestamp 1649977179
transform 1 0 62284 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_671
timestamp 1649977179
transform 1 0 62836 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_673
timestamp 1649977179
transform 1 0 63020 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_685
timestamp 1649977179
transform 1 0 64124 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_697
timestamp 1649977179
transform 1 0 65228 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_709
timestamp 1649977179
transform 1 0 66332 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_721
timestamp 1649977179
transform 1 0 67436 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_727
timestamp 1649977179
transform 1 0 67988 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_729
timestamp 1649977179
transform 1 0 68172 0 -1 44608
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_78_3
timestamp 1649977179
transform 1 0 1380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_15
timestamp 1649977179
transform 1 0 2484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 1649977179
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_29
timestamp 1649977179
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_41
timestamp 1649977179
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_53
timestamp 1649977179
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_65
timestamp 1649977179
transform 1 0 7084 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_77
timestamp 1649977179
transform 1 0 8188 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_83
timestamp 1649977179
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_85
timestamp 1649977179
transform 1 0 8924 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_97
timestamp 1649977179
transform 1 0 10028 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_109
timestamp 1649977179
transform 1 0 11132 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_121
timestamp 1649977179
transform 1 0 12236 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_133
timestamp 1649977179
transform 1 0 13340 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_139
timestamp 1649977179
transform 1 0 13892 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_141
timestamp 1649977179
transform 1 0 14076 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_153
timestamp 1649977179
transform 1 0 15180 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_165
timestamp 1649977179
transform 1 0 16284 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_177
timestamp 1649977179
transform 1 0 17388 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_189
timestamp 1649977179
transform 1 0 18492 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_195
timestamp 1649977179
transform 1 0 19044 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_197
timestamp 1649977179
transform 1 0 19228 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_209
timestamp 1649977179
transform 1 0 20332 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_221
timestamp 1649977179
transform 1 0 21436 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_233
timestamp 1649977179
transform 1 0 22540 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_245
timestamp 1649977179
transform 1 0 23644 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_251
timestamp 1649977179
transform 1 0 24196 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_253
timestamp 1649977179
transform 1 0 24380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_265
timestamp 1649977179
transform 1 0 25484 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_277
timestamp 1649977179
transform 1 0 26588 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_289
timestamp 1649977179
transform 1 0 27692 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_301
timestamp 1649977179
transform 1 0 28796 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_307
timestamp 1649977179
transform 1 0 29348 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_309
timestamp 1649977179
transform 1 0 29532 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_321
timestamp 1649977179
transform 1 0 30636 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_333
timestamp 1649977179
transform 1 0 31740 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_345
timestamp 1649977179
transform 1 0 32844 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_357
timestamp 1649977179
transform 1 0 33948 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_363
timestamp 1649977179
transform 1 0 34500 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_365
timestamp 1649977179
transform 1 0 34684 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_377
timestamp 1649977179
transform 1 0 35788 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_389
timestamp 1649977179
transform 1 0 36892 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_401
timestamp 1649977179
transform 1 0 37996 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_413
timestamp 1649977179
transform 1 0 39100 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_419
timestamp 1649977179
transform 1 0 39652 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_421
timestamp 1649977179
transform 1 0 39836 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_433
timestamp 1649977179
transform 1 0 40940 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_445
timestamp 1649977179
transform 1 0 42044 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_457
timestamp 1649977179
transform 1 0 43148 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_469
timestamp 1649977179
transform 1 0 44252 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_475
timestamp 1649977179
transform 1 0 44804 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_477
timestamp 1649977179
transform 1 0 44988 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_489
timestamp 1649977179
transform 1 0 46092 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_501
timestamp 1649977179
transform 1 0 47196 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_513
timestamp 1649977179
transform 1 0 48300 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_525
timestamp 1649977179
transform 1 0 49404 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_531
timestamp 1649977179
transform 1 0 49956 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_533
timestamp 1649977179
transform 1 0 50140 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_545
timestamp 1649977179
transform 1 0 51244 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_557
timestamp 1649977179
transform 1 0 52348 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_569
timestamp 1649977179
transform 1 0 53452 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_581
timestamp 1649977179
transform 1 0 54556 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_587
timestamp 1649977179
transform 1 0 55108 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_589
timestamp 1649977179
transform 1 0 55292 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_601
timestamp 1649977179
transform 1 0 56396 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_613
timestamp 1649977179
transform 1 0 57500 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_625
timestamp 1649977179
transform 1 0 58604 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_637
timestamp 1649977179
transform 1 0 59708 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_643
timestamp 1649977179
transform 1 0 60260 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_645
timestamp 1649977179
transform 1 0 60444 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_657
timestamp 1649977179
transform 1 0 61548 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_669
timestamp 1649977179
transform 1 0 62652 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_681
timestamp 1649977179
transform 1 0 63756 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_693
timestamp 1649977179
transform 1 0 64860 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_699
timestamp 1649977179
transform 1 0 65412 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_701
timestamp 1649977179
transform 1 0 65596 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_713
timestamp 1649977179
transform 1 0 66700 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_725
timestamp 1649977179
transform 1 0 67804 0 1 44608
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_79_3
timestamp 1649977179
transform 1 0 1380 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_15
timestamp 1649977179
transform 1 0 2484 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_27
timestamp 1649977179
transform 1 0 3588 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_39
timestamp 1649977179
transform 1 0 4692 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_51
timestamp 1649977179
transform 1 0 5796 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_55
timestamp 1649977179
transform 1 0 6164 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_57
timestamp 1649977179
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_69
timestamp 1649977179
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_81
timestamp 1649977179
transform 1 0 8556 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_93
timestamp 1649977179
transform 1 0 9660 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_105
timestamp 1649977179
transform 1 0 10764 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_111
timestamp 1649977179
transform 1 0 11316 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_113
timestamp 1649977179
transform 1 0 11500 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_125
timestamp 1649977179
transform 1 0 12604 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_137
timestamp 1649977179
transform 1 0 13708 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_149
timestamp 1649977179
transform 1 0 14812 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_161
timestamp 1649977179
transform 1 0 15916 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_167
timestamp 1649977179
transform 1 0 16468 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_169
timestamp 1649977179
transform 1 0 16652 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_181
timestamp 1649977179
transform 1 0 17756 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_193
timestamp 1649977179
transform 1 0 18860 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_205
timestamp 1649977179
transform 1 0 19964 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_217
timestamp 1649977179
transform 1 0 21068 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_223
timestamp 1649977179
transform 1 0 21620 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_225
timestamp 1649977179
transform 1 0 21804 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_237
timestamp 1649977179
transform 1 0 22908 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_249
timestamp 1649977179
transform 1 0 24012 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_261
timestamp 1649977179
transform 1 0 25116 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_273
timestamp 1649977179
transform 1 0 26220 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_279
timestamp 1649977179
transform 1 0 26772 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_281
timestamp 1649977179
transform 1 0 26956 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_293
timestamp 1649977179
transform 1 0 28060 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_305
timestamp 1649977179
transform 1 0 29164 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_317
timestamp 1649977179
transform 1 0 30268 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_329
timestamp 1649977179
transform 1 0 31372 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_335
timestamp 1649977179
transform 1 0 31924 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_337
timestamp 1649977179
transform 1 0 32108 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_349
timestamp 1649977179
transform 1 0 33212 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_361
timestamp 1649977179
transform 1 0 34316 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_373
timestamp 1649977179
transform 1 0 35420 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_385
timestamp 1649977179
transform 1 0 36524 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_391
timestamp 1649977179
transform 1 0 37076 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_393
timestamp 1649977179
transform 1 0 37260 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_405
timestamp 1649977179
transform 1 0 38364 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_417
timestamp 1649977179
transform 1 0 39468 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_429
timestamp 1649977179
transform 1 0 40572 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_441
timestamp 1649977179
transform 1 0 41676 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_447
timestamp 1649977179
transform 1 0 42228 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_449
timestamp 1649977179
transform 1 0 42412 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_461
timestamp 1649977179
transform 1 0 43516 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_473
timestamp 1649977179
transform 1 0 44620 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_485
timestamp 1649977179
transform 1 0 45724 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_497
timestamp 1649977179
transform 1 0 46828 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_503
timestamp 1649977179
transform 1 0 47380 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_505
timestamp 1649977179
transform 1 0 47564 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_517
timestamp 1649977179
transform 1 0 48668 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_529
timestamp 1649977179
transform 1 0 49772 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_541
timestamp 1649977179
transform 1 0 50876 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_553
timestamp 1649977179
transform 1 0 51980 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_559
timestamp 1649977179
transform 1 0 52532 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_561
timestamp 1649977179
transform 1 0 52716 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_573
timestamp 1649977179
transform 1 0 53820 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_585
timestamp 1649977179
transform 1 0 54924 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_597
timestamp 1649977179
transform 1 0 56028 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_609
timestamp 1649977179
transform 1 0 57132 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_615
timestamp 1649977179
transform 1 0 57684 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_617
timestamp 1649977179
transform 1 0 57868 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_629
timestamp 1649977179
transform 1 0 58972 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_641
timestamp 1649977179
transform 1 0 60076 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_653
timestamp 1649977179
transform 1 0 61180 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_665
timestamp 1649977179
transform 1 0 62284 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_671
timestamp 1649977179
transform 1 0 62836 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_673
timestamp 1649977179
transform 1 0 63020 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_685
timestamp 1649977179
transform 1 0 64124 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_697
timestamp 1649977179
transform 1 0 65228 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_709
timestamp 1649977179
transform 1 0 66332 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_721
timestamp 1649977179
transform 1 0 67436 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_727
timestamp 1649977179
transform 1 0 67988 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_729
timestamp 1649977179
transform 1 0 68172 0 -1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_80_3
timestamp 1649977179
transform 1 0 1380 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_15
timestamp 1649977179
transform 1 0 2484 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 1649977179
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_29
timestamp 1649977179
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_41
timestamp 1649977179
transform 1 0 4876 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_53
timestamp 1649977179
transform 1 0 5980 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_65
timestamp 1649977179
transform 1 0 7084 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_77
timestamp 1649977179
transform 1 0 8188 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_83
timestamp 1649977179
transform 1 0 8740 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_85
timestamp 1649977179
transform 1 0 8924 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_97
timestamp 1649977179
transform 1 0 10028 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_109
timestamp 1649977179
transform 1 0 11132 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_121
timestamp 1649977179
transform 1 0 12236 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_133
timestamp 1649977179
transform 1 0 13340 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_139
timestamp 1649977179
transform 1 0 13892 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_141
timestamp 1649977179
transform 1 0 14076 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_153
timestamp 1649977179
transform 1 0 15180 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_165
timestamp 1649977179
transform 1 0 16284 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_177
timestamp 1649977179
transform 1 0 17388 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_189
timestamp 1649977179
transform 1 0 18492 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_195
timestamp 1649977179
transform 1 0 19044 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_197
timestamp 1649977179
transform 1 0 19228 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_209
timestamp 1649977179
transform 1 0 20332 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_221
timestamp 1649977179
transform 1 0 21436 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_233
timestamp 1649977179
transform 1 0 22540 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_245
timestamp 1649977179
transform 1 0 23644 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_251
timestamp 1649977179
transform 1 0 24196 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_253
timestamp 1649977179
transform 1 0 24380 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_265
timestamp 1649977179
transform 1 0 25484 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_277
timestamp 1649977179
transform 1 0 26588 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_289
timestamp 1649977179
transform 1 0 27692 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_301
timestamp 1649977179
transform 1 0 28796 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_307
timestamp 1649977179
transform 1 0 29348 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_309
timestamp 1649977179
transform 1 0 29532 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_321
timestamp 1649977179
transform 1 0 30636 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_333
timestamp 1649977179
transform 1 0 31740 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_345
timestamp 1649977179
transform 1 0 32844 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_357
timestamp 1649977179
transform 1 0 33948 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_363
timestamp 1649977179
transform 1 0 34500 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_365
timestamp 1649977179
transform 1 0 34684 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_377
timestamp 1649977179
transform 1 0 35788 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_389
timestamp 1649977179
transform 1 0 36892 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_401
timestamp 1649977179
transform 1 0 37996 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_413
timestamp 1649977179
transform 1 0 39100 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_419
timestamp 1649977179
transform 1 0 39652 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_421
timestamp 1649977179
transform 1 0 39836 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_433
timestamp 1649977179
transform 1 0 40940 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_445
timestamp 1649977179
transform 1 0 42044 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_457
timestamp 1649977179
transform 1 0 43148 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_469
timestamp 1649977179
transform 1 0 44252 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_475
timestamp 1649977179
transform 1 0 44804 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_477
timestamp 1649977179
transform 1 0 44988 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_489
timestamp 1649977179
transform 1 0 46092 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_501
timestamp 1649977179
transform 1 0 47196 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_513
timestamp 1649977179
transform 1 0 48300 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_525
timestamp 1649977179
transform 1 0 49404 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_531
timestamp 1649977179
transform 1 0 49956 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_533
timestamp 1649977179
transform 1 0 50140 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_545
timestamp 1649977179
transform 1 0 51244 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_557
timestamp 1649977179
transform 1 0 52348 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_569
timestamp 1649977179
transform 1 0 53452 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_581
timestamp 1649977179
transform 1 0 54556 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_587
timestamp 1649977179
transform 1 0 55108 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_589
timestamp 1649977179
transform 1 0 55292 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_601
timestamp 1649977179
transform 1 0 56396 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_613
timestamp 1649977179
transform 1 0 57500 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_625
timestamp 1649977179
transform 1 0 58604 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_637
timestamp 1649977179
transform 1 0 59708 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_643
timestamp 1649977179
transform 1 0 60260 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_645
timestamp 1649977179
transform 1 0 60444 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_657
timestamp 1649977179
transform 1 0 61548 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_669
timestamp 1649977179
transform 1 0 62652 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_681
timestamp 1649977179
transform 1 0 63756 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_693
timestamp 1649977179
transform 1 0 64860 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_699
timestamp 1649977179
transform 1 0 65412 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_701
timestamp 1649977179
transform 1 0 65596 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_713
timestamp 1649977179
transform 1 0 66700 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_725
timestamp 1649977179
transform 1 0 67804 0 1 45696
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_81_3
timestamp 1649977179
transform 1 0 1380 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_15
timestamp 1649977179
transform 1 0 2484 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_27
timestamp 1649977179
transform 1 0 3588 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_39
timestamp 1649977179
transform 1 0 4692 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_51
timestamp 1649977179
transform 1 0 5796 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_55
timestamp 1649977179
transform 1 0 6164 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_57
timestamp 1649977179
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_69
timestamp 1649977179
transform 1 0 7452 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_81
timestamp 1649977179
transform 1 0 8556 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_93
timestamp 1649977179
transform 1 0 9660 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_105
timestamp 1649977179
transform 1 0 10764 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_111
timestamp 1649977179
transform 1 0 11316 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_113
timestamp 1649977179
transform 1 0 11500 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_125
timestamp 1649977179
transform 1 0 12604 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_137
timestamp 1649977179
transform 1 0 13708 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_149
timestamp 1649977179
transform 1 0 14812 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_161
timestamp 1649977179
transform 1 0 15916 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_167
timestamp 1649977179
transform 1 0 16468 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_169
timestamp 1649977179
transform 1 0 16652 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_181
timestamp 1649977179
transform 1 0 17756 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_193
timestamp 1649977179
transform 1 0 18860 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_205
timestamp 1649977179
transform 1 0 19964 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_217
timestamp 1649977179
transform 1 0 21068 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_223
timestamp 1649977179
transform 1 0 21620 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_225
timestamp 1649977179
transform 1 0 21804 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_237
timestamp 1649977179
transform 1 0 22908 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_249
timestamp 1649977179
transform 1 0 24012 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_261
timestamp 1649977179
transform 1 0 25116 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_273
timestamp 1649977179
transform 1 0 26220 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_279
timestamp 1649977179
transform 1 0 26772 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_281
timestamp 1649977179
transform 1 0 26956 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_293
timestamp 1649977179
transform 1 0 28060 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_305
timestamp 1649977179
transform 1 0 29164 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_317
timestamp 1649977179
transform 1 0 30268 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_329
timestamp 1649977179
transform 1 0 31372 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_335
timestamp 1649977179
transform 1 0 31924 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_337
timestamp 1649977179
transform 1 0 32108 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_349
timestamp 1649977179
transform 1 0 33212 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_361
timestamp 1649977179
transform 1 0 34316 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_373
timestamp 1649977179
transform 1 0 35420 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_385
timestamp 1649977179
transform 1 0 36524 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_391
timestamp 1649977179
transform 1 0 37076 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_393
timestamp 1649977179
transform 1 0 37260 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_405
timestamp 1649977179
transform 1 0 38364 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_417
timestamp 1649977179
transform 1 0 39468 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_429
timestamp 1649977179
transform 1 0 40572 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_441
timestamp 1649977179
transform 1 0 41676 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_447
timestamp 1649977179
transform 1 0 42228 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_449
timestamp 1649977179
transform 1 0 42412 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_461
timestamp 1649977179
transform 1 0 43516 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_473
timestamp 1649977179
transform 1 0 44620 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_485
timestamp 1649977179
transform 1 0 45724 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_497
timestamp 1649977179
transform 1 0 46828 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_503
timestamp 1649977179
transform 1 0 47380 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_505
timestamp 1649977179
transform 1 0 47564 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_517
timestamp 1649977179
transform 1 0 48668 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_529
timestamp 1649977179
transform 1 0 49772 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_541
timestamp 1649977179
transform 1 0 50876 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_553
timestamp 1649977179
transform 1 0 51980 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_559
timestamp 1649977179
transform 1 0 52532 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_561
timestamp 1649977179
transform 1 0 52716 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_573
timestamp 1649977179
transform 1 0 53820 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_585
timestamp 1649977179
transform 1 0 54924 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_597
timestamp 1649977179
transform 1 0 56028 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_609
timestamp 1649977179
transform 1 0 57132 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_615
timestamp 1649977179
transform 1 0 57684 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_617
timestamp 1649977179
transform 1 0 57868 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_629
timestamp 1649977179
transform 1 0 58972 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_641
timestamp 1649977179
transform 1 0 60076 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_653
timestamp 1649977179
transform 1 0 61180 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_665
timestamp 1649977179
transform 1 0 62284 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_671
timestamp 1649977179
transform 1 0 62836 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_673
timestamp 1649977179
transform 1 0 63020 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_685
timestamp 1649977179
transform 1 0 64124 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_697
timestamp 1649977179
transform 1 0 65228 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_709
timestamp 1649977179
transform 1 0 66332 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_721
timestamp 1649977179
transform 1 0 67436 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_727
timestamp 1649977179
transform 1 0 67988 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_729
timestamp 1649977179
transform 1 0 68172 0 -1 46784
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_82_3
timestamp 1649977179
transform 1 0 1380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_15
timestamp 1649977179
transform 1 0 2484 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 1649977179
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_29
timestamp 1649977179
transform 1 0 3772 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_41
timestamp 1649977179
transform 1 0 4876 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_53
timestamp 1649977179
transform 1 0 5980 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_65
timestamp 1649977179
transform 1 0 7084 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_77
timestamp 1649977179
transform 1 0 8188 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_83
timestamp 1649977179
transform 1 0 8740 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_85
timestamp 1649977179
transform 1 0 8924 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_97
timestamp 1649977179
transform 1 0 10028 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_109
timestamp 1649977179
transform 1 0 11132 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_121
timestamp 1649977179
transform 1 0 12236 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_133
timestamp 1649977179
transform 1 0 13340 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_139
timestamp 1649977179
transform 1 0 13892 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_141
timestamp 1649977179
transform 1 0 14076 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_153
timestamp 1649977179
transform 1 0 15180 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_165
timestamp 1649977179
transform 1 0 16284 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_177
timestamp 1649977179
transform 1 0 17388 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_189
timestamp 1649977179
transform 1 0 18492 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_195
timestamp 1649977179
transform 1 0 19044 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_197
timestamp 1649977179
transform 1 0 19228 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_209
timestamp 1649977179
transform 1 0 20332 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_221
timestamp 1649977179
transform 1 0 21436 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_233
timestamp 1649977179
transform 1 0 22540 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_245
timestamp 1649977179
transform 1 0 23644 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_251
timestamp 1649977179
transform 1 0 24196 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_253
timestamp 1649977179
transform 1 0 24380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_265
timestamp 1649977179
transform 1 0 25484 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_277
timestamp 1649977179
transform 1 0 26588 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_289
timestamp 1649977179
transform 1 0 27692 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_301
timestamp 1649977179
transform 1 0 28796 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_307
timestamp 1649977179
transform 1 0 29348 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_309
timestamp 1649977179
transform 1 0 29532 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_321
timestamp 1649977179
transform 1 0 30636 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_333
timestamp 1649977179
transform 1 0 31740 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_345
timestamp 1649977179
transform 1 0 32844 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_357
timestamp 1649977179
transform 1 0 33948 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_363
timestamp 1649977179
transform 1 0 34500 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_365
timestamp 1649977179
transform 1 0 34684 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_377
timestamp 1649977179
transform 1 0 35788 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_389
timestamp 1649977179
transform 1 0 36892 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_401
timestamp 1649977179
transform 1 0 37996 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_413
timestamp 1649977179
transform 1 0 39100 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_419
timestamp 1649977179
transform 1 0 39652 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_421
timestamp 1649977179
transform 1 0 39836 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_433
timestamp 1649977179
transform 1 0 40940 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_445
timestamp 1649977179
transform 1 0 42044 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_457
timestamp 1649977179
transform 1 0 43148 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_469
timestamp 1649977179
transform 1 0 44252 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_475
timestamp 1649977179
transform 1 0 44804 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_477
timestamp 1649977179
transform 1 0 44988 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_489
timestamp 1649977179
transform 1 0 46092 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_501
timestamp 1649977179
transform 1 0 47196 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_513
timestamp 1649977179
transform 1 0 48300 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_525
timestamp 1649977179
transform 1 0 49404 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_531
timestamp 1649977179
transform 1 0 49956 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_533
timestamp 1649977179
transform 1 0 50140 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_545
timestamp 1649977179
transform 1 0 51244 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_557
timestamp 1649977179
transform 1 0 52348 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_569
timestamp 1649977179
transform 1 0 53452 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_581
timestamp 1649977179
transform 1 0 54556 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_587
timestamp 1649977179
transform 1 0 55108 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_589
timestamp 1649977179
transform 1 0 55292 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_601
timestamp 1649977179
transform 1 0 56396 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_613
timestamp 1649977179
transform 1 0 57500 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_625
timestamp 1649977179
transform 1 0 58604 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_637
timestamp 1649977179
transform 1 0 59708 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_643
timestamp 1649977179
transform 1 0 60260 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_645
timestamp 1649977179
transform 1 0 60444 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_657
timestamp 1649977179
transform 1 0 61548 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_669
timestamp 1649977179
transform 1 0 62652 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_681
timestamp 1649977179
transform 1 0 63756 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_693
timestamp 1649977179
transform 1 0 64860 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_699
timestamp 1649977179
transform 1 0 65412 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_701
timestamp 1649977179
transform 1 0 65596 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_713
timestamp 1649977179
transform 1 0 66700 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_725
timestamp 1649977179
transform 1 0 67804 0 1 46784
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_83_3
timestamp 1649977179
transform 1 0 1380 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_15
timestamp 1649977179
transform 1 0 2484 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_27
timestamp 1649977179
transform 1 0 3588 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_39
timestamp 1649977179
transform 1 0 4692 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_51
timestamp 1649977179
transform 1 0 5796 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_55
timestamp 1649977179
transform 1 0 6164 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_57
timestamp 1649977179
transform 1 0 6348 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_69
timestamp 1649977179
transform 1 0 7452 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_81
timestamp 1649977179
transform 1 0 8556 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_93
timestamp 1649977179
transform 1 0 9660 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_105
timestamp 1649977179
transform 1 0 10764 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_111
timestamp 1649977179
transform 1 0 11316 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_113
timestamp 1649977179
transform 1 0 11500 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_125
timestamp 1649977179
transform 1 0 12604 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_137
timestamp 1649977179
transform 1 0 13708 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_149
timestamp 1649977179
transform 1 0 14812 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_161
timestamp 1649977179
transform 1 0 15916 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_167
timestamp 1649977179
transform 1 0 16468 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_169
timestamp 1649977179
transform 1 0 16652 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_181
timestamp 1649977179
transform 1 0 17756 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_193
timestamp 1649977179
transform 1 0 18860 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_205
timestamp 1649977179
transform 1 0 19964 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_217
timestamp 1649977179
transform 1 0 21068 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_223
timestamp 1649977179
transform 1 0 21620 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_225
timestamp 1649977179
transform 1 0 21804 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_237
timestamp 1649977179
transform 1 0 22908 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_249
timestamp 1649977179
transform 1 0 24012 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_261
timestamp 1649977179
transform 1 0 25116 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_273
timestamp 1649977179
transform 1 0 26220 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_279
timestamp 1649977179
transform 1 0 26772 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_281
timestamp 1649977179
transform 1 0 26956 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_293
timestamp 1649977179
transform 1 0 28060 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_305
timestamp 1649977179
transform 1 0 29164 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_317
timestamp 1649977179
transform 1 0 30268 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_329
timestamp 1649977179
transform 1 0 31372 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_335
timestamp 1649977179
transform 1 0 31924 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_337
timestamp 1649977179
transform 1 0 32108 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_349
timestamp 1649977179
transform 1 0 33212 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_361
timestamp 1649977179
transform 1 0 34316 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_373
timestamp 1649977179
transform 1 0 35420 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_385
timestamp 1649977179
transform 1 0 36524 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_391
timestamp 1649977179
transform 1 0 37076 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_393
timestamp 1649977179
transform 1 0 37260 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_405
timestamp 1649977179
transform 1 0 38364 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_417
timestamp 1649977179
transform 1 0 39468 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_429
timestamp 1649977179
transform 1 0 40572 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_441
timestamp 1649977179
transform 1 0 41676 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_447
timestamp 1649977179
transform 1 0 42228 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_449
timestamp 1649977179
transform 1 0 42412 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_461
timestamp 1649977179
transform 1 0 43516 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_473
timestamp 1649977179
transform 1 0 44620 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_485
timestamp 1649977179
transform 1 0 45724 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_497
timestamp 1649977179
transform 1 0 46828 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_503
timestamp 1649977179
transform 1 0 47380 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_505
timestamp 1649977179
transform 1 0 47564 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_517
timestamp 1649977179
transform 1 0 48668 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_529
timestamp 1649977179
transform 1 0 49772 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_541
timestamp 1649977179
transform 1 0 50876 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_553
timestamp 1649977179
transform 1 0 51980 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_559
timestamp 1649977179
transform 1 0 52532 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_561
timestamp 1649977179
transform 1 0 52716 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_573
timestamp 1649977179
transform 1 0 53820 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_585
timestamp 1649977179
transform 1 0 54924 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_597
timestamp 1649977179
transform 1 0 56028 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_609
timestamp 1649977179
transform 1 0 57132 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_615
timestamp 1649977179
transform 1 0 57684 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_617
timestamp 1649977179
transform 1 0 57868 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_629
timestamp 1649977179
transform 1 0 58972 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_641
timestamp 1649977179
transform 1 0 60076 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_653
timestamp 1649977179
transform 1 0 61180 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_665
timestamp 1649977179
transform 1 0 62284 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_671
timestamp 1649977179
transform 1 0 62836 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_673
timestamp 1649977179
transform 1 0 63020 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_685
timestamp 1649977179
transform 1 0 64124 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_697
timestamp 1649977179
transform 1 0 65228 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_709
timestamp 1649977179
transform 1 0 66332 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_721
timestamp 1649977179
transform 1 0 67436 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_727
timestamp 1649977179
transform 1 0 67988 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_83_729
timestamp 1649977179
transform 1 0 68172 0 -1 47872
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_84_3
timestamp 1649977179
transform 1 0 1380 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_15
timestamp 1649977179
transform 1 0 2484 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_84_27
timestamp 1649977179
transform 1 0 3588 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_29
timestamp 1649977179
transform 1 0 3772 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_41
timestamp 1649977179
transform 1 0 4876 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_53
timestamp 1649977179
transform 1 0 5980 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_65
timestamp 1649977179
transform 1 0 7084 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_77
timestamp 1649977179
transform 1 0 8188 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_83
timestamp 1649977179
transform 1 0 8740 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_85
timestamp 1649977179
transform 1 0 8924 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_97
timestamp 1649977179
transform 1 0 10028 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_109
timestamp 1649977179
transform 1 0 11132 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_121
timestamp 1649977179
transform 1 0 12236 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_133
timestamp 1649977179
transform 1 0 13340 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_139
timestamp 1649977179
transform 1 0 13892 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_141
timestamp 1649977179
transform 1 0 14076 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_153
timestamp 1649977179
transform 1 0 15180 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_165
timestamp 1649977179
transform 1 0 16284 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_177
timestamp 1649977179
transform 1 0 17388 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_189
timestamp 1649977179
transform 1 0 18492 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_195
timestamp 1649977179
transform 1 0 19044 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_197
timestamp 1649977179
transform 1 0 19228 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_209
timestamp 1649977179
transform 1 0 20332 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_221
timestamp 1649977179
transform 1 0 21436 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_233
timestamp 1649977179
transform 1 0 22540 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_245
timestamp 1649977179
transform 1 0 23644 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_251
timestamp 1649977179
transform 1 0 24196 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_253
timestamp 1649977179
transform 1 0 24380 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_265
timestamp 1649977179
transform 1 0 25484 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_277
timestamp 1649977179
transform 1 0 26588 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_289
timestamp 1649977179
transform 1 0 27692 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_301
timestamp 1649977179
transform 1 0 28796 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_307
timestamp 1649977179
transform 1 0 29348 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_309
timestamp 1649977179
transform 1 0 29532 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_321
timestamp 1649977179
transform 1 0 30636 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_333
timestamp 1649977179
transform 1 0 31740 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_345
timestamp 1649977179
transform 1 0 32844 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_357
timestamp 1649977179
transform 1 0 33948 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_363
timestamp 1649977179
transform 1 0 34500 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_365
timestamp 1649977179
transform 1 0 34684 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_377
timestamp 1649977179
transform 1 0 35788 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_389
timestamp 1649977179
transform 1 0 36892 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_401
timestamp 1649977179
transform 1 0 37996 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_413
timestamp 1649977179
transform 1 0 39100 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_419
timestamp 1649977179
transform 1 0 39652 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_421
timestamp 1649977179
transform 1 0 39836 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_433
timestamp 1649977179
transform 1 0 40940 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_445
timestamp 1649977179
transform 1 0 42044 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_457
timestamp 1649977179
transform 1 0 43148 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_469
timestamp 1649977179
transform 1 0 44252 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_475
timestamp 1649977179
transform 1 0 44804 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_477
timestamp 1649977179
transform 1 0 44988 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_489
timestamp 1649977179
transform 1 0 46092 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_501
timestamp 1649977179
transform 1 0 47196 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_513
timestamp 1649977179
transform 1 0 48300 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_525
timestamp 1649977179
transform 1 0 49404 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_531
timestamp 1649977179
transform 1 0 49956 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_533
timestamp 1649977179
transform 1 0 50140 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_545
timestamp 1649977179
transform 1 0 51244 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_557
timestamp 1649977179
transform 1 0 52348 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_569
timestamp 1649977179
transform 1 0 53452 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_581
timestamp 1649977179
transform 1 0 54556 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_587
timestamp 1649977179
transform 1 0 55108 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_589
timestamp 1649977179
transform 1 0 55292 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_601
timestamp 1649977179
transform 1 0 56396 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_613
timestamp 1649977179
transform 1 0 57500 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_625
timestamp 1649977179
transform 1 0 58604 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_637
timestamp 1649977179
transform 1 0 59708 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_643
timestamp 1649977179
transform 1 0 60260 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_645
timestamp 1649977179
transform 1 0 60444 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_657
timestamp 1649977179
transform 1 0 61548 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_669
timestamp 1649977179
transform 1 0 62652 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_681
timestamp 1649977179
transform 1 0 63756 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_693
timestamp 1649977179
transform 1 0 64860 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_699
timestamp 1649977179
transform 1 0 65412 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_701
timestamp 1649977179
transform 1 0 65596 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_713
timestamp 1649977179
transform 1 0 66700 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_84_725
timestamp 1649977179
transform 1 0 67804 0 1 47872
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_85_3
timestamp 1649977179
transform 1 0 1380 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_15
timestamp 1649977179
transform 1 0 2484 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_27
timestamp 1649977179
transform 1 0 3588 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_39
timestamp 1649977179
transform 1 0 4692 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_51
timestamp 1649977179
transform 1 0 5796 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_55
timestamp 1649977179
transform 1 0 6164 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_57
timestamp 1649977179
transform 1 0 6348 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_69
timestamp 1649977179
transform 1 0 7452 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_81
timestamp 1649977179
transform 1 0 8556 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_93
timestamp 1649977179
transform 1 0 9660 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_105
timestamp 1649977179
transform 1 0 10764 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_111
timestamp 1649977179
transform 1 0 11316 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_113
timestamp 1649977179
transform 1 0 11500 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_125
timestamp 1649977179
transform 1 0 12604 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_137
timestamp 1649977179
transform 1 0 13708 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_149
timestamp 1649977179
transform 1 0 14812 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_161
timestamp 1649977179
transform 1 0 15916 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_167
timestamp 1649977179
transform 1 0 16468 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_169
timestamp 1649977179
transform 1 0 16652 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_181
timestamp 1649977179
transform 1 0 17756 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_193
timestamp 1649977179
transform 1 0 18860 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_205
timestamp 1649977179
transform 1 0 19964 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_217
timestamp 1649977179
transform 1 0 21068 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_223
timestamp 1649977179
transform 1 0 21620 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_225
timestamp 1649977179
transform 1 0 21804 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_237
timestamp 1649977179
transform 1 0 22908 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_249
timestamp 1649977179
transform 1 0 24012 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_261
timestamp 1649977179
transform 1 0 25116 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_273
timestamp 1649977179
transform 1 0 26220 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_279
timestamp 1649977179
transform 1 0 26772 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_281
timestamp 1649977179
transform 1 0 26956 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_293
timestamp 1649977179
transform 1 0 28060 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_305
timestamp 1649977179
transform 1 0 29164 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_317
timestamp 1649977179
transform 1 0 30268 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_329
timestamp 1649977179
transform 1 0 31372 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_335
timestamp 1649977179
transform 1 0 31924 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_337
timestamp 1649977179
transform 1 0 32108 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_349
timestamp 1649977179
transform 1 0 33212 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_361
timestamp 1649977179
transform 1 0 34316 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_373
timestamp 1649977179
transform 1 0 35420 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_385
timestamp 1649977179
transform 1 0 36524 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_391
timestamp 1649977179
transform 1 0 37076 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_393
timestamp 1649977179
transform 1 0 37260 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_405
timestamp 1649977179
transform 1 0 38364 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_417
timestamp 1649977179
transform 1 0 39468 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_429
timestamp 1649977179
transform 1 0 40572 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_441
timestamp 1649977179
transform 1 0 41676 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_447
timestamp 1649977179
transform 1 0 42228 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_449
timestamp 1649977179
transform 1 0 42412 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_461
timestamp 1649977179
transform 1 0 43516 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_473
timestamp 1649977179
transform 1 0 44620 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_485
timestamp 1649977179
transform 1 0 45724 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_497
timestamp 1649977179
transform 1 0 46828 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_503
timestamp 1649977179
transform 1 0 47380 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_505
timestamp 1649977179
transform 1 0 47564 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_517
timestamp 1649977179
transform 1 0 48668 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_529
timestamp 1649977179
transform 1 0 49772 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_541
timestamp 1649977179
transform 1 0 50876 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_553
timestamp 1649977179
transform 1 0 51980 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_559
timestamp 1649977179
transform 1 0 52532 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_561
timestamp 1649977179
transform 1 0 52716 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_573
timestamp 1649977179
transform 1 0 53820 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_585
timestamp 1649977179
transform 1 0 54924 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_597
timestamp 1649977179
transform 1 0 56028 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_609
timestamp 1649977179
transform 1 0 57132 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_615
timestamp 1649977179
transform 1 0 57684 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_617
timestamp 1649977179
transform 1 0 57868 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_629
timestamp 1649977179
transform 1 0 58972 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_641
timestamp 1649977179
transform 1 0 60076 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_653
timestamp 1649977179
transform 1 0 61180 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_665
timestamp 1649977179
transform 1 0 62284 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_671
timestamp 1649977179
transform 1 0 62836 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_673
timestamp 1649977179
transform 1 0 63020 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_685
timestamp 1649977179
transform 1 0 64124 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_697
timestamp 1649977179
transform 1 0 65228 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_709
timestamp 1649977179
transform 1 0 66332 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_721
timestamp 1649977179
transform 1 0 67436 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_727
timestamp 1649977179
transform 1 0 67988 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_729
timestamp 1649977179
transform 1 0 68172 0 -1 48960
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_86_3
timestamp 1649977179
transform 1 0 1380 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_15
timestamp 1649977179
transform 1 0 2484 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_86_27
timestamp 1649977179
transform 1 0 3588 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_29
timestamp 1649977179
transform 1 0 3772 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_41
timestamp 1649977179
transform 1 0 4876 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_53
timestamp 1649977179
transform 1 0 5980 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_65
timestamp 1649977179
transform 1 0 7084 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_77
timestamp 1649977179
transform 1 0 8188 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_83
timestamp 1649977179
transform 1 0 8740 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_85
timestamp 1649977179
transform 1 0 8924 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_97
timestamp 1649977179
transform 1 0 10028 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_109
timestamp 1649977179
transform 1 0 11132 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_121
timestamp 1649977179
transform 1 0 12236 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_133
timestamp 1649977179
transform 1 0 13340 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_139
timestamp 1649977179
transform 1 0 13892 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_141
timestamp 1649977179
transform 1 0 14076 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_153
timestamp 1649977179
transform 1 0 15180 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_165
timestamp 1649977179
transform 1 0 16284 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_177
timestamp 1649977179
transform 1 0 17388 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_189
timestamp 1649977179
transform 1 0 18492 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_195
timestamp 1649977179
transform 1 0 19044 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_197
timestamp 1649977179
transform 1 0 19228 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_209
timestamp 1649977179
transform 1 0 20332 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_221
timestamp 1649977179
transform 1 0 21436 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_233
timestamp 1649977179
transform 1 0 22540 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_245
timestamp 1649977179
transform 1 0 23644 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_251
timestamp 1649977179
transform 1 0 24196 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_253
timestamp 1649977179
transform 1 0 24380 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_265
timestamp 1649977179
transform 1 0 25484 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_277
timestamp 1649977179
transform 1 0 26588 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_289
timestamp 1649977179
transform 1 0 27692 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_301
timestamp 1649977179
transform 1 0 28796 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_307
timestamp 1649977179
transform 1 0 29348 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_309
timestamp 1649977179
transform 1 0 29532 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_321
timestamp 1649977179
transform 1 0 30636 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_333
timestamp 1649977179
transform 1 0 31740 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_345
timestamp 1649977179
transform 1 0 32844 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_357
timestamp 1649977179
transform 1 0 33948 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_363
timestamp 1649977179
transform 1 0 34500 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_365
timestamp 1649977179
transform 1 0 34684 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_377
timestamp 1649977179
transform 1 0 35788 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_389
timestamp 1649977179
transform 1 0 36892 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_401
timestamp 1649977179
transform 1 0 37996 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_413
timestamp 1649977179
transform 1 0 39100 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_419
timestamp 1649977179
transform 1 0 39652 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_421
timestamp 1649977179
transform 1 0 39836 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_433
timestamp 1649977179
transform 1 0 40940 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_445
timestamp 1649977179
transform 1 0 42044 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_457
timestamp 1649977179
transform 1 0 43148 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_469
timestamp 1649977179
transform 1 0 44252 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_475
timestamp 1649977179
transform 1 0 44804 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_477
timestamp 1649977179
transform 1 0 44988 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_489
timestamp 1649977179
transform 1 0 46092 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_501
timestamp 1649977179
transform 1 0 47196 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_513
timestamp 1649977179
transform 1 0 48300 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_525
timestamp 1649977179
transform 1 0 49404 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_531
timestamp 1649977179
transform 1 0 49956 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_533
timestamp 1649977179
transform 1 0 50140 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_545
timestamp 1649977179
transform 1 0 51244 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_557
timestamp 1649977179
transform 1 0 52348 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_569
timestamp 1649977179
transform 1 0 53452 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_581
timestamp 1649977179
transform 1 0 54556 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_587
timestamp 1649977179
transform 1 0 55108 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_589
timestamp 1649977179
transform 1 0 55292 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_601
timestamp 1649977179
transform 1 0 56396 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_613
timestamp 1649977179
transform 1 0 57500 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_625
timestamp 1649977179
transform 1 0 58604 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_637
timestamp 1649977179
transform 1 0 59708 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_643
timestamp 1649977179
transform 1 0 60260 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_645
timestamp 1649977179
transform 1 0 60444 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_657
timestamp 1649977179
transform 1 0 61548 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_669
timestamp 1649977179
transform 1 0 62652 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_681
timestamp 1649977179
transform 1 0 63756 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_693
timestamp 1649977179
transform 1 0 64860 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_699
timestamp 1649977179
transform 1 0 65412 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_701
timestamp 1649977179
transform 1 0 65596 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_713
timestamp 1649977179
transform 1 0 66700 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_725
timestamp 1649977179
transform 1 0 67804 0 1 48960
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_87_3
timestamp 1649977179
transform 1 0 1380 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_15
timestamp 1649977179
transform 1 0 2484 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_27
timestamp 1649977179
transform 1 0 3588 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_39
timestamp 1649977179
transform 1 0 4692 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_51
timestamp 1649977179
transform 1 0 5796 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_55
timestamp 1649977179
transform 1 0 6164 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_57
timestamp 1649977179
transform 1 0 6348 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_69
timestamp 1649977179
transform 1 0 7452 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_81
timestamp 1649977179
transform 1 0 8556 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_93
timestamp 1649977179
transform 1 0 9660 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_105
timestamp 1649977179
transform 1 0 10764 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_111
timestamp 1649977179
transform 1 0 11316 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_113
timestamp 1649977179
transform 1 0 11500 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_125
timestamp 1649977179
transform 1 0 12604 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_137
timestamp 1649977179
transform 1 0 13708 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_149
timestamp 1649977179
transform 1 0 14812 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_161
timestamp 1649977179
transform 1 0 15916 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_167
timestamp 1649977179
transform 1 0 16468 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_169
timestamp 1649977179
transform 1 0 16652 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_181
timestamp 1649977179
transform 1 0 17756 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_193
timestamp 1649977179
transform 1 0 18860 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_205
timestamp 1649977179
transform 1 0 19964 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_217
timestamp 1649977179
transform 1 0 21068 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_223
timestamp 1649977179
transform 1 0 21620 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_225
timestamp 1649977179
transform 1 0 21804 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_237
timestamp 1649977179
transform 1 0 22908 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_249
timestamp 1649977179
transform 1 0 24012 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_261
timestamp 1649977179
transform 1 0 25116 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_273
timestamp 1649977179
transform 1 0 26220 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_279
timestamp 1649977179
transform 1 0 26772 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_281
timestamp 1649977179
transform 1 0 26956 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_293
timestamp 1649977179
transform 1 0 28060 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_305
timestamp 1649977179
transform 1 0 29164 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_317
timestamp 1649977179
transform 1 0 30268 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_329
timestamp 1649977179
transform 1 0 31372 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_335
timestamp 1649977179
transform 1 0 31924 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_337
timestamp 1649977179
transform 1 0 32108 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_349
timestamp 1649977179
transform 1 0 33212 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_361
timestamp 1649977179
transform 1 0 34316 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_373
timestamp 1649977179
transform 1 0 35420 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_385
timestamp 1649977179
transform 1 0 36524 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_391
timestamp 1649977179
transform 1 0 37076 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_393
timestamp 1649977179
transform 1 0 37260 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_405
timestamp 1649977179
transform 1 0 38364 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_417
timestamp 1649977179
transform 1 0 39468 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_429
timestamp 1649977179
transform 1 0 40572 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_441
timestamp 1649977179
transform 1 0 41676 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_447
timestamp 1649977179
transform 1 0 42228 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_449
timestamp 1649977179
transform 1 0 42412 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_461
timestamp 1649977179
transform 1 0 43516 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_473
timestamp 1649977179
transform 1 0 44620 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_485
timestamp 1649977179
transform 1 0 45724 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_497
timestamp 1649977179
transform 1 0 46828 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_503
timestamp 1649977179
transform 1 0 47380 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_505
timestamp 1649977179
transform 1 0 47564 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_517
timestamp 1649977179
transform 1 0 48668 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_529
timestamp 1649977179
transform 1 0 49772 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_541
timestamp 1649977179
transform 1 0 50876 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_553
timestamp 1649977179
transform 1 0 51980 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_559
timestamp 1649977179
transform 1 0 52532 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_561
timestamp 1649977179
transform 1 0 52716 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_573
timestamp 1649977179
transform 1 0 53820 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_585
timestamp 1649977179
transform 1 0 54924 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_597
timestamp 1649977179
transform 1 0 56028 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_609
timestamp 1649977179
transform 1 0 57132 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_615
timestamp 1649977179
transform 1 0 57684 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_617
timestamp 1649977179
transform 1 0 57868 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_629
timestamp 1649977179
transform 1 0 58972 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_641
timestamp 1649977179
transform 1 0 60076 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_653
timestamp 1649977179
transform 1 0 61180 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_665
timestamp 1649977179
transform 1 0 62284 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_671
timestamp 1649977179
transform 1 0 62836 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_673
timestamp 1649977179
transform 1 0 63020 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_685
timestamp 1649977179
transform 1 0 64124 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_697
timestamp 1649977179
transform 1 0 65228 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_709
timestamp 1649977179
transform 1 0 66332 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_721
timestamp 1649977179
transform 1 0 67436 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_727
timestamp 1649977179
transform 1 0 67988 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_87_729
timestamp 1649977179
transform 1 0 68172 0 -1 50048
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_88_3
timestamp 1649977179
transform 1 0 1380 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_15
timestamp 1649977179
transform 1 0 2484 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_88_27
timestamp 1649977179
transform 1 0 3588 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_29
timestamp 1649977179
transform 1 0 3772 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_41
timestamp 1649977179
transform 1 0 4876 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_53
timestamp 1649977179
transform 1 0 5980 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_65
timestamp 1649977179
transform 1 0 7084 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_77
timestamp 1649977179
transform 1 0 8188 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_83
timestamp 1649977179
transform 1 0 8740 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_85
timestamp 1649977179
transform 1 0 8924 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_97
timestamp 1649977179
transform 1 0 10028 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_109
timestamp 1649977179
transform 1 0 11132 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_121
timestamp 1649977179
transform 1 0 12236 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_133
timestamp 1649977179
transform 1 0 13340 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_139
timestamp 1649977179
transform 1 0 13892 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_141
timestamp 1649977179
transform 1 0 14076 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_153
timestamp 1649977179
transform 1 0 15180 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_165
timestamp 1649977179
transform 1 0 16284 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_177
timestamp 1649977179
transform 1 0 17388 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_189
timestamp 1649977179
transform 1 0 18492 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_195
timestamp 1649977179
transform 1 0 19044 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_197
timestamp 1649977179
transform 1 0 19228 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_209
timestamp 1649977179
transform 1 0 20332 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_221
timestamp 1649977179
transform 1 0 21436 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_233
timestamp 1649977179
transform 1 0 22540 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_245
timestamp 1649977179
transform 1 0 23644 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_251
timestamp 1649977179
transform 1 0 24196 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_253
timestamp 1649977179
transform 1 0 24380 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_265
timestamp 1649977179
transform 1 0 25484 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_277
timestamp 1649977179
transform 1 0 26588 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_289
timestamp 1649977179
transform 1 0 27692 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_301
timestamp 1649977179
transform 1 0 28796 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_307
timestamp 1649977179
transform 1 0 29348 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_309
timestamp 1649977179
transform 1 0 29532 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_321
timestamp 1649977179
transform 1 0 30636 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_333
timestamp 1649977179
transform 1 0 31740 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_345
timestamp 1649977179
transform 1 0 32844 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_357
timestamp 1649977179
transform 1 0 33948 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_363
timestamp 1649977179
transform 1 0 34500 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_365
timestamp 1649977179
transform 1 0 34684 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_377
timestamp 1649977179
transform 1 0 35788 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_389
timestamp 1649977179
transform 1 0 36892 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_401
timestamp 1649977179
transform 1 0 37996 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_413
timestamp 1649977179
transform 1 0 39100 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_419
timestamp 1649977179
transform 1 0 39652 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_421
timestamp 1649977179
transform 1 0 39836 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_433
timestamp 1649977179
transform 1 0 40940 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_445
timestamp 1649977179
transform 1 0 42044 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_457
timestamp 1649977179
transform 1 0 43148 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_469
timestamp 1649977179
transform 1 0 44252 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_475
timestamp 1649977179
transform 1 0 44804 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_477
timestamp 1649977179
transform 1 0 44988 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_489
timestamp 1649977179
transform 1 0 46092 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_501
timestamp 1649977179
transform 1 0 47196 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_513
timestamp 1649977179
transform 1 0 48300 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_525
timestamp 1649977179
transform 1 0 49404 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_531
timestamp 1649977179
transform 1 0 49956 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_533
timestamp 1649977179
transform 1 0 50140 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_545
timestamp 1649977179
transform 1 0 51244 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_557
timestamp 1649977179
transform 1 0 52348 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_569
timestamp 1649977179
transform 1 0 53452 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_581
timestamp 1649977179
transform 1 0 54556 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_587
timestamp 1649977179
transform 1 0 55108 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_589
timestamp 1649977179
transform 1 0 55292 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_601
timestamp 1649977179
transform 1 0 56396 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_613
timestamp 1649977179
transform 1 0 57500 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_625
timestamp 1649977179
transform 1 0 58604 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_637
timestamp 1649977179
transform 1 0 59708 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_643
timestamp 1649977179
transform 1 0 60260 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_645
timestamp 1649977179
transform 1 0 60444 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_657
timestamp 1649977179
transform 1 0 61548 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_669
timestamp 1649977179
transform 1 0 62652 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_681
timestamp 1649977179
transform 1 0 63756 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_693
timestamp 1649977179
transform 1 0 64860 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_699
timestamp 1649977179
transform 1 0 65412 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_701
timestamp 1649977179
transform 1 0 65596 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_713
timestamp 1649977179
transform 1 0 66700 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_88_725
timestamp 1649977179
transform 1 0 67804 0 1 50048
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_89_3
timestamp 1649977179
transform 1 0 1380 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_15
timestamp 1649977179
transform 1 0 2484 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_27
timestamp 1649977179
transform 1 0 3588 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_39
timestamp 1649977179
transform 1 0 4692 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_51
timestamp 1649977179
transform 1 0 5796 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_55
timestamp 1649977179
transform 1 0 6164 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_57
timestamp 1649977179
transform 1 0 6348 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_69
timestamp 1649977179
transform 1 0 7452 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_81
timestamp 1649977179
transform 1 0 8556 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_93
timestamp 1649977179
transform 1 0 9660 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_105
timestamp 1649977179
transform 1 0 10764 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_111
timestamp 1649977179
transform 1 0 11316 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_113
timestamp 1649977179
transform 1 0 11500 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_125
timestamp 1649977179
transform 1 0 12604 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_137
timestamp 1649977179
transform 1 0 13708 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_149
timestamp 1649977179
transform 1 0 14812 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_161
timestamp 1649977179
transform 1 0 15916 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_167
timestamp 1649977179
transform 1 0 16468 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_169
timestamp 1649977179
transform 1 0 16652 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_181
timestamp 1649977179
transform 1 0 17756 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_193
timestamp 1649977179
transform 1 0 18860 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_205
timestamp 1649977179
transform 1 0 19964 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_217
timestamp 1649977179
transform 1 0 21068 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_223
timestamp 1649977179
transform 1 0 21620 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_225
timestamp 1649977179
transform 1 0 21804 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_237
timestamp 1649977179
transform 1 0 22908 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_249
timestamp 1649977179
transform 1 0 24012 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_261
timestamp 1649977179
transform 1 0 25116 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_273
timestamp 1649977179
transform 1 0 26220 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_279
timestamp 1649977179
transform 1 0 26772 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_281
timestamp 1649977179
transform 1 0 26956 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_293
timestamp 1649977179
transform 1 0 28060 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_305
timestamp 1649977179
transform 1 0 29164 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_317
timestamp 1649977179
transform 1 0 30268 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_329
timestamp 1649977179
transform 1 0 31372 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_335
timestamp 1649977179
transform 1 0 31924 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_337
timestamp 1649977179
transform 1 0 32108 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_349
timestamp 1649977179
transform 1 0 33212 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_361
timestamp 1649977179
transform 1 0 34316 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_373
timestamp 1649977179
transform 1 0 35420 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_385
timestamp 1649977179
transform 1 0 36524 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_391
timestamp 1649977179
transform 1 0 37076 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_393
timestamp 1649977179
transform 1 0 37260 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_405
timestamp 1649977179
transform 1 0 38364 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_417
timestamp 1649977179
transform 1 0 39468 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_429
timestamp 1649977179
transform 1 0 40572 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_441
timestamp 1649977179
transform 1 0 41676 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_447
timestamp 1649977179
transform 1 0 42228 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_449
timestamp 1649977179
transform 1 0 42412 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_461
timestamp 1649977179
transform 1 0 43516 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_473
timestamp 1649977179
transform 1 0 44620 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_485
timestamp 1649977179
transform 1 0 45724 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_497
timestamp 1649977179
transform 1 0 46828 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_503
timestamp 1649977179
transform 1 0 47380 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_505
timestamp 1649977179
transform 1 0 47564 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_517
timestamp 1649977179
transform 1 0 48668 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_529
timestamp 1649977179
transform 1 0 49772 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_541
timestamp 1649977179
transform 1 0 50876 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_553
timestamp 1649977179
transform 1 0 51980 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_559
timestamp 1649977179
transform 1 0 52532 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_561
timestamp 1649977179
transform 1 0 52716 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_573
timestamp 1649977179
transform 1 0 53820 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_585
timestamp 1649977179
transform 1 0 54924 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_597
timestamp 1649977179
transform 1 0 56028 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_609
timestamp 1649977179
transform 1 0 57132 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_615
timestamp 1649977179
transform 1 0 57684 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_617
timestamp 1649977179
transform 1 0 57868 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_629
timestamp 1649977179
transform 1 0 58972 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_641
timestamp 1649977179
transform 1 0 60076 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_653
timestamp 1649977179
transform 1 0 61180 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_665
timestamp 1649977179
transform 1 0 62284 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_671
timestamp 1649977179
transform 1 0 62836 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_673
timestamp 1649977179
transform 1 0 63020 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_685
timestamp 1649977179
transform 1 0 64124 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_697
timestamp 1649977179
transform 1 0 65228 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_709
timestamp 1649977179
transform 1 0 66332 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_721
timestamp 1649977179
transform 1 0 67436 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_727
timestamp 1649977179
transform 1 0 67988 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_89_729
timestamp 1649977179
transform 1 0 68172 0 -1 51136
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_90_3
timestamp 1649977179
transform 1 0 1380 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_15
timestamp 1649977179
transform 1 0 2484 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_90_27
timestamp 1649977179
transform 1 0 3588 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_29
timestamp 1649977179
transform 1 0 3772 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_41
timestamp 1649977179
transform 1 0 4876 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_53
timestamp 1649977179
transform 1 0 5980 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_65
timestamp 1649977179
transform 1 0 7084 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_77
timestamp 1649977179
transform 1 0 8188 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_83
timestamp 1649977179
transform 1 0 8740 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_85
timestamp 1649977179
transform 1 0 8924 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_97
timestamp 1649977179
transform 1 0 10028 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_109
timestamp 1649977179
transform 1 0 11132 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_121
timestamp 1649977179
transform 1 0 12236 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_133
timestamp 1649977179
transform 1 0 13340 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_139
timestamp 1649977179
transform 1 0 13892 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_141
timestamp 1649977179
transform 1 0 14076 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_153
timestamp 1649977179
transform 1 0 15180 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_165
timestamp 1649977179
transform 1 0 16284 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_177
timestamp 1649977179
transform 1 0 17388 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_189
timestamp 1649977179
transform 1 0 18492 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_195
timestamp 1649977179
transform 1 0 19044 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_197
timestamp 1649977179
transform 1 0 19228 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_209
timestamp 1649977179
transform 1 0 20332 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_221
timestamp 1649977179
transform 1 0 21436 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_233
timestamp 1649977179
transform 1 0 22540 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_245
timestamp 1649977179
transform 1 0 23644 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_251
timestamp 1649977179
transform 1 0 24196 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_253
timestamp 1649977179
transform 1 0 24380 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_265
timestamp 1649977179
transform 1 0 25484 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_277
timestamp 1649977179
transform 1 0 26588 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_289
timestamp 1649977179
transform 1 0 27692 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_301
timestamp 1649977179
transform 1 0 28796 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_307
timestamp 1649977179
transform 1 0 29348 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_309
timestamp 1649977179
transform 1 0 29532 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_321
timestamp 1649977179
transform 1 0 30636 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_333
timestamp 1649977179
transform 1 0 31740 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_345
timestamp 1649977179
transform 1 0 32844 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_357
timestamp 1649977179
transform 1 0 33948 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_363
timestamp 1649977179
transform 1 0 34500 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_365
timestamp 1649977179
transform 1 0 34684 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_377
timestamp 1649977179
transform 1 0 35788 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_389
timestamp 1649977179
transform 1 0 36892 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_401
timestamp 1649977179
transform 1 0 37996 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_413
timestamp 1649977179
transform 1 0 39100 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_419
timestamp 1649977179
transform 1 0 39652 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_421
timestamp 1649977179
transform 1 0 39836 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_433
timestamp 1649977179
transform 1 0 40940 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_445
timestamp 1649977179
transform 1 0 42044 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_457
timestamp 1649977179
transform 1 0 43148 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_469
timestamp 1649977179
transform 1 0 44252 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_475
timestamp 1649977179
transform 1 0 44804 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_477
timestamp 1649977179
transform 1 0 44988 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_489
timestamp 1649977179
transform 1 0 46092 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_501
timestamp 1649977179
transform 1 0 47196 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_513
timestamp 1649977179
transform 1 0 48300 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_525
timestamp 1649977179
transform 1 0 49404 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_531
timestamp 1649977179
transform 1 0 49956 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_533
timestamp 1649977179
transform 1 0 50140 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_545
timestamp 1649977179
transform 1 0 51244 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_557
timestamp 1649977179
transform 1 0 52348 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_569
timestamp 1649977179
transform 1 0 53452 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_581
timestamp 1649977179
transform 1 0 54556 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_587
timestamp 1649977179
transform 1 0 55108 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_589
timestamp 1649977179
transform 1 0 55292 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_601
timestamp 1649977179
transform 1 0 56396 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_613
timestamp 1649977179
transform 1 0 57500 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_625
timestamp 1649977179
transform 1 0 58604 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_637
timestamp 1649977179
transform 1 0 59708 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_643
timestamp 1649977179
transform 1 0 60260 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_645
timestamp 1649977179
transform 1 0 60444 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_657
timestamp 1649977179
transform 1 0 61548 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_669
timestamp 1649977179
transform 1 0 62652 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_681
timestamp 1649977179
transform 1 0 63756 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_693
timestamp 1649977179
transform 1 0 64860 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_699
timestamp 1649977179
transform 1 0 65412 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_701
timestamp 1649977179
transform 1 0 65596 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_713
timestamp 1649977179
transform 1 0 66700 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_90_725
timestamp 1649977179
transform 1 0 67804 0 1 51136
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_91_3
timestamp 1649977179
transform 1 0 1380 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_15
timestamp 1649977179
transform 1 0 2484 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_27
timestamp 1649977179
transform 1 0 3588 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_39
timestamp 1649977179
transform 1 0 4692 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_91_51
timestamp 1649977179
transform 1 0 5796 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_91_55
timestamp 1649977179
transform 1 0 6164 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_57
timestamp 1649977179
transform 1 0 6348 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_69
timestamp 1649977179
transform 1 0 7452 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_81
timestamp 1649977179
transform 1 0 8556 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_93
timestamp 1649977179
transform 1 0 9660 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_105
timestamp 1649977179
transform 1 0 10764 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_111
timestamp 1649977179
transform 1 0 11316 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_113
timestamp 1649977179
transform 1 0 11500 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_125
timestamp 1649977179
transform 1 0 12604 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_137
timestamp 1649977179
transform 1 0 13708 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_149
timestamp 1649977179
transform 1 0 14812 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_161
timestamp 1649977179
transform 1 0 15916 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_167
timestamp 1649977179
transform 1 0 16468 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_169
timestamp 1649977179
transform 1 0 16652 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_181
timestamp 1649977179
transform 1 0 17756 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_193
timestamp 1649977179
transform 1 0 18860 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_205
timestamp 1649977179
transform 1 0 19964 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_217
timestamp 1649977179
transform 1 0 21068 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_223
timestamp 1649977179
transform 1 0 21620 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_225
timestamp 1649977179
transform 1 0 21804 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_237
timestamp 1649977179
transform 1 0 22908 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_249
timestamp 1649977179
transform 1 0 24012 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_261
timestamp 1649977179
transform 1 0 25116 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_273
timestamp 1649977179
transform 1 0 26220 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_279
timestamp 1649977179
transform 1 0 26772 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_281
timestamp 1649977179
transform 1 0 26956 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_293
timestamp 1649977179
transform 1 0 28060 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_305
timestamp 1649977179
transform 1 0 29164 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_317
timestamp 1649977179
transform 1 0 30268 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_329
timestamp 1649977179
transform 1 0 31372 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_335
timestamp 1649977179
transform 1 0 31924 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_337
timestamp 1649977179
transform 1 0 32108 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_349
timestamp 1649977179
transform 1 0 33212 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_361
timestamp 1649977179
transform 1 0 34316 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_373
timestamp 1649977179
transform 1 0 35420 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_385
timestamp 1649977179
transform 1 0 36524 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_391
timestamp 1649977179
transform 1 0 37076 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_393
timestamp 1649977179
transform 1 0 37260 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_405
timestamp 1649977179
transform 1 0 38364 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_417
timestamp 1649977179
transform 1 0 39468 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_429
timestamp 1649977179
transform 1 0 40572 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_441
timestamp 1649977179
transform 1 0 41676 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_447
timestamp 1649977179
transform 1 0 42228 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_449
timestamp 1649977179
transform 1 0 42412 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_461
timestamp 1649977179
transform 1 0 43516 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_473
timestamp 1649977179
transform 1 0 44620 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_485
timestamp 1649977179
transform 1 0 45724 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_497
timestamp 1649977179
transform 1 0 46828 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_503
timestamp 1649977179
transform 1 0 47380 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_505
timestamp 1649977179
transform 1 0 47564 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_517
timestamp 1649977179
transform 1 0 48668 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_529
timestamp 1649977179
transform 1 0 49772 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_541
timestamp 1649977179
transform 1 0 50876 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_553
timestamp 1649977179
transform 1 0 51980 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_559
timestamp 1649977179
transform 1 0 52532 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_561
timestamp 1649977179
transform 1 0 52716 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_573
timestamp 1649977179
transform 1 0 53820 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_585
timestamp 1649977179
transform 1 0 54924 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_597
timestamp 1649977179
transform 1 0 56028 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_609
timestamp 1649977179
transform 1 0 57132 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_615
timestamp 1649977179
transform 1 0 57684 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_617
timestamp 1649977179
transform 1 0 57868 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_629
timestamp 1649977179
transform 1 0 58972 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_641
timestamp 1649977179
transform 1 0 60076 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_653
timestamp 1649977179
transform 1 0 61180 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_665
timestamp 1649977179
transform 1 0 62284 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_671
timestamp 1649977179
transform 1 0 62836 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_673
timestamp 1649977179
transform 1 0 63020 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_685
timestamp 1649977179
transform 1 0 64124 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_697
timestamp 1649977179
transform 1 0 65228 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_709
timestamp 1649977179
transform 1 0 66332 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_721
timestamp 1649977179
transform 1 0 67436 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_727
timestamp 1649977179
transform 1 0 67988 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_91_729
timestamp 1649977179
transform 1 0 68172 0 -1 52224
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_92_3
timestamp 1649977179
transform 1 0 1380 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_15
timestamp 1649977179
transform 1 0 2484 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_92_27
timestamp 1649977179
transform 1 0 3588 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_29
timestamp 1649977179
transform 1 0 3772 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_41
timestamp 1649977179
transform 1 0 4876 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_53
timestamp 1649977179
transform 1 0 5980 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_65
timestamp 1649977179
transform 1 0 7084 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_77
timestamp 1649977179
transform 1 0 8188 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_83
timestamp 1649977179
transform 1 0 8740 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_85
timestamp 1649977179
transform 1 0 8924 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_97
timestamp 1649977179
transform 1 0 10028 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_109
timestamp 1649977179
transform 1 0 11132 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_121
timestamp 1649977179
transform 1 0 12236 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_133
timestamp 1649977179
transform 1 0 13340 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_139
timestamp 1649977179
transform 1 0 13892 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_141
timestamp 1649977179
transform 1 0 14076 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_153
timestamp 1649977179
transform 1 0 15180 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_165
timestamp 1649977179
transform 1 0 16284 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_177
timestamp 1649977179
transform 1 0 17388 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_189
timestamp 1649977179
transform 1 0 18492 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_195
timestamp 1649977179
transform 1 0 19044 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_197
timestamp 1649977179
transform 1 0 19228 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_209
timestamp 1649977179
transform 1 0 20332 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_221
timestamp 1649977179
transform 1 0 21436 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_233
timestamp 1649977179
transform 1 0 22540 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_245
timestamp 1649977179
transform 1 0 23644 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_251
timestamp 1649977179
transform 1 0 24196 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_253
timestamp 1649977179
transform 1 0 24380 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_265
timestamp 1649977179
transform 1 0 25484 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_277
timestamp 1649977179
transform 1 0 26588 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_289
timestamp 1649977179
transform 1 0 27692 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_301
timestamp 1649977179
transform 1 0 28796 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_307
timestamp 1649977179
transform 1 0 29348 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_309
timestamp 1649977179
transform 1 0 29532 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_321
timestamp 1649977179
transform 1 0 30636 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_333
timestamp 1649977179
transform 1 0 31740 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_345
timestamp 1649977179
transform 1 0 32844 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_357
timestamp 1649977179
transform 1 0 33948 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_363
timestamp 1649977179
transform 1 0 34500 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_365
timestamp 1649977179
transform 1 0 34684 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_377
timestamp 1649977179
transform 1 0 35788 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_389
timestamp 1649977179
transform 1 0 36892 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_401
timestamp 1649977179
transform 1 0 37996 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_413
timestamp 1649977179
transform 1 0 39100 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_419
timestamp 1649977179
transform 1 0 39652 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_421
timestamp 1649977179
transform 1 0 39836 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_433
timestamp 1649977179
transform 1 0 40940 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_445
timestamp 1649977179
transform 1 0 42044 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_457
timestamp 1649977179
transform 1 0 43148 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_469
timestamp 1649977179
transform 1 0 44252 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_475
timestamp 1649977179
transform 1 0 44804 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_477
timestamp 1649977179
transform 1 0 44988 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_489
timestamp 1649977179
transform 1 0 46092 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_501
timestamp 1649977179
transform 1 0 47196 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_513
timestamp 1649977179
transform 1 0 48300 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_525
timestamp 1649977179
transform 1 0 49404 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_531
timestamp 1649977179
transform 1 0 49956 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_533
timestamp 1649977179
transform 1 0 50140 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_545
timestamp 1649977179
transform 1 0 51244 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_557
timestamp 1649977179
transform 1 0 52348 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_569
timestamp 1649977179
transform 1 0 53452 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_581
timestamp 1649977179
transform 1 0 54556 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_587
timestamp 1649977179
transform 1 0 55108 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_589
timestamp 1649977179
transform 1 0 55292 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_601
timestamp 1649977179
transform 1 0 56396 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_613
timestamp 1649977179
transform 1 0 57500 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_625
timestamp 1649977179
transform 1 0 58604 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_637
timestamp 1649977179
transform 1 0 59708 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_643
timestamp 1649977179
transform 1 0 60260 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_645
timestamp 1649977179
transform 1 0 60444 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_657
timestamp 1649977179
transform 1 0 61548 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_669
timestamp 1649977179
transform 1 0 62652 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_681
timestamp 1649977179
transform 1 0 63756 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_693
timestamp 1649977179
transform 1 0 64860 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_699
timestamp 1649977179
transform 1 0 65412 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_701
timestamp 1649977179
transform 1 0 65596 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_713
timestamp 1649977179
transform 1 0 66700 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_92_725
timestamp 1649977179
transform 1 0 67804 0 1 52224
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_93_3
timestamp 1649977179
transform 1 0 1380 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_15
timestamp 1649977179
transform 1 0 2484 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_27
timestamp 1649977179
transform 1 0 3588 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_39
timestamp 1649977179
transform 1 0 4692 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_51
timestamp 1649977179
transform 1 0 5796 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_55
timestamp 1649977179
transform 1 0 6164 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_57
timestamp 1649977179
transform 1 0 6348 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_69
timestamp 1649977179
transform 1 0 7452 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_81
timestamp 1649977179
transform 1 0 8556 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_93
timestamp 1649977179
transform 1 0 9660 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_105
timestamp 1649977179
transform 1 0 10764 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_111
timestamp 1649977179
transform 1 0 11316 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_113
timestamp 1649977179
transform 1 0 11500 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_125
timestamp 1649977179
transform 1 0 12604 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_137
timestamp 1649977179
transform 1 0 13708 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_149
timestamp 1649977179
transform 1 0 14812 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_161
timestamp 1649977179
transform 1 0 15916 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_167
timestamp 1649977179
transform 1 0 16468 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_169
timestamp 1649977179
transform 1 0 16652 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_181
timestamp 1649977179
transform 1 0 17756 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_193
timestamp 1649977179
transform 1 0 18860 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_205
timestamp 1649977179
transform 1 0 19964 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_217
timestamp 1649977179
transform 1 0 21068 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_223
timestamp 1649977179
transform 1 0 21620 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_225
timestamp 1649977179
transform 1 0 21804 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_237
timestamp 1649977179
transform 1 0 22908 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_249
timestamp 1649977179
transform 1 0 24012 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_261
timestamp 1649977179
transform 1 0 25116 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_273
timestamp 1649977179
transform 1 0 26220 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_279
timestamp 1649977179
transform 1 0 26772 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_281
timestamp 1649977179
transform 1 0 26956 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_293
timestamp 1649977179
transform 1 0 28060 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_305
timestamp 1649977179
transform 1 0 29164 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_317
timestamp 1649977179
transform 1 0 30268 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_329
timestamp 1649977179
transform 1 0 31372 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_335
timestamp 1649977179
transform 1 0 31924 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_337
timestamp 1649977179
transform 1 0 32108 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_349
timestamp 1649977179
transform 1 0 33212 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_361
timestamp 1649977179
transform 1 0 34316 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_373
timestamp 1649977179
transform 1 0 35420 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_385
timestamp 1649977179
transform 1 0 36524 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_391
timestamp 1649977179
transform 1 0 37076 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_393
timestamp 1649977179
transform 1 0 37260 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_405
timestamp 1649977179
transform 1 0 38364 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_417
timestamp 1649977179
transform 1 0 39468 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_429
timestamp 1649977179
transform 1 0 40572 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_441
timestamp 1649977179
transform 1 0 41676 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_447
timestamp 1649977179
transform 1 0 42228 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_449
timestamp 1649977179
transform 1 0 42412 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_461
timestamp 1649977179
transform 1 0 43516 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_473
timestamp 1649977179
transform 1 0 44620 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_485
timestamp 1649977179
transform 1 0 45724 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_497
timestamp 1649977179
transform 1 0 46828 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_503
timestamp 1649977179
transform 1 0 47380 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_505
timestamp 1649977179
transform 1 0 47564 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_517
timestamp 1649977179
transform 1 0 48668 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_529
timestamp 1649977179
transform 1 0 49772 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_541
timestamp 1649977179
transform 1 0 50876 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_553
timestamp 1649977179
transform 1 0 51980 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_559
timestamp 1649977179
transform 1 0 52532 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_561
timestamp 1649977179
transform 1 0 52716 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_573
timestamp 1649977179
transform 1 0 53820 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_585
timestamp 1649977179
transform 1 0 54924 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_597
timestamp 1649977179
transform 1 0 56028 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_609
timestamp 1649977179
transform 1 0 57132 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_615
timestamp 1649977179
transform 1 0 57684 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_617
timestamp 1649977179
transform 1 0 57868 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_629
timestamp 1649977179
transform 1 0 58972 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_641
timestamp 1649977179
transform 1 0 60076 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_653
timestamp 1649977179
transform 1 0 61180 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_665
timestamp 1649977179
transform 1 0 62284 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_671
timestamp 1649977179
transform 1 0 62836 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_673
timestamp 1649977179
transform 1 0 63020 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_685
timestamp 1649977179
transform 1 0 64124 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_697
timestamp 1649977179
transform 1 0 65228 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_709
timestamp 1649977179
transform 1 0 66332 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_721
timestamp 1649977179
transform 1 0 67436 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_727
timestamp 1649977179
transform 1 0 67988 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_93_729
timestamp 1649977179
transform 1 0 68172 0 -1 53312
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_94_3
timestamp 1649977179
transform 1 0 1380 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_15
timestamp 1649977179
transform 1 0 2484 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_94_27
timestamp 1649977179
transform 1 0 3588 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_29
timestamp 1649977179
transform 1 0 3772 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_41
timestamp 1649977179
transform 1 0 4876 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_53
timestamp 1649977179
transform 1 0 5980 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_65
timestamp 1649977179
transform 1 0 7084 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_77
timestamp 1649977179
transform 1 0 8188 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_83
timestamp 1649977179
transform 1 0 8740 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_85
timestamp 1649977179
transform 1 0 8924 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_97
timestamp 1649977179
transform 1 0 10028 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_109
timestamp 1649977179
transform 1 0 11132 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_121
timestamp 1649977179
transform 1 0 12236 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_133
timestamp 1649977179
transform 1 0 13340 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_139
timestamp 1649977179
transform 1 0 13892 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_141
timestamp 1649977179
transform 1 0 14076 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_153
timestamp 1649977179
transform 1 0 15180 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_165
timestamp 1649977179
transform 1 0 16284 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_177
timestamp 1649977179
transform 1 0 17388 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_189
timestamp 1649977179
transform 1 0 18492 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_195
timestamp 1649977179
transform 1 0 19044 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_197
timestamp 1649977179
transform 1 0 19228 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_209
timestamp 1649977179
transform 1 0 20332 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_221
timestamp 1649977179
transform 1 0 21436 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_233
timestamp 1649977179
transform 1 0 22540 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_245
timestamp 1649977179
transform 1 0 23644 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_251
timestamp 1649977179
transform 1 0 24196 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_253
timestamp 1649977179
transform 1 0 24380 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_265
timestamp 1649977179
transform 1 0 25484 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_277
timestamp 1649977179
transform 1 0 26588 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_289
timestamp 1649977179
transform 1 0 27692 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_301
timestamp 1649977179
transform 1 0 28796 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_307
timestamp 1649977179
transform 1 0 29348 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_309
timestamp 1649977179
transform 1 0 29532 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_321
timestamp 1649977179
transform 1 0 30636 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_333
timestamp 1649977179
transform 1 0 31740 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_345
timestamp 1649977179
transform 1 0 32844 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_357
timestamp 1649977179
transform 1 0 33948 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_363
timestamp 1649977179
transform 1 0 34500 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_365
timestamp 1649977179
transform 1 0 34684 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_377
timestamp 1649977179
transform 1 0 35788 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_389
timestamp 1649977179
transform 1 0 36892 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_401
timestamp 1649977179
transform 1 0 37996 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_413
timestamp 1649977179
transform 1 0 39100 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_419
timestamp 1649977179
transform 1 0 39652 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_421
timestamp 1649977179
transform 1 0 39836 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_433
timestamp 1649977179
transform 1 0 40940 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_445
timestamp 1649977179
transform 1 0 42044 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_457
timestamp 1649977179
transform 1 0 43148 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_469
timestamp 1649977179
transform 1 0 44252 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_475
timestamp 1649977179
transform 1 0 44804 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_477
timestamp 1649977179
transform 1 0 44988 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_489
timestamp 1649977179
transform 1 0 46092 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_501
timestamp 1649977179
transform 1 0 47196 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_513
timestamp 1649977179
transform 1 0 48300 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_525
timestamp 1649977179
transform 1 0 49404 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_531
timestamp 1649977179
transform 1 0 49956 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_533
timestamp 1649977179
transform 1 0 50140 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_545
timestamp 1649977179
transform 1 0 51244 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_557
timestamp 1649977179
transform 1 0 52348 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_569
timestamp 1649977179
transform 1 0 53452 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_581
timestamp 1649977179
transform 1 0 54556 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_587
timestamp 1649977179
transform 1 0 55108 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_589
timestamp 1649977179
transform 1 0 55292 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_601
timestamp 1649977179
transform 1 0 56396 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_613
timestamp 1649977179
transform 1 0 57500 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_625
timestamp 1649977179
transform 1 0 58604 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_637
timestamp 1649977179
transform 1 0 59708 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_643
timestamp 1649977179
transform 1 0 60260 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_645
timestamp 1649977179
transform 1 0 60444 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_657
timestamp 1649977179
transform 1 0 61548 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_669
timestamp 1649977179
transform 1 0 62652 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_681
timestamp 1649977179
transform 1 0 63756 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_693
timestamp 1649977179
transform 1 0 64860 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_699
timestamp 1649977179
transform 1 0 65412 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_701
timestamp 1649977179
transform 1 0 65596 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_713
timestamp 1649977179
transform 1 0 66700 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_94_725
timestamp 1649977179
transform 1 0 67804 0 1 53312
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_95_3
timestamp 1649977179
transform 1 0 1380 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_15
timestamp 1649977179
transform 1 0 2484 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_27
timestamp 1649977179
transform 1 0 3588 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_39
timestamp 1649977179
transform 1 0 4692 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_95_51
timestamp 1649977179
transform 1 0 5796 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_55
timestamp 1649977179
transform 1 0 6164 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_57
timestamp 1649977179
transform 1 0 6348 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_69
timestamp 1649977179
transform 1 0 7452 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_81
timestamp 1649977179
transform 1 0 8556 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_93
timestamp 1649977179
transform 1 0 9660 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_105
timestamp 1649977179
transform 1 0 10764 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_111
timestamp 1649977179
transform 1 0 11316 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_113
timestamp 1649977179
transform 1 0 11500 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_125
timestamp 1649977179
transform 1 0 12604 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_137
timestamp 1649977179
transform 1 0 13708 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_149
timestamp 1649977179
transform 1 0 14812 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_161
timestamp 1649977179
transform 1 0 15916 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_167
timestamp 1649977179
transform 1 0 16468 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_169
timestamp 1649977179
transform 1 0 16652 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_181
timestamp 1649977179
transform 1 0 17756 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_193
timestamp 1649977179
transform 1 0 18860 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_205
timestamp 1649977179
transform 1 0 19964 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_217
timestamp 1649977179
transform 1 0 21068 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_223
timestamp 1649977179
transform 1 0 21620 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_225
timestamp 1649977179
transform 1 0 21804 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_237
timestamp 1649977179
transform 1 0 22908 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_249
timestamp 1649977179
transform 1 0 24012 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_261
timestamp 1649977179
transform 1 0 25116 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_273
timestamp 1649977179
transform 1 0 26220 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_279
timestamp 1649977179
transform 1 0 26772 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_281
timestamp 1649977179
transform 1 0 26956 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_293
timestamp 1649977179
transform 1 0 28060 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_305
timestamp 1649977179
transform 1 0 29164 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_317
timestamp 1649977179
transform 1 0 30268 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_329
timestamp 1649977179
transform 1 0 31372 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_335
timestamp 1649977179
transform 1 0 31924 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_337
timestamp 1649977179
transform 1 0 32108 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_349
timestamp 1649977179
transform 1 0 33212 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_361
timestamp 1649977179
transform 1 0 34316 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_373
timestamp 1649977179
transform 1 0 35420 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_385
timestamp 1649977179
transform 1 0 36524 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_391
timestamp 1649977179
transform 1 0 37076 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_393
timestamp 1649977179
transform 1 0 37260 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_405
timestamp 1649977179
transform 1 0 38364 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_417
timestamp 1649977179
transform 1 0 39468 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_429
timestamp 1649977179
transform 1 0 40572 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_441
timestamp 1649977179
transform 1 0 41676 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_447
timestamp 1649977179
transform 1 0 42228 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_449
timestamp 1649977179
transform 1 0 42412 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_461
timestamp 1649977179
transform 1 0 43516 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_473
timestamp 1649977179
transform 1 0 44620 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_485
timestamp 1649977179
transform 1 0 45724 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_497
timestamp 1649977179
transform 1 0 46828 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_503
timestamp 1649977179
transform 1 0 47380 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_505
timestamp 1649977179
transform 1 0 47564 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_517
timestamp 1649977179
transform 1 0 48668 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_529
timestamp 1649977179
transform 1 0 49772 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_541
timestamp 1649977179
transform 1 0 50876 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_553
timestamp 1649977179
transform 1 0 51980 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_559
timestamp 1649977179
transform 1 0 52532 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_561
timestamp 1649977179
transform 1 0 52716 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_573
timestamp 1649977179
transform 1 0 53820 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_585
timestamp 1649977179
transform 1 0 54924 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_597
timestamp 1649977179
transform 1 0 56028 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_609
timestamp 1649977179
transform 1 0 57132 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_615
timestamp 1649977179
transform 1 0 57684 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_617
timestamp 1649977179
transform 1 0 57868 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_629
timestamp 1649977179
transform 1 0 58972 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_641
timestamp 1649977179
transform 1 0 60076 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_653
timestamp 1649977179
transform 1 0 61180 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_665
timestamp 1649977179
transform 1 0 62284 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_671
timestamp 1649977179
transform 1 0 62836 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_673
timestamp 1649977179
transform 1 0 63020 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_685
timestamp 1649977179
transform 1 0 64124 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_697
timestamp 1649977179
transform 1 0 65228 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_709
timestamp 1649977179
transform 1 0 66332 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_721
timestamp 1649977179
transform 1 0 67436 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_727
timestamp 1649977179
transform 1 0 67988 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_95_729
timestamp 1649977179
transform 1 0 68172 0 -1 54400
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_96_3
timestamp 1649977179
transform 1 0 1380 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_15
timestamp 1649977179
transform 1 0 2484 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_96_27
timestamp 1649977179
transform 1 0 3588 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_29
timestamp 1649977179
transform 1 0 3772 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_41
timestamp 1649977179
transform 1 0 4876 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_53
timestamp 1649977179
transform 1 0 5980 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_65
timestamp 1649977179
transform 1 0 7084 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_77
timestamp 1649977179
transform 1 0 8188 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_83
timestamp 1649977179
transform 1 0 8740 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_85
timestamp 1649977179
transform 1 0 8924 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_97
timestamp 1649977179
transform 1 0 10028 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_109
timestamp 1649977179
transform 1 0 11132 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_121
timestamp 1649977179
transform 1 0 12236 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_133
timestamp 1649977179
transform 1 0 13340 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_139
timestamp 1649977179
transform 1 0 13892 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_141
timestamp 1649977179
transform 1 0 14076 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_153
timestamp 1649977179
transform 1 0 15180 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_165
timestamp 1649977179
transform 1 0 16284 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_177
timestamp 1649977179
transform 1 0 17388 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_189
timestamp 1649977179
transform 1 0 18492 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_195
timestamp 1649977179
transform 1 0 19044 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_197
timestamp 1649977179
transform 1 0 19228 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_209
timestamp 1649977179
transform 1 0 20332 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_221
timestamp 1649977179
transform 1 0 21436 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_233
timestamp 1649977179
transform 1 0 22540 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_245
timestamp 1649977179
transform 1 0 23644 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_251
timestamp 1649977179
transform 1 0 24196 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_253
timestamp 1649977179
transform 1 0 24380 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_265
timestamp 1649977179
transform 1 0 25484 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_277
timestamp 1649977179
transform 1 0 26588 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_289
timestamp 1649977179
transform 1 0 27692 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_301
timestamp 1649977179
transform 1 0 28796 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_307
timestamp 1649977179
transform 1 0 29348 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_309
timestamp 1649977179
transform 1 0 29532 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_321
timestamp 1649977179
transform 1 0 30636 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_333
timestamp 1649977179
transform 1 0 31740 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_345
timestamp 1649977179
transform 1 0 32844 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_357
timestamp 1649977179
transform 1 0 33948 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_363
timestamp 1649977179
transform 1 0 34500 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_365
timestamp 1649977179
transform 1 0 34684 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_377
timestamp 1649977179
transform 1 0 35788 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_389
timestamp 1649977179
transform 1 0 36892 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_401
timestamp 1649977179
transform 1 0 37996 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_413
timestamp 1649977179
transform 1 0 39100 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_419
timestamp 1649977179
transform 1 0 39652 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_421
timestamp 1649977179
transform 1 0 39836 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_433
timestamp 1649977179
transform 1 0 40940 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_445
timestamp 1649977179
transform 1 0 42044 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_457
timestamp 1649977179
transform 1 0 43148 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_469
timestamp 1649977179
transform 1 0 44252 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_475
timestamp 1649977179
transform 1 0 44804 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_477
timestamp 1649977179
transform 1 0 44988 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_489
timestamp 1649977179
transform 1 0 46092 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_501
timestamp 1649977179
transform 1 0 47196 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_513
timestamp 1649977179
transform 1 0 48300 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_525
timestamp 1649977179
transform 1 0 49404 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_531
timestamp 1649977179
transform 1 0 49956 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_533
timestamp 1649977179
transform 1 0 50140 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_545
timestamp 1649977179
transform 1 0 51244 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_557
timestamp 1649977179
transform 1 0 52348 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_569
timestamp 1649977179
transform 1 0 53452 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_581
timestamp 1649977179
transform 1 0 54556 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_587
timestamp 1649977179
transform 1 0 55108 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_589
timestamp 1649977179
transform 1 0 55292 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_601
timestamp 1649977179
transform 1 0 56396 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_613
timestamp 1649977179
transform 1 0 57500 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_625
timestamp 1649977179
transform 1 0 58604 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_637
timestamp 1649977179
transform 1 0 59708 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_643
timestamp 1649977179
transform 1 0 60260 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_645
timestamp 1649977179
transform 1 0 60444 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_657
timestamp 1649977179
transform 1 0 61548 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_669
timestamp 1649977179
transform 1 0 62652 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_681
timestamp 1649977179
transform 1 0 63756 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_693
timestamp 1649977179
transform 1 0 64860 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_699
timestamp 1649977179
transform 1 0 65412 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_701
timestamp 1649977179
transform 1 0 65596 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_713
timestamp 1649977179
transform 1 0 66700 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_96_725
timestamp 1649977179
transform 1 0 67804 0 1 54400
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_97_3
timestamp 1649977179
transform 1 0 1380 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_15
timestamp 1649977179
transform 1 0 2484 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_27
timestamp 1649977179
transform 1 0 3588 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_39
timestamp 1649977179
transform 1 0 4692 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_97_51
timestamp 1649977179
transform 1 0 5796 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_97_55
timestamp 1649977179
transform 1 0 6164 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_57
timestamp 1649977179
transform 1 0 6348 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_69
timestamp 1649977179
transform 1 0 7452 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_81
timestamp 1649977179
transform 1 0 8556 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_93
timestamp 1649977179
transform 1 0 9660 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_105
timestamp 1649977179
transform 1 0 10764 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_111
timestamp 1649977179
transform 1 0 11316 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_113
timestamp 1649977179
transform 1 0 11500 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_125
timestamp 1649977179
transform 1 0 12604 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_137
timestamp 1649977179
transform 1 0 13708 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_149
timestamp 1649977179
transform 1 0 14812 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_161
timestamp 1649977179
transform 1 0 15916 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_167
timestamp 1649977179
transform 1 0 16468 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_169
timestamp 1649977179
transform 1 0 16652 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_181
timestamp 1649977179
transform 1 0 17756 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_193
timestamp 1649977179
transform 1 0 18860 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_205
timestamp 1649977179
transform 1 0 19964 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_217
timestamp 1649977179
transform 1 0 21068 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_223
timestamp 1649977179
transform 1 0 21620 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_225
timestamp 1649977179
transform 1 0 21804 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_237
timestamp 1649977179
transform 1 0 22908 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_249
timestamp 1649977179
transform 1 0 24012 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_261
timestamp 1649977179
transform 1 0 25116 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_273
timestamp 1649977179
transform 1 0 26220 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_279
timestamp 1649977179
transform 1 0 26772 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_281
timestamp 1649977179
transform 1 0 26956 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_293
timestamp 1649977179
transform 1 0 28060 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_305
timestamp 1649977179
transform 1 0 29164 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_317
timestamp 1649977179
transform 1 0 30268 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_329
timestamp 1649977179
transform 1 0 31372 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_335
timestamp 1649977179
transform 1 0 31924 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_337
timestamp 1649977179
transform 1 0 32108 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_349
timestamp 1649977179
transform 1 0 33212 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_361
timestamp 1649977179
transform 1 0 34316 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_373
timestamp 1649977179
transform 1 0 35420 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_385
timestamp 1649977179
transform 1 0 36524 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_391
timestamp 1649977179
transform 1 0 37076 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_393
timestamp 1649977179
transform 1 0 37260 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_405
timestamp 1649977179
transform 1 0 38364 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_417
timestamp 1649977179
transform 1 0 39468 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_429
timestamp 1649977179
transform 1 0 40572 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_441
timestamp 1649977179
transform 1 0 41676 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_447
timestamp 1649977179
transform 1 0 42228 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_449
timestamp 1649977179
transform 1 0 42412 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_461
timestamp 1649977179
transform 1 0 43516 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_473
timestamp 1649977179
transform 1 0 44620 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_485
timestamp 1649977179
transform 1 0 45724 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_497
timestamp 1649977179
transform 1 0 46828 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_503
timestamp 1649977179
transform 1 0 47380 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_505
timestamp 1649977179
transform 1 0 47564 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_517
timestamp 1649977179
transform 1 0 48668 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_529
timestamp 1649977179
transform 1 0 49772 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_541
timestamp 1649977179
transform 1 0 50876 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_553
timestamp 1649977179
transform 1 0 51980 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_559
timestamp 1649977179
transform 1 0 52532 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_561
timestamp 1649977179
transform 1 0 52716 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_573
timestamp 1649977179
transform 1 0 53820 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_585
timestamp 1649977179
transform 1 0 54924 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_597
timestamp 1649977179
transform 1 0 56028 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_609
timestamp 1649977179
transform 1 0 57132 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_615
timestamp 1649977179
transform 1 0 57684 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_617
timestamp 1649977179
transform 1 0 57868 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_629
timestamp 1649977179
transform 1 0 58972 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_641
timestamp 1649977179
transform 1 0 60076 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_653
timestamp 1649977179
transform 1 0 61180 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_665
timestamp 1649977179
transform 1 0 62284 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_671
timestamp 1649977179
transform 1 0 62836 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_673
timestamp 1649977179
transform 1 0 63020 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_685
timestamp 1649977179
transform 1 0 64124 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_697
timestamp 1649977179
transform 1 0 65228 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_709
timestamp 1649977179
transform 1 0 66332 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_721
timestamp 1649977179
transform 1 0 67436 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_727
timestamp 1649977179
transform 1 0 67988 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_97_729
timestamp 1649977179
transform 1 0 68172 0 -1 55488
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_98_3
timestamp 1649977179
transform 1 0 1380 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_15
timestamp 1649977179
transform 1 0 2484 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_98_27
timestamp 1649977179
transform 1 0 3588 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_29
timestamp 1649977179
transform 1 0 3772 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_41
timestamp 1649977179
transform 1 0 4876 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_53
timestamp 1649977179
transform 1 0 5980 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_65
timestamp 1649977179
transform 1 0 7084 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_77
timestamp 1649977179
transform 1 0 8188 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_83
timestamp 1649977179
transform 1 0 8740 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_85
timestamp 1649977179
transform 1 0 8924 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_97
timestamp 1649977179
transform 1 0 10028 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_109
timestamp 1649977179
transform 1 0 11132 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_121
timestamp 1649977179
transform 1 0 12236 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_133
timestamp 1649977179
transform 1 0 13340 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_139
timestamp 1649977179
transform 1 0 13892 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_141
timestamp 1649977179
transform 1 0 14076 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_153
timestamp 1649977179
transform 1 0 15180 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_165
timestamp 1649977179
transform 1 0 16284 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_177
timestamp 1649977179
transform 1 0 17388 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_189
timestamp 1649977179
transform 1 0 18492 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_195
timestamp 1649977179
transform 1 0 19044 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_197
timestamp 1649977179
transform 1 0 19228 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_209
timestamp 1649977179
transform 1 0 20332 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_221
timestamp 1649977179
transform 1 0 21436 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_233
timestamp 1649977179
transform 1 0 22540 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_245
timestamp 1649977179
transform 1 0 23644 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_251
timestamp 1649977179
transform 1 0 24196 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_253
timestamp 1649977179
transform 1 0 24380 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_265
timestamp 1649977179
transform 1 0 25484 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_277
timestamp 1649977179
transform 1 0 26588 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_289
timestamp 1649977179
transform 1 0 27692 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_301
timestamp 1649977179
transform 1 0 28796 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_307
timestamp 1649977179
transform 1 0 29348 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_309
timestamp 1649977179
transform 1 0 29532 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_321
timestamp 1649977179
transform 1 0 30636 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_333
timestamp 1649977179
transform 1 0 31740 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_345
timestamp 1649977179
transform 1 0 32844 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_357
timestamp 1649977179
transform 1 0 33948 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_363
timestamp 1649977179
transform 1 0 34500 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_365
timestamp 1649977179
transform 1 0 34684 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_377
timestamp 1649977179
transform 1 0 35788 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_389
timestamp 1649977179
transform 1 0 36892 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_401
timestamp 1649977179
transform 1 0 37996 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_413
timestamp 1649977179
transform 1 0 39100 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_419
timestamp 1649977179
transform 1 0 39652 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_421
timestamp 1649977179
transform 1 0 39836 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_433
timestamp 1649977179
transform 1 0 40940 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_445
timestamp 1649977179
transform 1 0 42044 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_457
timestamp 1649977179
transform 1 0 43148 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_469
timestamp 1649977179
transform 1 0 44252 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_475
timestamp 1649977179
transform 1 0 44804 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_477
timestamp 1649977179
transform 1 0 44988 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_489
timestamp 1649977179
transform 1 0 46092 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_501
timestamp 1649977179
transform 1 0 47196 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_513
timestamp 1649977179
transform 1 0 48300 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_525
timestamp 1649977179
transform 1 0 49404 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_531
timestamp 1649977179
transform 1 0 49956 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_533
timestamp 1649977179
transform 1 0 50140 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_545
timestamp 1649977179
transform 1 0 51244 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_557
timestamp 1649977179
transform 1 0 52348 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_569
timestamp 1649977179
transform 1 0 53452 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_581
timestamp 1649977179
transform 1 0 54556 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_587
timestamp 1649977179
transform 1 0 55108 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_589
timestamp 1649977179
transform 1 0 55292 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_601
timestamp 1649977179
transform 1 0 56396 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_613
timestamp 1649977179
transform 1 0 57500 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_625
timestamp 1649977179
transform 1 0 58604 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_637
timestamp 1649977179
transform 1 0 59708 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_643
timestamp 1649977179
transform 1 0 60260 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_645
timestamp 1649977179
transform 1 0 60444 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_657
timestamp 1649977179
transform 1 0 61548 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_669
timestamp 1649977179
transform 1 0 62652 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_681
timestamp 1649977179
transform 1 0 63756 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_693
timestamp 1649977179
transform 1 0 64860 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_699
timestamp 1649977179
transform 1 0 65412 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_701
timestamp 1649977179
transform 1 0 65596 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_713
timestamp 1649977179
transform 1 0 66700 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_98_725
timestamp 1649977179
transform 1 0 67804 0 1 55488
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_99_3
timestamp 1649977179
transform 1 0 1380 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_15
timestamp 1649977179
transform 1 0 2484 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_27
timestamp 1649977179
transform 1 0 3588 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_39
timestamp 1649977179
transform 1 0 4692 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_99_51
timestamp 1649977179
transform 1 0 5796 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_99_55
timestamp 1649977179
transform 1 0 6164 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_57
timestamp 1649977179
transform 1 0 6348 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_69
timestamp 1649977179
transform 1 0 7452 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_81
timestamp 1649977179
transform 1 0 8556 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_93
timestamp 1649977179
transform 1 0 9660 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_105
timestamp 1649977179
transform 1 0 10764 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_111
timestamp 1649977179
transform 1 0 11316 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_113
timestamp 1649977179
transform 1 0 11500 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_125
timestamp 1649977179
transform 1 0 12604 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_137
timestamp 1649977179
transform 1 0 13708 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_149
timestamp 1649977179
transform 1 0 14812 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_161
timestamp 1649977179
transform 1 0 15916 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_167
timestamp 1649977179
transform 1 0 16468 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_169
timestamp 1649977179
transform 1 0 16652 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_181
timestamp 1649977179
transform 1 0 17756 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_193
timestamp 1649977179
transform 1 0 18860 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_205
timestamp 1649977179
transform 1 0 19964 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_217
timestamp 1649977179
transform 1 0 21068 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_223
timestamp 1649977179
transform 1 0 21620 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_225
timestamp 1649977179
transform 1 0 21804 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_237
timestamp 1649977179
transform 1 0 22908 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_249
timestamp 1649977179
transform 1 0 24012 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_261
timestamp 1649977179
transform 1 0 25116 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_273
timestamp 1649977179
transform 1 0 26220 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_279
timestamp 1649977179
transform 1 0 26772 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_281
timestamp 1649977179
transform 1 0 26956 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_293
timestamp 1649977179
transform 1 0 28060 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_305
timestamp 1649977179
transform 1 0 29164 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_317
timestamp 1649977179
transform 1 0 30268 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_329
timestamp 1649977179
transform 1 0 31372 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_335
timestamp 1649977179
transform 1 0 31924 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_337
timestamp 1649977179
transform 1 0 32108 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_349
timestamp 1649977179
transform 1 0 33212 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_361
timestamp 1649977179
transform 1 0 34316 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_373
timestamp 1649977179
transform 1 0 35420 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_385
timestamp 1649977179
transform 1 0 36524 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_391
timestamp 1649977179
transform 1 0 37076 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_393
timestamp 1649977179
transform 1 0 37260 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_405
timestamp 1649977179
transform 1 0 38364 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_417
timestamp 1649977179
transform 1 0 39468 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_429
timestamp 1649977179
transform 1 0 40572 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_441
timestamp 1649977179
transform 1 0 41676 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_447
timestamp 1649977179
transform 1 0 42228 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_449
timestamp 1649977179
transform 1 0 42412 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_461
timestamp 1649977179
transform 1 0 43516 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_473
timestamp 1649977179
transform 1 0 44620 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_485
timestamp 1649977179
transform 1 0 45724 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_497
timestamp 1649977179
transform 1 0 46828 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_503
timestamp 1649977179
transform 1 0 47380 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_505
timestamp 1649977179
transform 1 0 47564 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_517
timestamp 1649977179
transform 1 0 48668 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_529
timestamp 1649977179
transform 1 0 49772 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_541
timestamp 1649977179
transform 1 0 50876 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_553
timestamp 1649977179
transform 1 0 51980 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_559
timestamp 1649977179
transform 1 0 52532 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_561
timestamp 1649977179
transform 1 0 52716 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_573
timestamp 1649977179
transform 1 0 53820 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_585
timestamp 1649977179
transform 1 0 54924 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_597
timestamp 1649977179
transform 1 0 56028 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_609
timestamp 1649977179
transform 1 0 57132 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_615
timestamp 1649977179
transform 1 0 57684 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_617
timestamp 1649977179
transform 1 0 57868 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_629
timestamp 1649977179
transform 1 0 58972 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_641
timestamp 1649977179
transform 1 0 60076 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_653
timestamp 1649977179
transform 1 0 61180 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_665
timestamp 1649977179
transform 1 0 62284 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_671
timestamp 1649977179
transform 1 0 62836 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_673
timestamp 1649977179
transform 1 0 63020 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_685
timestamp 1649977179
transform 1 0 64124 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_697
timestamp 1649977179
transform 1 0 65228 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_709
timestamp 1649977179
transform 1 0 66332 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_721
timestamp 1649977179
transform 1 0 67436 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_727
timestamp 1649977179
transform 1 0 67988 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_99_729
timestamp 1649977179
transform 1 0 68172 0 -1 56576
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_100_3
timestamp 1649977179
transform 1 0 1380 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_15
timestamp 1649977179
transform 1 0 2484 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_100_27
timestamp 1649977179
transform 1 0 3588 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_29
timestamp 1649977179
transform 1 0 3772 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_41
timestamp 1649977179
transform 1 0 4876 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_53
timestamp 1649977179
transform 1 0 5980 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_65
timestamp 1649977179
transform 1 0 7084 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_77
timestamp 1649977179
transform 1 0 8188 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_83
timestamp 1649977179
transform 1 0 8740 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_85
timestamp 1649977179
transform 1 0 8924 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_97
timestamp 1649977179
transform 1 0 10028 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_109
timestamp 1649977179
transform 1 0 11132 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_121
timestamp 1649977179
transform 1 0 12236 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_133
timestamp 1649977179
transform 1 0 13340 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_139
timestamp 1649977179
transform 1 0 13892 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_141
timestamp 1649977179
transform 1 0 14076 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_153
timestamp 1649977179
transform 1 0 15180 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_165
timestamp 1649977179
transform 1 0 16284 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_177
timestamp 1649977179
transform 1 0 17388 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_189
timestamp 1649977179
transform 1 0 18492 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_195
timestamp 1649977179
transform 1 0 19044 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_197
timestamp 1649977179
transform 1 0 19228 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_209
timestamp 1649977179
transform 1 0 20332 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_100_221
timestamp 1649977179
transform 1 0 21436 0 1 56576
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_100_228
timestamp 1649977179
transform 1 0 22080 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_240
timestamp 1649977179
transform 1 0 23184 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_253
timestamp 1649977179
transform 1 0 24380 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_265
timestamp 1649977179
transform 1 0 25484 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_100_277
timestamp 1649977179
transform 1 0 26588 0 1 56576
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_100_282
timestamp 1649977179
transform 1 0 27048 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_294
timestamp 1649977179
transform 1 0 28152 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_100_306
timestamp 1649977179
transform 1 0 29256 0 1 56576
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_100_309
timestamp 1649977179
transform 1 0 29532 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_321
timestamp 1649977179
transform 1 0 30636 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_333
timestamp 1649977179
transform 1 0 31740 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_345
timestamp 1649977179
transform 1 0 32844 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_357
timestamp 1649977179
transform 1 0 33948 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_363
timestamp 1649977179
transform 1 0 34500 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_365
timestamp 1649977179
transform 1 0 34684 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_377
timestamp 1649977179
transform 1 0 35788 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_389
timestamp 1649977179
transform 1 0 36892 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_401
timestamp 1649977179
transform 1 0 37996 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_100_409
timestamp 1649977179
transform 1 0 38732 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_100_414
timestamp 1649977179
transform 1 0 39192 0 1 56576
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_100_421
timestamp 1649977179
transform 1 0 39836 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_433
timestamp 1649977179
transform 1 0 40940 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_445
timestamp 1649977179
transform 1 0 42044 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_457
timestamp 1649977179
transform 1 0 43148 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_469
timestamp 1649977179
transform 1 0 44252 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_475
timestamp 1649977179
transform 1 0 44804 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_477
timestamp 1649977179
transform 1 0 44988 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_489
timestamp 1649977179
transform 1 0 46092 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_501
timestamp 1649977179
transform 1 0 47196 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_513
timestamp 1649977179
transform 1 0 48300 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_525
timestamp 1649977179
transform 1 0 49404 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_531
timestamp 1649977179
transform 1 0 49956 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_533
timestamp 1649977179
transform 1 0 50140 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_545
timestamp 1649977179
transform 1 0 51244 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_557
timestamp 1649977179
transform 1 0 52348 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_569
timestamp 1649977179
transform 1 0 53452 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_581
timestamp 1649977179
transform 1 0 54556 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_587
timestamp 1649977179
transform 1 0 55108 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_589
timestamp 1649977179
transform 1 0 55292 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_601
timestamp 1649977179
transform 1 0 56396 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_613
timestamp 1649977179
transform 1 0 57500 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_625
timestamp 1649977179
transform 1 0 58604 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_637
timestamp 1649977179
transform 1 0 59708 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_643
timestamp 1649977179
transform 1 0 60260 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_645
timestamp 1649977179
transform 1 0 60444 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_657
timestamp 1649977179
transform 1 0 61548 0 1 56576
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_100_666
timestamp 1649977179
transform 1 0 62376 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_678
timestamp 1649977179
transform 1 0 63480 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_690
timestamp 1649977179
transform 1 0 64584 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_100_698
timestamp 1649977179
transform 1 0 65320 0 1 56576
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_100_701
timestamp 1649977179
transform 1 0 65596 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_713
timestamp 1649977179
transform 1 0 66700 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_725
timestamp 1649977179
transform 1 0 67804 0 1 56576
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_101_3
timestamp 1649977179
transform 1 0 1380 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_15
timestamp 1649977179
transform 1 0 2484 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_101_24
timestamp 1649977179
transform 1 0 3312 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_29
timestamp 1649977179
transform 1 0 3772 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_101_36
timestamp 1649977179
transform 1 0 4416 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_101_45
timestamp 1649977179
transform 1 0 5244 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_52
timestamp 1649977179
transform 1 0 5888 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_57
timestamp 1649977179
transform 1 0 6348 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_61
timestamp 1649977179
transform 1 0 6716 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_65
timestamp 1649977179
transform 1 0 7084 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_72
timestamp 1649977179
transform 1 0 7728 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_76
timestamp 1649977179
transform 1 0 8096 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_80
timestamp 1649977179
transform 1 0 8464 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_101_85
timestamp 1649977179
transform 1 0 8924 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_101_90
timestamp 1649977179
transform 1 0 9384 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_101_101
timestamp 1649977179
transform 1 0 10396 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_108
timestamp 1649977179
transform 1 0 11040 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_101_113
timestamp 1649977179
transform 1 0 11500 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_101_119
timestamp 1649977179
transform 1 0 12052 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_101_126
timestamp 1649977179
transform 1 0 12696 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_132
timestamp 1649977179
transform 1 0 13248 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_136
timestamp 1649977179
transform 1 0 13616 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_101_144
timestamp 1649977179
transform 1 0 14352 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_101_155
timestamp 1649977179
transform 1 0 15364 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_101_162
timestamp 1649977179
transform 1 0 16008 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_169
timestamp 1649977179
transform 1 0 16652 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_173
timestamp 1649977179
transform 1 0 17020 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_101_180
timestamp 1649977179
transform 1 0 17664 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_101_188
timestamp 1649977179
transform 1 0 18400 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_192
timestamp 1649977179
transform 1 0 18768 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_101_200
timestamp 1649977179
transform 1 0 19504 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_101_209
timestamp 1649977179
transform 1 0 20332 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_101_216
timestamp 1649977179
transform 1 0 20976 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_101_225
timestamp 1649977179
transform 1 0 21804 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_101_234
timestamp 1649977179
transform 1 0 22632 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_101_242
timestamp 1649977179
transform 1 0 23368 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_101_246
timestamp 1649977179
transform 1 0 23736 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_101_256
timestamp 1649977179
transform 1 0 24656 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_263
timestamp 1649977179
transform 1 0 25300 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_101_270
timestamp 1649977179
transform 1 0 25944 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_101_278
timestamp 1649977179
transform 1 0 26680 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_101_281
timestamp 1649977179
transform 1 0 26956 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_101_288
timestamp 1649977179
transform 1 0 27600 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_101_297
timestamp 1649977179
transform 1 0 28428 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_304
timestamp 1649977179
transform 1 0 29072 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_309
timestamp 1649977179
transform 1 0 29532 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_313
timestamp 1649977179
transform 1 0 29900 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_317
timestamp 1649977179
transform 1 0 30268 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_324
timestamp 1649977179
transform 1 0 30912 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_328
timestamp 1649977179
transform 1 0 31280 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_332
timestamp 1649977179
transform 1 0 31648 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_101_337
timestamp 1649977179
transform 1 0 32108 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_101_342
timestamp 1649977179
transform 1 0 32568 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_101_353
timestamp 1649977179
transform 1 0 33580 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_360
timestamp 1649977179
transform 1 0 34224 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_101_365
timestamp 1649977179
transform 1 0 34684 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_101_371
timestamp 1649977179
transform 1 0 35236 0 -1 57664
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_101_378
timestamp 1649977179
transform 1 0 35880 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_101_390
timestamp 1649977179
transform 1 0 36984 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_101_396
timestamp 1649977179
transform 1 0 37536 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_403
timestamp 1649977179
transform 1 0 38180 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_101_410
timestamp 1649977179
transform 1 0 38824 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_101_418
timestamp 1649977179
transform 1 0 39560 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_421
timestamp 1649977179
transform 1 0 39836 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_101_426
timestamp 1649977179
transform 1 0 40296 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_101_433
timestamp 1649977179
transform 1 0 40940 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_101_444
timestamp 1649977179
transform 1 0 41952 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_101_452
timestamp 1649977179
transform 1 0 42688 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_458
timestamp 1649977179
transform 1 0 43240 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_462
timestamp 1649977179
transform 1 0 43608 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_101_469
timestamp 1649977179
transform 1 0 44252 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_475
timestamp 1649977179
transform 1 0 44804 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_480
timestamp 1649977179
transform 1 0 45264 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_101_487
timestamp 1649977179
transform 1 0 45908 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_101_498
timestamp 1649977179
transform 1 0 46920 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_101_508
timestamp 1649977179
transform 1 0 47840 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_512
timestamp 1649977179
transform 1 0 48208 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_516
timestamp 1649977179
transform 1 0 48576 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_101_523
timestamp 1649977179
transform 1 0 49220 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_101_531
timestamp 1649977179
transform 1 0 49956 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_536
timestamp 1649977179
transform 1 0 50416 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_101_543
timestamp 1649977179
transform 1 0 51060 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_101_552
timestamp 1649977179
transform 1 0 51888 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_101_564
timestamp 1649977179
transform 1 0 52992 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_571
timestamp 1649977179
transform 1 0 53636 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_101_578
timestamp 1649977179
transform 1 0 54280 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_101_586
timestamp 1649977179
transform 1 0 55016 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_101_592
timestamp 1649977179
transform 1 0 55568 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_599
timestamp 1649977179
transform 1 0 56212 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_101_606
timestamp 1649977179
transform 1 0 56856 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_101_614
timestamp 1649977179
transform 1 0 57592 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_101_620
timestamp 1649977179
transform 1 0 58144 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_627
timestamp 1649977179
transform 1 0 58788 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_101_634
timestamp 1649977179
transform 1 0 59432 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_101_642
timestamp 1649977179
transform 1 0 60168 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_101_648
timestamp 1649977179
transform 1 0 60720 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_655
timestamp 1649977179
transform 1 0 61364 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_101_662
timestamp 1649977179
transform 1 0 62008 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_101_670
timestamp 1649977179
transform 1 0 62744 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_673
timestamp 1649977179
transform 1 0 63020 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_101_678
timestamp 1649977179
transform 1 0 63480 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_101_685
timestamp 1649977179
transform 1 0 64124 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_101_696
timestamp 1649977179
transform 1 0 65136 0 -1 57664
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_101_704
timestamp 1649977179
transform 1 0 65872 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_101_716
timestamp 1649977179
transform 1 0 66976 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_101_720
timestamp 1649977179
transform 1 0 67344 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_101_729
timestamp 1649977179
transform 1 0 68172 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1649977179
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1649977179
transform -1 0 68816 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1649977179
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1649977179
transform -1 0 68816 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1649977179
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1649977179
transform -1 0 68816 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1649977179
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1649977179
transform -1 0 68816 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1649977179
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1649977179
transform -1 0 68816 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1649977179
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1649977179
transform -1 0 68816 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1649977179
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1649977179
transform -1 0 68816 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1649977179
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1649977179
transform -1 0 68816 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1649977179
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1649977179
transform -1 0 68816 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1649977179
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1649977179
transform -1 0 68816 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1649977179
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1649977179
transform -1 0 68816 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1649977179
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1649977179
transform -1 0 68816 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1649977179
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1649977179
transform -1 0 68816 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1649977179
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1649977179
transform -1 0 68816 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1649977179
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1649977179
transform -1 0 68816 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1649977179
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1649977179
transform -1 0 68816 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1649977179
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1649977179
transform -1 0 68816 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1649977179
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1649977179
transform -1 0 68816 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1649977179
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1649977179
transform -1 0 68816 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1649977179
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1649977179
transform -1 0 68816 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1649977179
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1649977179
transform -1 0 68816 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1649977179
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1649977179
transform -1 0 68816 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1649977179
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1649977179
transform -1 0 68816 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1649977179
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1649977179
transform -1 0 68816 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1649977179
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1649977179
transform -1 0 68816 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1649977179
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1649977179
transform -1 0 68816 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1649977179
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1649977179
transform -1 0 68816 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1649977179
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1649977179
transform -1 0 68816 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1649977179
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1649977179
transform -1 0 68816 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1649977179
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1649977179
transform -1 0 68816 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1649977179
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1649977179
transform -1 0 68816 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1649977179
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1649977179
transform -1 0 68816 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1649977179
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1649977179
transform -1 0 68816 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1649977179
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1649977179
transform -1 0 68816 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1649977179
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1649977179
transform -1 0 68816 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1649977179
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1649977179
transform -1 0 68816 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1649977179
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1649977179
transform -1 0 68816 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1649977179
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1649977179
transform -1 0 68816 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1649977179
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1649977179
transform -1 0 68816 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1649977179
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1649977179
transform -1 0 68816 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1649977179
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1649977179
transform -1 0 68816 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1649977179
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1649977179
transform -1 0 68816 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1649977179
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1649977179
transform -1 0 68816 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1649977179
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1649977179
transform -1 0 68816 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1649977179
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1649977179
transform -1 0 68816 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1649977179
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1649977179
transform -1 0 68816 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1649977179
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1649977179
transform -1 0 68816 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1649977179
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1649977179
transform -1 0 68816 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1649977179
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1649977179
transform -1 0 68816 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1649977179
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1649977179
transform -1 0 68816 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1649977179
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1649977179
transform -1 0 68816 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1649977179
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1649977179
transform -1 0 68816 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1649977179
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1649977179
transform -1 0 68816 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1649977179
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1649977179
transform -1 0 68816 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1649977179
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1649977179
transform -1 0 68816 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1649977179
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1649977179
transform -1 0 68816 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1649977179
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1649977179
transform -1 0 68816 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1649977179
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1649977179
transform -1 0 68816 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1649977179
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1649977179
transform -1 0 68816 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1649977179
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1649977179
transform -1 0 68816 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1649977179
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1649977179
transform -1 0 68816 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1649977179
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1649977179
transform -1 0 68816 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1649977179
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1649977179
transform -1 0 68816 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1649977179
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1649977179
transform -1 0 68816 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1649977179
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1649977179
transform -1 0 68816 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1649977179
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1649977179
transform -1 0 68816 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1649977179
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1649977179
transform -1 0 68816 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1649977179
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1649977179
transform -1 0 68816 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1649977179
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1649977179
transform -1 0 68816 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1649977179
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1649977179
transform -1 0 68816 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1649977179
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1649977179
transform -1 0 68816 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1649977179
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1649977179
transform -1 0 68816 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1649977179
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1649977179
transform -1 0 68816 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1649977179
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1649977179
transform -1 0 68816 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1649977179
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1649977179
transform -1 0 68816 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1649977179
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1649977179
transform -1 0 68816 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1649977179
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1649977179
transform -1 0 68816 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1649977179
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1649977179
transform -1 0 68816 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1649977179
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1649977179
transform -1 0 68816 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1649977179
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1649977179
transform -1 0 68816 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1649977179
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1649977179
transform -1 0 68816 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1649977179
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1649977179
transform -1 0 68816 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1649977179
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1649977179
transform -1 0 68816 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_166
timestamp 1649977179
transform 1 0 1104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 1649977179
transform -1 0 68816 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_168
timestamp 1649977179
transform 1 0 1104 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_169
timestamp 1649977179
transform -1 0 68816 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_170
timestamp 1649977179
transform 1 0 1104 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_171
timestamp 1649977179
transform -1 0 68816 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_172
timestamp 1649977179
transform 1 0 1104 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_173
timestamp 1649977179
transform -1 0 68816 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_174
timestamp 1649977179
transform 1 0 1104 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_175
timestamp 1649977179
transform -1 0 68816 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_176
timestamp 1649977179
transform 1 0 1104 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_177
timestamp 1649977179
transform -1 0 68816 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_178
timestamp 1649977179
transform 1 0 1104 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_179
timestamp 1649977179
transform -1 0 68816 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_180
timestamp 1649977179
transform 1 0 1104 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_181
timestamp 1649977179
transform -1 0 68816 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_182
timestamp 1649977179
transform 1 0 1104 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_183
timestamp 1649977179
transform -1 0 68816 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_184
timestamp 1649977179
transform 1 0 1104 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_185
timestamp 1649977179
transform -1 0 68816 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_186
timestamp 1649977179
transform 1 0 1104 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_187
timestamp 1649977179
transform -1 0 68816 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_188
timestamp 1649977179
transform 1 0 1104 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_189
timestamp 1649977179
transform -1 0 68816 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_190
timestamp 1649977179
transform 1 0 1104 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_191
timestamp 1649977179
transform -1 0 68816 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_192
timestamp 1649977179
transform 1 0 1104 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_193
timestamp 1649977179
transform -1 0 68816 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_194
timestamp 1649977179
transform 1 0 1104 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_195
timestamp 1649977179
transform -1 0 68816 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_196
timestamp 1649977179
transform 1 0 1104 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_197
timestamp 1649977179
transform -1 0 68816 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_198
timestamp 1649977179
transform 1 0 1104 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_199
timestamp 1649977179
transform -1 0 68816 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_200
timestamp 1649977179
transform 1 0 1104 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_201
timestamp 1649977179
transform -1 0 68816 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_202
timestamp 1649977179
transform 1 0 1104 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_203
timestamp 1649977179
transform -1 0 68816 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1649977179
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1649977179
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1649977179
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1649977179
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1649977179
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1649977179
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1649977179
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1649977179
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1649977179
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1649977179
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1649977179
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1649977179
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1649977179
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1649977179
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1649977179
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1649977179
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1649977179
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1649977179
transform 1 0 50048 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1649977179
transform 1 0 52624 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1649977179
transform 1 0 55200 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1649977179
transform 1 0 57776 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1649977179
transform 1 0 60352 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1649977179
transform 1 0 62928 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1649977179
transform 1 0 65504 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1649977179
transform 1 0 68080 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1649977179
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1649977179
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1649977179
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1649977179
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1649977179
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1649977179
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1649977179
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1649977179
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1649977179
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1649977179
transform 1 0 52624 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1649977179
transform 1 0 57776 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1649977179
transform 1 0 62928 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1649977179
transform 1 0 68080 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1649977179
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1649977179
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1649977179
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1649977179
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1649977179
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1649977179
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1649977179
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1649977179
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1649977179
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1649977179
transform 1 0 50048 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1649977179
transform 1 0 55200 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1649977179
transform 1 0 60352 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1649977179
transform 1 0 65504 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1649977179
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1649977179
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1649977179
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1649977179
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1649977179
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1649977179
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1649977179
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1649977179
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1649977179
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1649977179
transform 1 0 52624 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1649977179
transform 1 0 57776 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1649977179
transform 1 0 62928 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1649977179
transform 1 0 68080 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1649977179
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1649977179
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1649977179
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1649977179
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1649977179
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1649977179
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1649977179
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1649977179
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1649977179
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1649977179
transform 1 0 50048 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1649977179
transform 1 0 55200 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1649977179
transform 1 0 60352 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1649977179
transform 1 0 65504 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1649977179
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1649977179
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1649977179
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1649977179
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1649977179
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1649977179
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1649977179
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1649977179
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1649977179
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1649977179
transform 1 0 52624 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1649977179
transform 1 0 57776 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1649977179
transform 1 0 62928 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1649977179
transform 1 0 68080 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1649977179
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1649977179
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1649977179
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1649977179
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1649977179
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1649977179
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1649977179
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1649977179
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1649977179
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1649977179
transform 1 0 50048 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1649977179
transform 1 0 55200 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1649977179
transform 1 0 60352 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1649977179
transform 1 0 65504 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1649977179
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1649977179
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1649977179
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1649977179
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1649977179
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1649977179
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1649977179
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1649977179
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1649977179
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1649977179
transform 1 0 52624 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1649977179
transform 1 0 57776 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1649977179
transform 1 0 62928 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1649977179
transform 1 0 68080 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1649977179
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1649977179
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1649977179
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1649977179
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1649977179
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1649977179
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1649977179
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1649977179
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1649977179
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1649977179
transform 1 0 50048 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1649977179
transform 1 0 55200 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1649977179
transform 1 0 60352 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1649977179
transform 1 0 65504 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1649977179
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1649977179
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1649977179
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1649977179
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1649977179
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1649977179
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1649977179
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1649977179
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1649977179
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1649977179
transform 1 0 52624 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1649977179
transform 1 0 57776 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1649977179
transform 1 0 62928 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1649977179
transform 1 0 68080 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1649977179
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1649977179
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1649977179
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1649977179
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1649977179
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1649977179
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1649977179
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1649977179
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1649977179
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1649977179
transform 1 0 50048 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1649977179
transform 1 0 55200 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1649977179
transform 1 0 60352 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1649977179
transform 1 0 65504 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1649977179
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1649977179
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1649977179
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1649977179
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1649977179
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1649977179
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1649977179
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1649977179
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1649977179
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1649977179
transform 1 0 52624 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1649977179
transform 1 0 57776 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1649977179
transform 1 0 62928 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1649977179
transform 1 0 68080 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1649977179
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1649977179
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1649977179
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1649977179
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1649977179
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1649977179
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1649977179
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1649977179
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1649977179
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1649977179
transform 1 0 50048 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1649977179
transform 1 0 55200 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1649977179
transform 1 0 60352 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1649977179
transform 1 0 65504 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1649977179
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1649977179
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1649977179
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1649977179
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1649977179
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1649977179
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1649977179
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1649977179
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1649977179
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1649977179
transform 1 0 52624 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1649977179
transform 1 0 57776 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1649977179
transform 1 0 62928 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1649977179
transform 1 0 68080 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1649977179
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1649977179
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1649977179
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1649977179
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1649977179
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1649977179
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1649977179
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1649977179
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1649977179
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1649977179
transform 1 0 50048 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1649977179
transform 1 0 55200 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1649977179
transform 1 0 60352 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1649977179
transform 1 0 65504 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1649977179
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1649977179
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1649977179
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1649977179
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1649977179
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1649977179
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1649977179
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1649977179
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1649977179
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1649977179
transform 1 0 52624 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1649977179
transform 1 0 57776 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1649977179
transform 1 0 62928 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1649977179
transform 1 0 68080 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1649977179
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1649977179
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1649977179
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1649977179
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1649977179
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1649977179
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1649977179
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1649977179
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1649977179
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1649977179
transform 1 0 50048 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1649977179
transform 1 0 55200 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1649977179
transform 1 0 60352 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1649977179
transform 1 0 65504 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1649977179
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1649977179
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1649977179
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1649977179
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1649977179
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1649977179
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1649977179
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1649977179
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1649977179
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1649977179
transform 1 0 52624 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1649977179
transform 1 0 57776 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1649977179
transform 1 0 62928 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1649977179
transform 1 0 68080 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1649977179
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1649977179
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1649977179
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1649977179
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1649977179
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1649977179
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1649977179
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1649977179
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1649977179
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1649977179
transform 1 0 50048 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1649977179
transform 1 0 55200 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1649977179
transform 1 0 60352 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1649977179
transform 1 0 65504 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1649977179
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1649977179
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1649977179
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1649977179
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1649977179
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1649977179
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1649977179
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1649977179
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1649977179
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1649977179
transform 1 0 52624 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1649977179
transform 1 0 57776 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1649977179
transform 1 0 62928 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1649977179
transform 1 0 68080 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1649977179
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1649977179
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1649977179
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1649977179
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1649977179
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1649977179
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1649977179
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1649977179
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1649977179
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1649977179
transform 1 0 50048 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1649977179
transform 1 0 55200 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1649977179
transform 1 0 60352 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1649977179
transform 1 0 65504 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1649977179
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1649977179
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1649977179
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1649977179
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1649977179
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1649977179
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1649977179
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1649977179
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1649977179
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1649977179
transform 1 0 52624 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1649977179
transform 1 0 57776 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1649977179
transform 1 0 62928 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1649977179
transform 1 0 68080 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1649977179
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1649977179
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1649977179
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1649977179
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1649977179
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1649977179
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1649977179
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1649977179
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1649977179
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1649977179
transform 1 0 50048 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1649977179
transform 1 0 55200 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1649977179
transform 1 0 60352 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1649977179
transform 1 0 65504 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1649977179
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1649977179
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1649977179
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1649977179
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1649977179
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1649977179
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1649977179
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1649977179
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1649977179
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1649977179
transform 1 0 52624 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1649977179
transform 1 0 57776 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1649977179
transform 1 0 62928 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1649977179
transform 1 0 68080 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1649977179
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1649977179
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1649977179
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1649977179
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1649977179
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1649977179
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1649977179
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1649977179
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1649977179
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1649977179
transform 1 0 50048 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1649977179
transform 1 0 55200 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1649977179
transform 1 0 60352 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1649977179
transform 1 0 65504 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1649977179
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1649977179
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1649977179
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1649977179
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1649977179
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1649977179
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1649977179
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1649977179
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1649977179
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1649977179
transform 1 0 52624 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1649977179
transform 1 0 57776 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1649977179
transform 1 0 62928 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1649977179
transform 1 0 68080 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1649977179
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1649977179
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1649977179
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1649977179
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1649977179
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1649977179
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1649977179
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1649977179
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1649977179
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1649977179
transform 1 0 50048 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1649977179
transform 1 0 55200 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1649977179
transform 1 0 60352 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1649977179
transform 1 0 65504 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1649977179
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1649977179
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1649977179
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1649977179
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1649977179
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1649977179
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1649977179
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1649977179
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1649977179
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1649977179
transform 1 0 52624 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1649977179
transform 1 0 57776 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1649977179
transform 1 0 62928 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1649977179
transform 1 0 68080 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1649977179
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1649977179
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1649977179
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1649977179
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1649977179
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1649977179
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1649977179
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1649977179
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1649977179
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1649977179
transform 1 0 50048 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1649977179
transform 1 0 55200 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1649977179
transform 1 0 60352 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1649977179
transform 1 0 65504 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1649977179
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1649977179
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1649977179
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1649977179
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1649977179
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1649977179
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1649977179
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1649977179
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1649977179
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1649977179
transform 1 0 52624 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1649977179
transform 1 0 57776 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1649977179
transform 1 0 62928 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1649977179
transform 1 0 68080 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1649977179
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1649977179
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1649977179
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1649977179
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1649977179
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1649977179
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1649977179
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1649977179
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1649977179
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1649977179
transform 1 0 50048 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1649977179
transform 1 0 55200 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1649977179
transform 1 0 60352 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1649977179
transform 1 0 65504 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1649977179
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1649977179
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1649977179
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1649977179
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1649977179
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1649977179
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1649977179
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1649977179
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1649977179
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1649977179
transform 1 0 52624 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1649977179
transform 1 0 57776 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1649977179
transform 1 0 62928 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1649977179
transform 1 0 68080 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1649977179
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1649977179
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1649977179
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1649977179
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1649977179
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1649977179
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1649977179
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1649977179
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1649977179
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1649977179
transform 1 0 50048 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1649977179
transform 1 0 55200 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1649977179
transform 1 0 60352 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1649977179
transform 1 0 65504 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1649977179
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1649977179
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1649977179
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1649977179
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1649977179
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1649977179
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1649977179
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1649977179
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1649977179
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1649977179
transform 1 0 52624 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1649977179
transform 1 0 57776 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1649977179
transform 1 0 62928 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1649977179
transform 1 0 68080 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1649977179
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1649977179
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1649977179
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1649977179
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1649977179
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1649977179
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1649977179
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1649977179
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1649977179
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1649977179
transform 1 0 50048 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1649977179
transform 1 0 55200 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1649977179
transform 1 0 60352 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1649977179
transform 1 0 65504 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1649977179
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1649977179
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1649977179
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1649977179
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1649977179
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1649977179
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1649977179
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1649977179
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1649977179
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1649977179
transform 1 0 52624 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1649977179
transform 1 0 57776 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1649977179
transform 1 0 62928 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1649977179
transform 1 0 68080 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1649977179
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1649977179
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1649977179
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1649977179
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1649977179
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1649977179
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1649977179
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1649977179
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1649977179
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1649977179
transform 1 0 50048 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1649977179
transform 1 0 55200 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1649977179
transform 1 0 60352 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1649977179
transform 1 0 65504 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1649977179
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1649977179
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1649977179
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1649977179
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1649977179
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1649977179
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1649977179
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1649977179
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1649977179
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1649977179
transform 1 0 52624 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1649977179
transform 1 0 57776 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1649977179
transform 1 0 62928 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1649977179
transform 1 0 68080 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1649977179
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1649977179
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1649977179
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1649977179
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1649977179
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1649977179
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1649977179
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1649977179
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1649977179
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1649977179
transform 1 0 50048 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1649977179
transform 1 0 55200 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1649977179
transform 1 0 60352 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1649977179
transform 1 0 65504 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1649977179
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1649977179
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1649977179
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1649977179
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1649977179
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1649977179
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1649977179
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1649977179
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1649977179
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1649977179
transform 1 0 52624 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1649977179
transform 1 0 57776 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1649977179
transform 1 0 62928 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1649977179
transform 1 0 68080 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1649977179
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1649977179
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1649977179
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1649977179
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1649977179
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1649977179
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1649977179
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1649977179
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1649977179
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1649977179
transform 1 0 50048 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1649977179
transform 1 0 55200 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1649977179
transform 1 0 60352 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1649977179
transform 1 0 65504 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1649977179
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1649977179
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1649977179
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1649977179
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1649977179
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1649977179
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1649977179
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1649977179
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1649977179
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1649977179
transform 1 0 52624 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1649977179
transform 1 0 57776 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1649977179
transform 1 0 62928 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1649977179
transform 1 0 68080 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1649977179
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1649977179
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1649977179
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1649977179
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1649977179
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1649977179
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1649977179
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1649977179
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1649977179
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1649977179
transform 1 0 50048 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1649977179
transform 1 0 55200 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1649977179
transform 1 0 60352 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1649977179
transform 1 0 65504 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1649977179
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1649977179
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1649977179
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1649977179
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1649977179
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1649977179
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1649977179
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1649977179
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1649977179
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1649977179
transform 1 0 52624 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1649977179
transform 1 0 57776 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1649977179
transform 1 0 62928 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1649977179
transform 1 0 68080 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1649977179
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1649977179
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1649977179
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1649977179
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1649977179
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1649977179
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1649977179
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1649977179
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1649977179
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1649977179
transform 1 0 50048 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1649977179
transform 1 0 55200 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1649977179
transform 1 0 60352 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1649977179
transform 1 0 65504 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1649977179
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1649977179
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1649977179
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1649977179
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1649977179
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1649977179
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1649977179
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1649977179
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1649977179
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1649977179
transform 1 0 52624 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1649977179
transform 1 0 57776 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1649977179
transform 1 0 62928 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1649977179
transform 1 0 68080 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1649977179
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1649977179
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1649977179
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1649977179
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1649977179
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1649977179
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1649977179
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1649977179
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1649977179
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1649977179
transform 1 0 50048 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1649977179
transform 1 0 55200 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1649977179
transform 1 0 60352 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1649977179
transform 1 0 65504 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1649977179
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1649977179
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1649977179
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1649977179
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1649977179
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1649977179
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1649977179
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1649977179
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1649977179
transform 1 0 47472 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1649977179
transform 1 0 52624 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1649977179
transform 1 0 57776 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1649977179
transform 1 0 62928 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1649977179
transform 1 0 68080 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1649977179
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1649977179
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1649977179
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1649977179
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1649977179
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1649977179
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1649977179
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1649977179
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1649977179
transform 1 0 44896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1649977179
transform 1 0 50048 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1649977179
transform 1 0 55200 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1649977179
transform 1 0 60352 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1649977179
transform 1 0 65504 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1649977179
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1649977179
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1649977179
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1649977179
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1649977179
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1649977179
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1649977179
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1649977179
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1649977179
transform 1 0 47472 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1649977179
transform 1 0 52624 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1649977179
transform 1 0 57776 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1649977179
transform 1 0 62928 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1649977179
transform 1 0 68080 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1649977179
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1649977179
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1649977179
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1649977179
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1649977179
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1649977179
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1649977179
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1649977179
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1649977179
transform 1 0 44896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1649977179
transform 1 0 50048 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1649977179
transform 1 0 55200 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1649977179
transform 1 0 60352 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1649977179
transform 1 0 65504 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1649977179
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1649977179
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1649977179
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1649977179
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1649977179
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1649977179
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1649977179
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1649977179
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1649977179
transform 1 0 47472 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1649977179
transform 1 0 52624 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1649977179
transform 1 0 57776 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1649977179
transform 1 0 62928 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1649977179
transform 1 0 68080 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1649977179
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1649977179
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1649977179
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1649977179
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1649977179
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1649977179
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1649977179
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1649977179
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1649977179
transform 1 0 44896 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1649977179
transform 1 0 50048 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1649977179
transform 1 0 55200 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1649977179
transform 1 0 60352 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1649977179
transform 1 0 65504 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1649977179
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1649977179
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1649977179
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1649977179
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1649977179
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1649977179
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1649977179
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1649977179
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1649977179
transform 1 0 47472 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1649977179
transform 1 0 52624 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1649977179
transform 1 0 57776 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1649977179
transform 1 0 62928 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1649977179
transform 1 0 68080 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_919
timestamp 1649977179
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_920
timestamp 1649977179
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_921
timestamp 1649977179
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_922
timestamp 1649977179
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_923
timestamp 1649977179
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_924
timestamp 1649977179
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_925
timestamp 1649977179
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_926
timestamp 1649977179
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_927
timestamp 1649977179
transform 1 0 44896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_928
timestamp 1649977179
transform 1 0 50048 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_929
timestamp 1649977179
transform 1 0 55200 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_930
timestamp 1649977179
transform 1 0 60352 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_931
timestamp 1649977179
transform 1 0 65504 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_932
timestamp 1649977179
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_933
timestamp 1649977179
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_934
timestamp 1649977179
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_935
timestamp 1649977179
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_936
timestamp 1649977179
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_937
timestamp 1649977179
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_938
timestamp 1649977179
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_939
timestamp 1649977179
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_940
timestamp 1649977179
transform 1 0 47472 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_941
timestamp 1649977179
transform 1 0 52624 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_942
timestamp 1649977179
transform 1 0 57776 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_943
timestamp 1649977179
transform 1 0 62928 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_944
timestamp 1649977179
transform 1 0 68080 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_945
timestamp 1649977179
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_946
timestamp 1649977179
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_947
timestamp 1649977179
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_948
timestamp 1649977179
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_949
timestamp 1649977179
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_950
timestamp 1649977179
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_951
timestamp 1649977179
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_952
timestamp 1649977179
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_953
timestamp 1649977179
transform 1 0 44896 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_954
timestamp 1649977179
transform 1 0 50048 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_955
timestamp 1649977179
transform 1 0 55200 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_956
timestamp 1649977179
transform 1 0 60352 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_957
timestamp 1649977179
transform 1 0 65504 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_958
timestamp 1649977179
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_959
timestamp 1649977179
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_960
timestamp 1649977179
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_961
timestamp 1649977179
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_962
timestamp 1649977179
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_963
timestamp 1649977179
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_964
timestamp 1649977179
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_965
timestamp 1649977179
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_966
timestamp 1649977179
transform 1 0 47472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_967
timestamp 1649977179
transform 1 0 52624 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_968
timestamp 1649977179
transform 1 0 57776 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_969
timestamp 1649977179
transform 1 0 62928 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_970
timestamp 1649977179
transform 1 0 68080 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_971
timestamp 1649977179
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_972
timestamp 1649977179
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_973
timestamp 1649977179
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_974
timestamp 1649977179
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_975
timestamp 1649977179
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_976
timestamp 1649977179
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_977
timestamp 1649977179
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_978
timestamp 1649977179
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_979
timestamp 1649977179
transform 1 0 44896 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_980
timestamp 1649977179
transform 1 0 50048 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_981
timestamp 1649977179
transform 1 0 55200 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_982
timestamp 1649977179
transform 1 0 60352 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_983
timestamp 1649977179
transform 1 0 65504 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_984
timestamp 1649977179
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_985
timestamp 1649977179
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_986
timestamp 1649977179
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_987
timestamp 1649977179
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_988
timestamp 1649977179
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_989
timestamp 1649977179
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_990
timestamp 1649977179
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_991
timestamp 1649977179
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_992
timestamp 1649977179
transform 1 0 47472 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_993
timestamp 1649977179
transform 1 0 52624 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_994
timestamp 1649977179
transform 1 0 57776 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_995
timestamp 1649977179
transform 1 0 62928 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_996
timestamp 1649977179
transform 1 0 68080 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_997
timestamp 1649977179
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_998
timestamp 1649977179
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_999
timestamp 1649977179
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1000
timestamp 1649977179
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1001
timestamp 1649977179
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1002
timestamp 1649977179
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1003
timestamp 1649977179
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1004
timestamp 1649977179
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1005
timestamp 1649977179
transform 1 0 44896 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1006
timestamp 1649977179
transform 1 0 50048 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1007
timestamp 1649977179
transform 1 0 55200 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1008
timestamp 1649977179
transform 1 0 60352 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1009
timestamp 1649977179
transform 1 0 65504 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1010
timestamp 1649977179
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1011
timestamp 1649977179
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1012
timestamp 1649977179
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1013
timestamp 1649977179
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1014
timestamp 1649977179
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1015
timestamp 1649977179
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1016
timestamp 1649977179
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1017
timestamp 1649977179
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1018
timestamp 1649977179
transform 1 0 47472 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1019
timestamp 1649977179
transform 1 0 52624 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1020
timestamp 1649977179
transform 1 0 57776 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1021
timestamp 1649977179
transform 1 0 62928 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1022
timestamp 1649977179
transform 1 0 68080 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1023
timestamp 1649977179
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1024
timestamp 1649977179
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1025
timestamp 1649977179
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1026
timestamp 1649977179
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1027
timestamp 1649977179
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1028
timestamp 1649977179
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1029
timestamp 1649977179
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1030
timestamp 1649977179
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1031
timestamp 1649977179
transform 1 0 44896 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1032
timestamp 1649977179
transform 1 0 50048 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1033
timestamp 1649977179
transform 1 0 55200 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1034
timestamp 1649977179
transform 1 0 60352 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1035
timestamp 1649977179
transform 1 0 65504 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1036
timestamp 1649977179
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1037
timestamp 1649977179
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1038
timestamp 1649977179
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1039
timestamp 1649977179
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1040
timestamp 1649977179
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1041
timestamp 1649977179
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1042
timestamp 1649977179
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1043
timestamp 1649977179
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1044
timestamp 1649977179
transform 1 0 47472 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1045
timestamp 1649977179
transform 1 0 52624 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1046
timestamp 1649977179
transform 1 0 57776 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1047
timestamp 1649977179
transform 1 0 62928 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1048
timestamp 1649977179
transform 1 0 68080 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1049
timestamp 1649977179
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1050
timestamp 1649977179
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1051
timestamp 1649977179
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1052
timestamp 1649977179
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1053
timestamp 1649977179
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1054
timestamp 1649977179
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1055
timestamp 1649977179
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1056
timestamp 1649977179
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1057
timestamp 1649977179
transform 1 0 44896 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1058
timestamp 1649977179
transform 1 0 50048 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1059
timestamp 1649977179
transform 1 0 55200 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1060
timestamp 1649977179
transform 1 0 60352 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1061
timestamp 1649977179
transform 1 0 65504 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1062
timestamp 1649977179
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1063
timestamp 1649977179
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1064
timestamp 1649977179
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1065
timestamp 1649977179
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1066
timestamp 1649977179
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1067
timestamp 1649977179
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1068
timestamp 1649977179
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1069
timestamp 1649977179
transform 1 0 42320 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1070
timestamp 1649977179
transform 1 0 47472 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1071
timestamp 1649977179
transform 1 0 52624 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1072
timestamp 1649977179
transform 1 0 57776 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1073
timestamp 1649977179
transform 1 0 62928 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1074
timestamp 1649977179
transform 1 0 68080 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1075
timestamp 1649977179
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1076
timestamp 1649977179
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1077
timestamp 1649977179
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1078
timestamp 1649977179
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1079
timestamp 1649977179
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1080
timestamp 1649977179
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1081
timestamp 1649977179
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1082
timestamp 1649977179
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1083
timestamp 1649977179
transform 1 0 44896 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1084
timestamp 1649977179
transform 1 0 50048 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1085
timestamp 1649977179
transform 1 0 55200 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1086
timestamp 1649977179
transform 1 0 60352 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1087
timestamp 1649977179
transform 1 0 65504 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1088
timestamp 1649977179
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1089
timestamp 1649977179
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1090
timestamp 1649977179
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1091
timestamp 1649977179
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1092
timestamp 1649977179
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1093
timestamp 1649977179
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1094
timestamp 1649977179
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1095
timestamp 1649977179
transform 1 0 42320 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1096
timestamp 1649977179
transform 1 0 47472 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1097
timestamp 1649977179
transform 1 0 52624 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1098
timestamp 1649977179
transform 1 0 57776 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1099
timestamp 1649977179
transform 1 0 62928 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1100
timestamp 1649977179
transform 1 0 68080 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1101
timestamp 1649977179
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1102
timestamp 1649977179
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1103
timestamp 1649977179
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1104
timestamp 1649977179
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1105
timestamp 1649977179
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1106
timestamp 1649977179
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1107
timestamp 1649977179
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1108
timestamp 1649977179
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1109
timestamp 1649977179
transform 1 0 44896 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1110
timestamp 1649977179
transform 1 0 50048 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1111
timestamp 1649977179
transform 1 0 55200 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1112
timestamp 1649977179
transform 1 0 60352 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1113
timestamp 1649977179
transform 1 0 65504 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1114
timestamp 1649977179
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1115
timestamp 1649977179
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1116
timestamp 1649977179
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1117
timestamp 1649977179
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1118
timestamp 1649977179
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1119
timestamp 1649977179
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1120
timestamp 1649977179
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1121
timestamp 1649977179
transform 1 0 42320 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1122
timestamp 1649977179
transform 1 0 47472 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1123
timestamp 1649977179
transform 1 0 52624 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1124
timestamp 1649977179
transform 1 0 57776 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1125
timestamp 1649977179
transform 1 0 62928 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1126
timestamp 1649977179
transform 1 0 68080 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1127
timestamp 1649977179
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1128
timestamp 1649977179
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1129
timestamp 1649977179
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1130
timestamp 1649977179
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1131
timestamp 1649977179
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1132
timestamp 1649977179
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1133
timestamp 1649977179
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1134
timestamp 1649977179
transform 1 0 39744 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1135
timestamp 1649977179
transform 1 0 44896 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1136
timestamp 1649977179
transform 1 0 50048 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1137
timestamp 1649977179
transform 1 0 55200 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1138
timestamp 1649977179
transform 1 0 60352 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1139
timestamp 1649977179
transform 1 0 65504 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1140
timestamp 1649977179
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1141
timestamp 1649977179
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1142
timestamp 1649977179
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1143
timestamp 1649977179
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1144
timestamp 1649977179
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1145
timestamp 1649977179
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1146
timestamp 1649977179
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1147
timestamp 1649977179
transform 1 0 42320 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1148
timestamp 1649977179
transform 1 0 47472 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1149
timestamp 1649977179
transform 1 0 52624 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1150
timestamp 1649977179
transform 1 0 57776 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1151
timestamp 1649977179
transform 1 0 62928 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1152
timestamp 1649977179
transform 1 0 68080 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1153
timestamp 1649977179
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1154
timestamp 1649977179
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1155
timestamp 1649977179
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1156
timestamp 1649977179
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1157
timestamp 1649977179
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1158
timestamp 1649977179
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1159
timestamp 1649977179
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1160
timestamp 1649977179
transform 1 0 39744 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1161
timestamp 1649977179
transform 1 0 44896 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1162
timestamp 1649977179
transform 1 0 50048 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1163
timestamp 1649977179
transform 1 0 55200 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1164
timestamp 1649977179
transform 1 0 60352 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1165
timestamp 1649977179
transform 1 0 65504 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1166
timestamp 1649977179
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1167
timestamp 1649977179
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1168
timestamp 1649977179
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1169
timestamp 1649977179
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1170
timestamp 1649977179
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1171
timestamp 1649977179
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1172
timestamp 1649977179
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1173
timestamp 1649977179
transform 1 0 42320 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1174
timestamp 1649977179
transform 1 0 47472 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1175
timestamp 1649977179
transform 1 0 52624 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1176
timestamp 1649977179
transform 1 0 57776 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1177
timestamp 1649977179
transform 1 0 62928 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1178
timestamp 1649977179
transform 1 0 68080 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1179
timestamp 1649977179
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1180
timestamp 1649977179
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1181
timestamp 1649977179
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1182
timestamp 1649977179
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1183
timestamp 1649977179
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1184
timestamp 1649977179
transform 1 0 29440 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1185
timestamp 1649977179
transform 1 0 34592 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1186
timestamp 1649977179
transform 1 0 39744 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1187
timestamp 1649977179
transform 1 0 44896 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1188
timestamp 1649977179
transform 1 0 50048 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1189
timestamp 1649977179
transform 1 0 55200 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1190
timestamp 1649977179
transform 1 0 60352 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1191
timestamp 1649977179
transform 1 0 65504 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1192
timestamp 1649977179
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1193
timestamp 1649977179
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1194
timestamp 1649977179
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1195
timestamp 1649977179
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1196
timestamp 1649977179
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1197
timestamp 1649977179
transform 1 0 32016 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1198
timestamp 1649977179
transform 1 0 37168 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1199
timestamp 1649977179
transform 1 0 42320 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1200
timestamp 1649977179
transform 1 0 47472 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1201
timestamp 1649977179
transform 1 0 52624 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1202
timestamp 1649977179
transform 1 0 57776 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1203
timestamp 1649977179
transform 1 0 62928 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1204
timestamp 1649977179
transform 1 0 68080 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1205
timestamp 1649977179
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1206
timestamp 1649977179
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1207
timestamp 1649977179
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1208
timestamp 1649977179
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1209
timestamp 1649977179
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1210
timestamp 1649977179
transform 1 0 29440 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1211
timestamp 1649977179
transform 1 0 34592 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1212
timestamp 1649977179
transform 1 0 39744 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1213
timestamp 1649977179
transform 1 0 44896 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1214
timestamp 1649977179
transform 1 0 50048 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1215
timestamp 1649977179
transform 1 0 55200 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1216
timestamp 1649977179
transform 1 0 60352 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1217
timestamp 1649977179
transform 1 0 65504 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1218
timestamp 1649977179
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1219
timestamp 1649977179
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1220
timestamp 1649977179
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1221
timestamp 1649977179
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1222
timestamp 1649977179
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1223
timestamp 1649977179
transform 1 0 32016 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1224
timestamp 1649977179
transform 1 0 37168 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1225
timestamp 1649977179
transform 1 0 42320 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1226
timestamp 1649977179
transform 1 0 47472 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1227
timestamp 1649977179
transform 1 0 52624 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1228
timestamp 1649977179
transform 1 0 57776 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1229
timestamp 1649977179
transform 1 0 62928 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1230
timestamp 1649977179
transform 1 0 68080 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1231
timestamp 1649977179
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1232
timestamp 1649977179
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1233
timestamp 1649977179
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1234
timestamp 1649977179
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1235
timestamp 1649977179
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1236
timestamp 1649977179
transform 1 0 29440 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1237
timestamp 1649977179
transform 1 0 34592 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1238
timestamp 1649977179
transform 1 0 39744 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1239
timestamp 1649977179
transform 1 0 44896 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1240
timestamp 1649977179
transform 1 0 50048 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1241
timestamp 1649977179
transform 1 0 55200 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1242
timestamp 1649977179
transform 1 0 60352 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1243
timestamp 1649977179
transform 1 0 65504 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1244
timestamp 1649977179
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1245
timestamp 1649977179
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1246
timestamp 1649977179
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1247
timestamp 1649977179
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1248
timestamp 1649977179
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1249
timestamp 1649977179
transform 1 0 32016 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1250
timestamp 1649977179
transform 1 0 37168 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1251
timestamp 1649977179
transform 1 0 42320 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1252
timestamp 1649977179
transform 1 0 47472 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1253
timestamp 1649977179
transform 1 0 52624 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1254
timestamp 1649977179
transform 1 0 57776 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1255
timestamp 1649977179
transform 1 0 62928 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1256
timestamp 1649977179
transform 1 0 68080 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1257
timestamp 1649977179
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1258
timestamp 1649977179
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1259
timestamp 1649977179
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1260
timestamp 1649977179
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1261
timestamp 1649977179
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1262
timestamp 1649977179
transform 1 0 29440 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1263
timestamp 1649977179
transform 1 0 34592 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1264
timestamp 1649977179
transform 1 0 39744 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1265
timestamp 1649977179
transform 1 0 44896 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1266
timestamp 1649977179
transform 1 0 50048 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1267
timestamp 1649977179
transform 1 0 55200 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1268
timestamp 1649977179
transform 1 0 60352 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1269
timestamp 1649977179
transform 1 0 65504 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1270
timestamp 1649977179
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1271
timestamp 1649977179
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1272
timestamp 1649977179
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1273
timestamp 1649977179
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1274
timestamp 1649977179
transform 1 0 26864 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1275
timestamp 1649977179
transform 1 0 32016 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1276
timestamp 1649977179
transform 1 0 37168 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1277
timestamp 1649977179
transform 1 0 42320 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1278
timestamp 1649977179
transform 1 0 47472 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1279
timestamp 1649977179
transform 1 0 52624 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1280
timestamp 1649977179
transform 1 0 57776 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1281
timestamp 1649977179
transform 1 0 62928 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1282
timestamp 1649977179
transform 1 0 68080 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1283
timestamp 1649977179
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1284
timestamp 1649977179
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1285
timestamp 1649977179
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1286
timestamp 1649977179
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1287
timestamp 1649977179
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1288
timestamp 1649977179
transform 1 0 29440 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1289
timestamp 1649977179
transform 1 0 34592 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1290
timestamp 1649977179
transform 1 0 39744 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1291
timestamp 1649977179
transform 1 0 44896 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1292
timestamp 1649977179
transform 1 0 50048 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1293
timestamp 1649977179
transform 1 0 55200 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1294
timestamp 1649977179
transform 1 0 60352 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1295
timestamp 1649977179
transform 1 0 65504 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1296
timestamp 1649977179
transform 1 0 6256 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1297
timestamp 1649977179
transform 1 0 11408 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1298
timestamp 1649977179
transform 1 0 16560 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1299
timestamp 1649977179
transform 1 0 21712 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1300
timestamp 1649977179
transform 1 0 26864 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1301
timestamp 1649977179
transform 1 0 32016 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1302
timestamp 1649977179
transform 1 0 37168 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1303
timestamp 1649977179
transform 1 0 42320 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1304
timestamp 1649977179
transform 1 0 47472 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1305
timestamp 1649977179
transform 1 0 52624 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1306
timestamp 1649977179
transform 1 0 57776 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1307
timestamp 1649977179
transform 1 0 62928 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1308
timestamp 1649977179
transform 1 0 68080 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1309
timestamp 1649977179
transform 1 0 3680 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1310
timestamp 1649977179
transform 1 0 8832 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1311
timestamp 1649977179
transform 1 0 13984 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1312
timestamp 1649977179
transform 1 0 19136 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1313
timestamp 1649977179
transform 1 0 24288 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1314
timestamp 1649977179
transform 1 0 29440 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1315
timestamp 1649977179
transform 1 0 34592 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1316
timestamp 1649977179
transform 1 0 39744 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1317
timestamp 1649977179
transform 1 0 44896 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1318
timestamp 1649977179
transform 1 0 50048 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1319
timestamp 1649977179
transform 1 0 55200 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1320
timestamp 1649977179
transform 1 0 60352 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1321
timestamp 1649977179
transform 1 0 65504 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1322
timestamp 1649977179
transform 1 0 6256 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1323
timestamp 1649977179
transform 1 0 11408 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1324
timestamp 1649977179
transform 1 0 16560 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1325
timestamp 1649977179
transform 1 0 21712 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1326
timestamp 1649977179
transform 1 0 26864 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1327
timestamp 1649977179
transform 1 0 32016 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1328
timestamp 1649977179
transform 1 0 37168 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1329
timestamp 1649977179
transform 1 0 42320 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1330
timestamp 1649977179
transform 1 0 47472 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1331
timestamp 1649977179
transform 1 0 52624 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1332
timestamp 1649977179
transform 1 0 57776 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1333
timestamp 1649977179
transform 1 0 62928 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1334
timestamp 1649977179
transform 1 0 68080 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1335
timestamp 1649977179
transform 1 0 3680 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1336
timestamp 1649977179
transform 1 0 8832 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1337
timestamp 1649977179
transform 1 0 13984 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1338
timestamp 1649977179
transform 1 0 19136 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1339
timestamp 1649977179
transform 1 0 24288 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1340
timestamp 1649977179
transform 1 0 29440 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1341
timestamp 1649977179
transform 1 0 34592 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1342
timestamp 1649977179
transform 1 0 39744 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1343
timestamp 1649977179
transform 1 0 44896 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1344
timestamp 1649977179
transform 1 0 50048 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1345
timestamp 1649977179
transform 1 0 55200 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1346
timestamp 1649977179
transform 1 0 60352 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1347
timestamp 1649977179
transform 1 0 65504 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1348
timestamp 1649977179
transform 1 0 6256 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1349
timestamp 1649977179
transform 1 0 11408 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1350
timestamp 1649977179
transform 1 0 16560 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1351
timestamp 1649977179
transform 1 0 21712 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1352
timestamp 1649977179
transform 1 0 26864 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1353
timestamp 1649977179
transform 1 0 32016 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1354
timestamp 1649977179
transform 1 0 37168 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1355
timestamp 1649977179
transform 1 0 42320 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1356
timestamp 1649977179
transform 1 0 47472 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1357
timestamp 1649977179
transform 1 0 52624 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1358
timestamp 1649977179
transform 1 0 57776 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1359
timestamp 1649977179
transform 1 0 62928 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1360
timestamp 1649977179
transform 1 0 68080 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1361
timestamp 1649977179
transform 1 0 3680 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1362
timestamp 1649977179
transform 1 0 8832 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1363
timestamp 1649977179
transform 1 0 13984 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1364
timestamp 1649977179
transform 1 0 19136 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1365
timestamp 1649977179
transform 1 0 24288 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1366
timestamp 1649977179
transform 1 0 29440 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1367
timestamp 1649977179
transform 1 0 34592 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1368
timestamp 1649977179
transform 1 0 39744 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1369
timestamp 1649977179
transform 1 0 44896 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1370
timestamp 1649977179
transform 1 0 50048 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1371
timestamp 1649977179
transform 1 0 55200 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1372
timestamp 1649977179
transform 1 0 60352 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1373
timestamp 1649977179
transform 1 0 65504 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1374
timestamp 1649977179
transform 1 0 6256 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1375
timestamp 1649977179
transform 1 0 11408 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1376
timestamp 1649977179
transform 1 0 16560 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1377
timestamp 1649977179
transform 1 0 21712 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1378
timestamp 1649977179
transform 1 0 26864 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1379
timestamp 1649977179
transform 1 0 32016 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1380
timestamp 1649977179
transform 1 0 37168 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1381
timestamp 1649977179
transform 1 0 42320 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1382
timestamp 1649977179
transform 1 0 47472 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1383
timestamp 1649977179
transform 1 0 52624 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1384
timestamp 1649977179
transform 1 0 57776 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1385
timestamp 1649977179
transform 1 0 62928 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1386
timestamp 1649977179
transform 1 0 68080 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1387
timestamp 1649977179
transform 1 0 3680 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1388
timestamp 1649977179
transform 1 0 8832 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1389
timestamp 1649977179
transform 1 0 13984 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1390
timestamp 1649977179
transform 1 0 19136 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1391
timestamp 1649977179
transform 1 0 24288 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1392
timestamp 1649977179
transform 1 0 29440 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1393
timestamp 1649977179
transform 1 0 34592 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1394
timestamp 1649977179
transform 1 0 39744 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1395
timestamp 1649977179
transform 1 0 44896 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1396
timestamp 1649977179
transform 1 0 50048 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1397
timestamp 1649977179
transform 1 0 55200 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1398
timestamp 1649977179
transform 1 0 60352 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1399
timestamp 1649977179
transform 1 0 65504 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1400
timestamp 1649977179
transform 1 0 6256 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1401
timestamp 1649977179
transform 1 0 11408 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1402
timestamp 1649977179
transform 1 0 16560 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1403
timestamp 1649977179
transform 1 0 21712 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1404
timestamp 1649977179
transform 1 0 26864 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1405
timestamp 1649977179
transform 1 0 32016 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1406
timestamp 1649977179
transform 1 0 37168 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1407
timestamp 1649977179
transform 1 0 42320 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1408
timestamp 1649977179
transform 1 0 47472 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1409
timestamp 1649977179
transform 1 0 52624 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1410
timestamp 1649977179
transform 1 0 57776 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1411
timestamp 1649977179
transform 1 0 62928 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1412
timestamp 1649977179
transform 1 0 68080 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1413
timestamp 1649977179
transform 1 0 3680 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1414
timestamp 1649977179
transform 1 0 8832 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1415
timestamp 1649977179
transform 1 0 13984 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1416
timestamp 1649977179
transform 1 0 19136 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1417
timestamp 1649977179
transform 1 0 24288 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1418
timestamp 1649977179
transform 1 0 29440 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1419
timestamp 1649977179
transform 1 0 34592 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1420
timestamp 1649977179
transform 1 0 39744 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1421
timestamp 1649977179
transform 1 0 44896 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1422
timestamp 1649977179
transform 1 0 50048 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1423
timestamp 1649977179
transform 1 0 55200 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1424
timestamp 1649977179
transform 1 0 60352 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1425
timestamp 1649977179
transform 1 0 65504 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1426
timestamp 1649977179
transform 1 0 6256 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1427
timestamp 1649977179
transform 1 0 11408 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1428
timestamp 1649977179
transform 1 0 16560 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1429
timestamp 1649977179
transform 1 0 21712 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1430
timestamp 1649977179
transform 1 0 26864 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1431
timestamp 1649977179
transform 1 0 32016 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1432
timestamp 1649977179
transform 1 0 37168 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1433
timestamp 1649977179
transform 1 0 42320 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1434
timestamp 1649977179
transform 1 0 47472 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1435
timestamp 1649977179
transform 1 0 52624 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1436
timestamp 1649977179
transform 1 0 57776 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1437
timestamp 1649977179
transform 1 0 62928 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1438
timestamp 1649977179
transform 1 0 68080 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1439
timestamp 1649977179
transform 1 0 3680 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1440
timestamp 1649977179
transform 1 0 8832 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1441
timestamp 1649977179
transform 1 0 13984 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1442
timestamp 1649977179
transform 1 0 19136 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1443
timestamp 1649977179
transform 1 0 24288 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1444
timestamp 1649977179
transform 1 0 29440 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1445
timestamp 1649977179
transform 1 0 34592 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1446
timestamp 1649977179
transform 1 0 39744 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1447
timestamp 1649977179
transform 1 0 44896 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1448
timestamp 1649977179
transform 1 0 50048 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1449
timestamp 1649977179
transform 1 0 55200 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1450
timestamp 1649977179
transform 1 0 60352 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1451
timestamp 1649977179
transform 1 0 65504 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1452
timestamp 1649977179
transform 1 0 6256 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1453
timestamp 1649977179
transform 1 0 11408 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1454
timestamp 1649977179
transform 1 0 16560 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1455
timestamp 1649977179
transform 1 0 21712 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1456
timestamp 1649977179
transform 1 0 26864 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1457
timestamp 1649977179
transform 1 0 32016 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1458
timestamp 1649977179
transform 1 0 37168 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1459
timestamp 1649977179
transform 1 0 42320 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1460
timestamp 1649977179
transform 1 0 47472 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1461
timestamp 1649977179
transform 1 0 52624 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1462
timestamp 1649977179
transform 1 0 57776 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1463
timestamp 1649977179
transform 1 0 62928 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1464
timestamp 1649977179
transform 1 0 68080 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1465
timestamp 1649977179
transform 1 0 3680 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1466
timestamp 1649977179
transform 1 0 8832 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1467
timestamp 1649977179
transform 1 0 13984 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1468
timestamp 1649977179
transform 1 0 19136 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1469
timestamp 1649977179
transform 1 0 24288 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1470
timestamp 1649977179
transform 1 0 29440 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1471
timestamp 1649977179
transform 1 0 34592 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1472
timestamp 1649977179
transform 1 0 39744 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1473
timestamp 1649977179
transform 1 0 44896 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1474
timestamp 1649977179
transform 1 0 50048 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1475
timestamp 1649977179
transform 1 0 55200 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1476
timestamp 1649977179
transform 1 0 60352 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1477
timestamp 1649977179
transform 1 0 65504 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1478
timestamp 1649977179
transform 1 0 6256 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1479
timestamp 1649977179
transform 1 0 11408 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1480
timestamp 1649977179
transform 1 0 16560 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1481
timestamp 1649977179
transform 1 0 21712 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1482
timestamp 1649977179
transform 1 0 26864 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1483
timestamp 1649977179
transform 1 0 32016 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1484
timestamp 1649977179
transform 1 0 37168 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1485
timestamp 1649977179
transform 1 0 42320 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1486
timestamp 1649977179
transform 1 0 47472 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1487
timestamp 1649977179
transform 1 0 52624 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1488
timestamp 1649977179
transform 1 0 57776 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1489
timestamp 1649977179
transform 1 0 62928 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1490
timestamp 1649977179
transform 1 0 68080 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1491
timestamp 1649977179
transform 1 0 3680 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1492
timestamp 1649977179
transform 1 0 8832 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1493
timestamp 1649977179
transform 1 0 13984 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1494
timestamp 1649977179
transform 1 0 19136 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1495
timestamp 1649977179
transform 1 0 24288 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1496
timestamp 1649977179
transform 1 0 29440 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1497
timestamp 1649977179
transform 1 0 34592 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1498
timestamp 1649977179
transform 1 0 39744 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1499
timestamp 1649977179
transform 1 0 44896 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1500
timestamp 1649977179
transform 1 0 50048 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1501
timestamp 1649977179
transform 1 0 55200 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1502
timestamp 1649977179
transform 1 0 60352 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1503
timestamp 1649977179
transform 1 0 65504 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1504
timestamp 1649977179
transform 1 0 6256 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1505
timestamp 1649977179
transform 1 0 11408 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1506
timestamp 1649977179
transform 1 0 16560 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1507
timestamp 1649977179
transform 1 0 21712 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1508
timestamp 1649977179
transform 1 0 26864 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1509
timestamp 1649977179
transform 1 0 32016 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1510
timestamp 1649977179
transform 1 0 37168 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1511
timestamp 1649977179
transform 1 0 42320 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1512
timestamp 1649977179
transform 1 0 47472 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1513
timestamp 1649977179
transform 1 0 52624 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1514
timestamp 1649977179
transform 1 0 57776 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1515
timestamp 1649977179
transform 1 0 62928 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1516
timestamp 1649977179
transform 1 0 68080 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1517
timestamp 1649977179
transform 1 0 3680 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1518
timestamp 1649977179
transform 1 0 8832 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1519
timestamp 1649977179
transform 1 0 13984 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1520
timestamp 1649977179
transform 1 0 19136 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1521
timestamp 1649977179
transform 1 0 24288 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1522
timestamp 1649977179
transform 1 0 29440 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1523
timestamp 1649977179
transform 1 0 34592 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1524
timestamp 1649977179
transform 1 0 39744 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1525
timestamp 1649977179
transform 1 0 44896 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1526
timestamp 1649977179
transform 1 0 50048 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1527
timestamp 1649977179
transform 1 0 55200 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1528
timestamp 1649977179
transform 1 0 60352 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1529
timestamp 1649977179
transform 1 0 65504 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1530
timestamp 1649977179
transform 1 0 3680 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1531
timestamp 1649977179
transform 1 0 6256 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1532
timestamp 1649977179
transform 1 0 8832 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1533
timestamp 1649977179
transform 1 0 11408 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1534
timestamp 1649977179
transform 1 0 13984 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1535
timestamp 1649977179
transform 1 0 16560 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1536
timestamp 1649977179
transform 1 0 19136 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1537
timestamp 1649977179
transform 1 0 21712 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1538
timestamp 1649977179
transform 1 0 24288 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1539
timestamp 1649977179
transform 1 0 26864 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1540
timestamp 1649977179
transform 1 0 29440 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1541
timestamp 1649977179
transform 1 0 32016 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1542
timestamp 1649977179
transform 1 0 34592 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1543
timestamp 1649977179
transform 1 0 37168 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1544
timestamp 1649977179
transform 1 0 39744 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1545
timestamp 1649977179
transform 1 0 42320 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1546
timestamp 1649977179
transform 1 0 44896 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1547
timestamp 1649977179
transform 1 0 47472 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1548
timestamp 1649977179
transform 1 0 50048 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1549
timestamp 1649977179
transform 1 0 52624 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1550
timestamp 1649977179
transform 1 0 55200 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1551
timestamp 1649977179
transform 1 0 57776 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1552
timestamp 1649977179
transform 1 0 60352 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1553
timestamp 1649977179
transform 1 0 62928 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1554
timestamp 1649977179
transform 1 0 65504 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1555
timestamp 1649977179
transform 1 0 68080 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__or4_1  _162_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 9200 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _163_
timestamp 1649977179
transform 1 0 10028 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nor4_2  _164_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 10856 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _165_
timestamp 1649977179
transform 1 0 19964 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _166_
timestamp 1649977179
transform 1 0 23184 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__nor4_1  _167_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 24288 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _168_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 12696 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _169_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 7820 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__or4bb_1  _170_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 21160 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _171_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 20700 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _172_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 5612 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _173_
timestamp 1649977179
transform -1 0 11040 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_2  _174_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2576 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _175_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 5336 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _176_
timestamp 1649977179
transform 1 0 8188 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _177_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 4416 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _178_
timestamp 1649977179
transform -1 0 20608 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _179_
timestamp 1649977179
transform 1 0 5244 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _180_
timestamp 1649977179
transform -1 0 3588 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _181_
timestamp 1649977179
transform 1 0 6348 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _182_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 4784 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _183_
timestamp 1649977179
transform -1 0 4876 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _184_
timestamp 1649977179
transform -1 0 5612 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _185_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 6624 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _186_
timestamp 1649977179
transform 1 0 4968 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _187_
timestamp 1649977179
transform -1 0 6440 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _188_
timestamp 1649977179
transform 1 0 4140 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _189_
timestamp 1649977179
transform -1 0 5428 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _190_
timestamp 1649977179
transform 1 0 4140 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _191_
timestamp 1649977179
transform -1 0 5428 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _192_
timestamp 1649977179
transform 1 0 5336 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _193_
timestamp 1649977179
transform -1 0 7084 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _194_
timestamp 1649977179
transform -1 0 6624 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _195_
timestamp 1649977179
transform -1 0 5796 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _196_
timestamp 1649977179
transform -1 0 5888 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _197_
timestamp 1649977179
transform -1 0 4324 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _198_
timestamp 1649977179
transform 1 0 5336 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _199_
timestamp 1649977179
transform -1 0 5152 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _200_
timestamp 1649977179
transform -1 0 6624 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _201_
timestamp 1649977179
transform 1 0 4692 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _202_
timestamp 1649977179
transform -1 0 6164 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _203_
timestamp 1649977179
transform 1 0 6348 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _204_
timestamp 1649977179
transform -1 0 7084 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _205_
timestamp 1649977179
transform 1 0 5428 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _206_
timestamp 1649977179
transform -1 0 6900 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _207_
timestamp 1649977179
transform 1 0 5244 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _208_
timestamp 1649977179
transform -1 0 7084 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _209_
timestamp 1649977179
transform -1 0 12880 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _210_
timestamp 1649977179
transform -1 0 9660 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _211_
timestamp 1649977179
transform -1 0 9752 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _212_
timestamp 1649977179
transform -1 0 10396 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _213_
timestamp 1649977179
transform -1 0 9752 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _214_
timestamp 1649977179
transform 1 0 12696 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _215_
timestamp 1649977179
transform -1 0 10764 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _216_
timestamp 1649977179
transform 1 0 10120 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _217_
timestamp 1649977179
transform 1 0 10120 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _218_
timestamp 1649977179
transform 1 0 11960 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _219_
timestamp 1649977179
transform -1 0 13616 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _220_
timestamp 1649977179
transform 1 0 11040 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _221_
timestamp 1649977179
transform -1 0 12972 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _222_
timestamp 1649977179
transform 1 0 11592 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _223_
timestamp 1649977179
transform -1 0 13248 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _224_
timestamp 1649977179
transform 1 0 16652 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _225_
timestamp 1649977179
transform -1 0 11868 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _226_
timestamp 1649977179
transform 1 0 20240 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _227_
timestamp 1649977179
transform -1 0 10396 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _228_
timestamp 1649977179
transform 1 0 17296 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _229_
timestamp 1649977179
transform 1 0 16652 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _230_
timestamp 1649977179
transform 1 0 16652 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _231_
timestamp 1649977179
transform 1 0 14536 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _232_
timestamp 1649977179
transform 1 0 14996 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _233_
timestamp 1649977179
transform 1 0 16376 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _234_
timestamp 1649977179
transform 1 0 16652 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _235_
timestamp 1649977179
transform 1 0 15272 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _236_
timestamp 1649977179
transform 1 0 15088 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _237_
timestamp 1649977179
transform 1 0 15456 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _238_
timestamp 1649977179
transform 1 0 16192 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _239_
timestamp 1649977179
transform -1 0 15916 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _240_
timestamp 1649977179
transform -1 0 21344 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _241_
timestamp 1649977179
transform 1 0 20424 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _242_
timestamp 1649977179
transform -1 0 9752 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _243_
timestamp 1649977179
transform -1 0 21436 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _244_
timestamp 1649977179
transform -1 0 16192 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _245_
timestamp 1649977179
transform 1 0 20424 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _246_
timestamp 1649977179
transform -1 0 20148 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _247_
timestamp 1649977179
transform 1 0 20148 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _248_
timestamp 1649977179
transform 1 0 21804 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _249_
timestamp 1649977179
transform -1 0 22908 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _250_
timestamp 1649977179
transform 1 0 21804 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _251_
timestamp 1649977179
transform 1 0 21068 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _252_
timestamp 1649977179
transform 1 0 20516 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _253_
timestamp 1649977179
transform 1 0 20608 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _254_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 4508 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _255_
timestamp 1649977179
transform 1 0 14720 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _256_
timestamp 1649977179
transform -1 0 7544 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _257_
timestamp 1649977179
transform -1 0 7544 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _258_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 8004 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _259_
timestamp 1649977179
transform 1 0 4140 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _260_
timestamp 1649977179
transform -1 0 12420 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _261_
timestamp 1649977179
transform 1 0 10304 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _262_
timestamp 1649977179
transform 1 0 7912 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _263_
timestamp 1649977179
transform 1 0 11592 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _264_
timestamp 1649977179
transform 1 0 8832 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _265_
timestamp 1649977179
transform 1 0 12512 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _266_
timestamp 1649977179
transform 1 0 9016 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _267_
timestamp 1649977179
transform 1 0 10304 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _268_
timestamp 1649977179
transform 1 0 8924 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _269_
timestamp 1649977179
transform -1 0 13800 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _270_
timestamp 1649977179
transform -1 0 5060 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _271_
timestamp 1649977179
transform -1 0 2944 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _272_
timestamp 1649977179
transform -1 0 3588 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _273_
timestamp 1649977179
transform 1 0 3496 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _274_
timestamp 1649977179
transform -1 0 5888 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _275_
timestamp 1649977179
transform -1 0 5980 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _276_
timestamp 1649977179
transform 1 0 3956 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _277_
timestamp 1649977179
transform -1 0 5888 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _278_
timestamp 1649977179
transform 1 0 3772 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _279_
timestamp 1649977179
transform -1 0 7084 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _280_
timestamp 1649977179
transform 1 0 3772 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _281_
timestamp 1649977179
transform -1 0 4784 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _282_
timestamp 1649977179
transform 1 0 3312 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _283_
timestamp 1649977179
transform -1 0 5888 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _284_
timestamp 1649977179
transform -1 0 13340 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _285_
timestamp 1649977179
transform -1 0 4692 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _286_
timestamp 1649977179
transform -1 0 14444 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _287_
timestamp 1649977179
transform 1 0 12328 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _288_
timestamp 1649977179
transform 1 0 13616 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _289_
timestamp 1649977179
transform 1 0 12512 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _290_
timestamp 1649977179
transform 1 0 11684 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _291_
timestamp 1649977179
transform -1 0 12788 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _292_
timestamp 1649977179
transform 1 0 14812 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _293_
timestamp 1649977179
transform -1 0 16468 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _294_
timestamp 1649977179
transform -1 0 15088 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _295_
timestamp 1649977179
transform -1 0 14260 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _296_
timestamp 1649977179
transform 1 0 14996 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _297_
timestamp 1649977179
transform -1 0 17388 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _298_
timestamp 1649977179
transform 1 0 21896 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _299_
timestamp 1649977179
transform 1 0 24380 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _300_
timestamp 1649977179
transform 1 0 21804 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _301_
timestamp 1649977179
transform -1 0 21068 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _302_
timestamp 1649977179
transform 1 0 22908 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _303_
timestamp 1649977179
transform 1 0 20976 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _304_
timestamp 1649977179
transform 1 0 21436 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _305_
timestamp 1649977179
transform 1 0 21804 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _306_
timestamp 1649977179
transform 1 0 22448 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _307_
timestamp 1649977179
transform 1 0 23276 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _308_
timestamp 1649977179
transform 1 0 24380 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _309_
timestamp 1649977179
transform 1 0 23092 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _310_
timestamp 1649977179
transform 1 0 23276 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _311_
timestamp 1649977179
transform 1 0 23000 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _312_
timestamp 1649977179
transform 1 0 21804 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _313_
timestamp 1649977179
transform -1 0 22080 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _314_
timestamp 1649977179
transform -1 0 21344 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _315_
timestamp 1649977179
transform 1 0 23460 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _316_
timestamp 1649977179
transform 1 0 21344 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _317_
timestamp 1649977179
transform 1 0 22724 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _318_
timestamp 1649977179
transform 1 0 22632 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _319_
timestamp 1649977179
transform 1 0 22724 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _320_
timestamp 1649977179
transform 1 0 23000 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _321_
timestamp 1649977179
transform -1 0 23920 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _322_
timestamp 1649977179
transform 1 0 22356 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _323_
timestamp 1649977179
transform 1 0 22632 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _324_
timestamp 1649977179
transform -1 0 22264 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _325_
timestamp 1649977179
transform 1 0 20240 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _326_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 6992 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _327_
timestamp 1649977179
transform 1 0 7176 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _328_
timestamp 1649977179
transform -1 0 10488 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _329_
timestamp 1649977179
transform 1 0 6992 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _330_
timestamp 1649977179
transform 1 0 7728 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _331_
timestamp 1649977179
transform 1 0 6992 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _332_
timestamp 1649977179
transform 1 0 6992 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _333_
timestamp 1649977179
transform 1 0 6992 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _334_
timestamp 1649977179
transform 1 0 6992 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _335_
timestamp 1649977179
transform 1 0 6532 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _336_
timestamp 1649977179
transform 1 0 10764 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _337_
timestamp 1649977179
transform 1 0 10304 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _338_
timestamp 1649977179
transform -1 0 15732 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _339_
timestamp 1649977179
transform 1 0 12880 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _340_
timestamp 1649977179
transform 1 0 14076 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _341_
timestamp 1649977179
transform 1 0 12972 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _342_
timestamp 1649977179
transform 1 0 13432 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _343_
timestamp 1649977179
transform 1 0 16100 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _344_
timestamp 1649977179
transform 1 0 14628 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _345_
timestamp 1649977179
transform 1 0 15364 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _346_
timestamp 1649977179
transform 1 0 18400 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _347_
timestamp 1649977179
transform 1 0 18124 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _348_
timestamp 1649977179
transform 1 0 15456 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _349_
timestamp 1649977179
transform 1 0 17296 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _350_
timestamp 1649977179
transform 1 0 19228 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _351_
timestamp 1649977179
transform 1 0 9568 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _352_
timestamp 1649977179
transform -1 0 11776 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _353_
timestamp 1649977179
transform 1 0 11960 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _354_
timestamp 1649977179
transform 1 0 10120 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _355_
timestamp 1649977179
transform -1 0 13616 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _356_
timestamp 1649977179
transform 1 0 8372 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _357_
timestamp 1649977179
transform 1 0 6992 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _358_
timestamp 1649977179
transform 1 0 7176 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _359_
timestamp 1649977179
transform 1 0 10304 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _360_
timestamp 1649977179
transform 1 0 9292 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _361_
timestamp 1649977179
transform 1 0 10120 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _362_
timestamp 1649977179
transform 1 0 13156 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _363_
timestamp 1649977179
transform -1 0 18676 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _364_
timestamp 1649977179
transform -1 0 16100 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _365_
timestamp 1649977179
transform -1 0 18492 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _366_
timestamp 1649977179
transform -1 0 18124 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _367_
timestamp 1649977179
transform -1 0 19596 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _368_
timestamp 1649977179
transform 1 0 17940 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _369_
timestamp 1649977179
transform 1 0 19228 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _370_
timestamp 1649977179
transform 1 0 18400 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _371_
timestamp 1649977179
transform 1 0 18124 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _372_
timestamp 1649977179
transform 1 0 17296 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _373_
timestamp 1649977179
transform 1 0 18124 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _374_
timestamp 1649977179
transform 1 0 19228 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _375_
timestamp 1649977179
transform 1 0 15916 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wb_clk_i dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 13340 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_wb_clk_i
timestamp 1649977179
transform -1 0 9660 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_wb_clk_i
timestamp 1649977179
transform -1 0 9660 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_wb_clk_i
timestamp 1649977179
transform 1 0 15640 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_wb_clk_i
timestamp 1649977179
transform 1 0 15640 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1649977179
transform -1 0 4140 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1649977179
transform -1 0 19872 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1649977179
transform -1 0 18032 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1649977179
transform 1 0 21804 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1649977179
transform -1 0 21344 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1649977179
transform -1 0 9568 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1649977179
transform 1 0 7728 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1649977179
transform 1 0 14996 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1649977179
transform -1 0 8464 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1649977179
transform 1 0 15456 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1649977179
transform 1 0 13340 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1649977179
transform 1 0 12236 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1649977179
transform -1 0 16192 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1649977179
transform 1 0 17848 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1649977179
transform -1 0 9752 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1649977179
transform 1 0 15916 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1649977179
transform 1 0 17480 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1649977179
transform 1 0 11408 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1649977179
transform -1 0 18768 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1649977179
transform -1 0 19504 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1649977179
transform -1 0 17112 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1649977179
transform -1 0 18768 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1649977179
transform -1 0 18124 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1649977179
transform 1 0 10764 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1649977179
transform 1 0 4508 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1649977179
transform 1 0 6532 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1649977179
transform 1 0 12696 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1649977179
transform 1 0 12052 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1649977179
transform 1 0 9476 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1649977179
transform 1 0 14352 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1649977179
transform 1 0 7544 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1649977179
transform 1 0 13616 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1649977179
transform -1 0 11868 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1649977179
transform 1 0 6348 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output35
timestamp 1649977179
transform 1 0 26128 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output36
timestamp 1649977179
transform 1 0 26956 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output37
timestamp 1649977179
transform 1 0 13156 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output38
timestamp 1649977179
transform 1 0 13248 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output39
timestamp 1649977179
transform 1 0 15824 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output40
timestamp 1649977179
transform -1 0 15364 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output41
timestamp 1649977179
transform 1 0 14352 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output42
timestamp 1649977179
transform 1 0 17204 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output43
timestamp 1649977179
transform -1 0 15456 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output44
timestamp 1649977179
transform -1 0 18584 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output45
timestamp 1649977179
transform -1 0 22172 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output46
timestamp 1649977179
transform -1 0 16192 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output47
timestamp 1649977179
transform -1 0 20332 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output48
timestamp 1649977179
transform -1 0 9568 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output49
timestamp 1649977179
transform -1 0 19596 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output50
timestamp 1649977179
transform -1 0 21252 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output51
timestamp 1649977179
transform -1 0 20608 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output52
timestamp 1649977179
transform -1 0 19780 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output53
timestamp 1649977179
transform -1 0 20516 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output54
timestamp 1649977179
transform 1 0 13248 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output55
timestamp 1649977179
transform -1 0 10304 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output56
timestamp 1649977179
transform -1 0 11040 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output57
timestamp 1649977179
transform 1 0 11960 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output58
timestamp 1649977179
transform 1 0 11776 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output59
timestamp 1649977179
transform 1 0 12512 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output60
timestamp 1649977179
transform 1 0 14260 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output61
timestamp 1649977179
transform 1 0 15088 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  pixel_macro_62 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 67344 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_63
timestamp 1649977179
transform 1 0 6348 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_64
timestamp 1649977179
transform 1 0 18952 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_65
timestamp 1649977179
transform -1 0 24288 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_66
timestamp 1649977179
transform -1 0 22724 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_67
timestamp 1649977179
transform -1 0 21528 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_68
timestamp 1649977179
transform 1 0 19780 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_69
timestamp 1649977179
transform -1 0 24656 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_70
timestamp 1649977179
transform -1 0 23644 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_71
timestamp 1649977179
transform -1 0 23000 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_72
timestamp 1649977179
transform -1 0 23092 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_73
timestamp 1649977179
transform 1 0 22356 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_74
timestamp 1649977179
transform 1 0 23000 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_75
timestamp 1649977179
transform -1 0 23920 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_76
timestamp 1649977179
transform 1 0 23000 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_77
timestamp 1649977179
transform 1 0 23644 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_78
timestamp 1649977179
transform 1 0 23644 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_79
timestamp 1649977179
transform 1 0 24288 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_80
timestamp 1649977179
transform 1 0 25576 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_81
timestamp 1649977179
transform -1 0 26404 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_82
timestamp 1649977179
transform -1 0 26496 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_83
timestamp 1649977179
transform 1 0 25484 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_84
timestamp 1649977179
transform 1 0 27048 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_85
timestamp 1649977179
transform -1 0 27968 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_86
timestamp 1649977179
transform 1 0 27508 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_87
timestamp 1649977179
transform -1 0 28612 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_88
timestamp 1649977179
transform 1 0 28152 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_89
timestamp 1649977179
transform 1 0 28152 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_90
timestamp 1649977179
transform 1 0 28796 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_91
timestamp 1649977179
transform -1 0 29808 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_92
timestamp 1649977179
transform 1 0 28796 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_93
timestamp 1649977179
transform 1 0 29440 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_94
timestamp 1649977179
transform -1 0 30544 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_95
timestamp 1649977179
transform 1 0 30084 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_96
timestamp 1649977179
transform 1 0 30084 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_97
timestamp 1649977179
transform 1 0 30728 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_98
timestamp 1649977179
transform -1 0 31648 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_99
timestamp 1649977179
transform 1 0 30728 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_100
timestamp 1649977179
transform 1 0 31372 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_101
timestamp 1649977179
transform -1 0 32476 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_102
timestamp 1649977179
transform 1 0 31372 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_103
timestamp 1649977179
transform 1 0 32292 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_104
timestamp 1649977179
transform -1 0 33304 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_105
timestamp 1649977179
transform 1 0 32936 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_106
timestamp 1649977179
transform 1 0 32660 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_107
timestamp 1649977179
transform 1 0 33580 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_108
timestamp 1649977179
transform 1 0 33304 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_109
timestamp 1649977179
transform -1 0 34500 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_110
timestamp 1649977179
transform 1 0 33948 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_111
timestamp 1649977179
transform -1 0 35144 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_112
timestamp 1649977179
transform 1 0 34776 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_113
timestamp 1649977179
transform -1 0 35788 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_114
timestamp 1649977179
transform 1 0 35420 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_115
timestamp 1649977179
transform -1 0 36340 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_116
timestamp 1649977179
transform -1 0 36616 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_117
timestamp 1649977179
transform -1 0 37536 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_118
timestamp 1649977179
transform -1 0 37536 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_119
timestamp 1649977179
transform -1 0 38180 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_120
timestamp 1649977179
transform -1 0 38180 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_121
timestamp 1649977179
transform -1 0 38824 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_122
timestamp 1649977179
transform -1 0 38824 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_123
timestamp 1649977179
transform -1 0 40112 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_124
timestamp 1649977179
transform -1 0 39468 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_125
timestamp 1649977179
transform -1 0 40756 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_126
timestamp 1649977179
transform -1 0 40112 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_127
timestamp 1649977179
transform -1 0 41400 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_128
timestamp 1649977179
transform -1 0 40756 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_129
timestamp 1649977179
transform -1 0 40204 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_130
timestamp 1649977179
transform -1 0 40848 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_131
timestamp 1649977179
transform -1 0 41400 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_132
timestamp 1649977179
transform -1 0 42688 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_133
timestamp 1649977179
transform -1 0 41492 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_134
timestamp 1649977179
transform -1 0 43332 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_135
timestamp 1649977179
transform -1 0 42688 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_136
timestamp 1649977179
transform -1 0 42136 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_137
timestamp 1649977179
transform -1 0 43976 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_138
timestamp 1649977179
transform -1 0 43332 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_139
timestamp 1649977179
transform -1 0 42964 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_140
timestamp 1649977179
transform -1 0 43976 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_141
timestamp 1649977179
transform -1 0 45264 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_142
timestamp 1649977179
transform -1 0 44620 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_143
timestamp 1649977179
transform -1 0 44068 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_144
timestamp 1649977179
transform -1 0 45908 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_145
timestamp 1649977179
transform -1 0 45264 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_146
timestamp 1649977179
transform -1 0 46552 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_147
timestamp 1649977179
transform -1 0 45908 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_148
timestamp 1649977179
transform -1 0 45448 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_149
timestamp 1649977179
transform -1 0 46552 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_150
timestamp 1649977179
transform -1 0 46092 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_151
timestamp 1649977179
transform -1 0 47840 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_152
timestamp 1649977179
transform -1 0 46736 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_153
timestamp 1649977179
transform -1 0 48484 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_154
timestamp 1649977179
transform -1 0 47840 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_155
timestamp 1649977179
transform -1 0 49128 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_156
timestamp 1649977179
transform -1 0 48484 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_157
timestamp 1649977179
transform -1 0 47932 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_158
timestamp 1649977179
transform -1 0 48576 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_159
timestamp 1649977179
transform -1 0 49128 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_160
timestamp 1649977179
transform -1 0 50416 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_161
timestamp 1649977179
transform -1 0 49772 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_162
timestamp 1649977179
transform -1 0 51060 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_163
timestamp 1649977179
transform -1 0 50416 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_164
timestamp 1649977179
transform -1 0 50416 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_165
timestamp 1649977179
transform -1 0 51704 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_166
timestamp 1649977179
transform -1 0 51060 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_167
timestamp 1649977179
transform -1 0 51060 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_168
timestamp 1649977179
transform -1 0 51704 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_169
timestamp 1649977179
transform -1 0 52992 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_170
timestamp 1649977179
transform -1 0 51704 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_171
timestamp 1649977179
transform -1 0 52348 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_172
timestamp 1649977179
transform -1 0 53636 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_173
timestamp 1649977179
transform -1 0 52992 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_174
timestamp 1649977179
transform -1 0 54280 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_175
timestamp 1649977179
transform -1 0 53636 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_176
timestamp 1649977179
transform -1 0 53176 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_177
timestamp 1649977179
transform -1 0 54280 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_178
timestamp 1649977179
transform -1 0 53820 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_179
timestamp 1649977179
transform -1 0 55568 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_180
timestamp 1649977179
transform -1 0 54924 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_181
timestamp 1649977179
transform -1 0 56212 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_182
timestamp 1649977179
transform -1 0 55568 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_183
timestamp 1649977179
transform -1 0 56856 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_184
timestamp 1649977179
transform -1 0 56212 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_185
timestamp 1649977179
transform -1 0 55660 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_186
timestamp 1649977179
transform -1 0 56304 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_187
timestamp 1649977179
transform -1 0 56856 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_188
timestamp 1649977179
transform -1 0 58144 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_189
timestamp 1649977179
transform -1 0 56948 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_190
timestamp 1649977179
transform -1 0 58788 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_191
timestamp 1649977179
transform -1 0 58144 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_192
timestamp 1649977179
transform -1 0 57592 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_193
timestamp 1649977179
transform -1 0 59432 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_194
timestamp 1649977179
transform -1 0 58236 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_195
timestamp 1649977179
transform -1 0 58788 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_196
timestamp 1649977179
transform -1 0 4416 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_197
timestamp 1649977179
transform -1 0 5888 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_198
timestamp 1649977179
transform -1 0 7728 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_199
timestamp 1649977179
transform -1 0 9384 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_200
timestamp 1649977179
transform -1 0 11040 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_201
timestamp 1649977179
transform -1 0 12696 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_202
timestamp 1649977179
transform -1 0 14352 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_203
timestamp 1649977179
transform -1 0 16008 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_204
timestamp 1649977179
transform -1 0 17664 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_205
timestamp 1649977179
transform -1 0 19504 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_206
timestamp 1649977179
transform -1 0 20976 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_207
timestamp 1649977179
transform -1 0 22632 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_208
timestamp 1649977179
transform -1 0 24656 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_209
timestamp 1649977179
transform -1 0 25944 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_210
timestamp 1649977179
transform -1 0 27600 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_211
timestamp 1649977179
transform -1 0 29072 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_212
timestamp 1649977179
transform -1 0 30912 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_213
timestamp 1649977179
transform -1 0 32568 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_214
timestamp 1649977179
transform -1 0 34224 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_215
timestamp 1649977179
transform -1 0 35880 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_216
timestamp 1649977179
transform -1 0 38180 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_217
timestamp 1649977179
transform -1 0 39192 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_218
timestamp 1649977179
transform -1 0 40940 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_219
timestamp 1649977179
transform -1 0 42688 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_220
timestamp 1649977179
transform -1 0 44252 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_221
timestamp 1649977179
transform -1 0 45908 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_222
timestamp 1649977179
transform -1 0 47840 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_223
timestamp 1649977179
transform -1 0 49220 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_224
timestamp 1649977179
transform -1 0 51060 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_225
timestamp 1649977179
transform -1 0 52992 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_226
timestamp 1649977179
transform -1 0 54280 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_227
timestamp 1649977179
transform -1 0 56212 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_228
timestamp 1649977179
transform -1 0 58144 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_229
timestamp 1649977179
transform -1 0 59432 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_230
timestamp 1649977179
transform -1 0 61364 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_231
timestamp 1649977179
transform -1 0 62376 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_232
timestamp 1649977179
transform -1 0 64124 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_233
timestamp 1649977179
transform -1 0 65872 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_234
timestamp 1649977179
transform 1 0 3036 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_235
timestamp 1649977179
transform 1 0 4968 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_236
timestamp 1649977179
transform -1 0 7084 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_237
timestamp 1649977179
transform 1 0 8188 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_238
timestamp 1649977179
transform -1 0 10396 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_239
timestamp 1649977179
transform -1 0 12052 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_240
timestamp 1649977179
transform -1 0 13616 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_241
timestamp 1649977179
transform -1 0 15364 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_242
timestamp 1649977179
transform -1 0 17020 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_243
timestamp 1649977179
transform -1 0 18768 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_244
timestamp 1649977179
transform -1 0 20332 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_245
timestamp 1649977179
transform -1 0 22080 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_246
timestamp 1649977179
transform -1 0 23736 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_247
timestamp 1649977179
transform -1 0 25300 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_248
timestamp 1649977179
transform -1 0 27048 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_249
timestamp 1649977179
transform 1 0 28152 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_250
timestamp 1649977179
transform -1 0 30268 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_251
timestamp 1649977179
transform 1 0 31372 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_252
timestamp 1649977179
transform -1 0 33580 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_253
timestamp 1649977179
transform -1 0 35236 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_254
timestamp 1649977179
transform -1 0 37536 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_255
timestamp 1649977179
transform -1 0 38824 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_256
timestamp 1649977179
transform -1 0 40296 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_257
timestamp 1649977179
transform -1 0 41952 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_258
timestamp 1649977179
transform -1 0 43608 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_259
timestamp 1649977179
transform -1 0 45264 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_260
timestamp 1649977179
transform -1 0 46920 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_261
timestamp 1649977179
transform -1 0 48576 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_262
timestamp 1649977179
transform -1 0 50416 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_263
timestamp 1649977179
transform -1 0 51888 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_264
timestamp 1649977179
transform -1 0 53636 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_265
timestamp 1649977179
transform -1 0 55568 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_266
timestamp 1649977179
transform -1 0 56856 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_267
timestamp 1649977179
transform -1 0 58788 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_268
timestamp 1649977179
transform -1 0 60720 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_269
timestamp 1649977179
transform -1 0 62008 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_270
timestamp 1649977179
transform -1 0 63480 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_271
timestamp 1649977179
transform -1 0 65136 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_272
timestamp 1649977179
transform -1 0 21344 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_273
timestamp 1649977179
transform 1 0 25024 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_274
timestamp 1649977179
transform -1 0 25208 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_275
timestamp 1649977179
transform -1 0 25116 0 1 2176
box -38 -48 314 592
<< labels >>
flabel metal2 s 2962 59200 3018 60000 0 FreeSans 224 90 0 0 io_in[0]
port 0 nsew signal input
flabel metal2 s 19522 59200 19578 60000 0 FreeSans 224 90 0 0 io_in[10]
port 1 nsew signal input
flabel metal2 s 21178 59200 21234 60000 0 FreeSans 224 90 0 0 io_in[11]
port 2 nsew signal input
flabel metal2 s 22834 59200 22890 60000 0 FreeSans 224 90 0 0 io_in[12]
port 3 nsew signal input
flabel metal2 s 24490 59200 24546 60000 0 FreeSans 224 90 0 0 io_in[13]
port 4 nsew signal input
flabel metal2 s 26146 59200 26202 60000 0 FreeSans 224 90 0 0 io_in[14]
port 5 nsew signal input
flabel metal2 s 27802 59200 27858 60000 0 FreeSans 224 90 0 0 io_in[15]
port 6 nsew signal input
flabel metal2 s 29458 59200 29514 60000 0 FreeSans 224 90 0 0 io_in[16]
port 7 nsew signal input
flabel metal2 s 31114 59200 31170 60000 0 FreeSans 224 90 0 0 io_in[17]
port 8 nsew signal input
flabel metal2 s 32770 59200 32826 60000 0 FreeSans 224 90 0 0 io_in[18]
port 9 nsew signal input
flabel metal2 s 34426 59200 34482 60000 0 FreeSans 224 90 0 0 io_in[19]
port 10 nsew signal input
flabel metal2 s 4618 59200 4674 60000 0 FreeSans 224 90 0 0 io_in[1]
port 11 nsew signal input
flabel metal2 s 36082 59200 36138 60000 0 FreeSans 224 90 0 0 io_in[20]
port 12 nsew signal input
flabel metal2 s 37738 59200 37794 60000 0 FreeSans 224 90 0 0 io_in[21]
port 13 nsew signal input
flabel metal2 s 39394 59200 39450 60000 0 FreeSans 224 90 0 0 io_in[22]
port 14 nsew signal input
flabel metal2 s 41050 59200 41106 60000 0 FreeSans 224 90 0 0 io_in[23]
port 15 nsew signal input
flabel metal2 s 42706 59200 42762 60000 0 FreeSans 224 90 0 0 io_in[24]
port 16 nsew signal input
flabel metal2 s 44362 59200 44418 60000 0 FreeSans 224 90 0 0 io_in[25]
port 17 nsew signal input
flabel metal2 s 46018 59200 46074 60000 0 FreeSans 224 90 0 0 io_in[26]
port 18 nsew signal input
flabel metal2 s 47674 59200 47730 60000 0 FreeSans 224 90 0 0 io_in[27]
port 19 nsew signal input
flabel metal2 s 49330 59200 49386 60000 0 FreeSans 224 90 0 0 io_in[28]
port 20 nsew signal input
flabel metal2 s 50986 59200 51042 60000 0 FreeSans 224 90 0 0 io_in[29]
port 21 nsew signal input
flabel metal2 s 6274 59200 6330 60000 0 FreeSans 224 90 0 0 io_in[2]
port 22 nsew signal input
flabel metal2 s 52642 59200 52698 60000 0 FreeSans 224 90 0 0 io_in[30]
port 23 nsew signal input
flabel metal2 s 54298 59200 54354 60000 0 FreeSans 224 90 0 0 io_in[31]
port 24 nsew signal input
flabel metal2 s 55954 59200 56010 60000 0 FreeSans 224 90 0 0 io_in[32]
port 25 nsew signal input
flabel metal2 s 57610 59200 57666 60000 0 FreeSans 224 90 0 0 io_in[33]
port 26 nsew signal input
flabel metal2 s 59266 59200 59322 60000 0 FreeSans 224 90 0 0 io_in[34]
port 27 nsew signal input
flabel metal2 s 60922 59200 60978 60000 0 FreeSans 224 90 0 0 io_in[35]
port 28 nsew signal input
flabel metal2 s 62578 59200 62634 60000 0 FreeSans 224 90 0 0 io_in[36]
port 29 nsew signal input
flabel metal2 s 64234 59200 64290 60000 0 FreeSans 224 90 0 0 io_in[37]
port 30 nsew signal input
flabel metal2 s 7930 59200 7986 60000 0 FreeSans 224 90 0 0 io_in[3]
port 31 nsew signal input
flabel metal2 s 9586 59200 9642 60000 0 FreeSans 224 90 0 0 io_in[4]
port 32 nsew signal input
flabel metal2 s 11242 59200 11298 60000 0 FreeSans 224 90 0 0 io_in[5]
port 33 nsew signal input
flabel metal2 s 12898 59200 12954 60000 0 FreeSans 224 90 0 0 io_in[6]
port 34 nsew signal input
flabel metal2 s 14554 59200 14610 60000 0 FreeSans 224 90 0 0 io_in[7]
port 35 nsew signal input
flabel metal2 s 16210 59200 16266 60000 0 FreeSans 224 90 0 0 io_in[8]
port 36 nsew signal input
flabel metal2 s 17866 59200 17922 60000 0 FreeSans 224 90 0 0 io_in[9]
port 37 nsew signal input
flabel metal2 s 3514 59200 3570 60000 0 FreeSans 224 90 0 0 io_oeb[0]
port 38 nsew signal tristate
flabel metal2 s 20074 59200 20130 60000 0 FreeSans 224 90 0 0 io_oeb[10]
port 39 nsew signal tristate
flabel metal2 s 21730 59200 21786 60000 0 FreeSans 224 90 0 0 io_oeb[11]
port 40 nsew signal tristate
flabel metal2 s 23386 59200 23442 60000 0 FreeSans 224 90 0 0 io_oeb[12]
port 41 nsew signal tristate
flabel metal2 s 25042 59200 25098 60000 0 FreeSans 224 90 0 0 io_oeb[13]
port 42 nsew signal tristate
flabel metal2 s 26698 59200 26754 60000 0 FreeSans 224 90 0 0 io_oeb[14]
port 43 nsew signal tristate
flabel metal2 s 28354 59200 28410 60000 0 FreeSans 224 90 0 0 io_oeb[15]
port 44 nsew signal tristate
flabel metal2 s 30010 59200 30066 60000 0 FreeSans 224 90 0 0 io_oeb[16]
port 45 nsew signal tristate
flabel metal2 s 31666 59200 31722 60000 0 FreeSans 224 90 0 0 io_oeb[17]
port 46 nsew signal tristate
flabel metal2 s 33322 59200 33378 60000 0 FreeSans 224 90 0 0 io_oeb[18]
port 47 nsew signal tristate
flabel metal2 s 34978 59200 35034 60000 0 FreeSans 224 90 0 0 io_oeb[19]
port 48 nsew signal tristate
flabel metal2 s 5170 59200 5226 60000 0 FreeSans 224 90 0 0 io_oeb[1]
port 49 nsew signal tristate
flabel metal2 s 36634 59200 36690 60000 0 FreeSans 224 90 0 0 io_oeb[20]
port 50 nsew signal tristate
flabel metal2 s 38290 59200 38346 60000 0 FreeSans 224 90 0 0 io_oeb[21]
port 51 nsew signal tristate
flabel metal2 s 39946 59200 40002 60000 0 FreeSans 224 90 0 0 io_oeb[22]
port 52 nsew signal tristate
flabel metal2 s 41602 59200 41658 60000 0 FreeSans 224 90 0 0 io_oeb[23]
port 53 nsew signal tristate
flabel metal2 s 43258 59200 43314 60000 0 FreeSans 224 90 0 0 io_oeb[24]
port 54 nsew signal tristate
flabel metal2 s 44914 59200 44970 60000 0 FreeSans 224 90 0 0 io_oeb[25]
port 55 nsew signal tristate
flabel metal2 s 46570 59200 46626 60000 0 FreeSans 224 90 0 0 io_oeb[26]
port 56 nsew signal tristate
flabel metal2 s 48226 59200 48282 60000 0 FreeSans 224 90 0 0 io_oeb[27]
port 57 nsew signal tristate
flabel metal2 s 49882 59200 49938 60000 0 FreeSans 224 90 0 0 io_oeb[28]
port 58 nsew signal tristate
flabel metal2 s 51538 59200 51594 60000 0 FreeSans 224 90 0 0 io_oeb[29]
port 59 nsew signal tristate
flabel metal2 s 6826 59200 6882 60000 0 FreeSans 224 90 0 0 io_oeb[2]
port 60 nsew signal tristate
flabel metal2 s 53194 59200 53250 60000 0 FreeSans 224 90 0 0 io_oeb[30]
port 61 nsew signal tristate
flabel metal2 s 54850 59200 54906 60000 0 FreeSans 224 90 0 0 io_oeb[31]
port 62 nsew signal tristate
flabel metal2 s 56506 59200 56562 60000 0 FreeSans 224 90 0 0 io_oeb[32]
port 63 nsew signal tristate
flabel metal2 s 58162 59200 58218 60000 0 FreeSans 224 90 0 0 io_oeb[33]
port 64 nsew signal tristate
flabel metal2 s 59818 59200 59874 60000 0 FreeSans 224 90 0 0 io_oeb[34]
port 65 nsew signal tristate
flabel metal2 s 61474 59200 61530 60000 0 FreeSans 224 90 0 0 io_oeb[35]
port 66 nsew signal tristate
flabel metal2 s 63130 59200 63186 60000 0 FreeSans 224 90 0 0 io_oeb[36]
port 67 nsew signal tristate
flabel metal2 s 64786 59200 64842 60000 0 FreeSans 224 90 0 0 io_oeb[37]
port 68 nsew signal tristate
flabel metal2 s 8482 59200 8538 60000 0 FreeSans 224 90 0 0 io_oeb[3]
port 69 nsew signal tristate
flabel metal2 s 10138 59200 10194 60000 0 FreeSans 224 90 0 0 io_oeb[4]
port 70 nsew signal tristate
flabel metal2 s 11794 59200 11850 60000 0 FreeSans 224 90 0 0 io_oeb[5]
port 71 nsew signal tristate
flabel metal2 s 13450 59200 13506 60000 0 FreeSans 224 90 0 0 io_oeb[6]
port 72 nsew signal tristate
flabel metal2 s 15106 59200 15162 60000 0 FreeSans 224 90 0 0 io_oeb[7]
port 73 nsew signal tristate
flabel metal2 s 16762 59200 16818 60000 0 FreeSans 224 90 0 0 io_oeb[8]
port 74 nsew signal tristate
flabel metal2 s 18418 59200 18474 60000 0 FreeSans 224 90 0 0 io_oeb[9]
port 75 nsew signal tristate
flabel metal2 s 4066 59200 4122 60000 0 FreeSans 224 90 0 0 io_out[0]
port 76 nsew signal tristate
flabel metal2 s 20626 59200 20682 60000 0 FreeSans 224 90 0 0 io_out[10]
port 77 nsew signal tristate
flabel metal2 s 22282 59200 22338 60000 0 FreeSans 224 90 0 0 io_out[11]
port 78 nsew signal tristate
flabel metal2 s 23938 59200 23994 60000 0 FreeSans 224 90 0 0 io_out[12]
port 79 nsew signal tristate
flabel metal2 s 25594 59200 25650 60000 0 FreeSans 224 90 0 0 io_out[13]
port 80 nsew signal tristate
flabel metal2 s 27250 59200 27306 60000 0 FreeSans 224 90 0 0 io_out[14]
port 81 nsew signal tristate
flabel metal2 s 28906 59200 28962 60000 0 FreeSans 224 90 0 0 io_out[15]
port 82 nsew signal tristate
flabel metal2 s 30562 59200 30618 60000 0 FreeSans 224 90 0 0 io_out[16]
port 83 nsew signal tristate
flabel metal2 s 32218 59200 32274 60000 0 FreeSans 224 90 0 0 io_out[17]
port 84 nsew signal tristate
flabel metal2 s 33874 59200 33930 60000 0 FreeSans 224 90 0 0 io_out[18]
port 85 nsew signal tristate
flabel metal2 s 35530 59200 35586 60000 0 FreeSans 224 90 0 0 io_out[19]
port 86 nsew signal tristate
flabel metal2 s 5722 59200 5778 60000 0 FreeSans 224 90 0 0 io_out[1]
port 87 nsew signal tristate
flabel metal2 s 37186 59200 37242 60000 0 FreeSans 224 90 0 0 io_out[20]
port 88 nsew signal tristate
flabel metal2 s 38842 59200 38898 60000 0 FreeSans 224 90 0 0 io_out[21]
port 89 nsew signal tristate
flabel metal2 s 40498 59200 40554 60000 0 FreeSans 224 90 0 0 io_out[22]
port 90 nsew signal tristate
flabel metal2 s 42154 59200 42210 60000 0 FreeSans 224 90 0 0 io_out[23]
port 91 nsew signal tristate
flabel metal2 s 43810 59200 43866 60000 0 FreeSans 224 90 0 0 io_out[24]
port 92 nsew signal tristate
flabel metal2 s 45466 59200 45522 60000 0 FreeSans 224 90 0 0 io_out[25]
port 93 nsew signal tristate
flabel metal2 s 47122 59200 47178 60000 0 FreeSans 224 90 0 0 io_out[26]
port 94 nsew signal tristate
flabel metal2 s 48778 59200 48834 60000 0 FreeSans 224 90 0 0 io_out[27]
port 95 nsew signal tristate
flabel metal2 s 50434 59200 50490 60000 0 FreeSans 224 90 0 0 io_out[28]
port 96 nsew signal tristate
flabel metal2 s 52090 59200 52146 60000 0 FreeSans 224 90 0 0 io_out[29]
port 97 nsew signal tristate
flabel metal2 s 7378 59200 7434 60000 0 FreeSans 224 90 0 0 io_out[2]
port 98 nsew signal tristate
flabel metal2 s 53746 59200 53802 60000 0 FreeSans 224 90 0 0 io_out[30]
port 99 nsew signal tristate
flabel metal2 s 55402 59200 55458 60000 0 FreeSans 224 90 0 0 io_out[31]
port 100 nsew signal tristate
flabel metal2 s 57058 59200 57114 60000 0 FreeSans 224 90 0 0 io_out[32]
port 101 nsew signal tristate
flabel metal2 s 58714 59200 58770 60000 0 FreeSans 224 90 0 0 io_out[33]
port 102 nsew signal tristate
flabel metal2 s 60370 59200 60426 60000 0 FreeSans 224 90 0 0 io_out[34]
port 103 nsew signal tristate
flabel metal2 s 62026 59200 62082 60000 0 FreeSans 224 90 0 0 io_out[35]
port 104 nsew signal tristate
flabel metal2 s 63682 59200 63738 60000 0 FreeSans 224 90 0 0 io_out[36]
port 105 nsew signal tristate
flabel metal2 s 65338 59200 65394 60000 0 FreeSans 224 90 0 0 io_out[37]
port 106 nsew signal tristate
flabel metal2 s 9034 59200 9090 60000 0 FreeSans 224 90 0 0 io_out[3]
port 107 nsew signal tristate
flabel metal2 s 10690 59200 10746 60000 0 FreeSans 224 90 0 0 io_out[4]
port 108 nsew signal tristate
flabel metal2 s 12346 59200 12402 60000 0 FreeSans 224 90 0 0 io_out[5]
port 109 nsew signal tristate
flabel metal2 s 14002 59200 14058 60000 0 FreeSans 224 90 0 0 io_out[6]
port 110 nsew signal tristate
flabel metal2 s 15658 59200 15714 60000 0 FreeSans 224 90 0 0 io_out[7]
port 111 nsew signal tristate
flabel metal2 s 17314 59200 17370 60000 0 FreeSans 224 90 0 0 io_out[8]
port 112 nsew signal tristate
flabel metal2 s 18970 59200 19026 60000 0 FreeSans 224 90 0 0 io_out[9]
port 113 nsew signal tristate
flabel metal2 s 57426 0 57482 800 0 FreeSans 224 90 0 0 irq[0]
port 114 nsew signal tristate
flabel metal2 s 57518 0 57574 800 0 FreeSans 224 90 0 0 irq[1]
port 115 nsew signal tristate
flabel metal2 s 57610 0 57666 800 0 FreeSans 224 90 0 0 irq[2]
port 116 nsew signal tristate
flabel metal2 s 22098 0 22154 800 0 FreeSans 224 90 0 0 la_data_in[0]
port 117 nsew signal input
flabel metal2 s 49698 0 49754 800 0 FreeSans 224 90 0 0 la_data_in[100]
port 118 nsew signal input
flabel metal2 s 49974 0 50030 800 0 FreeSans 224 90 0 0 la_data_in[101]
port 119 nsew signal input
flabel metal2 s 50250 0 50306 800 0 FreeSans 224 90 0 0 la_data_in[102]
port 120 nsew signal input
flabel metal2 s 50526 0 50582 800 0 FreeSans 224 90 0 0 la_data_in[103]
port 121 nsew signal input
flabel metal2 s 50802 0 50858 800 0 FreeSans 224 90 0 0 la_data_in[104]
port 122 nsew signal input
flabel metal2 s 51078 0 51134 800 0 FreeSans 224 90 0 0 la_data_in[105]
port 123 nsew signal input
flabel metal2 s 51354 0 51410 800 0 FreeSans 224 90 0 0 la_data_in[106]
port 124 nsew signal input
flabel metal2 s 51630 0 51686 800 0 FreeSans 224 90 0 0 la_data_in[107]
port 125 nsew signal input
flabel metal2 s 51906 0 51962 800 0 FreeSans 224 90 0 0 la_data_in[108]
port 126 nsew signal input
flabel metal2 s 52182 0 52238 800 0 FreeSans 224 90 0 0 la_data_in[109]
port 127 nsew signal input
flabel metal2 s 24858 0 24914 800 0 FreeSans 224 90 0 0 la_data_in[10]
port 128 nsew signal input
flabel metal2 s 52458 0 52514 800 0 FreeSans 224 90 0 0 la_data_in[110]
port 129 nsew signal input
flabel metal2 s 52734 0 52790 800 0 FreeSans 224 90 0 0 la_data_in[111]
port 130 nsew signal input
flabel metal2 s 53010 0 53066 800 0 FreeSans 224 90 0 0 la_data_in[112]
port 131 nsew signal input
flabel metal2 s 53286 0 53342 800 0 FreeSans 224 90 0 0 la_data_in[113]
port 132 nsew signal input
flabel metal2 s 53562 0 53618 800 0 FreeSans 224 90 0 0 la_data_in[114]
port 133 nsew signal input
flabel metal2 s 53838 0 53894 800 0 FreeSans 224 90 0 0 la_data_in[115]
port 134 nsew signal input
flabel metal2 s 54114 0 54170 800 0 FreeSans 224 90 0 0 la_data_in[116]
port 135 nsew signal input
flabel metal2 s 54390 0 54446 800 0 FreeSans 224 90 0 0 la_data_in[117]
port 136 nsew signal input
flabel metal2 s 54666 0 54722 800 0 FreeSans 224 90 0 0 la_data_in[118]
port 137 nsew signal input
flabel metal2 s 54942 0 54998 800 0 FreeSans 224 90 0 0 la_data_in[119]
port 138 nsew signal input
flabel metal2 s 25134 0 25190 800 0 FreeSans 224 90 0 0 la_data_in[11]
port 139 nsew signal input
flabel metal2 s 55218 0 55274 800 0 FreeSans 224 90 0 0 la_data_in[120]
port 140 nsew signal input
flabel metal2 s 55494 0 55550 800 0 FreeSans 224 90 0 0 la_data_in[121]
port 141 nsew signal input
flabel metal2 s 55770 0 55826 800 0 FreeSans 224 90 0 0 la_data_in[122]
port 142 nsew signal input
flabel metal2 s 56046 0 56102 800 0 FreeSans 224 90 0 0 la_data_in[123]
port 143 nsew signal input
flabel metal2 s 56322 0 56378 800 0 FreeSans 224 90 0 0 la_data_in[124]
port 144 nsew signal input
flabel metal2 s 56598 0 56654 800 0 FreeSans 224 90 0 0 la_data_in[125]
port 145 nsew signal input
flabel metal2 s 56874 0 56930 800 0 FreeSans 224 90 0 0 la_data_in[126]
port 146 nsew signal input
flabel metal2 s 57150 0 57206 800 0 FreeSans 224 90 0 0 la_data_in[127]
port 147 nsew signal input
flabel metal2 s 25410 0 25466 800 0 FreeSans 224 90 0 0 la_data_in[12]
port 148 nsew signal input
flabel metal2 s 25686 0 25742 800 0 FreeSans 224 90 0 0 la_data_in[13]
port 149 nsew signal input
flabel metal2 s 25962 0 26018 800 0 FreeSans 224 90 0 0 la_data_in[14]
port 150 nsew signal input
flabel metal2 s 26238 0 26294 800 0 FreeSans 224 90 0 0 la_data_in[15]
port 151 nsew signal input
flabel metal2 s 26514 0 26570 800 0 FreeSans 224 90 0 0 la_data_in[16]
port 152 nsew signal input
flabel metal2 s 26790 0 26846 800 0 FreeSans 224 90 0 0 la_data_in[17]
port 153 nsew signal input
flabel metal2 s 27066 0 27122 800 0 FreeSans 224 90 0 0 la_data_in[18]
port 154 nsew signal input
flabel metal2 s 27342 0 27398 800 0 FreeSans 224 90 0 0 la_data_in[19]
port 155 nsew signal input
flabel metal2 s 22374 0 22430 800 0 FreeSans 224 90 0 0 la_data_in[1]
port 156 nsew signal input
flabel metal2 s 27618 0 27674 800 0 FreeSans 224 90 0 0 la_data_in[20]
port 157 nsew signal input
flabel metal2 s 27894 0 27950 800 0 FreeSans 224 90 0 0 la_data_in[21]
port 158 nsew signal input
flabel metal2 s 28170 0 28226 800 0 FreeSans 224 90 0 0 la_data_in[22]
port 159 nsew signal input
flabel metal2 s 28446 0 28502 800 0 FreeSans 224 90 0 0 la_data_in[23]
port 160 nsew signal input
flabel metal2 s 28722 0 28778 800 0 FreeSans 224 90 0 0 la_data_in[24]
port 161 nsew signal input
flabel metal2 s 28998 0 29054 800 0 FreeSans 224 90 0 0 la_data_in[25]
port 162 nsew signal input
flabel metal2 s 29274 0 29330 800 0 FreeSans 224 90 0 0 la_data_in[26]
port 163 nsew signal input
flabel metal2 s 29550 0 29606 800 0 FreeSans 224 90 0 0 la_data_in[27]
port 164 nsew signal input
flabel metal2 s 29826 0 29882 800 0 FreeSans 224 90 0 0 la_data_in[28]
port 165 nsew signal input
flabel metal2 s 30102 0 30158 800 0 FreeSans 224 90 0 0 la_data_in[29]
port 166 nsew signal input
flabel metal2 s 22650 0 22706 800 0 FreeSans 224 90 0 0 la_data_in[2]
port 167 nsew signal input
flabel metal2 s 30378 0 30434 800 0 FreeSans 224 90 0 0 la_data_in[30]
port 168 nsew signal input
flabel metal2 s 30654 0 30710 800 0 FreeSans 224 90 0 0 la_data_in[31]
port 169 nsew signal input
flabel metal2 s 30930 0 30986 800 0 FreeSans 224 90 0 0 la_data_in[32]
port 170 nsew signal input
flabel metal2 s 31206 0 31262 800 0 FreeSans 224 90 0 0 la_data_in[33]
port 171 nsew signal input
flabel metal2 s 31482 0 31538 800 0 FreeSans 224 90 0 0 la_data_in[34]
port 172 nsew signal input
flabel metal2 s 31758 0 31814 800 0 FreeSans 224 90 0 0 la_data_in[35]
port 173 nsew signal input
flabel metal2 s 32034 0 32090 800 0 FreeSans 224 90 0 0 la_data_in[36]
port 174 nsew signal input
flabel metal2 s 32310 0 32366 800 0 FreeSans 224 90 0 0 la_data_in[37]
port 175 nsew signal input
flabel metal2 s 32586 0 32642 800 0 FreeSans 224 90 0 0 la_data_in[38]
port 176 nsew signal input
flabel metal2 s 32862 0 32918 800 0 FreeSans 224 90 0 0 la_data_in[39]
port 177 nsew signal input
flabel metal2 s 22926 0 22982 800 0 FreeSans 224 90 0 0 la_data_in[3]
port 178 nsew signal input
flabel metal2 s 33138 0 33194 800 0 FreeSans 224 90 0 0 la_data_in[40]
port 179 nsew signal input
flabel metal2 s 33414 0 33470 800 0 FreeSans 224 90 0 0 la_data_in[41]
port 180 nsew signal input
flabel metal2 s 33690 0 33746 800 0 FreeSans 224 90 0 0 la_data_in[42]
port 181 nsew signal input
flabel metal2 s 33966 0 34022 800 0 FreeSans 224 90 0 0 la_data_in[43]
port 182 nsew signal input
flabel metal2 s 34242 0 34298 800 0 FreeSans 224 90 0 0 la_data_in[44]
port 183 nsew signal input
flabel metal2 s 34518 0 34574 800 0 FreeSans 224 90 0 0 la_data_in[45]
port 184 nsew signal input
flabel metal2 s 34794 0 34850 800 0 FreeSans 224 90 0 0 la_data_in[46]
port 185 nsew signal input
flabel metal2 s 35070 0 35126 800 0 FreeSans 224 90 0 0 la_data_in[47]
port 186 nsew signal input
flabel metal2 s 35346 0 35402 800 0 FreeSans 224 90 0 0 la_data_in[48]
port 187 nsew signal input
flabel metal2 s 35622 0 35678 800 0 FreeSans 224 90 0 0 la_data_in[49]
port 188 nsew signal input
flabel metal2 s 23202 0 23258 800 0 FreeSans 224 90 0 0 la_data_in[4]
port 189 nsew signal input
flabel metal2 s 35898 0 35954 800 0 FreeSans 224 90 0 0 la_data_in[50]
port 190 nsew signal input
flabel metal2 s 36174 0 36230 800 0 FreeSans 224 90 0 0 la_data_in[51]
port 191 nsew signal input
flabel metal2 s 36450 0 36506 800 0 FreeSans 224 90 0 0 la_data_in[52]
port 192 nsew signal input
flabel metal2 s 36726 0 36782 800 0 FreeSans 224 90 0 0 la_data_in[53]
port 193 nsew signal input
flabel metal2 s 37002 0 37058 800 0 FreeSans 224 90 0 0 la_data_in[54]
port 194 nsew signal input
flabel metal2 s 37278 0 37334 800 0 FreeSans 224 90 0 0 la_data_in[55]
port 195 nsew signal input
flabel metal2 s 37554 0 37610 800 0 FreeSans 224 90 0 0 la_data_in[56]
port 196 nsew signal input
flabel metal2 s 37830 0 37886 800 0 FreeSans 224 90 0 0 la_data_in[57]
port 197 nsew signal input
flabel metal2 s 38106 0 38162 800 0 FreeSans 224 90 0 0 la_data_in[58]
port 198 nsew signal input
flabel metal2 s 38382 0 38438 800 0 FreeSans 224 90 0 0 la_data_in[59]
port 199 nsew signal input
flabel metal2 s 23478 0 23534 800 0 FreeSans 224 90 0 0 la_data_in[5]
port 200 nsew signal input
flabel metal2 s 38658 0 38714 800 0 FreeSans 224 90 0 0 la_data_in[60]
port 201 nsew signal input
flabel metal2 s 38934 0 38990 800 0 FreeSans 224 90 0 0 la_data_in[61]
port 202 nsew signal input
flabel metal2 s 39210 0 39266 800 0 FreeSans 224 90 0 0 la_data_in[62]
port 203 nsew signal input
flabel metal2 s 39486 0 39542 800 0 FreeSans 224 90 0 0 la_data_in[63]
port 204 nsew signal input
flabel metal2 s 39762 0 39818 800 0 FreeSans 224 90 0 0 la_data_in[64]
port 205 nsew signal input
flabel metal2 s 40038 0 40094 800 0 FreeSans 224 90 0 0 la_data_in[65]
port 206 nsew signal input
flabel metal2 s 40314 0 40370 800 0 FreeSans 224 90 0 0 la_data_in[66]
port 207 nsew signal input
flabel metal2 s 40590 0 40646 800 0 FreeSans 224 90 0 0 la_data_in[67]
port 208 nsew signal input
flabel metal2 s 40866 0 40922 800 0 FreeSans 224 90 0 0 la_data_in[68]
port 209 nsew signal input
flabel metal2 s 41142 0 41198 800 0 FreeSans 224 90 0 0 la_data_in[69]
port 210 nsew signal input
flabel metal2 s 23754 0 23810 800 0 FreeSans 224 90 0 0 la_data_in[6]
port 211 nsew signal input
flabel metal2 s 41418 0 41474 800 0 FreeSans 224 90 0 0 la_data_in[70]
port 212 nsew signal input
flabel metal2 s 41694 0 41750 800 0 FreeSans 224 90 0 0 la_data_in[71]
port 213 nsew signal input
flabel metal2 s 41970 0 42026 800 0 FreeSans 224 90 0 0 la_data_in[72]
port 214 nsew signal input
flabel metal2 s 42246 0 42302 800 0 FreeSans 224 90 0 0 la_data_in[73]
port 215 nsew signal input
flabel metal2 s 42522 0 42578 800 0 FreeSans 224 90 0 0 la_data_in[74]
port 216 nsew signal input
flabel metal2 s 42798 0 42854 800 0 FreeSans 224 90 0 0 la_data_in[75]
port 217 nsew signal input
flabel metal2 s 43074 0 43130 800 0 FreeSans 224 90 0 0 la_data_in[76]
port 218 nsew signal input
flabel metal2 s 43350 0 43406 800 0 FreeSans 224 90 0 0 la_data_in[77]
port 219 nsew signal input
flabel metal2 s 43626 0 43682 800 0 FreeSans 224 90 0 0 la_data_in[78]
port 220 nsew signal input
flabel metal2 s 43902 0 43958 800 0 FreeSans 224 90 0 0 la_data_in[79]
port 221 nsew signal input
flabel metal2 s 24030 0 24086 800 0 FreeSans 224 90 0 0 la_data_in[7]
port 222 nsew signal input
flabel metal2 s 44178 0 44234 800 0 FreeSans 224 90 0 0 la_data_in[80]
port 223 nsew signal input
flabel metal2 s 44454 0 44510 800 0 FreeSans 224 90 0 0 la_data_in[81]
port 224 nsew signal input
flabel metal2 s 44730 0 44786 800 0 FreeSans 224 90 0 0 la_data_in[82]
port 225 nsew signal input
flabel metal2 s 45006 0 45062 800 0 FreeSans 224 90 0 0 la_data_in[83]
port 226 nsew signal input
flabel metal2 s 45282 0 45338 800 0 FreeSans 224 90 0 0 la_data_in[84]
port 227 nsew signal input
flabel metal2 s 45558 0 45614 800 0 FreeSans 224 90 0 0 la_data_in[85]
port 228 nsew signal input
flabel metal2 s 45834 0 45890 800 0 FreeSans 224 90 0 0 la_data_in[86]
port 229 nsew signal input
flabel metal2 s 46110 0 46166 800 0 FreeSans 224 90 0 0 la_data_in[87]
port 230 nsew signal input
flabel metal2 s 46386 0 46442 800 0 FreeSans 224 90 0 0 la_data_in[88]
port 231 nsew signal input
flabel metal2 s 46662 0 46718 800 0 FreeSans 224 90 0 0 la_data_in[89]
port 232 nsew signal input
flabel metal2 s 24306 0 24362 800 0 FreeSans 224 90 0 0 la_data_in[8]
port 233 nsew signal input
flabel metal2 s 46938 0 46994 800 0 FreeSans 224 90 0 0 la_data_in[90]
port 234 nsew signal input
flabel metal2 s 47214 0 47270 800 0 FreeSans 224 90 0 0 la_data_in[91]
port 235 nsew signal input
flabel metal2 s 47490 0 47546 800 0 FreeSans 224 90 0 0 la_data_in[92]
port 236 nsew signal input
flabel metal2 s 47766 0 47822 800 0 FreeSans 224 90 0 0 la_data_in[93]
port 237 nsew signal input
flabel metal2 s 48042 0 48098 800 0 FreeSans 224 90 0 0 la_data_in[94]
port 238 nsew signal input
flabel metal2 s 48318 0 48374 800 0 FreeSans 224 90 0 0 la_data_in[95]
port 239 nsew signal input
flabel metal2 s 48594 0 48650 800 0 FreeSans 224 90 0 0 la_data_in[96]
port 240 nsew signal input
flabel metal2 s 48870 0 48926 800 0 FreeSans 224 90 0 0 la_data_in[97]
port 241 nsew signal input
flabel metal2 s 49146 0 49202 800 0 FreeSans 224 90 0 0 la_data_in[98]
port 242 nsew signal input
flabel metal2 s 49422 0 49478 800 0 FreeSans 224 90 0 0 la_data_in[99]
port 243 nsew signal input
flabel metal2 s 24582 0 24638 800 0 FreeSans 224 90 0 0 la_data_in[9]
port 244 nsew signal input
flabel metal2 s 22190 0 22246 800 0 FreeSans 224 90 0 0 la_data_out[0]
port 245 nsew signal tristate
flabel metal2 s 49790 0 49846 800 0 FreeSans 224 90 0 0 la_data_out[100]
port 246 nsew signal tristate
flabel metal2 s 50066 0 50122 800 0 FreeSans 224 90 0 0 la_data_out[101]
port 247 nsew signal tristate
flabel metal2 s 50342 0 50398 800 0 FreeSans 224 90 0 0 la_data_out[102]
port 248 nsew signal tristate
flabel metal2 s 50618 0 50674 800 0 FreeSans 224 90 0 0 la_data_out[103]
port 249 nsew signal tristate
flabel metal2 s 50894 0 50950 800 0 FreeSans 224 90 0 0 la_data_out[104]
port 250 nsew signal tristate
flabel metal2 s 51170 0 51226 800 0 FreeSans 224 90 0 0 la_data_out[105]
port 251 nsew signal tristate
flabel metal2 s 51446 0 51502 800 0 FreeSans 224 90 0 0 la_data_out[106]
port 252 nsew signal tristate
flabel metal2 s 51722 0 51778 800 0 FreeSans 224 90 0 0 la_data_out[107]
port 253 nsew signal tristate
flabel metal2 s 51998 0 52054 800 0 FreeSans 224 90 0 0 la_data_out[108]
port 254 nsew signal tristate
flabel metal2 s 52274 0 52330 800 0 FreeSans 224 90 0 0 la_data_out[109]
port 255 nsew signal tristate
flabel metal2 s 24950 0 25006 800 0 FreeSans 224 90 0 0 la_data_out[10]
port 256 nsew signal tristate
flabel metal2 s 52550 0 52606 800 0 FreeSans 224 90 0 0 la_data_out[110]
port 257 nsew signal tristate
flabel metal2 s 52826 0 52882 800 0 FreeSans 224 90 0 0 la_data_out[111]
port 258 nsew signal tristate
flabel metal2 s 53102 0 53158 800 0 FreeSans 224 90 0 0 la_data_out[112]
port 259 nsew signal tristate
flabel metal2 s 53378 0 53434 800 0 FreeSans 224 90 0 0 la_data_out[113]
port 260 nsew signal tristate
flabel metal2 s 53654 0 53710 800 0 FreeSans 224 90 0 0 la_data_out[114]
port 261 nsew signal tristate
flabel metal2 s 53930 0 53986 800 0 FreeSans 224 90 0 0 la_data_out[115]
port 262 nsew signal tristate
flabel metal2 s 54206 0 54262 800 0 FreeSans 224 90 0 0 la_data_out[116]
port 263 nsew signal tristate
flabel metal2 s 54482 0 54538 800 0 FreeSans 224 90 0 0 la_data_out[117]
port 264 nsew signal tristate
flabel metal2 s 54758 0 54814 800 0 FreeSans 224 90 0 0 la_data_out[118]
port 265 nsew signal tristate
flabel metal2 s 55034 0 55090 800 0 FreeSans 224 90 0 0 la_data_out[119]
port 266 nsew signal tristate
flabel metal2 s 25226 0 25282 800 0 FreeSans 224 90 0 0 la_data_out[11]
port 267 nsew signal tristate
flabel metal2 s 55310 0 55366 800 0 FreeSans 224 90 0 0 la_data_out[120]
port 268 nsew signal tristate
flabel metal2 s 55586 0 55642 800 0 FreeSans 224 90 0 0 la_data_out[121]
port 269 nsew signal tristate
flabel metal2 s 55862 0 55918 800 0 FreeSans 224 90 0 0 la_data_out[122]
port 270 nsew signal tristate
flabel metal2 s 56138 0 56194 800 0 FreeSans 224 90 0 0 la_data_out[123]
port 271 nsew signal tristate
flabel metal2 s 56414 0 56470 800 0 FreeSans 224 90 0 0 la_data_out[124]
port 272 nsew signal tristate
flabel metal2 s 56690 0 56746 800 0 FreeSans 224 90 0 0 la_data_out[125]
port 273 nsew signal tristate
flabel metal2 s 56966 0 57022 800 0 FreeSans 224 90 0 0 la_data_out[126]
port 274 nsew signal tristate
flabel metal2 s 57242 0 57298 800 0 FreeSans 224 90 0 0 la_data_out[127]
port 275 nsew signal tristate
flabel metal2 s 25502 0 25558 800 0 FreeSans 224 90 0 0 la_data_out[12]
port 276 nsew signal tristate
flabel metal2 s 25778 0 25834 800 0 FreeSans 224 90 0 0 la_data_out[13]
port 277 nsew signal tristate
flabel metal2 s 26054 0 26110 800 0 FreeSans 224 90 0 0 la_data_out[14]
port 278 nsew signal tristate
flabel metal2 s 26330 0 26386 800 0 FreeSans 224 90 0 0 la_data_out[15]
port 279 nsew signal tristate
flabel metal2 s 26606 0 26662 800 0 FreeSans 224 90 0 0 la_data_out[16]
port 280 nsew signal tristate
flabel metal2 s 26882 0 26938 800 0 FreeSans 224 90 0 0 la_data_out[17]
port 281 nsew signal tristate
flabel metal2 s 27158 0 27214 800 0 FreeSans 224 90 0 0 la_data_out[18]
port 282 nsew signal tristate
flabel metal2 s 27434 0 27490 800 0 FreeSans 224 90 0 0 la_data_out[19]
port 283 nsew signal tristate
flabel metal2 s 22466 0 22522 800 0 FreeSans 224 90 0 0 la_data_out[1]
port 284 nsew signal tristate
flabel metal2 s 27710 0 27766 800 0 FreeSans 224 90 0 0 la_data_out[20]
port 285 nsew signal tristate
flabel metal2 s 27986 0 28042 800 0 FreeSans 224 90 0 0 la_data_out[21]
port 286 nsew signal tristate
flabel metal2 s 28262 0 28318 800 0 FreeSans 224 90 0 0 la_data_out[22]
port 287 nsew signal tristate
flabel metal2 s 28538 0 28594 800 0 FreeSans 224 90 0 0 la_data_out[23]
port 288 nsew signal tristate
flabel metal2 s 28814 0 28870 800 0 FreeSans 224 90 0 0 la_data_out[24]
port 289 nsew signal tristate
flabel metal2 s 29090 0 29146 800 0 FreeSans 224 90 0 0 la_data_out[25]
port 290 nsew signal tristate
flabel metal2 s 29366 0 29422 800 0 FreeSans 224 90 0 0 la_data_out[26]
port 291 nsew signal tristate
flabel metal2 s 29642 0 29698 800 0 FreeSans 224 90 0 0 la_data_out[27]
port 292 nsew signal tristate
flabel metal2 s 29918 0 29974 800 0 FreeSans 224 90 0 0 la_data_out[28]
port 293 nsew signal tristate
flabel metal2 s 30194 0 30250 800 0 FreeSans 224 90 0 0 la_data_out[29]
port 294 nsew signal tristate
flabel metal2 s 22742 0 22798 800 0 FreeSans 224 90 0 0 la_data_out[2]
port 295 nsew signal tristate
flabel metal2 s 30470 0 30526 800 0 FreeSans 224 90 0 0 la_data_out[30]
port 296 nsew signal tristate
flabel metal2 s 30746 0 30802 800 0 FreeSans 224 90 0 0 la_data_out[31]
port 297 nsew signal tristate
flabel metal2 s 31022 0 31078 800 0 FreeSans 224 90 0 0 la_data_out[32]
port 298 nsew signal tristate
flabel metal2 s 31298 0 31354 800 0 FreeSans 224 90 0 0 la_data_out[33]
port 299 nsew signal tristate
flabel metal2 s 31574 0 31630 800 0 FreeSans 224 90 0 0 la_data_out[34]
port 300 nsew signal tristate
flabel metal2 s 31850 0 31906 800 0 FreeSans 224 90 0 0 la_data_out[35]
port 301 nsew signal tristate
flabel metal2 s 32126 0 32182 800 0 FreeSans 224 90 0 0 la_data_out[36]
port 302 nsew signal tristate
flabel metal2 s 32402 0 32458 800 0 FreeSans 224 90 0 0 la_data_out[37]
port 303 nsew signal tristate
flabel metal2 s 32678 0 32734 800 0 FreeSans 224 90 0 0 la_data_out[38]
port 304 nsew signal tristate
flabel metal2 s 32954 0 33010 800 0 FreeSans 224 90 0 0 la_data_out[39]
port 305 nsew signal tristate
flabel metal2 s 23018 0 23074 800 0 FreeSans 224 90 0 0 la_data_out[3]
port 306 nsew signal tristate
flabel metal2 s 33230 0 33286 800 0 FreeSans 224 90 0 0 la_data_out[40]
port 307 nsew signal tristate
flabel metal2 s 33506 0 33562 800 0 FreeSans 224 90 0 0 la_data_out[41]
port 308 nsew signal tristate
flabel metal2 s 33782 0 33838 800 0 FreeSans 224 90 0 0 la_data_out[42]
port 309 nsew signal tristate
flabel metal2 s 34058 0 34114 800 0 FreeSans 224 90 0 0 la_data_out[43]
port 310 nsew signal tristate
flabel metal2 s 34334 0 34390 800 0 FreeSans 224 90 0 0 la_data_out[44]
port 311 nsew signal tristate
flabel metal2 s 34610 0 34666 800 0 FreeSans 224 90 0 0 la_data_out[45]
port 312 nsew signal tristate
flabel metal2 s 34886 0 34942 800 0 FreeSans 224 90 0 0 la_data_out[46]
port 313 nsew signal tristate
flabel metal2 s 35162 0 35218 800 0 FreeSans 224 90 0 0 la_data_out[47]
port 314 nsew signal tristate
flabel metal2 s 35438 0 35494 800 0 FreeSans 224 90 0 0 la_data_out[48]
port 315 nsew signal tristate
flabel metal2 s 35714 0 35770 800 0 FreeSans 224 90 0 0 la_data_out[49]
port 316 nsew signal tristate
flabel metal2 s 23294 0 23350 800 0 FreeSans 224 90 0 0 la_data_out[4]
port 317 nsew signal tristate
flabel metal2 s 35990 0 36046 800 0 FreeSans 224 90 0 0 la_data_out[50]
port 318 nsew signal tristate
flabel metal2 s 36266 0 36322 800 0 FreeSans 224 90 0 0 la_data_out[51]
port 319 nsew signal tristate
flabel metal2 s 36542 0 36598 800 0 FreeSans 224 90 0 0 la_data_out[52]
port 320 nsew signal tristate
flabel metal2 s 36818 0 36874 800 0 FreeSans 224 90 0 0 la_data_out[53]
port 321 nsew signal tristate
flabel metal2 s 37094 0 37150 800 0 FreeSans 224 90 0 0 la_data_out[54]
port 322 nsew signal tristate
flabel metal2 s 37370 0 37426 800 0 FreeSans 224 90 0 0 la_data_out[55]
port 323 nsew signal tristate
flabel metal2 s 37646 0 37702 800 0 FreeSans 224 90 0 0 la_data_out[56]
port 324 nsew signal tristate
flabel metal2 s 37922 0 37978 800 0 FreeSans 224 90 0 0 la_data_out[57]
port 325 nsew signal tristate
flabel metal2 s 38198 0 38254 800 0 FreeSans 224 90 0 0 la_data_out[58]
port 326 nsew signal tristate
flabel metal2 s 38474 0 38530 800 0 FreeSans 224 90 0 0 la_data_out[59]
port 327 nsew signal tristate
flabel metal2 s 23570 0 23626 800 0 FreeSans 224 90 0 0 la_data_out[5]
port 328 nsew signal tristate
flabel metal2 s 38750 0 38806 800 0 FreeSans 224 90 0 0 la_data_out[60]
port 329 nsew signal tristate
flabel metal2 s 39026 0 39082 800 0 FreeSans 224 90 0 0 la_data_out[61]
port 330 nsew signal tristate
flabel metal2 s 39302 0 39358 800 0 FreeSans 224 90 0 0 la_data_out[62]
port 331 nsew signal tristate
flabel metal2 s 39578 0 39634 800 0 FreeSans 224 90 0 0 la_data_out[63]
port 332 nsew signal tristate
flabel metal2 s 39854 0 39910 800 0 FreeSans 224 90 0 0 la_data_out[64]
port 333 nsew signal tristate
flabel metal2 s 40130 0 40186 800 0 FreeSans 224 90 0 0 la_data_out[65]
port 334 nsew signal tristate
flabel metal2 s 40406 0 40462 800 0 FreeSans 224 90 0 0 la_data_out[66]
port 335 nsew signal tristate
flabel metal2 s 40682 0 40738 800 0 FreeSans 224 90 0 0 la_data_out[67]
port 336 nsew signal tristate
flabel metal2 s 40958 0 41014 800 0 FreeSans 224 90 0 0 la_data_out[68]
port 337 nsew signal tristate
flabel metal2 s 41234 0 41290 800 0 FreeSans 224 90 0 0 la_data_out[69]
port 338 nsew signal tristate
flabel metal2 s 23846 0 23902 800 0 FreeSans 224 90 0 0 la_data_out[6]
port 339 nsew signal tristate
flabel metal2 s 41510 0 41566 800 0 FreeSans 224 90 0 0 la_data_out[70]
port 340 nsew signal tristate
flabel metal2 s 41786 0 41842 800 0 FreeSans 224 90 0 0 la_data_out[71]
port 341 nsew signal tristate
flabel metal2 s 42062 0 42118 800 0 FreeSans 224 90 0 0 la_data_out[72]
port 342 nsew signal tristate
flabel metal2 s 42338 0 42394 800 0 FreeSans 224 90 0 0 la_data_out[73]
port 343 nsew signal tristate
flabel metal2 s 42614 0 42670 800 0 FreeSans 224 90 0 0 la_data_out[74]
port 344 nsew signal tristate
flabel metal2 s 42890 0 42946 800 0 FreeSans 224 90 0 0 la_data_out[75]
port 345 nsew signal tristate
flabel metal2 s 43166 0 43222 800 0 FreeSans 224 90 0 0 la_data_out[76]
port 346 nsew signal tristate
flabel metal2 s 43442 0 43498 800 0 FreeSans 224 90 0 0 la_data_out[77]
port 347 nsew signal tristate
flabel metal2 s 43718 0 43774 800 0 FreeSans 224 90 0 0 la_data_out[78]
port 348 nsew signal tristate
flabel metal2 s 43994 0 44050 800 0 FreeSans 224 90 0 0 la_data_out[79]
port 349 nsew signal tristate
flabel metal2 s 24122 0 24178 800 0 FreeSans 224 90 0 0 la_data_out[7]
port 350 nsew signal tristate
flabel metal2 s 44270 0 44326 800 0 FreeSans 224 90 0 0 la_data_out[80]
port 351 nsew signal tristate
flabel metal2 s 44546 0 44602 800 0 FreeSans 224 90 0 0 la_data_out[81]
port 352 nsew signal tristate
flabel metal2 s 44822 0 44878 800 0 FreeSans 224 90 0 0 la_data_out[82]
port 353 nsew signal tristate
flabel metal2 s 45098 0 45154 800 0 FreeSans 224 90 0 0 la_data_out[83]
port 354 nsew signal tristate
flabel metal2 s 45374 0 45430 800 0 FreeSans 224 90 0 0 la_data_out[84]
port 355 nsew signal tristate
flabel metal2 s 45650 0 45706 800 0 FreeSans 224 90 0 0 la_data_out[85]
port 356 nsew signal tristate
flabel metal2 s 45926 0 45982 800 0 FreeSans 224 90 0 0 la_data_out[86]
port 357 nsew signal tristate
flabel metal2 s 46202 0 46258 800 0 FreeSans 224 90 0 0 la_data_out[87]
port 358 nsew signal tristate
flabel metal2 s 46478 0 46534 800 0 FreeSans 224 90 0 0 la_data_out[88]
port 359 nsew signal tristate
flabel metal2 s 46754 0 46810 800 0 FreeSans 224 90 0 0 la_data_out[89]
port 360 nsew signal tristate
flabel metal2 s 24398 0 24454 800 0 FreeSans 224 90 0 0 la_data_out[8]
port 361 nsew signal tristate
flabel metal2 s 47030 0 47086 800 0 FreeSans 224 90 0 0 la_data_out[90]
port 362 nsew signal tristate
flabel metal2 s 47306 0 47362 800 0 FreeSans 224 90 0 0 la_data_out[91]
port 363 nsew signal tristate
flabel metal2 s 47582 0 47638 800 0 FreeSans 224 90 0 0 la_data_out[92]
port 364 nsew signal tristate
flabel metal2 s 47858 0 47914 800 0 FreeSans 224 90 0 0 la_data_out[93]
port 365 nsew signal tristate
flabel metal2 s 48134 0 48190 800 0 FreeSans 224 90 0 0 la_data_out[94]
port 366 nsew signal tristate
flabel metal2 s 48410 0 48466 800 0 FreeSans 224 90 0 0 la_data_out[95]
port 367 nsew signal tristate
flabel metal2 s 48686 0 48742 800 0 FreeSans 224 90 0 0 la_data_out[96]
port 368 nsew signal tristate
flabel metal2 s 48962 0 49018 800 0 FreeSans 224 90 0 0 la_data_out[97]
port 369 nsew signal tristate
flabel metal2 s 49238 0 49294 800 0 FreeSans 224 90 0 0 la_data_out[98]
port 370 nsew signal tristate
flabel metal2 s 49514 0 49570 800 0 FreeSans 224 90 0 0 la_data_out[99]
port 371 nsew signal tristate
flabel metal2 s 24674 0 24730 800 0 FreeSans 224 90 0 0 la_data_out[9]
port 372 nsew signal tristate
flabel metal2 s 22282 0 22338 800 0 FreeSans 224 90 0 0 la_oenb[0]
port 373 nsew signal input
flabel metal2 s 49882 0 49938 800 0 FreeSans 224 90 0 0 la_oenb[100]
port 374 nsew signal input
flabel metal2 s 50158 0 50214 800 0 FreeSans 224 90 0 0 la_oenb[101]
port 375 nsew signal input
flabel metal2 s 50434 0 50490 800 0 FreeSans 224 90 0 0 la_oenb[102]
port 376 nsew signal input
flabel metal2 s 50710 0 50766 800 0 FreeSans 224 90 0 0 la_oenb[103]
port 377 nsew signal input
flabel metal2 s 50986 0 51042 800 0 FreeSans 224 90 0 0 la_oenb[104]
port 378 nsew signal input
flabel metal2 s 51262 0 51318 800 0 FreeSans 224 90 0 0 la_oenb[105]
port 379 nsew signal input
flabel metal2 s 51538 0 51594 800 0 FreeSans 224 90 0 0 la_oenb[106]
port 380 nsew signal input
flabel metal2 s 51814 0 51870 800 0 FreeSans 224 90 0 0 la_oenb[107]
port 381 nsew signal input
flabel metal2 s 52090 0 52146 800 0 FreeSans 224 90 0 0 la_oenb[108]
port 382 nsew signal input
flabel metal2 s 52366 0 52422 800 0 FreeSans 224 90 0 0 la_oenb[109]
port 383 nsew signal input
flabel metal2 s 25042 0 25098 800 0 FreeSans 224 90 0 0 la_oenb[10]
port 384 nsew signal input
flabel metal2 s 52642 0 52698 800 0 FreeSans 224 90 0 0 la_oenb[110]
port 385 nsew signal input
flabel metal2 s 52918 0 52974 800 0 FreeSans 224 90 0 0 la_oenb[111]
port 386 nsew signal input
flabel metal2 s 53194 0 53250 800 0 FreeSans 224 90 0 0 la_oenb[112]
port 387 nsew signal input
flabel metal2 s 53470 0 53526 800 0 FreeSans 224 90 0 0 la_oenb[113]
port 388 nsew signal input
flabel metal2 s 53746 0 53802 800 0 FreeSans 224 90 0 0 la_oenb[114]
port 389 nsew signal input
flabel metal2 s 54022 0 54078 800 0 FreeSans 224 90 0 0 la_oenb[115]
port 390 nsew signal input
flabel metal2 s 54298 0 54354 800 0 FreeSans 224 90 0 0 la_oenb[116]
port 391 nsew signal input
flabel metal2 s 54574 0 54630 800 0 FreeSans 224 90 0 0 la_oenb[117]
port 392 nsew signal input
flabel metal2 s 54850 0 54906 800 0 FreeSans 224 90 0 0 la_oenb[118]
port 393 nsew signal input
flabel metal2 s 55126 0 55182 800 0 FreeSans 224 90 0 0 la_oenb[119]
port 394 nsew signal input
flabel metal2 s 25318 0 25374 800 0 FreeSans 224 90 0 0 la_oenb[11]
port 395 nsew signal input
flabel metal2 s 55402 0 55458 800 0 FreeSans 224 90 0 0 la_oenb[120]
port 396 nsew signal input
flabel metal2 s 55678 0 55734 800 0 FreeSans 224 90 0 0 la_oenb[121]
port 397 nsew signal input
flabel metal2 s 55954 0 56010 800 0 FreeSans 224 90 0 0 la_oenb[122]
port 398 nsew signal input
flabel metal2 s 56230 0 56286 800 0 FreeSans 224 90 0 0 la_oenb[123]
port 399 nsew signal input
flabel metal2 s 56506 0 56562 800 0 FreeSans 224 90 0 0 la_oenb[124]
port 400 nsew signal input
flabel metal2 s 56782 0 56838 800 0 FreeSans 224 90 0 0 la_oenb[125]
port 401 nsew signal input
flabel metal2 s 57058 0 57114 800 0 FreeSans 224 90 0 0 la_oenb[126]
port 402 nsew signal input
flabel metal2 s 57334 0 57390 800 0 FreeSans 224 90 0 0 la_oenb[127]
port 403 nsew signal input
flabel metal2 s 25594 0 25650 800 0 FreeSans 224 90 0 0 la_oenb[12]
port 404 nsew signal input
flabel metal2 s 25870 0 25926 800 0 FreeSans 224 90 0 0 la_oenb[13]
port 405 nsew signal input
flabel metal2 s 26146 0 26202 800 0 FreeSans 224 90 0 0 la_oenb[14]
port 406 nsew signal input
flabel metal2 s 26422 0 26478 800 0 FreeSans 224 90 0 0 la_oenb[15]
port 407 nsew signal input
flabel metal2 s 26698 0 26754 800 0 FreeSans 224 90 0 0 la_oenb[16]
port 408 nsew signal input
flabel metal2 s 26974 0 27030 800 0 FreeSans 224 90 0 0 la_oenb[17]
port 409 nsew signal input
flabel metal2 s 27250 0 27306 800 0 FreeSans 224 90 0 0 la_oenb[18]
port 410 nsew signal input
flabel metal2 s 27526 0 27582 800 0 FreeSans 224 90 0 0 la_oenb[19]
port 411 nsew signal input
flabel metal2 s 22558 0 22614 800 0 FreeSans 224 90 0 0 la_oenb[1]
port 412 nsew signal input
flabel metal2 s 27802 0 27858 800 0 FreeSans 224 90 0 0 la_oenb[20]
port 413 nsew signal input
flabel metal2 s 28078 0 28134 800 0 FreeSans 224 90 0 0 la_oenb[21]
port 414 nsew signal input
flabel metal2 s 28354 0 28410 800 0 FreeSans 224 90 0 0 la_oenb[22]
port 415 nsew signal input
flabel metal2 s 28630 0 28686 800 0 FreeSans 224 90 0 0 la_oenb[23]
port 416 nsew signal input
flabel metal2 s 28906 0 28962 800 0 FreeSans 224 90 0 0 la_oenb[24]
port 417 nsew signal input
flabel metal2 s 29182 0 29238 800 0 FreeSans 224 90 0 0 la_oenb[25]
port 418 nsew signal input
flabel metal2 s 29458 0 29514 800 0 FreeSans 224 90 0 0 la_oenb[26]
port 419 nsew signal input
flabel metal2 s 29734 0 29790 800 0 FreeSans 224 90 0 0 la_oenb[27]
port 420 nsew signal input
flabel metal2 s 30010 0 30066 800 0 FreeSans 224 90 0 0 la_oenb[28]
port 421 nsew signal input
flabel metal2 s 30286 0 30342 800 0 FreeSans 224 90 0 0 la_oenb[29]
port 422 nsew signal input
flabel metal2 s 22834 0 22890 800 0 FreeSans 224 90 0 0 la_oenb[2]
port 423 nsew signal input
flabel metal2 s 30562 0 30618 800 0 FreeSans 224 90 0 0 la_oenb[30]
port 424 nsew signal input
flabel metal2 s 30838 0 30894 800 0 FreeSans 224 90 0 0 la_oenb[31]
port 425 nsew signal input
flabel metal2 s 31114 0 31170 800 0 FreeSans 224 90 0 0 la_oenb[32]
port 426 nsew signal input
flabel metal2 s 31390 0 31446 800 0 FreeSans 224 90 0 0 la_oenb[33]
port 427 nsew signal input
flabel metal2 s 31666 0 31722 800 0 FreeSans 224 90 0 0 la_oenb[34]
port 428 nsew signal input
flabel metal2 s 31942 0 31998 800 0 FreeSans 224 90 0 0 la_oenb[35]
port 429 nsew signal input
flabel metal2 s 32218 0 32274 800 0 FreeSans 224 90 0 0 la_oenb[36]
port 430 nsew signal input
flabel metal2 s 32494 0 32550 800 0 FreeSans 224 90 0 0 la_oenb[37]
port 431 nsew signal input
flabel metal2 s 32770 0 32826 800 0 FreeSans 224 90 0 0 la_oenb[38]
port 432 nsew signal input
flabel metal2 s 33046 0 33102 800 0 FreeSans 224 90 0 0 la_oenb[39]
port 433 nsew signal input
flabel metal2 s 23110 0 23166 800 0 FreeSans 224 90 0 0 la_oenb[3]
port 434 nsew signal input
flabel metal2 s 33322 0 33378 800 0 FreeSans 224 90 0 0 la_oenb[40]
port 435 nsew signal input
flabel metal2 s 33598 0 33654 800 0 FreeSans 224 90 0 0 la_oenb[41]
port 436 nsew signal input
flabel metal2 s 33874 0 33930 800 0 FreeSans 224 90 0 0 la_oenb[42]
port 437 nsew signal input
flabel metal2 s 34150 0 34206 800 0 FreeSans 224 90 0 0 la_oenb[43]
port 438 nsew signal input
flabel metal2 s 34426 0 34482 800 0 FreeSans 224 90 0 0 la_oenb[44]
port 439 nsew signal input
flabel metal2 s 34702 0 34758 800 0 FreeSans 224 90 0 0 la_oenb[45]
port 440 nsew signal input
flabel metal2 s 34978 0 35034 800 0 FreeSans 224 90 0 0 la_oenb[46]
port 441 nsew signal input
flabel metal2 s 35254 0 35310 800 0 FreeSans 224 90 0 0 la_oenb[47]
port 442 nsew signal input
flabel metal2 s 35530 0 35586 800 0 FreeSans 224 90 0 0 la_oenb[48]
port 443 nsew signal input
flabel metal2 s 35806 0 35862 800 0 FreeSans 224 90 0 0 la_oenb[49]
port 444 nsew signal input
flabel metal2 s 23386 0 23442 800 0 FreeSans 224 90 0 0 la_oenb[4]
port 445 nsew signal input
flabel metal2 s 36082 0 36138 800 0 FreeSans 224 90 0 0 la_oenb[50]
port 446 nsew signal input
flabel metal2 s 36358 0 36414 800 0 FreeSans 224 90 0 0 la_oenb[51]
port 447 nsew signal input
flabel metal2 s 36634 0 36690 800 0 FreeSans 224 90 0 0 la_oenb[52]
port 448 nsew signal input
flabel metal2 s 36910 0 36966 800 0 FreeSans 224 90 0 0 la_oenb[53]
port 449 nsew signal input
flabel metal2 s 37186 0 37242 800 0 FreeSans 224 90 0 0 la_oenb[54]
port 450 nsew signal input
flabel metal2 s 37462 0 37518 800 0 FreeSans 224 90 0 0 la_oenb[55]
port 451 nsew signal input
flabel metal2 s 37738 0 37794 800 0 FreeSans 224 90 0 0 la_oenb[56]
port 452 nsew signal input
flabel metal2 s 38014 0 38070 800 0 FreeSans 224 90 0 0 la_oenb[57]
port 453 nsew signal input
flabel metal2 s 38290 0 38346 800 0 FreeSans 224 90 0 0 la_oenb[58]
port 454 nsew signal input
flabel metal2 s 38566 0 38622 800 0 FreeSans 224 90 0 0 la_oenb[59]
port 455 nsew signal input
flabel metal2 s 23662 0 23718 800 0 FreeSans 224 90 0 0 la_oenb[5]
port 456 nsew signal input
flabel metal2 s 38842 0 38898 800 0 FreeSans 224 90 0 0 la_oenb[60]
port 457 nsew signal input
flabel metal2 s 39118 0 39174 800 0 FreeSans 224 90 0 0 la_oenb[61]
port 458 nsew signal input
flabel metal2 s 39394 0 39450 800 0 FreeSans 224 90 0 0 la_oenb[62]
port 459 nsew signal input
flabel metal2 s 39670 0 39726 800 0 FreeSans 224 90 0 0 la_oenb[63]
port 460 nsew signal input
flabel metal2 s 39946 0 40002 800 0 FreeSans 224 90 0 0 la_oenb[64]
port 461 nsew signal input
flabel metal2 s 40222 0 40278 800 0 FreeSans 224 90 0 0 la_oenb[65]
port 462 nsew signal input
flabel metal2 s 40498 0 40554 800 0 FreeSans 224 90 0 0 la_oenb[66]
port 463 nsew signal input
flabel metal2 s 40774 0 40830 800 0 FreeSans 224 90 0 0 la_oenb[67]
port 464 nsew signal input
flabel metal2 s 41050 0 41106 800 0 FreeSans 224 90 0 0 la_oenb[68]
port 465 nsew signal input
flabel metal2 s 41326 0 41382 800 0 FreeSans 224 90 0 0 la_oenb[69]
port 466 nsew signal input
flabel metal2 s 23938 0 23994 800 0 FreeSans 224 90 0 0 la_oenb[6]
port 467 nsew signal input
flabel metal2 s 41602 0 41658 800 0 FreeSans 224 90 0 0 la_oenb[70]
port 468 nsew signal input
flabel metal2 s 41878 0 41934 800 0 FreeSans 224 90 0 0 la_oenb[71]
port 469 nsew signal input
flabel metal2 s 42154 0 42210 800 0 FreeSans 224 90 0 0 la_oenb[72]
port 470 nsew signal input
flabel metal2 s 42430 0 42486 800 0 FreeSans 224 90 0 0 la_oenb[73]
port 471 nsew signal input
flabel metal2 s 42706 0 42762 800 0 FreeSans 224 90 0 0 la_oenb[74]
port 472 nsew signal input
flabel metal2 s 42982 0 43038 800 0 FreeSans 224 90 0 0 la_oenb[75]
port 473 nsew signal input
flabel metal2 s 43258 0 43314 800 0 FreeSans 224 90 0 0 la_oenb[76]
port 474 nsew signal input
flabel metal2 s 43534 0 43590 800 0 FreeSans 224 90 0 0 la_oenb[77]
port 475 nsew signal input
flabel metal2 s 43810 0 43866 800 0 FreeSans 224 90 0 0 la_oenb[78]
port 476 nsew signal input
flabel metal2 s 44086 0 44142 800 0 FreeSans 224 90 0 0 la_oenb[79]
port 477 nsew signal input
flabel metal2 s 24214 0 24270 800 0 FreeSans 224 90 0 0 la_oenb[7]
port 478 nsew signal input
flabel metal2 s 44362 0 44418 800 0 FreeSans 224 90 0 0 la_oenb[80]
port 479 nsew signal input
flabel metal2 s 44638 0 44694 800 0 FreeSans 224 90 0 0 la_oenb[81]
port 480 nsew signal input
flabel metal2 s 44914 0 44970 800 0 FreeSans 224 90 0 0 la_oenb[82]
port 481 nsew signal input
flabel metal2 s 45190 0 45246 800 0 FreeSans 224 90 0 0 la_oenb[83]
port 482 nsew signal input
flabel metal2 s 45466 0 45522 800 0 FreeSans 224 90 0 0 la_oenb[84]
port 483 nsew signal input
flabel metal2 s 45742 0 45798 800 0 FreeSans 224 90 0 0 la_oenb[85]
port 484 nsew signal input
flabel metal2 s 46018 0 46074 800 0 FreeSans 224 90 0 0 la_oenb[86]
port 485 nsew signal input
flabel metal2 s 46294 0 46350 800 0 FreeSans 224 90 0 0 la_oenb[87]
port 486 nsew signal input
flabel metal2 s 46570 0 46626 800 0 FreeSans 224 90 0 0 la_oenb[88]
port 487 nsew signal input
flabel metal2 s 46846 0 46902 800 0 FreeSans 224 90 0 0 la_oenb[89]
port 488 nsew signal input
flabel metal2 s 24490 0 24546 800 0 FreeSans 224 90 0 0 la_oenb[8]
port 489 nsew signal input
flabel metal2 s 47122 0 47178 800 0 FreeSans 224 90 0 0 la_oenb[90]
port 490 nsew signal input
flabel metal2 s 47398 0 47454 800 0 FreeSans 224 90 0 0 la_oenb[91]
port 491 nsew signal input
flabel metal2 s 47674 0 47730 800 0 FreeSans 224 90 0 0 la_oenb[92]
port 492 nsew signal input
flabel metal2 s 47950 0 48006 800 0 FreeSans 224 90 0 0 la_oenb[93]
port 493 nsew signal input
flabel metal2 s 48226 0 48282 800 0 FreeSans 224 90 0 0 la_oenb[94]
port 494 nsew signal input
flabel metal2 s 48502 0 48558 800 0 FreeSans 224 90 0 0 la_oenb[95]
port 495 nsew signal input
flabel metal2 s 48778 0 48834 800 0 FreeSans 224 90 0 0 la_oenb[96]
port 496 nsew signal input
flabel metal2 s 49054 0 49110 800 0 FreeSans 224 90 0 0 la_oenb[97]
port 497 nsew signal input
flabel metal2 s 49330 0 49386 800 0 FreeSans 224 90 0 0 la_oenb[98]
port 498 nsew signal input
flabel metal2 s 49606 0 49662 800 0 FreeSans 224 90 0 0 la_oenb[99]
port 499 nsew signal input
flabel metal2 s 24766 0 24822 800 0 FreeSans 224 90 0 0 la_oenb[9]
port 500 nsew signal input
flabel metal2 s 66994 59200 67050 60000 0 FreeSans 224 90 0 0 pxl_done
port 501 nsew signal tristate
flabel metal2 s 65890 59200 65946 60000 0 FreeSans 224 90 0 0 pxl_start_in_ext
port 502 nsew signal input
flabel metal2 s 66442 59200 66498 60000 0 FreeSans 224 90 0 0 pxl_start_out
port 503 nsew signal input
flabel metal4 s 4208 2128 4528 57712 0 FreeSans 1920 90 0 0 vccd1
port 504 nsew power bidirectional
flabel metal4 s 34928 2128 35248 57712 0 FreeSans 1920 90 0 0 vccd1
port 504 nsew power bidirectional
flabel metal4 s 65648 2128 65968 57712 0 FreeSans 1920 90 0 0 vccd1
port 504 nsew power bidirectional
flabel metal4 s 19568 2128 19888 57712 0 FreeSans 1920 90 0 0 vssd1
port 505 nsew ground bidirectional
flabel metal4 s 50288 2128 50608 57712 0 FreeSans 1920 90 0 0 vssd1
port 505 nsew ground bidirectional
flabel metal2 s 12346 0 12402 800 0 FreeSans 224 90 0 0 wb_clk_i
port 506 nsew signal input
flabel metal2 s 12438 0 12494 800 0 FreeSans 224 90 0 0 wb_rst_i
port 507 nsew signal input
flabel metal2 s 12530 0 12586 800 0 FreeSans 224 90 0 0 wbs_ack_o
port 508 nsew signal tristate
flabel metal2 s 12898 0 12954 800 0 FreeSans 224 90 0 0 wbs_adr_i[0]
port 509 nsew signal input
flabel metal2 s 16026 0 16082 800 0 FreeSans 224 90 0 0 wbs_adr_i[10]
port 510 nsew signal input
flabel metal2 s 16302 0 16358 800 0 FreeSans 224 90 0 0 wbs_adr_i[11]
port 511 nsew signal input
flabel metal2 s 16578 0 16634 800 0 FreeSans 224 90 0 0 wbs_adr_i[12]
port 512 nsew signal input
flabel metal2 s 16854 0 16910 800 0 FreeSans 224 90 0 0 wbs_adr_i[13]
port 513 nsew signal input
flabel metal2 s 17130 0 17186 800 0 FreeSans 224 90 0 0 wbs_adr_i[14]
port 514 nsew signal input
flabel metal2 s 17406 0 17462 800 0 FreeSans 224 90 0 0 wbs_adr_i[15]
port 515 nsew signal input
flabel metal2 s 17682 0 17738 800 0 FreeSans 224 90 0 0 wbs_adr_i[16]
port 516 nsew signal input
flabel metal2 s 17958 0 18014 800 0 FreeSans 224 90 0 0 wbs_adr_i[17]
port 517 nsew signal input
flabel metal2 s 18234 0 18290 800 0 FreeSans 224 90 0 0 wbs_adr_i[18]
port 518 nsew signal input
flabel metal2 s 18510 0 18566 800 0 FreeSans 224 90 0 0 wbs_adr_i[19]
port 519 nsew signal input
flabel metal2 s 13266 0 13322 800 0 FreeSans 224 90 0 0 wbs_adr_i[1]
port 520 nsew signal input
flabel metal2 s 18786 0 18842 800 0 FreeSans 224 90 0 0 wbs_adr_i[20]
port 521 nsew signal input
flabel metal2 s 19062 0 19118 800 0 FreeSans 224 90 0 0 wbs_adr_i[21]
port 522 nsew signal input
flabel metal2 s 19338 0 19394 800 0 FreeSans 224 90 0 0 wbs_adr_i[22]
port 523 nsew signal input
flabel metal2 s 19614 0 19670 800 0 FreeSans 224 90 0 0 wbs_adr_i[23]
port 524 nsew signal input
flabel metal2 s 19890 0 19946 800 0 FreeSans 224 90 0 0 wbs_adr_i[24]
port 525 nsew signal input
flabel metal2 s 20166 0 20222 800 0 FreeSans 224 90 0 0 wbs_adr_i[25]
port 526 nsew signal input
flabel metal2 s 20442 0 20498 800 0 FreeSans 224 90 0 0 wbs_adr_i[26]
port 527 nsew signal input
flabel metal2 s 20718 0 20774 800 0 FreeSans 224 90 0 0 wbs_adr_i[27]
port 528 nsew signal input
flabel metal2 s 20994 0 21050 800 0 FreeSans 224 90 0 0 wbs_adr_i[28]
port 529 nsew signal input
flabel metal2 s 21270 0 21326 800 0 FreeSans 224 90 0 0 wbs_adr_i[29]
port 530 nsew signal input
flabel metal2 s 13634 0 13690 800 0 FreeSans 224 90 0 0 wbs_adr_i[2]
port 531 nsew signal input
flabel metal2 s 21546 0 21602 800 0 FreeSans 224 90 0 0 wbs_adr_i[30]
port 532 nsew signal input
flabel metal2 s 21822 0 21878 800 0 FreeSans 224 90 0 0 wbs_adr_i[31]
port 533 nsew signal input
flabel metal2 s 14002 0 14058 800 0 FreeSans 224 90 0 0 wbs_adr_i[3]
port 534 nsew signal input
flabel metal2 s 14370 0 14426 800 0 FreeSans 224 90 0 0 wbs_adr_i[4]
port 535 nsew signal input
flabel metal2 s 14646 0 14702 800 0 FreeSans 224 90 0 0 wbs_adr_i[5]
port 536 nsew signal input
flabel metal2 s 14922 0 14978 800 0 FreeSans 224 90 0 0 wbs_adr_i[6]
port 537 nsew signal input
flabel metal2 s 15198 0 15254 800 0 FreeSans 224 90 0 0 wbs_adr_i[7]
port 538 nsew signal input
flabel metal2 s 15474 0 15530 800 0 FreeSans 224 90 0 0 wbs_adr_i[8]
port 539 nsew signal input
flabel metal2 s 15750 0 15806 800 0 FreeSans 224 90 0 0 wbs_adr_i[9]
port 540 nsew signal input
flabel metal2 s 12622 0 12678 800 0 FreeSans 224 90 0 0 wbs_cyc_i
port 541 nsew signal input
flabel metal2 s 12990 0 13046 800 0 FreeSans 224 90 0 0 wbs_dat_i[0]
port 542 nsew signal input
flabel metal2 s 16118 0 16174 800 0 FreeSans 224 90 0 0 wbs_dat_i[10]
port 543 nsew signal input
flabel metal2 s 16394 0 16450 800 0 FreeSans 224 90 0 0 wbs_dat_i[11]
port 544 nsew signal input
flabel metal2 s 16670 0 16726 800 0 FreeSans 224 90 0 0 wbs_dat_i[12]
port 545 nsew signal input
flabel metal2 s 16946 0 17002 800 0 FreeSans 224 90 0 0 wbs_dat_i[13]
port 546 nsew signal input
flabel metal2 s 17222 0 17278 800 0 FreeSans 224 90 0 0 wbs_dat_i[14]
port 547 nsew signal input
flabel metal2 s 17498 0 17554 800 0 FreeSans 224 90 0 0 wbs_dat_i[15]
port 548 nsew signal input
flabel metal2 s 17774 0 17830 800 0 FreeSans 224 90 0 0 wbs_dat_i[16]
port 549 nsew signal input
flabel metal2 s 18050 0 18106 800 0 FreeSans 224 90 0 0 wbs_dat_i[17]
port 550 nsew signal input
flabel metal2 s 18326 0 18382 800 0 FreeSans 224 90 0 0 wbs_dat_i[18]
port 551 nsew signal input
flabel metal2 s 18602 0 18658 800 0 FreeSans 224 90 0 0 wbs_dat_i[19]
port 552 nsew signal input
flabel metal2 s 13358 0 13414 800 0 FreeSans 224 90 0 0 wbs_dat_i[1]
port 553 nsew signal input
flabel metal2 s 18878 0 18934 800 0 FreeSans 224 90 0 0 wbs_dat_i[20]
port 554 nsew signal input
flabel metal2 s 19154 0 19210 800 0 FreeSans 224 90 0 0 wbs_dat_i[21]
port 555 nsew signal input
flabel metal2 s 19430 0 19486 800 0 FreeSans 224 90 0 0 wbs_dat_i[22]
port 556 nsew signal input
flabel metal2 s 19706 0 19762 800 0 FreeSans 224 90 0 0 wbs_dat_i[23]
port 557 nsew signal input
flabel metal2 s 19982 0 20038 800 0 FreeSans 224 90 0 0 wbs_dat_i[24]
port 558 nsew signal input
flabel metal2 s 20258 0 20314 800 0 FreeSans 224 90 0 0 wbs_dat_i[25]
port 559 nsew signal input
flabel metal2 s 20534 0 20590 800 0 FreeSans 224 90 0 0 wbs_dat_i[26]
port 560 nsew signal input
flabel metal2 s 20810 0 20866 800 0 FreeSans 224 90 0 0 wbs_dat_i[27]
port 561 nsew signal input
flabel metal2 s 21086 0 21142 800 0 FreeSans 224 90 0 0 wbs_dat_i[28]
port 562 nsew signal input
flabel metal2 s 21362 0 21418 800 0 FreeSans 224 90 0 0 wbs_dat_i[29]
port 563 nsew signal input
flabel metal2 s 13726 0 13782 800 0 FreeSans 224 90 0 0 wbs_dat_i[2]
port 564 nsew signal input
flabel metal2 s 21638 0 21694 800 0 FreeSans 224 90 0 0 wbs_dat_i[30]
port 565 nsew signal input
flabel metal2 s 21914 0 21970 800 0 FreeSans 224 90 0 0 wbs_dat_i[31]
port 566 nsew signal input
flabel metal2 s 14094 0 14150 800 0 FreeSans 224 90 0 0 wbs_dat_i[3]
port 567 nsew signal input
flabel metal2 s 14462 0 14518 800 0 FreeSans 224 90 0 0 wbs_dat_i[4]
port 568 nsew signal input
flabel metal2 s 14738 0 14794 800 0 FreeSans 224 90 0 0 wbs_dat_i[5]
port 569 nsew signal input
flabel metal2 s 15014 0 15070 800 0 FreeSans 224 90 0 0 wbs_dat_i[6]
port 570 nsew signal input
flabel metal2 s 15290 0 15346 800 0 FreeSans 224 90 0 0 wbs_dat_i[7]
port 571 nsew signal input
flabel metal2 s 15566 0 15622 800 0 FreeSans 224 90 0 0 wbs_dat_i[8]
port 572 nsew signal input
flabel metal2 s 15842 0 15898 800 0 FreeSans 224 90 0 0 wbs_dat_i[9]
port 573 nsew signal input
flabel metal2 s 13082 0 13138 800 0 FreeSans 224 90 0 0 wbs_dat_o[0]
port 574 nsew signal tristate
flabel metal2 s 16210 0 16266 800 0 FreeSans 224 90 0 0 wbs_dat_o[10]
port 575 nsew signal tristate
flabel metal2 s 16486 0 16542 800 0 FreeSans 224 90 0 0 wbs_dat_o[11]
port 576 nsew signal tristate
flabel metal2 s 16762 0 16818 800 0 FreeSans 224 90 0 0 wbs_dat_o[12]
port 577 nsew signal tristate
flabel metal2 s 17038 0 17094 800 0 FreeSans 224 90 0 0 wbs_dat_o[13]
port 578 nsew signal tristate
flabel metal2 s 17314 0 17370 800 0 FreeSans 224 90 0 0 wbs_dat_o[14]
port 579 nsew signal tristate
flabel metal2 s 17590 0 17646 800 0 FreeSans 224 90 0 0 wbs_dat_o[15]
port 580 nsew signal tristate
flabel metal2 s 17866 0 17922 800 0 FreeSans 224 90 0 0 wbs_dat_o[16]
port 581 nsew signal tristate
flabel metal2 s 18142 0 18198 800 0 FreeSans 224 90 0 0 wbs_dat_o[17]
port 582 nsew signal tristate
flabel metal2 s 18418 0 18474 800 0 FreeSans 224 90 0 0 wbs_dat_o[18]
port 583 nsew signal tristate
flabel metal2 s 18694 0 18750 800 0 FreeSans 224 90 0 0 wbs_dat_o[19]
port 584 nsew signal tristate
flabel metal2 s 13450 0 13506 800 0 FreeSans 224 90 0 0 wbs_dat_o[1]
port 585 nsew signal tristate
flabel metal2 s 18970 0 19026 800 0 FreeSans 224 90 0 0 wbs_dat_o[20]
port 586 nsew signal tristate
flabel metal2 s 19246 0 19302 800 0 FreeSans 224 90 0 0 wbs_dat_o[21]
port 587 nsew signal tristate
flabel metal2 s 19522 0 19578 800 0 FreeSans 224 90 0 0 wbs_dat_o[22]
port 588 nsew signal tristate
flabel metal2 s 19798 0 19854 800 0 FreeSans 224 90 0 0 wbs_dat_o[23]
port 589 nsew signal tristate
flabel metal2 s 20074 0 20130 800 0 FreeSans 224 90 0 0 wbs_dat_o[24]
port 590 nsew signal tristate
flabel metal2 s 20350 0 20406 800 0 FreeSans 224 90 0 0 wbs_dat_o[25]
port 591 nsew signal tristate
flabel metal2 s 20626 0 20682 800 0 FreeSans 224 90 0 0 wbs_dat_o[26]
port 592 nsew signal tristate
flabel metal2 s 20902 0 20958 800 0 FreeSans 224 90 0 0 wbs_dat_o[27]
port 593 nsew signal tristate
flabel metal2 s 21178 0 21234 800 0 FreeSans 224 90 0 0 wbs_dat_o[28]
port 594 nsew signal tristate
flabel metal2 s 21454 0 21510 800 0 FreeSans 224 90 0 0 wbs_dat_o[29]
port 595 nsew signal tristate
flabel metal2 s 13818 0 13874 800 0 FreeSans 224 90 0 0 wbs_dat_o[2]
port 596 nsew signal tristate
flabel metal2 s 21730 0 21786 800 0 FreeSans 224 90 0 0 wbs_dat_o[30]
port 597 nsew signal tristate
flabel metal2 s 22006 0 22062 800 0 FreeSans 224 90 0 0 wbs_dat_o[31]
port 598 nsew signal tristate
flabel metal2 s 14186 0 14242 800 0 FreeSans 224 90 0 0 wbs_dat_o[3]
port 599 nsew signal tristate
flabel metal2 s 14554 0 14610 800 0 FreeSans 224 90 0 0 wbs_dat_o[4]
port 600 nsew signal tristate
flabel metal2 s 14830 0 14886 800 0 FreeSans 224 90 0 0 wbs_dat_o[5]
port 601 nsew signal tristate
flabel metal2 s 15106 0 15162 800 0 FreeSans 224 90 0 0 wbs_dat_o[6]
port 602 nsew signal tristate
flabel metal2 s 15382 0 15438 800 0 FreeSans 224 90 0 0 wbs_dat_o[7]
port 603 nsew signal tristate
flabel metal2 s 15658 0 15714 800 0 FreeSans 224 90 0 0 wbs_dat_o[8]
port 604 nsew signal tristate
flabel metal2 s 15934 0 15990 800 0 FreeSans 224 90 0 0 wbs_dat_o[9]
port 605 nsew signal tristate
flabel metal2 s 13174 0 13230 800 0 FreeSans 224 90 0 0 wbs_sel_i[0]
port 606 nsew signal input
flabel metal2 s 13542 0 13598 800 0 FreeSans 224 90 0 0 wbs_sel_i[1]
port 607 nsew signal input
flabel metal2 s 13910 0 13966 800 0 FreeSans 224 90 0 0 wbs_sel_i[2]
port 608 nsew signal input
flabel metal2 s 14278 0 14334 800 0 FreeSans 224 90 0 0 wbs_sel_i[3]
port 609 nsew signal input
flabel metal2 s 12714 0 12770 800 0 FreeSans 224 90 0 0 wbs_stb_i
port 610 nsew signal input
flabel metal2 s 12806 0 12862 800 0 FreeSans 224 90 0 0 wbs_we_i
port 611 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 70000 60000
<< end >>
